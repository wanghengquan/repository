// Library - ice8chip, Cell - fabric_buf_ice8p, View - schematic
// LAST TIME SAVED: Aug 13 15:11:11 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module fabric_buf_ice8p ( f_out, f_in );
output  f_out;

input  f_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I_inv_lvt_2 ( .A(net6), .Y(f_out));
inv_lvt I_inv_lvt_1 ( .A(f_in), .Y(net6));

endmodule
// Library - io, Cell - cebdffrqn, View - schematic
// LAST TIME SAVED: Apr 27 16:16:03 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module cebdffrqn ( q, qn, ceb, clk, d, r );
output  q, qn;

input  ceb, clk, d, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I43 ( .A(so), .Y(low_s));
inv_lvt I50 ( .A(clkb), .Y(clkd));
inv_lvt Iinv_ckfb ( .A(clatb), .Y(net50));
inv_lvt I40 ( .A(r), .Y(rstb));
inv_lvt I_q_inv ( .A(qn), .Y(q));
inv_lvt I39 ( .A(net77), .Y(qn));
txgate_lvt I52 ( .in(so), .out(mi), .pp(clkb), .nn(clkd));
txgate_lvt I44 ( .in(d), .out(si), .pp(clkd), .nn(clkb));
txgate_lvt I51 ( .in(si), .out(low_s), .pp(clkb), .nn(clkd));
txgate_lvt I53 ( .in(mi), .out(qn), .pp(clkd), .nn(clkb));
nand2_lvt I290 ( .A(clk), .Y(clkb), .B(clatb));
nand2_lvt I42 ( .A(si), .Y(so), .B(rstb));
nor2_lvt INAND2_m ( .A(r), .B(mi), .Y(net77));
anor21_lvt I54 ( .A(net50), .B(clk), .Y(clatb), .C(ceb));

endmodule
// Library - io, Cell - dffrckb, View - schematic
// LAST TIME SAVED: Aug 12 13:15:42 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module dffrckb ( q, qn, clk, d, e, r );
output  q, qn;

input  clk, d, e, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



oai21x2_lvt I57 ( .A1(clk), .Y(clat), .A0(clatb), .B0(e));
nor2_lvt I48 ( .B(clat), .A(clk), .Y(clkb));
nand2_lvt I54 ( .A(rstb), .Y(qn), .B(q));
nand2_lvt I42 ( .A(si), .B(rstb), .Y(so));
txgate_lvt I59 ( .in(d), .out(si), .pp(clkb), .nn(clkd));
txgate_lvt I64 ( .in(low_s), .out(si), .pp(clkd), .nn(clkb));
txgate_lvt I62 ( .in(qn), .out(mi), .pp(clkb), .nn(clkd));
txgate_lvt I60 ( .in(so), .out(mi), .pp(clkd), .nn(clkb));
inv_lvt I55 ( .A(mi), .Y(q));
inv_lvt I50 ( .A(clkb), .Y(clkd));
inv_lvt I56 ( .A(clat), .Y(clatb));
inv_lvt I43 ( .A(so), .Y(low_s));
inv_lvt I40 ( .A(r), .Y(rstb));

endmodule
// Library - io, Cell - in_logic_v1_imp, View - schematic
// LAST TIME SAVED: Jun 24 11:06:20 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module in_logic_v1_imp ( dout0, dout1, sdo, bs_en, cbit, cbitb, ceb,
     clk, cntl, din, mode, rstio, sdi, shift, tclk, ud );
output  dout0, dout1, sdo;

input  bs_en, ceb, clk, cntl, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbitb;
input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



insel1_lvt_imp I_insel1 ( .in1(dinb), .in0(regb), .out(reg_),
     .sb({cbit1b, cbitb[0]}), .sel({cbit1, cbit[0]}), .in2(net037),
     .in3(net037));
mux2x1_hvt I_mux_mode ( .sel(mode), .in1(udd), .in0(reg_),
     .out(doutb));
mux2x1_hvt I_mux_clk ( .in1(tclk), .in0(clk), .out(ck2r0),
     .sel(bs_en));
mux2x1_hvt I_mux_data ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
mux2x1_hvt I_mux2_btw ( .in1(sdo), .in0(din), .out(net056),
     .sel(bs_en));
nand2_lvt I188 ( .A(cntl), .Y(cbit1b), .B(cbit[1]));
inv_lvt I_inv_dout0 ( .A(doutb), .Y(dout0));
inv_lvt I_inv_dout1 ( .A(udd), .Y(dout1));
inv_lvt I185 ( .A(cbit1b), .Y(cbit1));
inv_lvt I186 ( .A(dout0), .Y(net037));
inv_lvt I172 ( .A(din), .Y(dinb));
cebdffrqn I_dff0 ( .ceb(ceb), .clk(ck2r0), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff1 ( .e(ud), .clk(ck2r0), .qn(udd), .r(rstio), .q(net060),
     .d(net056));

endmodule
// Library - io, Cell - in_logic_v3_imp, View - schematic
// LAST TIME SAVED: Aug  9 13:26:43 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module in_logic_v3_imp ( dout0, dout1, sdo, sp12, bl, bs_en, ceb, clk,
     cntl, din, mode, pgate, prog, reset, rstio, sdi, shift, slfop,
     tclk, ud, vdd_cntl, wl );
output  dout0, dout1, sdo, sp12;


input  bs_en, ceb, clk, cntl, din, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
in_logic_v1_imp I_in_logic ( .ceb(ceb), .rstio(rstio), .din(din),
     .cntl(cntl), .dout1(dout1), .dout0(dout0), .shift(shift), .ud(ud),
     .clk(clk), .sdo(sdo), .sdi(sdi), .cbit({cbit[0], cbit[1]}),
     .cbitb({cbitb[0], cbitb[1]}), .tclk(tclk), .bs_en(bs_en),
     .mode(mode));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[3]), .sp12(sp12),
     .prog(prog));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - outsel1_lvt, View - schematic
// LAST TIME SAVED: Nov 22 19:11:18 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module outsel1_lvt ( out, clk, in0, in1, in2, sb, sel );
output  out;

input  clk, in0, in1, in2;

input [1:0]  sel;
input [1:0]  sb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I41 ( .A(in1), .Y(net036));
inv_lvt I40 ( .A(clk), .Y(clkb));
txgate_lvt I33 ( .in(whatever), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_lvt I_txgate1 ( .in(net036), .out(whatever), .pp(sb[0]),
     .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(whatever), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(ddr), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_lvt I38 ( .in(in2), .out(ddr), .pp(clkb), .nn(clk));
txgate_lvt I39 ( .in(in1), .out(ddr), .pp(clk), .nn(clkb));

endmodule
// Library - io, Cell - out_logic_v1, View - schematic
// LAST TIME SAVED: Aug 13 11:02:21 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module out_logic_v1 ( dout, sdo, bs_en, cbit, cbitb, ceb, clk, ddr0,
     ddr1, mode, rstio, sdi, shift, tclk, ud );
output  dout, sdo;

input  bs_en, ceb, clk, ddr0, ddr1, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



outsel1_lvt I169 ( .clk(ddrclk), .in2(udb), .sb(cbitb[1:0]),
     .sel(cbit[1:0]), .in1(net094), .in0(dinb), .out(muxob));
mux2x1_hvt I170 ( .sel(mode), .in1(udb), .in0(muxob), .out(doutb));
mux2x1_hvt I177 ( .in1(tclk), .in0(clk), .out(mux4clk), .sel(bs_en));
mux2x1_hvt I173 ( .in1(sdi), .in0(ddr0), .out(dd), .sel(shift));
mux2x1_hvt I176 ( .in1(sdo), .in0(ddr1), .out(mux4d), .sel(bs_en));
nor2_lvt I179 ( .A(mux4clk), .B(cbit[0]), .Y(ddrclk));
inv_lvt I171 ( .A(doutb), .Y(dout));
inv_lvt I172 ( .A(ddr0), .Y(dinb));
cebdffrqn I_reg0 ( .ceb(ceb), .clk(mux4clk), .qn(net094), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_reg1 ( .e(ud), .clk(mux4clk), .qn(udb), .r(rstio), .q(net44),
     .d(mux4d));

endmodule
// Library - io, Cell - out_logic_v3, View - schematic
// LAST TIME SAVED: Aug  9 13:26:57 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module out_logic_v3 ( dout, sdo, sp12, bl, bs_en, ceb, clk, ddr0, ddr1,
     mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk, ud,
     vdd_cntl, wl );
output  dout, sdo, sp12;


input  bs_en, ceb, clk, ddr0, ddr1, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;

wire  [3:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
out_logic_v1 I_outlogic_v1 ( .shift(shift), .ud(ud), .clk(clk),
     .sdo(sdo), .sdi(sdi), .ceb(ceb), .cbit({cbit[2], cbit[3]}),
     .cbitb({cbitb[2], cbitb[3]}), .dout(dout), .ddr0(ddr0),
     .tclk(tclk), .bs_en(bs_en), .rstio(rstio), .ddr1(ddr1),
     .mode(mode));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
odrv12 I_odrv12 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp12(sp12));

endmodule
// Library - io, Cell - ioesel_lvt, View - schematic
// LAST TIME SAVED: Dec  1 14:31:52 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioesel_lvt ( out, in0, in1, sb, sel );
output  out;

input  in0, in1;

input [1:0]  sb;
input [1:0]  sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I38 ( .A(sel[0]), .Y(net017));
txgate_lvt I33 ( .in(mid), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_lvt I_txgate1 ( .in(in1), .out(mid), .pp(sb[0]), .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(mid), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(net017), .out(out), .pp(sel[1]), .nn(sb[1]));

endmodule
// Library - io, Cell - ioe_logic_v1, View - schematic
// LAST TIME SAVED: Aug 13 14:52:51 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioe_logic_v1 ( outb, sdo, bs_en, cbit, cbitb, ceb, clk, din,
     mode, rstio, sdi, shift, tclk, ud );
output  outb, sdo;

input  bs_en, ceb, clk, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ioesel_lvt I_ioe_mux2 ( .sb(cbitb[1:0]), .sel(cbit[1:0]), .in1(regb),
     .in0(dinb), .out(regmuxb));
mux2x1_hvt I175 ( .in1(tclk), .in0(clk), .out(net039), .sel(bs_en));
mux2x1_hvt I170 ( .sel(mode), .in1(udd), .in0(regmuxb), .out(outb));
mux2x1_hvt I173 ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
inv_lvt I172 ( .A(din), .Y(dinb));
cebdffrqn I_dff_1 ( .ceb(ceb), .clk(net039), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff_2 ( .e(ud), .clk(net039), .qn(udd), .r(rstio), .q(net44),
     .d(sdo));

endmodule
// Library - io, Cell - ioe_logic_v3, View - schematic
// LAST TIME SAVED: Aug 12 13:29:42 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioe_logic_v3 ( padeb, sdo, sp12, bl, bs_en, ceb, clk, din,
     hiz_b, mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk,
     ud, vdd_cntl, wl );
output  padeb, sdo, sp12;


input  bs_en, ceb, clk, din, hiz_b, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbit;

wire  [3:0]  cbitb;



inv_lvt I_inv ( .A(oeb), .Y(oed));
nand2_lvt I_nand2 ( .A(oed), .Y(padeb), .B(hiz_b));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
ioe_logic_v1 I_ioe_logic ( .shift(shift), .ud(ud), .clk(clk),
     .sdo(sdo), .sdi(sdi), .cbit(cbit[3:2]), .din(din),
     .cbitb(cbitb[3:2]), .ceb(ceb), .rstio(rstio), .bs_en(bs_en),
     .tclk(tclk), .outb(oeb), .mode(mode));
odrv12 I_odrv12x2 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp12(sp12));

endmodule
// Library - leafcell, Cell - dffs, View - schematic
// LAST TIME SAVED: Dec  3 13:08:03 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module dffs ( Q, QN, CLK, D, S );
output  Q, QN;

input  CLK, D, S;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net45), .Y(net38));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net42));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net49), .Y(net42));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net49), .Y(net38));
nand2_hvt I5 ( .A(net38), .Y(net45), .B(net26));
nand2_hvt I125 ( .A(net42), .Y(net49), .B(net26));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));
inv_hvt I146 ( .A(net38), .Y(Q));
inv_hvt I147 ( .A(net45), .Y(QN));
inv_hvt I2 ( .A(S), .Y(net26));
inv_hvt I131 ( .A(CLK), .Y(clk_b));

endmodule
// Library - io, Cell - odrv12x3, View - schematic
// LAST TIME SAVED: Aug  9 13:26:19 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module odrv12x3 ( sp12, bl, pgate, prog, reset, slfop, vdd_cntl, wl );


input  prog;

output [2:0]  sp12;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  reset;
input [2:0]  slfop;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12_2_ ( .slfop(slfop[2]), .cbitb(cbitb[2]),
     .sp12(sp12[2]), .prog(prog));
odrv12 I_odrv12_1_ ( .slfop(slfop[1]), .cbitb(cbitb[1]),
     .sp12(sp12[1]), .prog(prog));
odrv12 I_odrv12_0_ ( .slfop(slfop[0]), .cbitb(cbitb[0]),
     .sp12(sp12[0]), .prog(prog));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioe_col2_v3, View - schematic
// LAST TIME SAVED: May 12 17:42:20 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioe_col2_v3 ( dout, padeb, pado, sdo, sp12_h_l, bl, bs_en, ceb,
     hiz_b, hold, inclk, mode, outclk, padin, pgate, prog, reset,
     rstio, sdi, shift, tclk, ti, update, vdd_cntl, wl );
output  sdo;


input  bs_en, ceb, hiz_b, hold, inclk, mode, outclk, prog, rstio, sdi,
     shift, tclk, update;

output [1:0]  pado;
output [23:0]  sp12_h_l;
output [3:0]  dout;
output [1:0]  padeb;

inout [1:0]  bl;

input [1:0]  padin;
input [5:0]  ti;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



in_logic_v3_imp I_in1 ( .slfop(dout[3]), .shift(shift),
     .dout1(dout[3]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[2]), .sp12(sp12_h_l[14]), .wl(wl[13:12]),
     .ceb(ceb), .reset(reset[13:12]), .sdo(s4), .sdi(s3),
     .vdd_cntl(vdd_cntl[13:12]), .pgate(pgate[13:12]), .din(padin[1]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode),
     .rstio(rstio));
in_logic_v3_imp I_in0 ( .slfop(dout[0]), .shift(shift),
     .dout1(dout[1]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[0]), .sp12(sp12_h_l[8]), .wl(wl[3:2]),
     .ceb(ceb), .reset(reset[3:2]), .sdo(s1), .sdi(s0),
     .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]), .din(padin[0]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode),
     .rstio(rstio));
out_logic_v3 I_out1 ( .shift(shift), .slfop(dout[3]), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .sp12(sp12_h_l[6]),
     .wl(wl[11:10]), .ceb(ceb), .reset(reset[11:10]), .sdo(s3),
     .sdi(s2), .vdd_cntl(vdd_cntl[11:10]), .pgate(pgate[11:10]),
     .dout(pado[1]), .tclk(tclk), .bs_en(bs_en), .rstio(rstio),
     .ddr1(ti[5]), .mode(mode), .ddr0(ti[4]));
out_logic_v3 I_out0 ( .shift(shift), .slfop(dout[0]), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .sp12(sp12_h_l[0]),
     .wl(wl[1:0]), .ceb(ceb), .reset(reset[1:0]), .sdo(s0), .sdi(sdi),
     .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]), .dout(pado[0]),
     .tclk(tclk), .bs_en(bs_en), .rstio(rstio), .ddr1(ti[2]),
     .mode(mode), .ddr0(ti[1]));
ioe_logic_v3 I_ioe0 ( .shift(shift), .hiz_b(hiz_b), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .padeb(padeb[0]),
     .slfop(dout[0]), .sp12(sp12_h_l[16]), .wl(wl[5:4]), .ceb(ceb),
     .reset(reset[5:4]), .sdo(s2), .sdi(s1), .pgate(pgate[5:4]),
     .din(ti[0]), .tclk(tclk), .vdd_cntl(vdd_cntl[5:4]), .bs_en(bs_en),
     .mode(mode), .rstio(rstio));
ioe_logic_v3 I_ioe1 ( .shift(shift), .hiz_b(hiz_b), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .padeb(padeb[1]),
     .slfop(dout[3]), .sp12(sp12_h_l[22]), .wl(wl[15:14]), .ceb(ceb),
     .reset(reset[15:14]), .sdo(sdo), .sdi(s4), .pgate(pgate[15:14]),
     .din(ti[3]), .tclk(tclk), .vdd_cntl(vdd_cntl[15:14]),
     .bs_en(bs_en), .mode(mode), .rstio(rstio));
odrv12x3 I_odrv12x3_1 ( .bl(bl[1:0]), .wl(wl[7:6]), .reset(reset[7:6]),
     .pgate(pgate[7:6]), .slfop({dout[1], dout[1], dout[1]}),
     .sp12({sp12_h_l[18], sp12_h_l[10], sp12_h_l[2]}),
     .vdd_cntl(vdd_cntl[7:6]), .prog(prog));
odrv12x3 I_odrv12x3_2 ( .bl(bl[1:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]), .slfop({dout[2], dout[2], dout[2]}),
     .sp12({sp12_h_l[20], sp12_h_l[12], sp12_h_l[4]}),
     .vdd_cntl(vdd_cntl[9:8]), .prog(prog));

endmodule
// Library - io, Cell - io_odrv4x5, View - schematic
// LAST TIME SAVED: Aug  9 13:55:12 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_odrv4x5 ( cbit, sp4_out, bl, pgate, prog,
     reset, slfop, vdd_cntl, wl );


input  prog, slfop;

output [4:0]  sp4_out;
output [7:5]  cbit;

inout [3:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
/* //////////////wire vddp_ = test.cds_globalsInst.vddp_; */ supply1 vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  cbitb;

wire  [1:0]  r_vdd;

wire [7:0] cbit_int;
assign cbit[7:5] = cbit_int[7:5];



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv4 I_odrv_4_ ( .cbitb(cbitb[4]), .sp4(sp4_out[4]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_3_ ( .cbitb(cbitb[3]), .sp4(sp4_out[3]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_2_ ( .cbitb(cbitb[2]), .sp4(sp4_out[2]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_1_ ( .cbitb(cbitb[1]), .sp4(sp4_out[1]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_0_ ( .cbitb(cbitb[0]), .sp4(sp4_out[0]), .slfop(slfop),
     .prog(prog));
cram2x2 Icram2x2_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset[1:0]), .q(cbit_int[7:4]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));
cram2x2 Icram2x2_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset[1:0]), .q(cbit_int[3:0]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - io_col_odrv4_x40bare_v3, View - schematic
// LAST TIME SAVED: Jun  2 10:03:19 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_col_odrv4_x40bare_v3 ( cf, bl, sp4_h_l,
     sp4_v_b, dout0, dout1,
     pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [23:0]  cf;

inout [3:0]  bl;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_b;

input [0:1]  dout1;
input [0:1]  dout0;
input [15:0]  wl;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
/* //////////////wire vddp_ = test.cds_globalsInst.vddp_; */ supply1 vddp_;
supply0 GND_;
supply1 VDD_;



io_odrv4x5 I_io_odrv4x5_6 ( cf[20:18], {sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6]}, bl[3:0], pgate[13:12],
     prog, reset[13:12], dout1[1], vdd_cntl[13:12], wl[13:12]);
io_odrv4x5 I_io_odrv4x5_4 ( cf[14:12], {sp4_h_l[36], sp4_h_l[28],
     sp4_h_l[20], sp4_h_l[12], sp4_h_l[4]}, bl[3:0], pgate[9:8], prog,
     reset[9:8], dout0[1], vdd_cntl[9:8], wl[9:8]);
io_odrv4x5 I_io_odrv4x5_7 ( cf[23:21], {sp4_v_b[15], sp4_v_b[11],
     sp4_v_b[7], sp4_v_b[3], sp4_h_l[46]}, bl[3:0], pgate[15:14], prog,
     reset[15:14], dout1[1], vdd_cntl[15:14], wl[15:14]);
io_odrv4x5 I_io_odrv4x5_3 ( cf[11:9], {sp4_v_b[13], sp4_v_b[9],
     sp4_v_b[5], sp4_v_b[1], sp4_h_l[42]}, bl[3:0], pgate[7:6], prog,
     reset[7:6], dout1[0], vdd_cntl[7:6], wl[7:6]);
io_odrv4x5 I_io_odrv4x5_2 ( cf[8:6], {sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2]}, bl[3:0], pgate[5:4], prog,
     reset[5:4], dout1[0], vdd_cntl[5:4], wl[5:4]);
io_odrv4x5 I_io_odrv4x5_0 ( cf[2:0], {sp4_h_l[32], sp4_h_l[24],
     sp4_h_l[16], sp4_h_l[8], sp4_h_l[0]}, bl[3:0], pgate[1:0], prog,
     reset[1:0], dout0[0], vdd_cntl[1:0], wl[1:0]);
io_odrv4x5 I_io_odrv4x5_1 ( cf[5:3], {sp4_v_b[12], sp4_v_b[8],
     sp4_v_b[4], sp4_v_b[0], sp4_h_l[40]}, bl[3:0], pgate[3:2], prog,
     reset[3:2], dout0[0], vdd_cntl[3:2], wl[3:2]);
io_odrv4x5 I_io_odrv4x5_5 ( cf[17:15], {sp4_v_b[14], sp4_v_b[10],
     sp4_v_b[6], sp4_v_b[2], sp4_h_l[44]}, bl[3:0], pgate[11:10], prog,
     reset[11:10], dout0[1], vdd_cntl[11:10], wl[11:10]);

endmodule
// Library - ice8chip, Cell - io_col4_rgt_ice8p_v2, View - schematic
// LAST TIME SAVED: Jan 12 14:59:31 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_col4_rgt_ice8p_v2 ( cbit_colcntl, cf, fabric_out, padeb,
     pado, sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t,
     sp12_h_l, bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold,
     lft_op, mode, padin, pgate, prog, r, reset, sdi, shift, spioeb,
     spiout, tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [23:0]  cf;
output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;
output [7:0]  cbit_colcntl;

inout [15:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;
inout [15:0]  sp4_v_t;
inout [23:0]  sp12_h_l;

input [1:0]  spioeb;
input [1:0]  spiout;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [15:0]  wl;
input [15:0]  reset;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [7:0]  glb_netwk;
input [1:0]  padin;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



rm7w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
sbox1_colbdlc_v4 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_gmux_x16bare_v4 I_io_gmux_x16bare_v4 (
     .cbit_colcntl(cbit_colcntl[7:0]), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});

endmodule
// Library - ice8chip, Cell - tckbufx32_ice8p, View - schematic
// LAST TIME SAVED: Aug 13 15:04:42 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module tckbufx32_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I_inv_lvt_1 ( .A(in), .Y(net4));
inv_lvt Iinv_lvt_2 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - tielo4x, View - schematic
// LAST TIME SAVED: May 18 10:31:28 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module tielo4x ( tielo );
output  tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - tiehi4x, View - schematic
// LAST TIME SAVED: May 18 10:33:00 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module tiehi4x ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - ice1chip, Cell - io_rgt_top_1x8_ice1f, View - schematic
// LAST TIME SAVED: Mar  4 20:34:44 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_rgt_top_1x8_ice1f ( cf_r, fabric_out_09, fabric_out_10,
     padeb, pado, sdo, slf_op_01, slf_op_02, slf_op_03, slf_op_04,
     slf_op_05, slf_op_06, slf_op_07, slf_op_08, tclk_o, SP4_h_l_01,
     SP4_h_l_02, SP4_h_l_03, SP4_h_l_04, SP4_h_l_05, SP4_h_l_06,
     SP4_h_l_07, SP4_h_l_08, SP12_h_l_01, SP12_h_l_02, SP12_h_l_03,
     SP12_h_l_04, SP12_h_l_05, SP12_h_l_06, SP12_h_l_07, SP12_h_l_08,
     bl, pgate, reset_b, sp4_v_b_13_09, sp4_v_t_08, vdd_cntl, wl,
     bnl_op_13_09, bs_en, ceb, glb_netwk_col, hiz_b, hold, lft_op_01,
     lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06, lft_op_07,
     lft_op_08, mode, padin, prog, r, sdi, shift, tclk, tnl_op_08,
     update );
output  fabric_out_09, fabric_out_10, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_03;
output [3:0]  slf_op_08;
output [3:0]  slf_op_06;
output [3:0]  slf_op_02;
output [24:13]  padeb;
output [24:13]  pado;
output [3:0]  slf_op_05;
output [3:0]  slf_op_07;
output [3:0]  slf_op_04;
output [191:0]  cf_r;
output [3:0]  slf_op_01;

inout [23:0]  SP12_h_l_08;
inout [47:0]  SP4_h_l_07;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_01;
inout [23:0]  SP12_h_l_03;
inout [23:0]  SP12_h_l_02;
inout [47:0]  SP4_h_l_03;
inout [15:0]  sp4_v_t_08;
inout [47:0]  SP4_h_l_02;
inout [127:0]  vdd_cntl;
inout [127:0]  reset_b;
inout [127:0]  pgate;
inout [23:0]  SP12_h_l_06;
inout [23:0]  SP12_h_l_01;
inout [23:0]  SP12_h_l_07;
inout [47:0]  SP4_h_l_04;
inout [23:0]  SP12_h_l_04;
inout [127:0]  wl;
inout [47:0]  SP4_h_l_08;
inout [47:0]  SP4_h_l_06;
inout [23:0]  SP12_h_l_05;
inout [15:0]  sp4_v_b_13_09;
inout [47:0]  SP4_h_l_05;

input [7:0]  lft_op_07;
input [7:0]  lft_op_02;
input [7:0]  bnl_op_13_09;
input [7:0]  tnl_op_08;
input [24:13]  padin;
input [7:0]  lft_op_03;
input [7:0]  lft_op_01;
input [7:0]  lft_op_05;
input [7:0]  lft_op_08;
input [7:0]  lft_op_04;
input [7:0]  glb_netwk_col;
input [7:0]  lft_op_06;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net632;

wire  [0:15]  net478;

wire  [7:0]  colbuf_cntl_t;

wire  [7:0]  colbuf_cntl_b;

wire  [7:0]  glb_netwk_b;

wire  [7:0]  glb_netwk_t;

wire  [0:15]  net586;

wire  [0:1]  net618;

wire  [0:1]  net630;

wire  [0:15]  net442;

wire  [0:7]  net633;

wire  [0:7]  net317;

wire  [0:7]  net461;

wire  [0:1]  net590;

wire  [0:1]  net624;

wire  [0:7]  net497;

wire  [0:1]  net625;

wire  [0:1]  net620;

wire  [0:15]  net370;

wire  [0:1]  net628;

wire  [0:1]  net476;

wire  [0:7]  net623;

wire  [0:1]  net616;

wire  [0:15]  net514;

wire  [0:1]  net477;

wire  [0:1]  net332;

wire  [0:1]  net629;

wire  [0:15]  net550;

wire  [0:15]  net406;



io_col4_rgt_ice8p_v2 I_io_00_08 ( .cbit_colcntl(net317[0:7]),
     .ceb(ceb), .sdo(sdo), .sdi(net355), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(net332[0:1]), .pado(net332[0:1]),
     .padeb(net616[0:1]), .sp4_v_t(sp4_v_t_08[15:0]),
     .sp4_h_l(SP4_h_l_08[47:0]), .sp12_h_l(SP12_h_l_08[23:0]),
     .prog(prog), .spi_ss_in_b(net628[0:1]), .tnl_op(tnl_op_08[7:0]),
     .lft_op(lft_op_08[7:0]), .bnl_op(lft_op_07[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net370[0:15]), .wl(wl[127:112]), .cf(cf_r[191:168]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_08[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net352));
io_col4_rgt_ice8p_v2 I_io_00_07 ( .cbit_colcntl(net632[0:7]),
     .ceb(ceb), .sdo(net355), .sdi(net427), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[24:23]), .pado(pado[24:23]),
     .padeb(padeb[24:23]), .sp4_v_t(net370[0:15]),
     .sp4_h_l(SP4_h_l_07[47:0]), .sp12_h_l(SP12_h_l_07[23:0]),
     .prog(prog), .spi_ss_in_b(net629[0:1]), .tnl_op(lft_op_08[7:0]),
     .lft_op(lft_op_07[7:0]), .bnl_op(lft_op_06[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net442[0:15]), .wl(wl[111:96]), .cf(cf_r[167:144]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_07[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net388));
io_col4_rgt_ice8p_v2 I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net391), .sdi(net571), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[20:19]), .pado(pado[20:19]),
     .padeb(padeb[20:19]), .sp4_v_t(net406[0:15]),
     .sp4_h_l(SP4_h_l_05[47:0]), .sp12_h_l(SP12_h_l_05[23:0]),
     .prog(prog), .spi_ss_in_b(net618[0:1]), .tnl_op(lft_op_06[7:0]),
     .lft_op(lft_op_05[7:0]), .bnl_op(lft_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net586[0:15]), .wl(wl[79:64]), .cf(cf_r[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net424));
io_col4_rgt_ice8p_v2 I_io_00_06 ( .cbit_colcntl(net633[0:7]),
     .ceb(ceb), .sdo(net427), .sdi(net391), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[22:21]), .pado(pado[22:21]),
     .padeb(padeb[22:21]), .sp4_v_t(net442[0:15]),
     .sp4_h_l(SP4_h_l_06[47:0]), .sp12_h_l(SP12_h_l_06[23:0]),
     .prog(prog), .spi_ss_in_b(net625[0:1]), .tnl_op(lft_op_07[7:0]),
     .lft_op(lft_op_06[7:0]), .bnl_op(lft_op_05[7:0]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net406[0:15]), .wl(wl[95:80]), .cf(cf_r[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net460));
io_col4_rgt_ice8p_v2 I_io_00_02 ( .cbit_colcntl(net461[0:7]),
     .ceb(ceb), .sdo(net463), .sdi(net499), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(net476[0:1]), .pado(net476[0:1]),
     .padeb(net477[0:1]), .sp4_v_t(net478[0:15]),
     .sp4_h_l(SP4_h_l_02[47:0]), .sp12_h_l(SP12_h_l_02[23:0]),
     .prog(prog), .spi_ss_in_b(net630[0:1]), .tnl_op(lft_op_03[7:0]),
     .lft_op(lft_op_02[7:0]), .bnl_op(lft_op_01[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(net514[0:15]), .wl(wl[31:16]), .cf(cf_r[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_10));
io_col4_rgt_ice8p_v2 I_io_00_01 ( .cbit_colcntl(net497[0:7]),
     .ceb(ceb), .sdo(net499), .sdi(sdi), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[14:13]), .pado(pado[14:13]),
     .padeb(padeb[14:13]), .sp4_v_t(net514[0:15]),
     .sp4_h_l(SP4_h_l_01[47:0]), .sp12_h_l(SP12_h_l_01[23:0]),
     .prog(prog), .spi_ss_in_b(net620[0:1]), .tnl_op(lft_op_02[7:0]),
     .lft_op(lft_op_01[7:0]), .bnl_op(bnl_op_13_09[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_v_b_13_09[15:0]), .wl(wl[15:0]), .cf(cf_r[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_09));
io_col4_rgt_ice8p_v2 I_io_00_03 ( .cbit_colcntl(net623[0:7]),
     .ceb(ceb), .sdo(net535), .sdi(net463), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[16:15]), .pado(pado[16:15]),
     .padeb(padeb[16:15]), .sp4_v_t(net550[0:15]),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b(net624[0:1]), .tnl_op(lft_op_04[7:0]),
     .lft_op(lft_op_03[7:0]), .bnl_op(lft_op_02[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net478[0:15]), .wl(wl[47:32]), .cf(cf_r[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net568));
io_col4_rgt_ice8p_v2 I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net571), .sdi(net535), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[18:17]), .pado(pado[18:17]),
     .padeb(padeb[18:17]), .sp4_v_t(net586[0:15]),
     .sp4_h_l(SP4_h_l_04[47:0]), .sp12_h_l(SP12_h_l_04[23:0]),
     .prog(prog), .spi_ss_in_b(net590[0:1]), .tnl_op(lft_op_05[7:0]),
     .lft_op(lft_op_04[7:0]), .bnl_op(lft_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net550[0:15]), .wl(wl[63:48]), .cf(cf_r[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net604));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - bram_bufferx4x6, View - schematic
// LAST TIME SAVED: Sep 15 13:53:57 2008
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_bufferx4x6 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I4 ( .in(d1), .out(d2));
bram_bufferx4 I5 ( .in(d2), .out(d3));
bram_bufferx4 I6 ( .in(d3), .out(d4));
bram_bufferx4 I7 ( .in(d4), .out(out));
bram_bufferx4 I3 ( .in(d0), .out(d1));
bram_bufferx4 I0 ( .in(in), .out(d0));

endmodule
// Library - leafcell, Cell - pllphase_sr_40lp, View - schematic
// LAST TIME SAVED: Jun  6 17:32:49 2011
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pllphase_sr_40lp ( f_dvd2, f_dvd4_p0, f_dvd4_p90, f_out, CLK,
     cbit, sr, tiehi, tielo );
output  f_dvd2, f_dvd4_p0, f_dvd4_p90, f_out;

input  CLK, cbit, sr, tiehi, tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  qn;



mux2_hvt I_MUX4DIV7 ( .in1(net077), .in0(net051), .out(net038),
     .sel(cbit));
inv_tri_2_hvt I21 ( .Tb(net0136), .T(net0136), .A(net0136),
     .Y(net0113));
nor2_hvt I22 ( .A(net0113), .B(tielo), .Y(net0116));
inv_hvt I26 ( .A(net089), .Y(net086));
inv_hvt I27 ( .A(CLK), .Y(net089));
inv_hvt I23 ( .A(net0116), .Y(net044));
inv_hvt I20 ( .A(net0138), .Y(net0136));
inv_hvt I19 ( .A(net0101), .Y(net0138));
inv_hvt I28 ( .A(net086), .Y(net057));
inv_hvt I29 ( .A(net057), .Y(net080));
inv_hvt I30 ( .A(net080), .Y(net088));
inv_hvt I31 ( .A(net088), .Y(net0101));
inv_hvt I8 ( .A(qn[1]), .Y(f_dvd4_p90));
inv_hvt I7 ( .A(net0100), .Y(f_dvd2));
inv_hvt I6 ( .A(net044), .Y(f_out));
inv_hvt I5 ( .A(qn[0]), .Y(f_dvd4_p0));
pll_ml_dff I2 ( .R(sr), .D(net056), .CLK(CLK), .QN(qn[1]), .Q(net051));
pll_ml_dff I0 ( .R(sr), .D(net054), .CLK(CLK), .QN(qn[0]), .Q(net056));
pll_ml_dff I3 ( .R(sr), .D(net051), .CLK(CLK), .QN(net061),
     .Q(net040));
pll_ml_dff I12 ( .R(sr), .D(net0100), .CLK(CLK), .QN(net0100),
     .Q(net067));
dffs I10 ( .D(net082), .QN(net071), .Q(net054), .CLK(CLK), .S(sr));
dffs I9 ( .D(net053), .QN(net076), .Q(net077), .CLK(CLK), .S(sr));
dffs I11 ( .D(net038), .QN(net081), .Q(net082), .CLK(CLK), .S(sr));
dffs I4 ( .D(net040), .CLK(CLK), .QN(net087), .Q(net053), .S(sr));

endmodule
// Library - leafcell, Cell - lowla_modified, View - schematic
// LAST TIME SAVED: Aug 12 09:10:07 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module lowla_modified ( lao, clk, min );
output  lao;

input  clk, min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I249 ( .in(lao), .out(st2), .pp(cbitb), .nn(clkd));
txgate_hvt I248 ( .in(min), .out(st2), .pp(clkd), .nn(cbitb));
inv_hvt I289 ( .A(net29), .Y(lao));
inv_hvt I290 ( .A(st2), .Y(net29));
inv_hvt I_inv ( .A(clk), .Y(cbitb));
inv_hvt I_inv3 ( .A(cbitb), .Y(clkd));

endmodule
// Library - ice8chip, Cell - scan_buf_ice8p, View - schematic
// LAST TIME SAVED: Jun 28 09:23:39 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module scan_buf_ice8p ( bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo,
     shift_o, tclk_o, update_o, bs_en_i, ceb_i, hiz_b_i, mode_i, r_i,
     sdi, shift_i, tclk_i, update_i );
output  bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo, shift_o, tclk_o,
     update_o;

input  bs_en_i, ceb_i, hiz_b_i, mode_i, r_i, sdi, shift_i, tclk_i,
     update_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



tckbufx32_ice8p I_tclkbuf ( .in(tclk_i), .out(tclk_o));
bram_bufferx4 I_bs_enbuf ( .in(bs_en_i), .out(bs_en_o));
bram_bufferx4 I_cebbuf ( .in(ceb_i), .out(ceb_o));
bram_bufferx4 I_modebuf ( .in(mode_i), .out(mode_o));
bram_bufferx4 I_hiz_bbuf ( .in(hiz_b_i), .out(hiz_b_o));
bram_bufferx4 I_updatebuf ( .in(update_i), .out(update_o));
bram_bufferx4 I_shiftbuf ( .in(shift_i), .out(shift_o));
bram_bufferx4 I_rbuf ( .in(r_i), .out(r_o));
bram_bufferx4x6 I_sdibuf ( .in(sdi), .out(sdi_2));
lowla_modified I_lowla ( .clk(tclk_i), .min(sdi_2), .lao(sdo));

endmodule
// Library - io, Cell - ioinmx1mux2_imp, View - schematic
// LAST TIME SAVED: Aug 13 14:11:56 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioinmx1mux2_imp ( clk, mo, ti, bl, cdone_in, ce, ceb, in, min,
     pgate, prog, reset, spi, vdd_cntl, wl );
output  clk, ti;


input  cdone_in, ceb, prog;

output [1:0]  mo;

inout [5:0]  bl;

input [1:0]  spi;
input [11:0]  ce;
input [1:0]  in;
input [7:0]  min;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  moo;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  mob;

wire  [1:0]  r_vdd;



mux2x1_hvt I_emux_1_ ( .in1(in[1]), .in0(spi[1]), .out(moo[1]),
     .sel(cdone_in));
mux2x1_hvt I_emux_0_ ( .in1(in[0]), .in0(spi[0]), .out(moo[0]),
     .sel(cdone_in));
inv_lvt inv_1_1_ ( .A(moo[1]), .Y(mob[1]));
inv_lvt inv_1_0_ ( .A(moo[0]), .Y(mob[0]));
inv_lvt I_inv_2_1_ ( .A(mob[1]), .Y(mo[1]));
inv_lvt I_inv_2_0_ ( .A(mob[0]), .Y(mo[0]));
ioin_mux_v2 I_ioin_mux ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clk_mux12to1 I_clk_mux12to1 ( .prog(prog), .min(ce[11:0]), .clk(clk),
     .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7], cbitb[10],
     cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7], cbit[10],
     cbit[6], cbit[4]}), .cenb(ceb));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc, View - schematic
// LAST TIME SAVED: Aug 12 13:51:42 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  spi;
output [1:0]  ti;

inout [5:0]  bl;

input [7:0]  min1;
input [7:0]  min0;
input [1:0]  padin;
input [1:0]  pgate;
input [7:0]  min2;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



inv_lvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_lvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
nor2_lvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_lvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
ioin_mux_v2 I_ioin_mux_bankcntl ( bankcntl, {cbit[11], cbit[8], cbit[9],
     cbit[10]}, {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0],
     prog);
ioin_mux_v2 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v2 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nand2inv, View - schematic
// LAST TIME SAVED: Oct  8 16:13:18 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioinmx2nand2inv ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [7:0]  min0;
input [7:0]  ce;
input [1:0]  reset;
input [1:0]  wl;
input [7:0]  min1;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



nand2_lvt I180 ( .A(update_b), .Y(updt), .B(bs_en));
inv_lvt I181 ( .A(update), .Y(update_b));
ioin_mux_v2 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v2 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc_v3, View - schematic
// LAST TIME SAVED: May 12 17:30:59 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox1_colbdlc_v3 ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  spi_ss_in_b;
output [1:0]  padeb;
output [5:0]  ti;
output [1:0]  pado;

inout [5:0]  bl;
inout [3:0]  t_mid;
inout [3:0]  sp4_v_b;
inout [3:0]  l;
inout [3:0]  r;

input [1:0]  out;
input [1:0]  padin;
input [11:0]  clk_in;
input [7:0]  min5;
input [1:0]  spiout;
input [7:0]  ceb_in;
input [7:0]  min4;
input [11:0]  inclk_in;
input [7:0]  min2;
input [1:0]  oeb;
input [7:0]  min1;
input [1:0]  spioeb;
input [7:0]  min3;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  min0;
input [7:0]  min6;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ioinmx1mux2_imp I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .in(out[1:0]), .ti(ti[2]), .min(min2[7:0]), .spi(spiout[1:0]),
     .wl(wl[9:8]), .reset(reset[9:8]), .pgate(pgate[9:8]),
     .cdone_in(cdone_in), .mo(pado[1:0]));
ioinmx1mux2_imp I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .in(oeb[1:0]), .ti(ti[5]), .min(min5[7:0]), .spi(spioeb[1:0]),
     .wl(wl[15:14]), .reset(reset[15:14]), .pgate(pgate[15:14]),
     .cdone_in(cdone_in), .mo(padeb[1:0]));
ioinmx2nor2invx2bdlc I5 ( .vdd_cntl(vdd_cntl[5:4]), .min2(min6[7:0]),
     .bankcntl(fabric_out), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx2nand2inv I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - io, Cell - io_gmux_x2v2, View - schematic
// LAST TIME SAVED: Jun  1 11:08:17 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_gmux_x2v2 ( .cbitb_colcntl({cbitb[11], cbitb[9]}), gout, bl,
     min0, min1, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [1:0]  gout;
output [11:0]  cbitb;

inout [5:0]  bl;

input [15:0]  min0;
input [1:0]  vdd_cntl;
input [15:0]  min1;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux I_g_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux I_g_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare_v3, View - schematic
// LAST TIME SAVED: Jun  2 10:52:40 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_gmux_x16bare_v3 ( cbitb_colcntl, lc_trk_g0, lc_trk_g1, bl,
     min0, min1, min2, min3, min4, min5, min6, min7, min8, min9, min10,
     min11, min12, min13, min14, min15, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  cbitb_colcntl;

inout [5:0]  bl;

input [15:0]  min7;
input [15:0]  min0;
input [15:0]  min9;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min15;
input [15:0]  min3;
input [15:0]  min14;
input [15:0]  min12;
input [15:0]  min6;
input [15:0]  min8;
input [15:0]  min5;
input [15:0]  min4;
input [15:0]  min11;
input [15:0]  min10;
input [15:0]  vdd_cntl;
input [15:0]  min2;
input [15:0]  reset;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net114;

wire  [0:1]  net187;

wire  [0:1]  net188;

wire  [0:1]  net124;



io_gmux_x2v2 I_io_gmux_x2_7 ( .cbitb_colcntl(net114[0:1]),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[15:14]));
io_gmux_x2v2 I_io_gmux_x2_6 ( .cbitb_colcntl(net124[0:1]),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[13:12]));
io_gmux_x2v2 I_io_gmux_x2_2 ( .cbitb_colcntl(cbitb_colcntl[5:4]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[5:4]));
io_gmux_x2v2 I_io_gmux_x2_0 ( .cbitb_colcntl(cbitb_colcntl[1:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[1:0]));
io_gmux_x2v2 _io_gmux_x2_1 ( .cbitb_colcntl(cbitb_colcntl[3:2]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[3:2]));
io_gmux_x2v2 I_io_gmux_x2_4 ( .cbitb_colcntl(net187[0:1]),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[9:8]));
io_gmux_x2v2 I_io_gmux_x2_5 ( .cbitb_colcntl(net188[0:1]),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[11:10]));
io_gmux_x2v2 I_io_gmux_x2_3 ( .cbitb_colcntl(cbitb_colcntl[7:6]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[7:6]));

endmodule
// Library - ice8chip, Cell - io_col4_top_ice8p, View - schematic
// LAST TIME SAVED: Jan 12 15:49:45 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_col4_top_ice8p ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  padeb;
output [1:0]  pado;
output [23:0]  cf;
output [3:0]  slf_op;
output [1:0]  spi_ss_in_b;

inout [15:0]  sp4_v_t;
inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [15:0]  sp4_v_b;
inout [47:0]  sp4_h_l;

input [1:0]  spioeb;
input [15:0]  wl;
input [7:0]  lft_op;
input [15:0]  reset;
input [1:0]  spiout;
input [15:0]  vdd_cntl;
input [7:0]  bnl_op;
input [15:0]  pgate;
input [7:0]  tnl_op;
input [1:0]  padin;
input [7:0]  glb_netwk;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  ti;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  om;

wire  [1:0]  oenm;

wire  [0:7]  net0100;



rm6w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
sbox1_colbdlc_v3 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
io_gmux_x16bare_v3 I_io_gmux_x16bare_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .cbitb_colcntl(net0100[0:7]), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29],
     sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13],
     sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5],
     tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));

endmodule
// Library - ice1chip, Cell - io_top_rgt_1x6_ice1f, View - schematic
// LAST TIME SAVED: Mar  8 10:17:00 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_top_rgt_1x6_ice1f ( bs_en_o, ceb_o, cf_t, fabric_out_07_17,
     fabric_out_08_17, hiz_b_o, mode_o, padeb_t_r, pado_t_r, r_o, sdo,
     shift_o, slf_op_01_17, slf_op_02_17, slf_op_03_17, slf_op_04_17,
     slf_op_05_17, slf_op_06_17, tclk_o, update_o, bl_01, bl_02, bl_03,
     bl_04, bl_05, bl_06, sp4_h_l_07_17, sp4_h_r_12_17, sp4_v_b_01_17,
     sp4_v_b_02_17, sp4_v_b_03_17, sp4_v_b_04_17, sp4_v_b_05_17,
     sp4_v_b_06_17, sp12_v_b_01_17, sp12_v_b_02_17, sp12_v_b_03_17,
     sp12_v_b_04_17, sp12_v_b_05_17, sp12_v_b_06_17, bnl_op_07_17,
     bnr_op_12_17, bs_en_i, ceb_i, glb_net_01, glb_net_02, glb_net_03,
     glb_net_04, glb_net_05, glb_net_06, hiz_b_i, hold_t_r,
     lft_op_01_17, lft_op_02_17, lft_op_03_17, lft_op_04_17,
     lft_op_05_17, lft_op_06_17, mode_i, padin_t_r, pgate_l, prog, r_i,
     reset_l, sdi, shift_i, tclk_i, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_07_17, fabric_out_08_17, hiz_b_o,
     mode_o, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_r, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_02_17;
output [3:0]  slf_op_06_17;
output [3:0]  slf_op_03_17;
output [143:0]  cf_t;
output [23:12]  padeb_t_r;
output [23:12]  pado_t_r;
output [3:0]  slf_op_04_17;
output [3:0]  slf_op_01_17;
output [3:0]  slf_op_05_17;

inout [47:0]  sp4_v_b_06_17;
inout [23:0]  sp12_v_b_06_17;
inout [23:0]  sp12_v_b_05_17;
inout [47:0]  sp4_v_b_05_17;
inout [47:0]  sp4_v_b_03_17;
inout [47:0]  sp4_v_b_01_17;
inout [23:0]  sp12_v_b_03_17;
inout [47:0]  sp4_v_b_02_17;
inout [47:0]  sp4_v_b_04_17;
inout [15:0]  sp4_h_l_07_17;
inout [23:0]  sp12_v_b_04_17;
inout [53:0]  bl_05;
inout [53:0]  bl_06;
inout [23:0]  sp12_v_b_02_17;
inout [41:0]  bl_04;
inout [53:0]  bl_03;
inout [15:0]  sp4_h_r_12_17;
inout [53:0]  bl_02;
inout [53:0]  bl_01;
inout [23:0]  sp12_v_b_01_17;

input [7:0]  bnr_op_12_17;
input [7:0]  glb_net_03;
input [7:0]  glb_net_01;
input [7:0]  lft_op_05_17;
input [7:0]  bnl_op_07_17;
input [7:0]  lft_op_03_17;
input [7:0]  lft_op_04_17;
input [7:0]  glb_net_06;
input [7:0]  lft_op_06_17;
input [7:0]  glb_net_02;
input [7:0]  glb_net_04;
input [23:12]  padin_t_r;
input [7:0]  lft_op_01_17;
input [15:0]  reset_l;
input [15:0]  wl_l;
input [7:0]  lft_op_02_17;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_05;
input [15:0]  pgate_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net433;

wire  [0:1]  net472;

wire  [0:15]  net363;

wire  [0:1]  net290;

wire  [0:15]  net503;

wire  [0:1]  net507;

wire  [0:15]  net328;

wire  [0:15]  net398;

wire  [0:1]  net402;

wire  [0:1]  net332;

wire  [0:1]  net289;



tckbufx32_ice8p I_tck_halfbankcenter ( .in(net273), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));
scan_buf_ice8p I345 ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net273), .shift_o(shift_o),
     .sdo(net453), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_top_ice8p I_IO_08_17 ( .sdo(net383), .sdi(net313),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net398[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_r[15:14]),
     .pado(pado_t_r[15:14]), .padeb(padeb_t_r[15:14]),
     .sp4_v_b(net328[0:15]), .sp4_h_l(sp4_v_b_02_17[47:0]),
     .sp12_h_l(sp12_v_b_02_17[23:0]), .prog(prog),
     .spi_ss_in_b(net332[0:1]), .tnl_op(lft_op_01_17[7:0]),
     .lft_op(lft_op_02_17[7:0]), .bnl_op(lft_op_03_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_02[5],
     bl_02[4], bl_02[37], bl_02[36], bl_02[35], bl_02[34], bl_02[33],
     bl_02[32], bl_02[14], bl_02[20], bl_02[19], bl_02[18], bl_02[17],
     bl_02[16], bl_02[27], bl_02[26], bl_02[25], bl_02[23]}),
     .wl(wl_l[15:0]), .cf(cf_t[47:24]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_02_17[3:0]),
     .glb_netwk(glb_net_02[7:0]), .hold(hold_t_r),
     .fabric_out(fabric_out_08_17));
io_col4_top_ice8p I_IO_10_17_bram ( .sdo(net488), .sdi(net348),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net503[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_r[19:18]),
     .pado(pado_t_r[19:18]), .padeb(padeb_t_r[19:18]),
     .sp4_v_b(net363[0:15]), .sp4_h_l(sp4_v_b_04_17[47:0]),
     .sp12_h_l(sp12_v_b_04_17[23:0]), .prog(prog),
     .spi_ss_in_b(net289[0:1]), .tnl_op(lft_op_03_17[7:0]),
     .lft_op(lft_op_04_17[7:0]), .bnl_op(lft_op_05_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_04[5],
     bl_04[4], bl_04[37], bl_04[36], bl_04[35], bl_04[34], bl_04[33],
     bl_04[32], bl_04[14], bl_04[20], bl_04[19], bl_04[18], bl_04[17],
     bl_04[16], bl_04[27], bl_04[26], bl_04[25], bl_04[23]}),
     .wl(wl_l[15:0]), .cf(cf_t[71:48]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_04_17[3:0]),
     .glb_netwk(glb_net_04[7:0]), .hold(hold_t_r),
     .fabric_out(net381));
io_col4_top_ice8p I_IO_07_17 ( .sdo(sdo), .sdi(net383),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_07_17[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_r[13:12]),
     .pado(pado_t_r[13:12]), .padeb(padeb_t_r[13:12]),
     .sp4_v_b(net398[0:15]), .sp4_h_l(sp4_v_b_01_17[47:0]),
     .sp12_h_l(sp12_v_b_01_17[23:0]), .prog(prog),
     .spi_ss_in_b(net402[0:1]), .tnl_op(bnl_op_07_17[7:0]),
     .lft_op(lft_op_01_17[7:0]), .bnl_op(lft_op_02_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_01[5],
     bl_01[4], bl_01[37], bl_01[36], bl_01[35], bl_01[34], bl_01[33],
     bl_01[32], bl_01[14], bl_01[20], bl_01[19], bl_01[18], bl_01[17],
     bl_01[16], bl_01[27], bl_01[26], bl_01[25], bl_01[23]}),
     .wl(wl_l[15:0]), .cf(cf_t[23:0]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_01_17[3:0]),
     .glb_netwk(glb_net_01[7:0]), .hold(hold_t_r),
     .fabric_out(fabric_out_07_17));
io_col4_top_ice8p I_IO_11_17 ( .sdo(net348), .sdi(net418),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net363[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_r[21:20]),
     .pado(pado_t_r[21:20]), .padeb(padeb_t_r[21:20]),
     .sp4_v_b(net433[0:15]), .sp4_h_l(sp4_v_b_05_17[47:0]),
     .sp12_h_l(sp12_v_b_05_17[23:0]), .prog(prog),
     .spi_ss_in_b(net290[0:1]), .tnl_op(lft_op_04_17[7:0]),
     .lft_op(lft_op_05_17[7:0]), .bnl_op(lft_op_06_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_05[5],
     bl_05[4], bl_05[37], bl_05[36], bl_05[35], bl_05[34], bl_05[33],
     bl_05[32], bl_05[14], bl_05[20], bl_05[19], bl_05[18], bl_05[17],
     bl_05[16], bl_05[27], bl_05[26], bl_05[25], bl_05[23]}),
     .wl(wl_l[15:0]), .cf(cf_t[119:96]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_05_17[3:0]),
     .glb_netwk(glb_net_05[7:0]), .hold(hold_t_r),
     .fabric_out(net451));
io_col4_top_ice8p I_IO_12_17 ( .sdo(net418), .sdi(net453),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net433[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_r[23:22]),
     .pado(pado_t_r[23:22]), .padeb(padeb_t_r[23:22]),
     .sp4_v_b(sp4_h_r_12_17[15:0]), .sp4_h_l(sp4_v_b_06_17[47:0]),
     .sp12_h_l(sp12_v_b_06_17[23:0]), .prog(prog),
     .spi_ss_in_b(net472[0:1]), .tnl_op(lft_op_05_17[7:0]),
     .lft_op(lft_op_06_17[7:0]), .bnl_op(bnr_op_12_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_l[15:0]), .cf(cf_t[143:120]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_06_17[3:0]),
     .glb_netwk(glb_net_06[7:0]), .hold(hold_t_r),
     .fabric_out(net486));
io_col4_top_ice8p I_IO_09_17 ( .sdo(net313), .sdi(net488),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net328[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_r[17:16]),
     .pado(pado_t_r[17:16]), .padeb(padeb_t_r[17:16]),
     .sp4_v_b(net503[0:15]), .sp4_h_l(sp4_v_b_03_17[47:0]),
     .sp12_h_l(sp12_v_b_03_17[23:0]), .prog(prog),
     .spi_ss_in_b(net507[0:1]), .tnl_op(lft_op_02_17[7:0]),
     .lft_op(lft_op_03_17[7:0]), .bnl_op(lft_op_04_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_03[5],
     bl_03[4], bl_03[37], bl_03[36], bl_03[35], bl_03[34], bl_03[33],
     bl_03[32], bl_03[14], bl_03[20], bl_03[19], bl_03[18], bl_03[17],
     bl_03[16], bl_03[27], bl_03[26], bl_03[25], bl_03[23]}),
     .wl(wl_l[15:0]), .cf(cf_t[95:72]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_03_17[3:0]),
     .glb_netwk(glb_net_03[7:0]), .hold(hold_t_r),
     .fabric_out(net521));

endmodule
// Library - leafcell, Cell - clkmux2buffer, View - schematic
// LAST TIME SAVED: Jun 29 15:54:22 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module clkmux2buffer ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate Itg20 ( .in(in1), .out(net16), .pp(net10), .nn(sel));
txgate I31 ( .in(in0), .out(net16), .pp(sel), .nn(net10));
inv I_inv1 ( .A(net16), .Y(outb));
inv I_inv2 ( .A(outb), .Y(out));
inv I1 ( .A(sel), .Y(net10));

endmodule
// Library - ice8chip, Cell - clk_quad_buf_ice8p, View - schematic
// LAST TIME SAVED: Aug 12 09:03:48 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module clk_quad_buf_ice8p ( clko, clki );
output  clko;

input  clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I19 ( .A(clkb), .Y(clko));
inv_lvt I22 ( .A(clki), .Y(clkb));

endmodule
// Library - ice8chip, Cell - clk_quad_buf_x8_ice8p, View - schematic
// LAST TIME SAVED: Jun 24 14:46:09 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module clk_quad_buf_x8_ice8p ( clko, clki );


output [7:0]  clko;

input [7:0]  clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_quad_buf_ice8p I_clk_quad_buf_ice8p_7_ ( .clki(clki[7]),
     .clko(clko[7]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_6_ ( .clki(clki[6]),
     .clko(clko[6]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_5_ ( .clki(clki[5]),
     .clko(clko[5]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_4_ ( .clki(clki[4]),
     .clko(clko[4]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_3_ ( .clki(clki[3]),
     .clko(clko[3]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_2_ ( .clki(clki[2]),
     .clko(clko[2]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_1_ ( .clki(clki[1]),
     .clko(clko[1]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_0_ ( .clki(clki[0]),
     .clko(clko[0]));

endmodule
// Library - leafcell, Cell - misc_module4_v3, View - schematic
// LAST TIME SAVED: Mar 21 13:25:15 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module misc_module4_v3 ( S_R, cbit, cbitb, clk, clkb, glb2local, sp4,
     bl, b, glb_netwk, l, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3,
     m, min0, min1, min2, min3, pgate, prog, r, reset_b, sp12,
     vdd_cntl, wl );
output  S_R, clk, clkb;


input  prog;

output [7:0]  sp4;
output [3:0]  glb2local;
output [63:0]  cbit;
output [63:0]  cbitb;

inout [3:0]  bl;

input [15:0]  pgate;
input [5:0]  lc_trk_g1;
input [15:0]  vdd_cntl;
input [5:0]  lc_trk_g3;
input [7:0]  min1;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g0;
input [15:0]  wl;
input [7:0]  min0;
input [7:0]  min2;
input [1:0]  r;
input [1:0]  l;
input [1:0]  m;
input [1:0]  b;
input [5:0]  lc_trk_g2;
input [15:0]  reset_b;
input [7:0]  sp12;
input [7:0]  min3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  r_vdd;



inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
pch_hvt  M0_15_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[15]), .S(r_vdd[15]));
pch_hvt  M0_14_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[14]), .S(r_vdd[14]));
pch_hvt  M0_13_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[13]), .S(r_vdd[13]));
pch_hvt  M0_12_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[12]), .S(r_vdd[12]));
pch_hvt  M0_11_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[11]), .S(r_vdd[11]));
pch_hvt  M0_10_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[10]), .S(r_vdd[10]));
pch_hvt  M0_9_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[9]), .S(r_vdd[9]));
pch_hvt  M0_8_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[8]), .S(r_vdd[8]));
pch_hvt  M0_7_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[7]), .S(r_vdd[7]));
pch_hvt  M0_6_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[6]), .S(r_vdd[6]));
pch_hvt  M0_5_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[5]), .S(r_vdd[5]));
pch_hvt  M0_4_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[4]), .S(r_vdd[4]));
pch_hvt  M0_3_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[3]), .S(r_vdd[3]));
pch_hvt  M0_2_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[2]), .S(r_vdd[2]));
pch_hvt  M0_1_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[1]), .S(r_vdd[1]));
pch_hvt  M0_0_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[0]), .S(r_vdd[0]));
clkmandcmuxrev0 I_clkmandcmuxrev0 ( .prog(progd),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]), .clk(clk),
     .clkb(clkb), .glb_netwk(glb_netwk[7:0]), .s_r(S_R),
     .glb2local(glb2local[3:0]), .cbit({cbit[2], cbit[1], cbit[0],
     cbit[27], cbit[25], cbit[26], cbit[24], cbit[23], cbit[21],
     cbit[22], cbit[20], cbit[19], cbit[17], cbit[18], cbit[16],
     cbit[15], cbit[13], cbit[14], cbit[12], cbit[31], cbit[29],
     cbit[30], cbit[28], cbit[11], cbit[9], cbit[10], cbit[8],
     cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}), .min2(min2[7:0]),
     .min1(min1[7:0]), .min0(min0[7:0]), .min3(min3[7:0]),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}));
sp12to4 I_sp12to4_7_ ( .prog(progd), .triout(sp4[7]),
     .cbitb(cbitb[62]), .drv(sp12[7]));
sp12to4 I_sp12to4_6_ ( .prog(progd), .triout(sp4[6]),
     .cbitb(cbitb[58]), .drv(sp12[6]));
sp12to4 I_sp12to4_5_ ( .prog(progd), .triout(sp4[5]),
     .cbitb(cbitb[54]), .drv(sp12[5]));
sp12to4 I_sp12to4_4_ ( .prog(progd), .triout(sp4[4]),
     .cbitb(cbitb[50]), .drv(sp12[4]));
sp12to4 I_sp12to4_3_ ( .prog(progd), .triout(sp4[3]),
     .cbitb(cbitb[46]), .drv(sp12[3]));
sp12to4 I_sp12to4_2_ ( .prog(progd), .triout(sp4[2]),
     .cbitb(cbitb[42]), .drv(sp12[2]));
sp12to4 I_sp12to4_1_ ( .prog(progd), .triout(sp4[1]), .cbitb(cbitb[5]),
     .drv(sp12[1]));
sp12to4 I_sp12to4_0_ ( .prog(progd), .triout(sp4[0]),
     .cbitb(cbitb[34]), .drv(sp12[0]));
sbox1 I_sbox1_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(progd));
sbox1 I_sbox1_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(progd));
cram16x4 I_cram16x4 ( .q(cbit[63:0]), .r_gnd(r_vdd[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));

endmodule
// Library - xpmem, Cell - cram_2x28, View - schematic
// LAST TIME SAVED: Jun 24 18:02:26 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module cram_2x28 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [55:0]  q;
output [55:0]  q_b;

inout [27:0]  bl;

input [1:0]  r_vdd;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 I_mstake_13_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[27:26]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[1:0]));
cram2x2 I_mstake_12_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[25:24]), .q_b(q_b[51:48]),
     .q(q[51:48]), .wl(wl[1:0]));
cram2x2 I_mstake_11_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[23:22]), .q_b(q_b[47:44]),
     .q(q[47:44]), .wl(wl[1:0]));
cram2x2 I_mstake_10_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[21:20]), .q_b(q_b[43:40]),
     .q(q[43:40]), .wl(wl[1:0]));
cram2x2 I_mstake_9_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[19:18]), .q_b(q_b[39:36]),
     .q(q[39:36]), .wl(wl[1:0]));
cram2x2 I_mstake_8_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[17:16]), .q_b(q_b[35:32]),
     .q(q[35:32]), .wl(wl[1:0]));
cram2x2 I_mstake_7_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[15:14]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[1:0]));
cram2x2 I_mstake_6_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[13:12]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[1:0]));
cram2x2 I_mstake_5_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 I_mstake_4_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 I_mstake_3_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 I_mstake_2_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 I_mstake_1_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 I_mstake_0_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - logic_cell_rev, View - schematic
// LAST TIME SAVED: Sep  3 10:41:29 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module logic_cell_rev ( carry_out, out, out_vic, carry_in, cbit, clk,
     clkb, in0, in1, in2, in3, prog, purst, s_r );
output  carry_out, out, out_vic;

input  carry_in, clk, clkb, in0, in1, in2, in3, prog, purst, s_r;

input [20:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clut4vic I_clut4 ( .lut4vic(out_vic), .in3b(in3b), .in3(in3),
     .in2b(in2b), .in2(in2), .in1b(in1b), .in1(in1), .in0b(in0b),
     .in0(in0), .cbit(cbit[15:0]), .lut4(LUT4_outd));
o_mux I_o_mux ( .prog(prog), .in1(rego), .in0(LUT4_outd),
     .cbit(cbit[19]), .out(out));
inv_lvt I196 ( .A(in3), .Y(in3b));
inv_lvt I189 ( .A(in0), .Y(in0b));
inv_lvt I194 ( .A(in1), .Y(in1b));
inv_lvt I195 ( .A(in2), .Y(in2b));
carry_logic_nand I_carry_logic ( .vg_en(cbit[20]), .carry_in(carry_in),
     .b_bar(in1b), .b(in1), .a_bar(in2b), .a(in2), .cout(carry_out));
coredffr I_coredffr ( .purst(purst), .d(LUT4_outd), .clkb(clkb),
     .clk(clk), .cbit(cbit[17:16]), .S_R(s_r), .q(rego));

endmodule
// Library - leafcell, Cell - lcmuxod3_0_0, View - schematic
// LAST TIME SAVED: Jun 24 17:41:19 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module lcmuxod3_0_0 ( carry_out, cbit, cbitb, op, op_vic, sp4_h_r,
     sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb,
     min0, min1, min2, min3, op_bot, pgate, prog, purst, reset_b, s_r,
     vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_h_r;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [1:0]  sp12_v_b;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [55:0]  cbit;
output [55:0]  cbitb;
output [2:0]  sp4_v_b;

input [15:0]  min2;
input [1:0]  pgate;
input [15:0]  min0;
input [15:0]  min1;
input [1:0]  reset_b;
input [15:0]  min3;
input [27:0]  bl;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



in_mux_nand_icc I_in2mux_nand ( .cbitb({cbitb[50], cbitb[12],
     cbitb[13], cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50],
     cbit[12], cbit[13], cbit[16], cbit[19], cbit[17]}),
     .op_bot(op_bot), .prog(prog), .inmuxo(in2), .min(min2[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_30 I_odrv30 ( .slfop(op), .prog(prog),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53], cbitb[55],
     cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44], cbitb[46],
     cbitb[43], cbitb[41], cbitb[42], cbitb[40]}), .sp12_h_r(sp12_h_r),
     .sp12_v_b(sp12_v_b[1:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));

endmodule
// Library - leafcell, Cell - lcmuxod3_0, View - schematic
// LAST TIME SAVED: Jun 23 08:18:57 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module lcmuxod3_0 ( carry_out, op, op_vic, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, op_bot, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_h_r;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [1:0]  sp12_v_b;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [2:0]  sp4_v_b;

input [1:0]  wl;
input [15:0]  min0;
input [1:0]  pgate;
input [15:0]  min1;
input [27:0]  bl;
input [1:0]  vdd_cntl;
input [15:0]  min3;
input [15:0]  min2;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [55:0]  cbitb;

wire  [55:0]  cbit;



in_mux_nand_icc I_in2mux_nand ( .cbitb({cbitb[50], cbitb[12],
     cbitb[13], cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50],
     cbit[12], cbit[13], cbit[16], cbit[19], cbit[17]}),
     .op_bot(op_bot), .prog(prog), .inmuxo(in2), .min(min2[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_30 I_odrv30 ( .slfop(op), .prog(prog),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53], cbitb[55],
     cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44], cbitb[46],
     cbitb[43], cbitb[41], cbitb[42], cbitb[40]}), .sp12_h_r(sp12_h_r),
     .sp12_v_b(sp12_v_b[1:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));

endmodule
// Library - leafcell, Cell - lcmuxod7_4, View - schematic
// LAST TIME SAVED: Jun 23 08:19:59 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module lcmuxod7_4 ( carry_out, op, op_vic, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, op_bot, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_v_b;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_h_r;

input [27:0]  bl;
input [15:0]  min1;
input [1:0]  reset_b;
input [15:0]  min0;
input [15:0]  min3;
input [1:0]  pgate;
input [15:0]  min2;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [55:0]  cbitb;

wire  [55:0]  cbit;



in_mux_nand_icc I_in2mux ( .cbitb({cbitb[50], cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50], cbit[12],
     cbit[13], cbit[16], cbit[19], cbit[17]}), .op_bot(op_bot),
     .prog(prog), .inmuxo(in2), .min(min2[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_74 I_odrv74 ( .slfop(op), .prog(prog), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));

endmodule
// Library - leafcell, Cell - lccol_rev0, View - schematic
// LAST TIME SAVED: Oct 18 13:49:45 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module lccol_rev0 ( carry_out, op_vic, slf_op, bl, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, cin2local, clk, clkb, lc_trk_g0,
     lc_trk_g1, lc_trk_g2, lc_trk_g3, op_bot, pgate, prog, purst,
     reset_b, s_r, vdd_cntl, wl );
output  carry_out, op_vic;


input  cin2local, clk, clkb, op_bot, prog, purst, s_r;

output [7:0]  slf_op;

inout [27:0]  bl;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;

input [15:0]  reset_b;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g2;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  wl;
input [7:0]  lc_trk_g3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbitb;

wire  [55:0]  cbit;



lcmuxod3_0_0 I_LC_00 ( .cbitb(cbitb[55:0]), .cbit(cbit[55:0]),
     .op_bot(op_bot), .op_vic(net0118), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .carry_out(c_01),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], cin}),
     .reset_b(reset_b[1:0]), .vdd_cntl(vdd_cntl[1:0]), .wl(wl[1:0]),
     .op(slf_op[0]), .s_r(s_r), .sp4_h_r({sp4_h_r[32], sp4_h_r[16],
     sp4_h_r[0]}), .sp12_v_b({sp12_v_b[16], sp12_v_b[0]}),
     .sp4_r_v_b({sp4_r_v_b[33], sp4_r_v_b[17], sp4_r_v_b[1]}),
     .sp4_v_b({sp4_v_b[32], sp4_v_b[16], sp4_v_b[0]}), .carry_in(cin),
     .sp12_h_r(sp12_h_r[8]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[1:0]), .prog(prog));
lcmuxod3_0 I_LC_02 ( .op_bot(net0166), .op_vic(net094),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .carry_out(c_23), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_12}),
     .reset_b(reset_b[5:4]), .vdd_cntl(vdd_cntl[5:4]), .wl(wl[5:4]),
     .op(slf_op[2]), .s_r(s_r), .sp4_h_r({sp4_h_r[36], sp4_h_r[20],
     sp4_h_r[4]}), .sp12_v_b({sp12_v_b[20], sp12_v_b[4]}),
     .sp4_r_v_b({sp4_r_v_b[37], sp4_r_v_b[21], sp4_r_v_b[5]}),
     .sp4_v_b({sp4_v_b[36], sp4_v_b[20], sp4_v_b[4]}), .carry_in(c_12),
     .sp12_h_r(sp12_h_r[12]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[5:4]), .prog(prog));
lcmuxod3_0 I_LC_03 ( .op_bot(net094), .op_vic(net0142),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .carry_out(c_34), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_23}),
     .reset_b(reset_b[7:6]), .vdd_cntl(vdd_cntl[7:6]), .wl(wl[7:6]),
     .op(slf_op[3]), .s_r(s_r), .sp4_h_r({sp4_h_r[38], sp4_h_r[22],
     sp4_h_r[6]}), .sp12_v_b({sp12_v_b[22], sp12_v_b[6]}),
     .sp4_r_v_b({sp4_r_v_b[39], sp4_r_v_b[23], sp4_r_v_b[7]}),
     .sp4_v_b({sp4_v_b[38], sp4_v_b[22], sp4_v_b[6]}), .carry_in(c_23),
     .sp12_h_r(sp12_h_r[14]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[7:6]), .prog(prog));
lcmuxod3_0 I_LC_01 ( .op_bot(net0118), .op_vic(net0166),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .carry_out(c_12), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_01}),
     .reset_b(reset_b[3:2]), .vdd_cntl(vdd_cntl[3:2]), .wl(wl[3:2]),
     .op(slf_op[1]), .s_r(s_r), .sp4_h_r({sp4_h_r[34], sp4_h_r[18],
     sp4_h_r[2]}), .sp12_v_b({sp12_v_b[18], sp12_v_b[2]}),
     .sp4_r_v_b({sp4_r_v_b[35], sp4_r_v_b[19], sp4_r_v_b[3]}),
     .sp4_v_b({sp4_v_b[34], sp4_v_b[18], sp4_v_b[2]}), .carry_in(c_01),
     .sp12_h_r(sp12_h_r[10]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[3:2]), .prog(prog));
lcmuxod7_4 I_LC_07 ( .op_vic(op_vic), .op_bot(net0261), .bl(bl[27:0]),
     .reset_b(reset_b[15:14]), .purst(purst), .wl(wl[15:14]),
     .vdd_cntl(vdd_cntl[15:14]), .sp4_r_v_b({sp4_r_v_b[47],
     sp4_r_v_b[31], sp4_r_v_b[15]}), .sp4_h_r({sp4_h_r[46],
     sp4_h_r[30], sp4_h_r[14]}), .sp4_v_b({sp4_v_b[46], sp4_v_b[30],
     sp4_v_b[14]}), .pgate(pgate[15:14]), .sp12_h_r({sp12_h_r[22],
     sp12_h_r[6]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_67}),
     .carry_out(carry_out), .op(slf_op[7]), .s_r(s_r),
     .sp12_v_b(sp12_v_b[14]), .clk(clk), .carry_in(c_67),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clkb(clkb), .prog(prog));
lcmuxod7_4 I_LC_04 ( .op_vic(net0213), .op_bot(net0142), .prog(prog),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_34}), .clkb(clkb),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .purst(purst),
     .sp4_h_r({sp4_h_r[40], sp4_h_r[24], sp4_h_r[8]}),
     .sp4_r_v_b({sp4_r_v_b[41], sp4_r_v_b[25], sp4_r_v_b[9]}),
     .sp12_v_b(sp12_v_b[8]), .reset_b(reset_b[9:8]),
     .vdd_cntl(vdd_cntl[9:8]), .bl(bl[27:0]), .pgate(pgate[9:8]),
     .wl(wl[9:8]), .sp4_v_b({sp4_v_b[40], sp4_v_b[24], sp4_v_b[8]}),
     .sp12_h_r({sp12_h_r[16], sp12_h_r[0]}), .carry_out(c_45),
     .carry_in(c_34), .op(slf_op[4]));
lcmuxod7_4 I_LC_05 ( .op_vic(net0237), .op_bot(net0213), .prog(prog),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_45}), .clkb(clkb),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .purst(purst),
     .sp4_h_r({sp4_h_r[42], sp4_h_r[26], sp4_h_r[10]}),
     .sp4_r_v_b({sp4_r_v_b[43], sp4_r_v_b[27], sp4_r_v_b[11]}),
     .sp12_v_b(sp12_v_b[10]), .reset_b(reset_b[11:10]),
     .vdd_cntl(vdd_cntl[11:10]), .bl(bl[27:0]), .pgate(pgate[11:10]),
     .wl(wl[11:10]), .sp4_v_b({sp4_v_b[42], sp4_v_b[26], sp4_v_b[10]}),
     .sp12_h_r({sp12_h_r[18], sp12_h_r[2]}), .carry_out(c_56),
     .carry_in(c_45), .op(slf_op[5]));
lcmuxod7_4 I_LC_06 ( .op_vic(net0261), .op_bot(net0237), .prog(prog),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_56}), .clkb(clkb),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .purst(purst),
     .sp4_h_r({sp4_h_r[44], sp4_h_r[28], sp4_h_r[12]}),
     .sp4_r_v_b({sp4_r_v_b[45], sp4_r_v_b[29], sp4_r_v_b[13]}),
     .sp12_v_b(sp12_v_b[12]), .reset_b(reset_b[13:12]),
     .vdd_cntl(vdd_cntl[13:12]), .bl(bl[27:0]), .pgate(pgate[13:12]),
     .wl(wl[13:12]), .sp4_v_b({sp4_v_b[44], sp4_v_b[28], sp4_v_b[12]}),
     .sp12_h_r({sp12_h_r[20], sp12_h_r[4]}), .carry_out(c_67),
     .carry_in(c_56), .op(slf_op[6]));
mux_4carry I_carry_cnt ( .cin(cin2local), .lcl_cin(cin),
     .cbitb({cbitb[45], cbitb[48]}), .prog(prog), .cbit({cbit[45],
     cbit[48]}));

endmodule
// Library - ice1chip, Cell - ltile4_ice1f, View - schematic
// LAST TIME SAVED: Mar 31 17:35:26 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ltile4_ice1f ( carry_out, cntl_cbit, op_vic, slf_op, bl,
     sp4_h_l, sp4_h_r, sp4_r_v_b, sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r,
     sp12_v_b, sp12_v_t, bnl_op, bnr_op, bot_op, carry_in, glb_netwk,
     lft_op, op_bot, pgate, prog, purst, reset_b, rgt_op, tnl_op,
     tnr_op, top_op, vdd_cntl, wl );
output  carry_out, op_vic;


input  carry_in, op_bot, prog, purst;

output [7:0]  slf_op;
output [7:0]  cntl_cbit;

inout [47:0]  sp4_v_t;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [23:0]  sp12_v_t;
inout [47:0]  sp4_h_r;
inout [53:0]  bl;

input [7:0]  bnl_op;
input [7:0]  tnl_op;
input [7:0]  glb_netwk;
input [7:0]  tnr_op;
input [7:0]  lft_op;
input [7:0]  bnr_op;
input [15:0]  pgate;
input [7:0]  bot_op;
input [15:0]  reset_b;
input [7:0]  top_op;
input [15:0]  vdd_cntl;
input [7:0]  rgt_op;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  lc_trk_g0;

wire  [1:0]  sp12_h_r_mid;

wire  [7:0]  lc_trk_g1;

wire  [3:0]  net_glb2local;

wire  [63:0]  cbitb_c;

wire  [1:0]  sp12_v_b_mid;

wire  [7:0]  lc_trk_g3;

wire  [7:0]  lc_trk_g2;

wire  [63:0]  cbit_c;

wire  [0:7]  net187;

wire  [0:7]  net188;



inv_hvt I97 ( .A(purst), .Y(purstb));
inv_hvt I98 ( .A(purstb), .Y(purstd));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(progd));
rm8y  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm8y  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm8y  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm8y  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm8y  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm8y  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm8y  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm8y  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm8y  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm8y  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm8y  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm8y  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm8y  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm8y  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm8y  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm8y  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm8y  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm8y  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm8y  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm8y  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm8y  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm8y  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm8y  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm8y  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
span4_ice8p I_sp4_sw ( .bram_cbit(net188[0:7]),
     .ccntrl_cbit(net187[0:7]), .sp4_h_l(sp4_h_l[47:0]), .bl(bl[13:4]),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_t(sp4_v_t[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .reset_b({reset_b[14], reset_b[15],
     reset_b[12], reset_b[13], reset_b[10], reset_b[11], reset_b[8],
     reset_b[9], reset_b[6], reset_b[7], reset_b[4], reset_b[5],
     reset_b[2], reset_b[3], reset_b[0], reset_b[1]}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .prog(progd));
misc_module4_v3 I_misc ( .cbitb(cbitb_c[63:0]), .cbit({cbit_c[63:61],
     cntl_cbit[7], cbit_c[59:57], cntl_cbit[6], cbit_c[55:53],
     cntl_cbit[5], cbit_c[51:49], cntl_cbit[4], cbit_c[47:45],
     cntl_cbit[3], cbit_c[43:41], cntl_cbit[2], cbit_c[39:33],
     cntl_cbit[1], cbit_c[31:4], cntl_cbit[0], cbit_c[2:0]}),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .lc_trk_g1(lc_trk_g1[5:0]), .glb2local(net_glb2local[3:0]),
     .clkb(clkb), .bl(bl[3:0]), .min2(glb_netwk[7:0]),
     .min3(glb_netwk[7:0]), .min1(glb_netwk[7:0]),
     .min0(glb_netwk[7:0]), .glb_netwk(glb_netwk[7:0]),
     .lc_trk_g0(lc_trk_g0[5:0]), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .sp4(sp4_h_r[23:16]), .l(sp12_h_r_mid[1:0]),
     .S_R(s_r), .clk(clk), .b(sp12_v_b[1:0]), .r(sp12_h_r[1:0]),
     .m(sp12_v_b_mid[1:0]), .prog(progd), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18],
     sp12_h_r[16], sp12_h_r[14], sp12_h_r[12], sp12_h_r[10],
     sp12_h_r[8]}), .reset_b({reset_b[14], reset_b[15], reset_b[12],
     reset_b[13], reset_b[10], reset_b[11], reset_b[8], reset_b[9],
     reset_b[6], reset_b[7], reset_b[4], reset_b[5], reset_b[2],
     reset_b[3], reset_b[0], reset_b[1]}), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}));
gmux_sp12to4 I_gmux_sp12to4 ( .reset_b({reset_b[14], reset_b[15],
     reset_b[12], reset_b[13], reset_b[10], reset_b[11], reset_b[8],
     reset_b[9], reset_b[6], reset_b[7], reset_b[4], reset_b[5],
     reset_b[2], reset_b[3], reset_b[0], reset_b[1]}),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .lft_op(lft_op[7:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .glb2local(net_glb2local[3:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .bnr_op(bnr_op[7:0]), .lc_trk_g2(lc_trk_g2[7:0]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .bl(bl[25:14]), .lc_trk_g3(lc_trk_g3[7:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .prog(progd));
rm7y  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7y  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7y  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7y  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7y  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7y  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7y  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7y  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7y  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7y  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7y  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7y  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7y  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7y  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7y  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7y  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7y  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7y  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7y  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7y  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7y  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7y  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7y  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7y  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
lccol_rev0 I_lccol_rev0 ( .op_bot(op_bot), .op_vic(op_vic),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .wl({wl[14], wl[15], wl[12], wl[13],
     wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2],
     wl[3], wl[0], wl[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .s_r(s_r), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .prog(progd), .purst(purstd), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .clkb(clkb), .clk(clk),
     .cin2local(carry_in), .slf_op(slf_op[7:0]), .carry_out(carry_out),
     .sp12_v_b(sp12_v_b[23:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .bl(bl[53:26]));

endmodule
// Library - leafcell, Cell - clkbuffer500um, View - schematic
// LAST TIME SAVED: May 13 10:52:41 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module clkbuffer500um ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I4 ( .A(net6), .Y(out));
inv I3 ( .A(in), .Y(net6));

endmodule
// Library - ice1chip, Cell - lt_1x8_top_ice1f, View - schematic
// LAST TIME SAVED: Jun  6 13:23:14 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module lt_1x8_top_ice1f ( carry_out, glb_netwk_b, glb_netwk_t, op_vic,
     slf_op_01, slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06,
     slf_op_07, slf_op_08, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02,
     sp4_h_l_03, sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07,
     sp4_h_l_08, sp4_h_r_01, sp4_h_r_02, sp4_h_r_03, sp4_h_r_04,
     sp4_h_r_05, sp4_h_r_06, sp4_h_r_07, sp4_h_r_08, sp4_r_v_b_01,
     sp4_r_v_b_02, sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05,
     sp4_r_v_b_06, sp4_r_v_b_07, sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02,
     sp4_v_b_03, sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07,
     sp4_v_b_08, sp4_v_t_08, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03,
     sp12_h_l_04, sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08,
     sp12_h_r_01, sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_h_r_05,
     sp12_h_r_06, sp12_h_r_07, sp12_h_r_08, sp12_v_b_01, sp12_v_t_08,
     vdd_cntl, wl, bnl_op_01, bnr_op_01, bot_op_01, carry_in,
     glb_netwk_col, lc_bot, lft_op_01, lft_op_02, lft_op_03, lft_op_04,
     lft_op_05, lft_op_06, lft_op_07, lft_op_08, prog, purst,
     rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04, rgt_op_05, rgt_op_06,
     rgt_op_07, rgt_op_08, tnl_op_08, tnr_op_08, top_op_08 );
output  carry_out, op_vic;


input  carry_in, lc_bot, prog, purst;

output [7:0]  slf_op_05;
output [7:0]  slf_op_07;
output [7:0]  slf_op_06;
output [7:0]  slf_op_08;
output [7:0]  slf_op_01;
output [7:0]  glb_netwk_t;
output [7:0]  glb_netwk_b;
output [7:0]  slf_op_04;
output [7:0]  slf_op_02;
output [7:0]  slf_op_03;

inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_r_08;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_h_r_06;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_v_b_05;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_r_08;
inout [23:0]  sp12_h_l_01;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_r_v_b_07;
inout [53:0]  bl;
inout [23:0]  sp12_h_r_05;
inout [23:0]  sp12_h_l_05;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_h_l_05;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_v_b_06;
inout [47:0]  sp4_h_l_01;
inout [23:0]  sp12_v_t_08;
inout [23:0]  sp12_h_l_04;
inout [23:0]  sp12_v_b_01;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_v_t_08;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_v_b_03;
inout [23:0]  sp12_h_r_02;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_l_06;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_r_v_b_05;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_h_r_07;
inout [127:0]  reset_b;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_r_v_b_04;
inout [127:0]  pgate;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_h_l_04;
inout [127:0]  vdd_cntl;
inout [127:0]  wl;

input [7:0]  rgt_op_05;
input [7:0]  rgt_op_07;
input [7:0]  lft_op_03;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_02;
input [7:0]  lft_op_04;
input [7:0]  bnr_op_01;
input [7:0]  lft_op_05;
input [7:0]  lft_op_01;
input [7:0]  rgt_op_01;
input [7:0]  lft_op_02;
input [7:0]  rgt_op_06;
input [7:0]  lft_op_07;
input [7:0]  lft_op_06;
input [7:0]  bnl_op_01;
input [7:0]  top_op_08;
input [7:0]  rgt_op_04;
input [7:0]  tnr_op_08;
input [7:0]  tnl_op_08;
input [7:0]  lft_op_08;
input [7:0]  rgt_op_08;
input [7:0]  glb_netwk_col;
input [7:0]  bot_op_01;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net0754;

wire  [0:23]  net711;

wire  [7:0]  colbuf_cntl_b;

wire  [0:7]  net947;

wire  [0:23]  net1083;

wire  [0:23]  net990;

wire  [0:23]  net959;

wire  [0:7]  net668;

wire  [0:23]  net680;

wire  [7:0]  colbuf_cntl_t;

wire  [0:23]  net742;

wire  [0:7]  net978;

wire  [0:7]  net637;

wire  [0:23]  net649;

wire  [0:7]  net1071;



ltile4_ice1f I_LT06 ( .cntl_cbit(net637[0:7]), .op_bot(net732),
     .op_vic(net639), .prog(prog), .carry_out(net641),
     .lft_op(lft_op_06[7:0]), .sp12_h_l(sp12_h_l_06[23:0]),
     .sp4_h_l(sp4_h_l_06[47:0]), .sp4_v_b(sp4_v_b_06[47:0]),
     .sp12_v_b(net742[0:23]), .sp12_h_r(sp12_h_r_06[23:0]),
     .sp4_h_r(sp4_h_r_06[47:0]), .sp12_v_t(net649[0:23]),
     .sp4_v_t(sp4_v_b_07[47:0]), .sp4_r_v_b(sp4_r_v_b_06[47:0]),
     .wl(wl[95:80]), .top_op(slf_op_07[7:0]), .rgt_op(rgt_op_06[7:0]),
     .bot_op(slf_op_05[7:0]), .bl(bl[53:0]), .reset_b(reset_b[95:80]),
     .vdd_cntl(vdd_cntl[95:80]), .glb_netwk(glb_netwk_t[7:0]),
     .carry_in(net734), .purst(purst), .slf_op(slf_op_06[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_05[7:0]),
     .bnl_op(lft_op_05[7:0]), .tnr_op(rgt_op_07[7:0]),
     .tnl_op(lft_op_07[7:0]));
ltile4_ice1f I_LT03 ( .cntl_cbit(net668[0:7]), .op_bot(net980),
     .op_vic(net670), .prog(prog), .carry_out(net672),
     .lft_op(lft_op_03[7:0]), .sp12_h_l(sp12_h_l_03[23:0]),
     .sp4_h_l(sp4_h_l_03[47:0]), .sp4_v_b(sp4_v_b_03[47:0]),
     .sp12_v_b(net990[0:23]), .sp12_h_r(sp12_h_r_03[23:0]),
     .sp4_h_r(sp4_h_r_03[47:0]), .sp12_v_t(net680[0:23]),
     .sp4_v_t(sp4_v_b_04[47:0]), .sp4_r_v_b(sp4_r_v_b_03[47:0]),
     .wl(wl[47:32]), .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(net982), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4_ice1f I_LT04 ( .cntl_cbit(colbuf_cntl_b[7:0]), .op_bot(net670),
     .op_vic(net701), .prog(prog), .carry_out(net703),
     .lft_op(lft_op_04[7:0]), .sp12_h_l(sp12_h_l_04[23:0]),
     .sp4_h_l(sp4_h_l_04[47:0]), .sp4_v_b(sp4_v_b_04[47:0]),
     .sp12_v_b(net680[0:23]), .sp12_h_r(sp12_h_r_04[23:0]),
     .sp4_h_r(sp4_h_r_04[47:0]), .sp12_v_t(net711[0:23]),
     .sp4_v_t(sp4_v_b_05[47:0]), .sp4_r_v_b(sp4_r_v_b_04[47:0]),
     .wl(wl[63:48]), .top_op(slf_op_05[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(net672), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(rgt_op_05[7:0]),
     .tnl_op(lft_op_05[7:0]));
ltile4_ice1f I_LT05 ( .cntl_cbit(colbuf_cntl_t[7:0]), .op_bot(net701),
     .op_vic(net732), .prog(prog), .carry_out(net734),
     .lft_op(lft_op_05[7:0]), .sp12_h_l(sp12_h_l_05[23:0]),
     .sp4_h_l(sp4_h_l_05[47:0]), .sp4_v_b(sp4_v_b_05[47:0]),
     .sp12_v_b(net711[0:23]), .sp12_h_r(sp12_h_r_05[23:0]),
     .sp4_h_r(sp4_h_r_05[47:0]), .sp12_v_t(net742[0:23]),
     .sp4_v_t(sp4_v_b_06[47:0]), .sp4_r_v_b(sp4_r_v_b_05[47:0]),
     .wl(wl[79:64]), .top_op(slf_op_06[7:0]), .rgt_op(rgt_op_05[7:0]),
     .bot_op(slf_op_04[7:0]), .bl(bl[53:0]), .reset_b(reset_b[79:64]),
     .vdd_cntl(vdd_cntl[79:64]), .glb_netwk(glb_netwk_t[7:0]),
     .carry_in(net703), .purst(purst), .slf_op(slf_op_05[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_04[7:0]),
     .bnl_op(lft_op_04[7:0]), .tnr_op(rgt_op_06[7:0]),
     .tnl_op(lft_op_06[7:0]));
ltile4_ice1f I_LT01 ( .cntl_cbit(net947[0:7]), .op_bot(lc_bot),
     .op_vic(net949), .prog(prog), .carry_out(net951),
     .lft_op(lft_op_01[7:0]), .sp12_h_l(sp12_h_l_01[23:0]),
     .sp4_h_l(sp4_h_l_01[47:0]), .sp4_v_b(sp4_v_b_01[47:0]),
     .sp12_v_b(sp12_v_b_01[23:0]), .sp12_h_r(sp12_h_r_01[23:0]),
     .sp4_h_r(sp4_h_r_01[47:0]), .sp12_v_t(net959[0:23]),
     .sp4_v_t(sp4_v_b_02[47:0]), .sp4_r_v_b(sp4_r_v_b_01[47:0]),
     .wl(wl[15:0]), .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4_ice1f I_LT02 ( .cntl_cbit(net978[0:7]), .op_bot(net949),
     .op_vic(net980), .prog(prog), .carry_out(net982),
     .lft_op(lft_op_02[7:0]), .sp12_h_l(sp12_h_l_02[23:0]),
     .sp4_h_l(sp4_h_l_02[47:0]), .sp4_v_b(sp4_v_b_02[47:0]),
     .sp12_v_b(net959[0:23]), .sp12_h_r(sp12_h_r_02[23:0]),
     .sp4_h_r(sp4_h_r_02[47:0]), .sp12_v_t(net990[0:23]),
     .sp4_v_t(sp4_v_b_03[47:0]), .sp4_r_v_b(sp4_r_v_b_02[47:0]),
     .wl(wl[31:16]), .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(net951), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));
ltile4_ice1f I_LT08 ( .cntl_cbit(net0754[0:7]), .op_bot(net1073),
     .op_vic(op_vic), .prog(prog), .carry_out(carry_out),
     .lft_op(lft_op_08[7:0]), .sp12_h_l(sp12_h_l_08[23:0]),
     .sp4_h_l(sp4_h_l_08[47:0]), .sp4_v_b(sp4_v_b_08[47:0]),
     .sp12_v_b(net1083[0:23]), .sp12_h_r(sp12_h_r_08[23:0]),
     .sp4_h_r(sp4_h_r_08[47:0]), .sp12_v_t(sp12_v_t_08[23:0]),
     .sp4_v_t(sp4_v_t_08[47:0]), .sp4_r_v_b(sp4_r_v_b_08[47:0]),
     .wl(wl[127:112]), .top_op(top_op_08[7:0]),
     .rgt_op(rgt_op_08[7:0]), .bot_op(slf_op_07[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[127:112]), .vdd_cntl(vdd_cntl[127:112]),
     .glb_netwk(glb_netwk_t[7:0]), .carry_in(net1075), .purst(purst),
     .slf_op(slf_op_08[7:0]), .pgate(pgate[127:112]),
     .bnr_op(rgt_op_07[7:0]), .bnl_op(lft_op_07[7:0]),
     .tnr_op(tnr_op_08[7:0]), .tnl_op(tnl_op_08[7:0]));
ltile4_ice1f I_LT07 ( .cntl_cbit(net1071[0:7]), .op_bot(net639),
     .op_vic(net1073), .prog(prog), .carry_out(net1075),
     .lft_op(lft_op_07[7:0]), .sp12_h_l(sp12_h_l_07[23:0]),
     .sp4_h_l(sp4_h_l_07[47:0]), .sp4_v_b(sp4_v_b_07[47:0]),
     .sp12_v_b(net649[0:23]), .sp12_h_r(sp12_h_r_07[23:0]),
     .sp4_h_r(sp4_h_r_07[47:0]), .sp12_v_t(net1083[0:23]),
     .sp4_v_t(sp4_v_b_08[47:0]), .sp4_r_v_b(sp4_r_v_b_07[47:0]),
     .wl(wl[111:96]), .top_op(slf_op_08[7:0]), .rgt_op(rgt_op_07[7:0]),
     .bot_op(slf_op_06[7:0]), .bl(bl[53:0]), .reset_b(reset_b[111:96]),
     .vdd_cntl(vdd_cntl[111:96]), .glb_netwk(glb_netwk_t[7:0]),
     .carry_in(net641), .purst(purst), .slf_op(slf_op_07[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_06[7:0]),
     .bnl_op(lft_op_06[7:0]), .tnr_op(rgt_op_08[7:0]),
     .tnl_op(lft_op_08[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - ice1chip, Cell - quad_tr_ice1, View - schematic
// LAST TIME SAVED: Apr 26 17:01:49 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module quad_tr_ice1 ( bm_aa_2bot, bm_ab_2bot, bm_sdo_o, bs_en_o, ceb_o,
     cf_r, cf_t, fabric_out_07_17, fabric_out_08_17, fabric_out_13_09,
     fabric_out_13_10, hiz_b_o, mode_o, padeb_r, padeb_t_r,
     padin_07_17a, padin_13_09a, pado_r, pado_t_r, r_o, sdo, shift_o,
     slf_op_07_09, slf_op_07_10, slf_op_07_11, slf_op_07_12,
     slf_op_07_13, slf_op_07_14, slf_op_07_15, slf_op_07_16,
     slf_op_07_17, slf_op_08_09, slf_op_09_09, slf_op_10_09,
     slf_op_11_09, slf_op_12_09, slf_op_13_09, tclk_o, update_o, bl,
     pgate_r, reset_b_r, sp4_h_l_07_09, sp4_h_l_07_10, sp4_h_l_07_11,
     sp4_h_l_07_12, sp4_h_l_07_13, sp4_h_l_07_14, sp4_h_l_07_15,
     sp4_h_l_07_16, sp4_h_l_07_17, sp4_h_r_13_09, sp4_v_b_07_09,
     sp4_v_b_07_10, sp4_v_b_07_11, sp4_v_b_07_12, sp4_v_b_07_13,
     sp4_v_b_07_14, sp4_v_b_07_15, sp4_v_b_07_16, sp4_v_b_08_09,
     sp4_v_b_09_09, sp4_v_b_10_09, sp4_v_b_11_09, sp4_v_b_12_09,
     sp12_h_l_07_09, sp12_h_l_07_10, sp12_h_l_07_11, sp12_h_l_07_12,
     sp12_h_l_07_13, sp12_h_l_07_14, sp12_h_l_07_15, sp12_h_l_07_16,
     sp12_v_b_07_09, sp12_v_b_08_09, sp12_v_b_09_09, sp12_v_b_10_09,
     sp12_v_b_11_09, sp12_v_b_12_09, vdd_cntl_r, wl_r, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_07_09,
     bnl_op_08_09, bnl_op_09_09, bnl_op_10_09, bnl_op_11_09,
     bnl_op_12_09, bnl_op_13_09, bnr_op_07_09, bnr_op_08_09,
     bnr_op_09_09, bnr_op_10_09, bnr_op_11_09, bnr_op_12_09,
     bot_op_07_09, bot_op_08_09, bot_op_09_09, bot_op_10_09,
     bot_op_11_09, bot_op_12_09, bs_en_i, carry_in_07_09,
     carry_in_08_09, carry_in_09_09, carry_in_11_09, carry_in_12_09,
     ceb_i, glb_in, hiz_b_i, hold_r_t, hold_t_r, lc_bot_07_09,
     lc_bot_08_09, lc_bot_09_09, lc_bot_11_09, lc_bot_12_09,
     lft_op_07_09, lft_op_07_10, lft_op_07_11, lft_op_07_12,
     lft_op_07_13, lft_op_07_14, lft_op_07_15, lft_op_07_16, mode_i,
     padin_r, padin_t_r, prog, purst, r_i, sdi, shift_i, tclk_i,
     tnl_op_07_16, update_i );
output  bs_en_o, ceb_o, fabric_out_07_17, fabric_out_08_17,
     fabric_out_13_09, fabric_out_13_10, hiz_b_o, mode_o, padin_07_17a,
     padin_13_09a, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, carry_in_07_09, carry_in_08_09,
     carry_in_09_09, carry_in_11_09, carry_in_12_09, ceb_i, hiz_b_i,
     hold_r_t, hold_t_r, lc_bot_07_09, lc_bot_08_09, lc_bot_09_09,
     lc_bot_11_09, lc_bot_12_09, mode_i, prog, purst, r_i, sdi,
     shift_i, tclk_i, update_i;

output [23:12]  pado_t_r;
output [7:0]  slf_op_07_15;
output [7:0]  slf_op_08_09;
output [143:0]  cf_t;
output [191:0]  cf_r;
output [3:0]  slf_op_07_17;
output [23:12]  padeb_t_r;
output [3:0]  slf_op_13_09;
output [7:0]  slf_op_07_10;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_12_09;
output [7:0]  slf_op_07_11;
output [7:0]  slf_op_07_09;
output [7:0]  slf_op_07_12;
output [24:13]  padeb_r;
output [10:0]  bm_ab_2bot;
output [24:13]  pado_r;
output [7:0]  slf_op_07_13;
output [7:0]  slf_op_10_09;
output [10:0]  bm_aa_2bot;
output [7:0]  slf_op_07_16;
output [7:0]  slf_op_11_09;
output [7:0]  slf_op_09_09;
output [7:0]  slf_op_07_14;

inout [23:0]  sp12_v_b_11_09;
inout [47:0]  sp4_v_b_11_09;
inout [23:0]  sp12_h_l_07_15;
inout [47:0]  sp4_v_b_07_16;
inout [47:0]  sp4_h_l_07_09;
inout [47:0]  sp4_h_l_07_12;
inout [47:0]  sp4_h_l_07_13;
inout [47:0]  sp4_h_l_07_14;
inout [23:0]  sp12_v_b_10_09;
inout [23:0]  sp12_h_l_07_16;
inout [23:0]  sp12_v_b_07_09;
inout [47:0]  sp4_v_b_09_09;
inout [47:0]  sp4_v_b_07_10;
inout [47:0]  sp4_v_b_10_09;
inout [23:0]  sp12_v_b_09_09;
inout [23:0]  sp12_h_l_07_14;
inout [143:0]  wl_r;
inout [143:0]  vdd_cntl_r;
inout [23:0]  sp12_v_b_12_09;
inout [47:0]  sp4_v_b_07_12;
inout [15:0]  sp4_h_l_07_17;
inout [47:0]  sp4_h_l_07_16;
inout [47:0]  sp4_v_b_07_14;
inout [23:0]  sp12_h_l_07_10;
inout [47:0]  sp4_v_b_07_11;
inout [47:0]  sp4_v_b_07_15;
inout [23:0]  sp12_h_l_07_11;
inout [47:0]  sp4_h_l_07_15;
inout [143:0]  pgate_r;
inout [143:0]  reset_b_r;
inout [23:0]  sp12_h_l_07_12;
inout [47:0]  sp4_v_b_12_09;
inout [23:0]  sp12_h_l_07_09;
inout [47:0]  sp4_h_l_07_10;
inout [15:0]  sp4_h_r_13_09;
inout [23:0]  sp12_v_b_08_09;
inout [47:0]  sp4_v_b_07_09;
inout [23:0]  sp12_h_l_07_13;
inout [47:0]  sp4_h_l_07_11;
inout [47:0]  sp4_v_b_07_13;
inout [47:0]  sp4_v_b_08_09;
inout [329:0]  bl;

input [7:0]  bnl_op_13_09;
input [1:0]  bm_sweb_i;
input [7:0]  bnl_op_12_09;
input [7:0]  bnr_op_08_09;
input [7:0]  bot_op_12_09;
input [1:0]  bm_sclkrw_i;
input [7:0]  bm_sa_i;
input [7:0]  bnr_op_07_09;
input [7:0]  bnr_op_12_09;
input [7:0]  lft_op_07_13;
input [1:0]  bm_sdi_i;
input [7:0]  bnl_op_11_09;
input [7:0]  bnl_op_07_09;
input [7:0]  bnr_op_10_09;
input [7:0]  bot_op_09_09;
input [24:13]  padin_r;
input [7:0]  bot_op_11_09;
input [7:0]  bot_op_10_09;
input [7:0]  lft_op_07_15;
input [7:0]  lft_op_07_11;
input [7:0]  lft_op_07_16;
input [7:0]  lft_op_07_14;
input [7:0]  bot_op_08_09;
input [7:0]  bnr_op_09_09;
input [7:0]  bnl_op_08_09;
input [7:0]  lft_op_07_09;
input [23:12]  padin_t_r;
input [7:0]  bnl_op_09_09;
input [7:0]  lft_op_07_10;
input [7:0]  bnr_op_11_09;
input [3:0]  tnl_op_07_16;
input [7:0]  lft_op_07_12;
input [7:0]  glb_in;
input [7:0]  bot_op_07_09;
input [7:0]  bnl_op_10_09;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:23]  net1153;

wire  [3:0]  slf_op_13_16;

wire  [3:0]  slf_op_13_12;

wire  [3:0]  slf_op_13_14;

wire  [0:0]  padinlat_t_r;

wire  [0:23]  net1014;

wire  [3:0]  slf_op_13_15;

wire  [0:47]  net1114;

wire  [3:0]  slf_op_13_10;

wire  [3:0]  slf_op_10_17;

wire  [3:0]  slf_op_08_17;

wire  [7:0]  clk_center;

wire  [7:0]  clk_tree_drv_tr;

wire  [3:0]  slf_op_12_17;

wire  [3:0]  slf_op_09_17;

wire  [1:0]  bm_sdi_b1_o;

wire  [3:0]  slf_op_11_17;

wire  [3:0]  slf_op_13_11;

wire  [3:0]  slf_op_13_13;

wire  [0:7]  net1224;

wire  [0:47]  net1111;

wire  [0:47]  net1365;

wire  [0:47]  net1400;

wire  [0:23]  net870;

wire  [0:7]  net1004;

wire  [0:47]  net938;

wire  [0:47]  net1157;

wire  [0:47]  net1402;

wire  [0:7]  net1405;

wire  [0:7]  net1190;

wire  [0:23]  net921;

wire  [0:47]  net996;

wire  [0:47]  net1067;

wire  [0:47]  net1220;

wire  [0:47]  net1032;

wire  [0:7]  net943;

wire  [0:23]  net1056;

wire  [0:23]  net1200;

wire  [0:47]  net1183;

wire  [0:47]  net1369;

wire  [0:7]  net1141;

wire  [0:47]  net1184;

wire  [0:23]  net1341;

wire  [0:47]  net879;

wire  [0:23]  net1107;

wire  [0:47]  net1430;

wire  [0:7]  net1407;

wire  [0:23]  net1150;

wire  [0:23]  net1297;

wire  [0:23]  net1109;

wire  [0:47]  net1252;

wire  [0:7]  net1284;

wire  [0:23]  net1108;

wire  [0:7]  net1130;

wire  [0:47]  net1368;

wire  [0:47]  net1062;

wire  [0:7]  net1227;

wire  [0:47]  net1090;

wire  [0:47]  net994;

wire  [0:47]  net1088;

wire  [0:47]  net1257;

wire  [0:47]  net1158;

wire  [0:47]  net1314;

wire  [0:23]  net965;

wire  [0:47]  net1069;

wire  [0:47]  net899;

wire  [0:47]  net1301;

wire  [0:47]  net973;

wire  [0:7]  net1131;

wire  [0:47]  net1431;

wire  [0:23]  net1377;

wire  [0:7]  net1097;

wire  [0:47]  net1020;

wire  [0:7]  net1225;

wire  [0:7]  net1191;

wire  [0:7]  net1098;

wire  [0:47]  net822;

wire  [0:47]  net1063;

wire  [0:47]  net1255;

wire  [0:47]  net1156;

wire  [0:7]  net813;

wire  [0:7]  net1192;

wire  [0:1]  net1387;

wire  [0:47]  net1019;

wire  [0:23]  net1013;

wire  [0:7]  net1095;

wire  [0:47]  net975;

wire  [0:47]  net817;

wire  [0:23]  net963;

wire  [0:7]  net1003;

wire  [0:7]  net1133;

wire  [0:47]  net1383;

wire  [0:47]  net1163;

wire  [0:23]  net934;

wire  [0:47]  net1432;

wire  [0:47]  net900;

wire  [0:47]  net824;

wire  [0:47]  net974;

wire  [0:23]  net918;

wire  [0:47]  net1256;

wire  [0:7]  net1408;

wire  [0:7]  net01228;

wire  [0:7]  net1047;

wire  [0:23]  net1151;

wire  [0:47]  net968;

wire  [0:47]  net995;

wire  [0:23]  net1393;

wire  [0:7]  net0848;

wire  [0:47]  net1361;

wire  [0:47]  net1428;

wire  [0:23]  net1216;

wire  [0:47]  net1207;

wire  [0:47]  net1161;

wire  [0:47]  net993;

wire  [0:47]  net972;

wire  [0:47]  net1087;

wire  [0:23]  net1244;

wire  [0:47]  net881;

wire  [0:23]  net868;

wire  [0:47]  net902;

wire  [0:47]  net1113;

wire  [0:7]  net953;

wire  [0:23]  net1294;

wire  [0:23]  net1201;

wire  [0:47]  net1371;

wire  [0:23]  net1386;

wire  [0:7]  net1039;

wire  [0:23]  net1106;

wire  [0:23]  net1059;

wire  [0:23]  net1245;

wire  [0:47]  net1182;

wire  [0:7]  net1318;

wire  [0:47]  net970;

wire  [0:7]  net1189;

wire  [0:47]  net1278;

wire  [0:47]  net0885;

wire  [0:47]  net1300;

wire  [0:7]  net1410;

wire  [0:47]  net878;

wire  [0:47]  net1160;

wire  [0:47]  net1018;

wire  [0:23]  net1203;

wire  [0:7]  net1285;

wire  [0:47]  net1427;

wire  [0:47]  net0882;

wire  [0:23]  net1355;

wire  [0:47]  net1089;

wire  [0:1]  net1380;

wire  [0:7]  net1404;

wire  [0:23]  net964;

wire  [0:47]  net1162;

wire  [0:23]  net1246;

wire  [0:47]  net1068;

wire  [0:23]  net1353;

wire  [0:23]  net1015;

wire  [0:47]  net1299;

wire  [0:7]  net01133;

wire  [0:7]  net1096;

wire  [0:23]  net1122;

wire  [0:47]  net820;

wire  [0:7]  net1036;

wire  [0:23]  net869;

wire  [0:47]  net1302;

wire  [0:15]  net793;

wire  [0:47]  net1254;

wire  [0:7]  net942;

wire  [0:47]  net821;

wire  [0:7]  net1001;

wire  [0:7]  net1409;

wire  [0:47]  net1372;

wire  [0:47]  net1205;

wire  [0:47]  net1275;

wire  [0:23]  net1385;

wire  [0:23]  net1295;

wire  [0:47]  net880;

wire  [0:7]  net1283;

wire  [0:47]  net1401;

wire  [0:23]  net1058;

wire  [0:47]  net1276;

wire  [0:47]  net1206;

wire  [0:7]  net01038;

wire  [0:7]  net1037;

wire  [0:47]  net1181;

wire  [0:23]  net919;

wire  [0:23]  net1202;

wire  [0:47]  net1017;

wire  [0:7]  net1423;

wire  [0:23]  net1152;

wire  [0:47]  net1064;

wire  [0:47]  net901;

wire  [0:7]  net1286;

wire  [0:7]  net1406;

wire  [0:47]  net1429;

wire  [0:7]  net1002;

wire  [0:23]  net1310;

wire  [0:23]  net1358;

wire  [0:47]  net1208;

wire  [0:47]  net969;

wire  [0:47]  net1250;

wire  [0:23]  net871;

wire  [0:47]  net1251;

wire  [0:23]  net1296;

wire  [0:7]  net1235;

wire  [0:23]  net1012;

wire  [0:47]  net1126;

wire  [0:23]  net1057;

wire  [0:7]  net1422;

wire  [0:23]  net1357;

wire  [0:7]  net0943;

wire  [0:23]  net1247;

wire  [0:23]  net1028;

wire  [0:23]  net920;

wire  [0:47]  net1066;

wire  [0:23]  net962;

wire  [0:47]  net823;

wire  [0:7]  net945;

wire  [0:47]  net1112;

wire  [0:47]  net1277;



bram1x4_ice1f I_lt_col_t10 ( .glb_netwk_top(net1423[0:7]), .prog(prog),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .reset_b(reset_b_r[127:0]), .bm_wdummymux_en_o(net1328),
     .bm_sreb_o(net1329), .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(net809),
     .bm_sa_o(net813[0:7]), .bm_rcapmux_en_o(net1333),
     .bm_init_o(net814), .lft_op_05(net1192[0:7]), .bl(bl[203:162]),
     .sp4_h_l_06(net995[0:47]), .sp12_h_l_02(net964[0:23]),
     .lft_op_06(net1191[0:7]), .sp12_h_l_03(net963[0:23]),
     .sp12_h_r_03(net1341[0:23]), .sp12_h_l_01(net965[0:23]),
     .sp4_v_b_04(net968[0:47]), .sp4_v_b_05(net1017[0:47]),
     .lft_op_07(net1190[0:7]), .sp4_v_b_06(net1018[0:47]),
     .sp4_v_b_08(net1020[0:47]), .sp4_v_b_07(net1019[0:47]),
     .lft_op_03(net1131[0:7]), .lft_op_01(slf_op_09_09[7:0]),
     .sp4_h_l_02(net974[0:47]), .sp12_h_l_06(net1013[0:23]),
     .sp12_h_r_07(net1353[0:23]), .sp12_h_l_05(net1012[0:23]),
     .sp12_h_r_06(net1355[0:23]), .sp12_h_l_04(net962[0:23]),
     .sp12_h_r_05(net1357[0:23]), .sp12_h_r_08(net1358[0:23]),
     .sp12_h_l_07(net1014[0:23]), .sp12_h_l_08(net1015[0:23]),
     .sp4_r_v_b_03(net1361[0:47]), .vdd_cntl(vdd_cntl_r[127:0]),
     .pgate(pgate_r[127:0]), .bot_op_01(bot_op_10_09[7:0]),
     .sp4_r_v_b_04(net1365[0:47]), .sp4_v_b_01(sp4_v_b_10_09[47:0]),
     .sp4_v_b_03(net969[0:47]), .sp4_h_r_08(net1368[0:47]),
     .sp4_r_v_b_05(net1369[0:47]), .sp4_v_b_02(net970[0:47]),
     .sp4_v_t_08(net1371[0:47]), .sp4_r_v_b_02(net1372[0:47]),
     .bnr_op_01(bnr_op_10_09[7:0]), .bm_sdi_o(bm_sdi_b1_o[1:0]),
     .sp4_h_l_04(net972[0:47]), .lft_op_08(net1189[0:7]),
     .sp12_h_r_01(net1377[0:23]), .bm_sdo_i({tiegnd_bram_t,
     bm_sdi_b1_o[0]}), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sweb_o(net1380[0:1]), .sp4_h_l_03(net973[0:47]),
     .sp4_h_l_01(net975[0:47]), .sp4_h_r_01(net1383[0:47]),
     .tnr_op_08({slf_op_11_17[3], slf_op_11_17[2], slf_op_11_17[1],
     slf_op_11_17[0], slf_op_11_17[3], slf_op_11_17[2],
     slf_op_11_17[1], slf_op_11_17[0]}), .sp12_h_r_02(net1385[0:23]),
     .sp12_h_r_04(net1386[0:23]), .bm_sclkrw_o(net1387[0:1]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .lft_op_02(net1133[0:7]),
     .lft_op_04(net1141[0:7]), .bm_sweb_i(bm_sweb_i[1:0]),
     .bnl_op_01(bnl_op_10_09[7:0]), .sp12_v_t_08(net1393[0:23]),
     .wl(wl_r[127:0]), .tnl_op_08({slf_op_09_17[3], slf_op_09_17[2],
     slf_op_09_17[1], slf_op_09_17[0], slf_op_09_17[3],
     slf_op_09_17[2], slf_op_09_17[1], slf_op_09_17[0]}),
     .top_op_08({slf_op_10_17[3], slf_op_10_17[2], slf_op_10_17[1],
     slf_op_10_17[0], slf_op_10_17[3], slf_op_10_17[2],
     slf_op_10_17[1], slf_op_10_17[0]}), .bm_ab_2bot(bm_ab_2bot[10:0]),
     .bm_aa_2bot(bm_aa_2bot[10:0]), .sp12_v_b_01(sp12_v_b_10_09[23:0]),
     .sp4_r_v_b_08(net1400[0:47]), .sp4_r_v_b_07(net1401[0:47]),
     .sp4_r_v_b_06(net1402[0:47]), .sp4_r_v_b_01(sp4_v_b_11_09[47:0]),
     .rgt_op_08(net1404[0:7]), .rgt_op_07(net1405[0:7]),
     .rgt_op_06(net1406[0:7]), .rgt_op_05(net1407[0:7]),
     .rgt_op_04(net1408[0:7]), .rgt_op_03(net1409[0:7]),
     .rgt_op_02(net1410[0:7]), .rgt_op_01(slf_op_11_09[7:0]),
     .slf_op_02(net945[0:7]), .slf_op_01(slf_op_10_09[7:0]),
     .slf_op_03(net943[0:7]), .slf_op_04(net953[0:7]),
     .slf_op_05(net1004[0:7]), .slf_op_06(net1003[0:7]),
     .slf_op_07(net1002[0:7]), .slf_op_08(net1001[0:7]),
     .bm_ab_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .bm_aa_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .glb_netwk_bot(net1422[0:7]), .sp4_h_l_08(net993[0:47]),
     .sp4_h_l_07(net994[0:47]), .sp4_h_l_05(net996[0:47]),
     .sp4_h_r_02(net1427[0:47]), .sp4_h_r_03(net1428[0:47]),
     .sp4_h_r_04(net1429[0:47]), .sp4_h_r_05(net1430[0:47]),
     .sp4_h_r_06(net1431[0:47]), .sp4_h_r_07(net1432[0:47]));
fabric_buf_ice8p I461 ( .f_in(net01448), .f_out(padin_13_09a));
fabric_buf_ice8p I_fabric_buf_8p_r_32 ( .f_in(net_fabric_out_13_09),
     .f_out(fabric_out_13_09));
fabric_buf_ice8p I451 ( .f_in(net_fabric_out_13_10),
     .f_out(fabric_out_13_10));
fabric_buf_ice8p I453 ( .f_in(net_fabric_out_07_17),
     .f_out(fabric_out_07_17));
fabric_buf_ice8p I454 ( .f_in(padinlat_t_r[0]), .f_out(padin_07_17a));
fabric_buf_ice8p I452 ( .f_in(net_fabric_out_08_17),
     .f_out(fabric_out_08_17));
io_rgt_top_1x8_ice1f I_lt_col_t13 ( .cf_r(cf_r[191:0]),
     .shift(shift_i), .bs_en(bs_en_i), .mode(mode_i), .sdi(sdi),
     .hiz_b(hiz_b_i), .prog(prog), .hold(hold_r_t), .update(update_i),
     .r(r_i), .SP4_h_l_05(net902[0:47]), .slf_op_05(slf_op_13_13[3:0]),
     .slf_op_01(slf_op_13_09[3:0]), .slf_op_06(slf_op_13_14[3:0]),
     .slf_op_02(slf_op_13_10[3:0]), .sdo(net680), .bl(bl[329:312]),
     .tclk(tclk_i), .reset_b(reset_b_r[127:0]),
     .lft_op_07(net1096[0:7]), .SP4_h_l_06(net901[0:47]),
     .sp4_v_t_08(net793[0:15]), .slf_op_04(slf_op_13_12[3:0]),
     .slf_op_03(slf_op_13_11[3:0]), .slf_op_07(slf_op_13_15[3:0]),
     .slf_op_08(slf_op_13_16[3:0]), .SP4_h_l_08(net899[0:47]),
     .SP4_h_l_07(net900[0:47]), .SP4_h_l_03(net879[0:47]),
     .SP4_h_l_04(net878[0:47]), .SP4_h_l_02(net880[0:47]),
     .SP4_h_l_01(net881[0:47]), .lft_op_04(net1047[0:7]),
     .lft_op_06(net1097[0:7]), .lft_op_01(slf_op_12_09[7:0]),
     .lft_op_08(net1095[0:7]), .lft_op_02(net1039[0:7]),
     .pgate(pgate_r[127:0]), .vdd_cntl(vdd_cntl_r[127:0]),
     .tnl_op_08({slf_op_12_17[3], slf_op_12_17[2], slf_op_12_17[1],
     slf_op_12_17[0], slf_op_12_17[3], slf_op_12_17[2],
     slf_op_12_17[1], slf_op_12_17[0]}), .wl(wl_r[127:0]),
     .tclk_o(net707), .ceb(ceb_i),
     .fabric_out_09(net_fabric_out_13_09), .SP12_h_l_02(net870[0:23]),
     .SP12_h_l_04(net868[0:23]), .SP12_h_l_08(net921[0:23]),
     .SP12_h_l_06(net919[0:23]), .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .SP12_h_l_05(net918[0:23]), .SP12_h_l_01(net871[0:23]),
     .SP12_h_l_03(net869[0:23]), .SP12_h_l_07(net920[0:23]),
     .fabric_out_10(net_fabric_out_13_10), .padin(padin_r[24:13]),
     .pado(pado_r[24:13]), .padeb(padeb_r[24:13]),
     .lft_op_03(net1037[0:7]), .bnl_op_13_09(bnl_op_13_09[7:0]),
     .lft_op_05(net1098[0:7]), .sp4_v_b_13_09(sp4_h_r_13_09[15:0]));
io_top_rgt_1x6_ice1f I_preio_top_l ( .pado_t_r(pado_t_r[23:12]),
     .padeb_t_r(padeb_t_r[23:12]), .padin_t_r(padin_t_r[23:12]),
     .cf_t(cf_t[143:0]), .fabric_out_08_17(net_fabric_out_08_17),
     .hold_t_r(hold_t_r), .wl_l({wl_r[142], wl_r[143], wl_r[141],
     wl_r[140], wl_r[138], wl_r[139], wl_r[137], wl_r[136], wl_r[134],
     wl_r[135], wl_r[133], wl_r[132], wl_r[130], wl_r[131], wl_r[129],
     wl_r[128]}), .lft_op_01_17(slf_op_07_16[7:0]),
     .vdd_cntl_l({vdd_cntl_r[142], vdd_cntl_r[143], vdd_cntl_r[141],
     vdd_cntl_r[140], vdd_cntl_r[138], vdd_cntl_r[139],
     vdd_cntl_r[137], vdd_cntl_r[136], vdd_cntl_r[134],
     vdd_cntl_r[135], vdd_cntl_r[133], vdd_cntl_r[132],
     vdd_cntl_r[130], vdd_cntl_r[131], vdd_cntl_r[129],
     vdd_cntl_r[128]}), .update_i(net736), .tclk_i(net737),
     .shift_i(net738), .sdi(net739), .reset_l({reset_b_r[142],
     reset_b_r[143], reset_b_r[141], reset_b_r[140], reset_b_r[138],
     reset_b_r[139], reset_b_r[137], reset_b_r[136], reset_b_r[134],
     reset_b_r[135], reset_b_r[133], reset_b_r[132], reset_b_r[130],
     reset_b_r[131], reset_b_r[129], reset_b_r[128]}), .r_i(net741),
     .prog(prog), .pgate_l({pgate_r[142], pgate_r[143], pgate_r[141],
     pgate_r[140], pgate_r[138], pgate_r[139], pgate_r[137],
     pgate_r[136], pgate_r[134], pgate_r[135], pgate_r[133],
     pgate_r[132], pgate_r[130], pgate_r[131], pgate_r[129],
     pgate_r[128]}), .mode_i(net744), .hiz_b_i(net745),
     .bs_en_i(net746), .update_o(update_o), .tclk_o(tclk_o),
     .shift_o(shift_o), .sdo(sdo), .r_o(r_o), .mode_o(mode_o),
     .hiz_b_o(hiz_b_o), .glb_net_06(net942[0:7]),
     .glb_net_05(net1130[0:7]), .glb_net_04(net1423[0:7]),
     .glb_net_03(net1036[0:7]), .glb_net_02(net1224[0:7]),
     .glb_net_01(net1318[0:7]), .bs_en_o(bs_en_o), .bl_06(bl[311:258]),
     .bl_05(bl[257:204]), .bl_02(bl[107:54]), .bl_01(bl[53:0]),
     .lft_op_03_17(net1189[0:7]), .sp4_v_b_04_17(net1371[0:47]),
     .lft_op_02_17(net1283[0:7]), .lft_op_04_17(net1001[0:7]),
     .sp4_v_b_06_17(net938[0:47]), .sp12_v_b_04_17(net1393[0:23]),
     .sp4_v_b_02_17(net1220[0:47]), .sp12_v_b_05_17(net1122[0:23]),
     .lft_op_06_17(net1095[0:7]), .slf_op_04_17(slf_op_10_17[3:0]),
     .sp4_v_b_05_17(net1126[0:47]), .sp12_v_b_03_17(net1028[0:23]),
     .slf_op_01_17(slf_op_07_17[3:0]), .sp4_v_b_01_17(net1314[0:47]),
     .sp4_v_b_03_17(net1032[0:47]), .slf_op_03_17(slf_op_09_17[3:0]),
     .lft_op_05_17(net1404[0:7]), .sp12_v_b_01_17(net1310[0:23]),
     .slf_op_06_17(slf_op_12_17[3:0]), .sp12_v_b_06_17(net934[0:23]),
     .slf_op_02_17(slf_op_08_17[3:0]), .sp12_v_b_02_17(net1216[0:23]),
     .bl_03(bl[161:108]), .bl_04(bl[203:162]), .ceb_o(ceb_o),
     .slf_op_05_17(slf_op_11_17[3:0]), .ceb_i(net791),
     .fabric_out_07_17(net_fabric_out_07_17),
     .sp4_h_r_12_17(net793[0:15]), .bnr_op_12_17({slf_op_13_16[3],
     slf_op_13_16[2], slf_op_13_16[1], slf_op_13_16[0],
     slf_op_13_16[3], slf_op_13_16[2], slf_op_13_16[1],
     slf_op_13_16[0]}), .sp4_h_l_07_17(sp4_h_l_07_17[15:0]),
     .bnl_op_07_17(lft_op_07_16[7:0]));
clk_quad_buf_x8_ice8p I428 ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));
clk_quad_buf_x8_ice8p I427 ( .clko(clk_tree_drv_tr[7:0]),
     .clki(clk_center[7:0]));
scan_buf_ice8p I446 ( .update_i(update_i), .tclk_i(net707),
     .shift_i(shift_i), .sdi(net680), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net736), .tclk_o(net737), .shift_o(net738),
     .sdo(net739), .r_o(net741), .mode_o(net744), .hiz_b_o(net745),
     .ceb_o(net791), .bs_en_o(net746));
tielo I430 ( .tielo(tiegnd_bram_t));
tielo I450 ( .tielo(net848));
lt_1x8_top_ice1f I_lt_col_t12 ( .glb_netwk_b(net0848[0:7]),
     .rgt_op_03({slf_op_13_11[3], slf_op_13_11[2], slf_op_13_11[1],
     slf_op_13_11[0], slf_op_13_11[3], slf_op_13_11[2],
     slf_op_13_11[1], slf_op_13_11[0]}), .slf_op_02(net1039[0:7]),
     .rgt_op_02({slf_op_13_10[3], slf_op_13_10[2], slf_op_13_10[1],
     slf_op_13_10[0], slf_op_13_10[3], slf_op_13_10[2],
     slf_op_13_10[1], slf_op_13_10[0]}), .rgt_op_01({slf_op_13_09[3],
     slf_op_13_09[2], slf_op_13_09[1], slf_op_13_09[0],
     slf_op_13_09[3], slf_op_13_09[2], slf_op_13_09[1],
     slf_op_13_09[0]}), .purst(purst), .prog(prog),
     .lft_op_04(net1408[0:7]), .lft_op_03(net1409[0:7]),
     .lft_op_02(net1410[0:7]), .lft_op_01(slf_op_11_09[7:0]),
     .rgt_op_04({slf_op_13_12[3], slf_op_13_12[2], slf_op_13_12[1],
     slf_op_13_12[0], slf_op_13_12[3], slf_op_13_12[2],
     slf_op_13_12[1], slf_op_13_12[0]}), .carry_in(carry_in_12_09),
     .bnl_op_01(bnl_op_12_09[7:0]), .slf_op_04(net1047[0:7]),
     .slf_op_03(net1037[0:7]), .slf_op_01(slf_op_12_09[7:0]),
     .sp4_h_l_04(net1066[0:47]), .carry_out(net866),
     .vdd_cntl(vdd_cntl_r[127:0]), .sp12_h_r_04(net868[0:23]),
     .sp12_h_r_03(net869[0:23]), .sp12_h_r_02(net870[0:23]),
     .sp12_h_r_01(net871[0:23]), .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_12_09[47:0]), .sp4_r_v_b_04(net0882[0:47]),
     .sp4_r_v_b_03(net820[0:47]), .sp4_r_v_b_02(net817[0:47]),
     .sp4_r_v_b_01(net0885[0:47]), .sp4_h_r_04(net878[0:47]),
     .sp4_h_r_03(net879[0:47]), .sp4_h_r_02(net880[0:47]),
     .sp4_h_r_01(net881[0:47]), .sp4_h_l_03(net1067[0:47]),
     .sp4_h_l_02(net1068[0:47]), .sp4_h_l_01(net1069[0:47]),
     .bl(bl[311:258]), .bot_op_01(bot_op_12_09[7:0]),
     .sp12_h_l_01(net1059[0:23]), .sp12_h_l_02(net1058[0:23]),
     .sp12_h_l_03(net1057[0:23]), .sp12_h_l_04(net1056[0:23]),
     .sp4_v_b_04(net1062[0:47]), .sp4_v_b_03(net1063[0:47]),
     .sp4_v_b_02(net1064[0:47]), .bnr_op_01(bnr_op_12_09[7:0]),
     .sp4_h_l_05(net1090[0:47]), .sp4_h_l_06(net1089[0:47]),
     .sp4_h_l_07(net1088[0:47]), .sp4_h_l_08(net1087[0:47]),
     .sp4_h_r_08(net899[0:47]), .sp4_h_r_07(net900[0:47]),
     .sp4_h_r_06(net901[0:47]), .sp4_h_r_05(net902[0:47]),
     .slf_op_05(net1098[0:7]), .slf_op_06(net1097[0:7]),
     .slf_op_07(net1096[0:7]), .slf_op_08(net1095[0:7]),
     .rgt_op_08({slf_op_13_16[3], slf_op_13_16[2], slf_op_13_16[1],
     slf_op_13_16[0], slf_op_13_16[3], slf_op_13_16[2],
     slf_op_13_16[1], slf_op_13_16[0]}), .rgt_op_07({slf_op_13_15[3],
     slf_op_13_15[2], slf_op_13_15[1], slf_op_13_15[0],
     slf_op_13_15[3], slf_op_13_15[2], slf_op_13_15[1],
     slf_op_13_15[0]}), .rgt_op_06({slf_op_13_14[3], slf_op_13_14[2],
     slf_op_13_14[1], slf_op_13_14[0], slf_op_13_14[3],
     slf_op_13_14[2], slf_op_13_14[1], slf_op_13_14[0]}),
     .rgt_op_05({slf_op_13_13[3], slf_op_13_13[2], slf_op_13_13[1],
     slf_op_13_13[0], slf_op_13_13[3], slf_op_13_13[2],
     slf_op_13_13[1], slf_op_13_13[0]}), .lft_op_08(net1404[0:7]),
     .lft_op_07(net1405[0:7]), .lft_op_06(net1406[0:7]),
     .lft_op_05(net1407[0:7]), .sp12_h_l_08(net1109[0:23]),
     .sp12_h_l_07(net1108[0:23]), .sp12_h_l_06(net1107[0:23]),
     .sp12_h_r_05(net918[0:23]), .sp12_h_r_06(net919[0:23]),
     .sp12_h_r_07(net920[0:23]), .sp12_h_r_08(net921[0:23]),
     .sp12_h_l_05(net1106[0:23]), .sp4_r_v_b_05(net824[0:47]),
     .sp4_r_v_b_06(net823[0:47]), .sp4_r_v_b_07(net821[0:47]),
     .sp4_r_v_b_08(net822[0:47]), .sp4_v_b_08(net1114[0:47]),
     .sp4_v_b_07(net1113[0:47]), .sp4_v_b_06(net1112[0:47]),
     .sp4_v_b_05(net1111[0:47]), .pgate(pgate_r[127:0]),
     .reset_b(reset_b_r[127:0]), .wl(wl_r[127:0]),
     .sp12_v_t_08(net934[0:23]), .tnr_op_08({net848, net848, net848,
     net848, net848, net848, net848, net848}),
     .top_op_08({slf_op_12_17[3], slf_op_12_17[2], slf_op_12_17[1],
     slf_op_12_17[0], slf_op_12_17[3], slf_op_12_17[2],
     slf_op_12_17[1], slf_op_12_17[0]}), .tnl_op_08({slf_op_11_17[3],
     slf_op_11_17[2], slf_op_11_17[1], slf_op_11_17[0],
     slf_op_11_17[3], slf_op_11_17[2], slf_op_11_17[1],
     slf_op_11_17[0]}), .sp4_v_t_08(net938[0:47]),
     .lc_bot(lc_bot_12_09), .op_vic(net940),
     .sp12_v_b_01(sp12_v_b_12_09[23:0]), .glb_netwk_t(net942[0:7]));
lt_1x8_top_ice1f I_lt_col_t09 ( .glb_netwk_b(net0943[0:7]),
     .rgt_op_03(net943[0:7]), .slf_op_02(net1133[0:7]),
     .rgt_op_02(net945[0:7]), .rgt_op_01(slf_op_10_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net1235[0:7]),
     .lft_op_03(net1225[0:7]), .lft_op_02(net1227[0:7]),
     .lft_op_01(slf_op_08_09[7:0]), .rgt_op_04(net953[0:7]),
     .carry_in(carry_in_09_09), .bnl_op_01(bnl_op_09_09[7:0]),
     .slf_op_04(net1141[0:7]), .slf_op_03(net1131[0:7]),
     .slf_op_01(slf_op_09_09[7:0]), .sp4_h_l_04(net1160[0:47]),
     .carry_out(net960), .vdd_cntl(vdd_cntl_r[127:0]),
     .sp12_h_r_04(net962[0:23]), .sp12_h_r_03(net963[0:23]),
     .sp12_h_r_02(net964[0:23]), .sp12_h_r_01(net965[0:23]),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_09_09[47:0]), .sp4_r_v_b_04(net968[0:47]),
     .sp4_r_v_b_03(net969[0:47]), .sp4_r_v_b_02(net970[0:47]),
     .sp4_r_v_b_01(sp4_v_b_10_09[47:0]), .sp4_h_r_04(net972[0:47]),
     .sp4_h_r_03(net973[0:47]), .sp4_h_r_02(net974[0:47]),
     .sp4_h_r_01(net975[0:47]), .sp4_h_l_03(net1161[0:47]),
     .sp4_h_l_02(net1162[0:47]), .sp4_h_l_01(net1163[0:47]),
     .bl(bl[161:108]), .bot_op_01(bot_op_09_09[7:0]),
     .sp12_h_l_01(net1153[0:23]), .sp12_h_l_02(net1152[0:23]),
     .sp12_h_l_03(net1151[0:23]), .sp12_h_l_04(net1150[0:23]),
     .sp4_v_b_04(net1156[0:47]), .sp4_v_b_03(net1157[0:47]),
     .sp4_v_b_02(net1158[0:47]), .bnr_op_01(bnr_op_09_09[7:0]),
     .sp4_h_l_05(net1184[0:47]), .sp4_h_l_06(net1183[0:47]),
     .sp4_h_l_07(net1182[0:47]), .sp4_h_l_08(net1181[0:47]),
     .sp4_h_r_08(net993[0:47]), .sp4_h_r_07(net994[0:47]),
     .sp4_h_r_06(net995[0:47]), .sp4_h_r_05(net996[0:47]),
     .slf_op_05(net1192[0:7]), .slf_op_06(net1191[0:7]),
     .slf_op_07(net1190[0:7]), .slf_op_08(net1189[0:7]),
     .rgt_op_08(net1001[0:7]), .rgt_op_07(net1002[0:7]),
     .rgt_op_06(net1003[0:7]), .rgt_op_05(net1004[0:7]),
     .lft_op_08(net1283[0:7]), .lft_op_07(net1284[0:7]),
     .lft_op_06(net1285[0:7]), .lft_op_05(net1286[0:7]),
     .sp12_h_l_08(net1203[0:23]), .sp12_h_l_07(net1202[0:23]),
     .sp12_h_l_06(net1201[0:23]), .sp12_h_r_05(net1012[0:23]),
     .sp12_h_r_06(net1013[0:23]), .sp12_h_r_07(net1014[0:23]),
     .sp12_h_r_08(net1015[0:23]), .sp12_h_l_05(net1200[0:23]),
     .sp4_r_v_b_05(net1017[0:47]), .sp4_r_v_b_06(net1018[0:47]),
     .sp4_r_v_b_07(net1019[0:47]), .sp4_r_v_b_08(net1020[0:47]),
     .sp4_v_b_08(net1208[0:47]), .sp4_v_b_07(net1207[0:47]),
     .sp4_v_b_06(net1206[0:47]), .sp4_v_b_05(net1205[0:47]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .wl(wl_r[127:0]), .sp12_v_t_08(net1028[0:23]),
     .tnr_op_08({slf_op_10_17[3], slf_op_10_17[2], slf_op_10_17[1],
     slf_op_10_17[0], slf_op_10_17[3], slf_op_10_17[2],
     slf_op_10_17[1], slf_op_10_17[0]}), .top_op_08({slf_op_09_17[3],
     slf_op_09_17[2], slf_op_09_17[1], slf_op_09_17[0],
     slf_op_09_17[3], slf_op_09_17[2], slf_op_09_17[1],
     slf_op_09_17[0]}), .tnl_op_08({slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0], slf_op_08_17[3],
     slf_op_08_17[2], slf_op_08_17[1], slf_op_08_17[0]}),
     .sp4_v_t_08(net1032[0:47]), .lc_bot(lc_bot_09_09),
     .op_vic(net1034), .sp12_v_b_01(sp12_v_b_09_09[23:0]),
     .glb_netwk_t(net1036[0:7]));
lt_1x8_top_ice1f I_lt_col_t11 ( .glb_netwk_b(net01038[0:7]),
     .rgt_op_03(net1037[0:7]), .slf_op_02(net1410[0:7]),
     .rgt_op_02(net1039[0:7]), .rgt_op_01(slf_op_12_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net953[0:7]),
     .lft_op_03(net943[0:7]), .lft_op_02(net945[0:7]),
     .lft_op_01(slf_op_10_09[7:0]), .rgt_op_04(net1047[0:7]),
     .carry_in(carry_in_11_09), .bnl_op_01(bnl_op_11_09[7:0]),
     .slf_op_04(net1408[0:7]), .slf_op_03(net1409[0:7]),
     .slf_op_01(slf_op_11_09[7:0]), .sp4_h_l_04(net1429[0:47]),
     .carry_out(net1054), .vdd_cntl(vdd_cntl_r[127:0]),
     .sp12_h_r_04(net1056[0:23]), .sp12_h_r_03(net1057[0:23]),
     .sp12_h_r_02(net1058[0:23]), .sp12_h_r_01(net1059[0:23]),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_11_09[47:0]), .sp4_r_v_b_04(net1062[0:47]),
     .sp4_r_v_b_03(net1063[0:47]), .sp4_r_v_b_02(net1064[0:47]),
     .sp4_r_v_b_01(sp4_v_b_12_09[47:0]), .sp4_h_r_04(net1066[0:47]),
     .sp4_h_r_03(net1067[0:47]), .sp4_h_r_02(net1068[0:47]),
     .sp4_h_r_01(net1069[0:47]), .sp4_h_l_03(net1428[0:47]),
     .sp4_h_l_02(net1427[0:47]), .sp4_h_l_01(net1383[0:47]),
     .bl(bl[257:204]), .bot_op_01(bot_op_11_09[7:0]),
     .sp12_h_l_01(net1377[0:23]), .sp12_h_l_02(net1385[0:23]),
     .sp12_h_l_03(net1341[0:23]), .sp12_h_l_04(net1386[0:23]),
     .sp4_v_b_04(net1365[0:47]), .sp4_v_b_03(net1361[0:47]),
     .sp4_v_b_02(net1372[0:47]), .bnr_op_01(bnr_op_11_09[7:0]),
     .sp4_h_l_05(net1430[0:47]), .sp4_h_l_06(net1431[0:47]),
     .sp4_h_l_07(net1432[0:47]), .sp4_h_l_08(net1368[0:47]),
     .sp4_h_r_08(net1087[0:47]), .sp4_h_r_07(net1088[0:47]),
     .sp4_h_r_06(net1089[0:47]), .sp4_h_r_05(net1090[0:47]),
     .slf_op_05(net1407[0:7]), .slf_op_06(net1406[0:7]),
     .slf_op_07(net1405[0:7]), .slf_op_08(net1404[0:7]),
     .rgt_op_08(net1095[0:7]), .rgt_op_07(net1096[0:7]),
     .rgt_op_06(net1097[0:7]), .rgt_op_05(net1098[0:7]),
     .lft_op_08(net1001[0:7]), .lft_op_07(net1002[0:7]),
     .lft_op_06(net1003[0:7]), .lft_op_05(net1004[0:7]),
     .sp12_h_l_08(net1358[0:23]), .sp12_h_l_07(net1353[0:23]),
     .sp12_h_l_06(net1355[0:23]), .sp12_h_r_05(net1106[0:23]),
     .sp12_h_r_06(net1107[0:23]), .sp12_h_r_07(net1108[0:23]),
     .sp12_h_r_08(net1109[0:23]), .sp12_h_l_05(net1357[0:23]),
     .sp4_r_v_b_05(net1111[0:47]), .sp4_r_v_b_06(net1112[0:47]),
     .sp4_r_v_b_07(net1113[0:47]), .sp4_r_v_b_08(net1114[0:47]),
     .sp4_v_b_08(net1400[0:47]), .sp4_v_b_07(net1401[0:47]),
     .sp4_v_b_06(net1402[0:47]), .sp4_v_b_05(net1369[0:47]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .wl(wl_r[127:0]), .sp12_v_t_08(net1122[0:23]),
     .tnr_op_08({slf_op_12_17[3], slf_op_12_17[2], slf_op_12_17[1],
     slf_op_12_17[0], slf_op_12_17[3], slf_op_12_17[2],
     slf_op_12_17[1], slf_op_12_17[0]}), .top_op_08({slf_op_11_17[3],
     slf_op_11_17[2], slf_op_11_17[1], slf_op_11_17[0],
     slf_op_11_17[3], slf_op_11_17[2], slf_op_11_17[1],
     slf_op_11_17[0]}), .tnl_op_08({slf_op_10_17[3], slf_op_10_17[2],
     slf_op_10_17[1], slf_op_10_17[0], slf_op_10_17[3],
     slf_op_10_17[2], slf_op_10_17[1], slf_op_10_17[0]}),
     .sp4_v_t_08(net1126[0:47]), .lc_bot(lc_bot_11_09),
     .op_vic(net1128), .sp12_v_b_01(sp12_v_b_11_09[23:0]),
     .glb_netwk_t(net1130[0:7]));
lt_1x8_top_ice1f I_lt_col_t08 ( .glb_netwk_b(net01133[0:7]),
     .rgt_op_03(net1131[0:7]), .slf_op_02(net1227[0:7]),
     .rgt_op_02(net1133[0:7]), .rgt_op_01(slf_op_09_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(slf_op_07_12[7:0]),
     .lft_op_03(slf_op_07_11[7:0]), .lft_op_02(slf_op_07_10[7:0]),
     .lft_op_01(slf_op_07_09[7:0]), .rgt_op_04(net1141[0:7]),
     .carry_in(carry_in_08_09), .bnl_op_01(bnl_op_08_09[7:0]),
     .slf_op_04(net1235[0:7]), .slf_op_03(net1225[0:7]),
     .slf_op_01(slf_op_08_09[7:0]), .sp4_h_l_04(net1254[0:47]),
     .carry_out(net1148), .vdd_cntl(vdd_cntl_r[127:0]),
     .sp12_h_r_04(net1150[0:23]), .sp12_h_r_03(net1151[0:23]),
     .sp12_h_r_02(net1152[0:23]), .sp12_h_r_01(net1153[0:23]),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_08_09[47:0]), .sp4_r_v_b_04(net1156[0:47]),
     .sp4_r_v_b_03(net1157[0:47]), .sp4_r_v_b_02(net1158[0:47]),
     .sp4_r_v_b_01(sp4_v_b_09_09[47:0]), .sp4_h_r_04(net1160[0:47]),
     .sp4_h_r_03(net1161[0:47]), .sp4_h_r_02(net1162[0:47]),
     .sp4_h_r_01(net1163[0:47]), .sp4_h_l_03(net1255[0:47]),
     .sp4_h_l_02(net1256[0:47]), .sp4_h_l_01(net1257[0:47]),
     .bl(bl[107:54]), .bot_op_01(bot_op_08_09[7:0]),
     .sp12_h_l_01(net1247[0:23]), .sp12_h_l_02(net1246[0:23]),
     .sp12_h_l_03(net1245[0:23]), .sp12_h_l_04(net1244[0:23]),
     .sp4_v_b_04(net1250[0:47]), .sp4_v_b_03(net1251[0:47]),
     .sp4_v_b_02(net1252[0:47]), .bnr_op_01(bnr_op_08_09[7:0]),
     .sp4_h_l_05(net1278[0:47]), .sp4_h_l_06(net1277[0:47]),
     .sp4_h_l_07(net1276[0:47]), .sp4_h_l_08(net1275[0:47]),
     .sp4_h_r_08(net1181[0:47]), .sp4_h_r_07(net1182[0:47]),
     .sp4_h_r_06(net1183[0:47]), .sp4_h_r_05(net1184[0:47]),
     .slf_op_05(net1286[0:7]), .slf_op_06(net1285[0:7]),
     .slf_op_07(net1284[0:7]), .slf_op_08(net1283[0:7]),
     .rgt_op_08(net1189[0:7]), .rgt_op_07(net1190[0:7]),
     .rgt_op_06(net1191[0:7]), .rgt_op_05(net1192[0:7]),
     .lft_op_08(slf_op_07_16[7:0]), .lft_op_07(slf_op_07_15[7:0]),
     .lft_op_06(slf_op_07_14[7:0]), .lft_op_05(slf_op_07_13[7:0]),
     .sp12_h_l_08(net1297[0:23]), .sp12_h_l_07(net1296[0:23]),
     .sp12_h_l_06(net1295[0:23]), .sp12_h_r_05(net1200[0:23]),
     .sp12_h_r_06(net1201[0:23]), .sp12_h_r_07(net1202[0:23]),
     .sp12_h_r_08(net1203[0:23]), .sp12_h_l_05(net1294[0:23]),
     .sp4_r_v_b_05(net1205[0:47]), .sp4_r_v_b_06(net1206[0:47]),
     .sp4_r_v_b_07(net1207[0:47]), .sp4_r_v_b_08(net1208[0:47]),
     .sp4_v_b_08(net1302[0:47]), .sp4_v_b_07(net1301[0:47]),
     .sp4_v_b_06(net1300[0:47]), .sp4_v_b_05(net1299[0:47]),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .wl(wl_r[127:0]), .sp12_v_t_08(net1216[0:23]),
     .tnr_op_08({slf_op_09_17[3], slf_op_09_17[2], slf_op_09_17[1],
     slf_op_09_17[0], slf_op_09_17[3], slf_op_09_17[2],
     slf_op_09_17[1], slf_op_09_17[0]}), .top_op_08({slf_op_08_17[3],
     slf_op_08_17[2], slf_op_08_17[1], slf_op_08_17[0],
     slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0]}), .tnl_op_08({slf_op_07_17[3], slf_op_07_17[2],
     slf_op_07_17[1], slf_op_07_17[0], slf_op_07_17[3],
     slf_op_07_17[2], slf_op_07_17[1], slf_op_07_17[0]}),
     .sp4_v_t_08(net1220[0:47]), .lc_bot(lc_bot_08_09),
     .op_vic(net1222), .sp12_v_b_01(sp12_v_b_08_09[23:0]),
     .glb_netwk_t(net1224[0:7]));
lt_1x8_top_ice1f I_lt_col_t07 ( .glb_netwk_b(net01228[0:7]),
     .rgt_op_03(net1225[0:7]), .slf_op_02(slf_op_07_10[7:0]),
     .rgt_op_02(net1227[0:7]), .rgt_op_01(slf_op_08_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(lft_op_07_12[7:0]),
     .lft_op_03(lft_op_07_11[7:0]), .lft_op_02(lft_op_07_10[7:0]),
     .lft_op_01(lft_op_07_09[7:0]), .rgt_op_04(net1235[0:7]),
     .carry_in(carry_in_07_09), .bnl_op_01(bnl_op_07_09[7:0]),
     .slf_op_04(slf_op_07_12[7:0]), .slf_op_03(slf_op_07_11[7:0]),
     .slf_op_01(slf_op_07_09[7:0]), .sp4_h_l_04(sp4_h_l_07_12[47:0]),
     .carry_out(net1242), .vdd_cntl(vdd_cntl_r[127:0]),
     .sp12_h_r_04(net1244[0:23]), .sp12_h_r_03(net1245[0:23]),
     .sp12_h_r_02(net1246[0:23]), .sp12_h_r_01(net1247[0:23]),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_07_09[47:0]), .sp4_r_v_b_04(net1250[0:47]),
     .sp4_r_v_b_03(net1251[0:47]), .sp4_r_v_b_02(net1252[0:47]),
     .sp4_r_v_b_01(sp4_v_b_08_09[47:0]), .sp4_h_r_04(net1254[0:47]),
     .sp4_h_r_03(net1255[0:47]), .sp4_h_r_02(net1256[0:47]),
     .sp4_h_r_01(net1257[0:47]), .sp4_h_l_03(sp4_h_l_07_11[47:0]),
     .sp4_h_l_02(sp4_h_l_07_10[47:0]),
     .sp4_h_l_01(sp4_h_l_07_09[47:0]), .bl(bl[53:0]),
     .bot_op_01(bot_op_07_09[7:0]), .sp12_h_l_01(sp12_h_l_07_09[23:0]),
     .sp12_h_l_02(sp12_h_l_07_10[23:0]),
     .sp12_h_l_03(sp12_h_l_07_11[23:0]),
     .sp12_h_l_04(sp12_h_l_07_12[23:0]),
     .sp4_v_b_04(sp4_v_b_07_12[47:0]),
     .sp4_v_b_03(sp4_v_b_07_11[47:0]),
     .sp4_v_b_02(sp4_v_b_07_10[47:0]), .bnr_op_01(bnr_op_07_09[7:0]),
     .sp4_h_l_05(sp4_h_l_07_13[47:0]),
     .sp4_h_l_06(sp4_h_l_07_14[47:0]),
     .sp4_h_l_07(sp4_h_l_07_15[47:0]),
     .sp4_h_l_08(sp4_h_l_07_16[47:0]), .sp4_h_r_08(net1275[0:47]),
     .sp4_h_r_07(net1276[0:47]), .sp4_h_r_06(net1277[0:47]),
     .sp4_h_r_05(net1278[0:47]), .slf_op_05(slf_op_07_13[7:0]),
     .slf_op_06(slf_op_07_14[7:0]), .slf_op_07(slf_op_07_15[7:0]),
     .slf_op_08(slf_op_07_16[7:0]), .rgt_op_08(net1283[0:7]),
     .rgt_op_07(net1284[0:7]), .rgt_op_06(net1285[0:7]),
     .rgt_op_05(net1286[0:7]), .lft_op_08(lft_op_07_16[7:0]),
     .lft_op_07(lft_op_07_15[7:0]), .lft_op_06(lft_op_07_14[7:0]),
     .lft_op_05(lft_op_07_13[7:0]), .sp12_h_l_08(sp12_h_l_07_16[23:0]),
     .sp12_h_l_07(sp12_h_l_07_15[23:0]),
     .sp12_h_l_06(sp12_h_l_07_14[23:0]), .sp12_h_r_05(net1294[0:23]),
     .sp12_h_r_06(net1295[0:23]), .sp12_h_r_07(net1296[0:23]),
     .sp12_h_r_08(net1297[0:23]), .sp12_h_l_05(sp12_h_l_07_13[23:0]),
     .sp4_r_v_b_05(net1299[0:47]), .sp4_r_v_b_06(net1300[0:47]),
     .sp4_r_v_b_07(net1301[0:47]), .sp4_r_v_b_08(net1302[0:47]),
     .sp4_v_b_08(sp4_v_b_07_16[47:0]),
     .sp4_v_b_07(sp4_v_b_07_15[47:0]),
     .sp4_v_b_06(sp4_v_b_07_14[47:0]),
     .sp4_v_b_05(sp4_v_b_07_13[47:0]), .pgate(pgate_r[127:0]),
     .reset_b(reset_b_r[127:0]), .wl(wl_r[127:0]),
     .sp12_v_t_08(net1310[0:23]), .tnr_op_08({slf_op_08_17[3],
     slf_op_08_17[2], slf_op_08_17[1], slf_op_08_17[0],
     slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0]}), .top_op_08({slf_op_07_17[3], slf_op_07_17[2],
     slf_op_07_17[1], slf_op_07_17[0], slf_op_07_17[3],
     slf_op_07_17[2], slf_op_07_17[1], slf_op_07_17[0]}),
     .tnl_op_08({tnl_op_07_16[3], tnl_op_07_16[2], tnl_op_07_16[1],
     tnl_op_07_16[0], tnl_op_07_16[3], tnl_op_07_16[2],
     tnl_op_07_16[1], tnl_op_07_16[0]}), .sp4_v_t_08(net1314[0:47]),
     .lc_bot(lc_bot_07_09), .op_vic(net1316),
     .sp12_v_b_01(sp12_v_b_07_09[23:0]), .glb_netwk_t(net1318[0:7]));
pinlatbuf12p I_pinlatbuf12p_r ( .pad_in(padin_r[13]),
     .icegate(hold_r_t), .cbit(cf_r[15]), .cout(net01448),
     .prog(prog));
pinlatbuf12p I_pinlatbuf12p ( .pad_in(padin_t_r[12]),
     .icegate(hold_t_r), .cbit(cf_t[15]), .cout(padinlat_t_r[0]),
     .prog(prog));

endmodule
// Library - ice8chip, Cell - io_col4_lft_ice8p_v2, View - schematic
// LAST TIME SAVED: Jan 12 15:05:42 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_col4_lft_ice8p_v2 ( cbit_colcntl, cf, fabric_out, padeb,
     pado, sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t,
     sp12_h_l, bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold,
     lft_op, mode, padin, pgate, prog, r, reset, sdi, shift, spioeb,
     spiout, tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [7:0]  cbit_colcntl;
output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;
output [23:0]  cf;

inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;

input [7:0]  glb_netwk;
input [1:0]  padin;
input [15:0]  wl;
input [15:0]  reset;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [1:0]  spiout;
input [1:0]  spioeb;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  tnl_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [1:0]  om;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [3:0]  t_mid;



rm7w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
sbox1_colbdlc_v4 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_gmux_x16bare_v4 I_io_gmux_x16bare_v4 (
     .cbit_colcntl(cbit_colcntl[7:0]), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));

endmodule
// Library - ice1chip, Cell - io_lft_top_1x8_ice1f, View - schematic
// LAST TIME SAVED: Apr 11 16:00:35 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_lft_top_1x8_ice1f ( cf_l, fabric_out_09, fo_dlyadj, padeb,
     pado, sdo, slf_op_01, slf_op_02, slf_op_03, slf_op_04, slf_op_05,
     slf_op_06, slf_op_07, slf_op_08, tclk_o, SP4_h_l_01, SP4_h_l_02,
     SP4_h_l_03, SP4_h_l_04, SP4_h_l_05, SP4_h_l_06, SP4_h_l_07,
     SP4_h_l_08, SP12_h_l_01, SP12_h_l_02, SP12_h_l_03, SP12_h_l_04,
     SP12_h_l_05, SP12_h_l_06, SP12_h_l_07, SP12_h_l_08, bl, pgate,
     reset_b, sp4_v_b_00_09, sp4_v_t_08, vdd_cntl, wl, bnr_op_00_09,
     bs_en, ceb, glb_netwk_col, hiz_b, hold, jtag_rowtest_mode_rowu1_b,
     last_rsr, mode, padin, prog, r, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, sdi, shift,
     tclk, tnr_op_08, update );
output  fabric_out_09, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu1_b, mode, prog,
     r, sdi, shift, tclk, update;

output [3:0]  slf_op_03;
output [3:0]  slf_op_01;
output [3:0]  slf_op_02;
output [3:0]  slf_op_06;
output [3:0]  slf_op_07;
output [3:0]  slf_op_08;
output [3:0]  slf_op_05;
output [191:0]  cf_l;
output [3:0]  slf_op_04;
output [7:3]  fo_dlyadj;
output [23:12]  padeb;
output [23:12]  pado;

inout [47:0]  SP4_h_l_02;
inout [47:0]  SP4_h_l_08;
inout [23:0]  SP12_h_l_02;
inout [23:0]  SP12_h_l_08;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_06;
inout [23:0]  SP12_h_l_03;
inout [23:0]  SP12_h_l_07;
inout [47:0]  SP4_h_l_04;
inout [47:0]  SP4_h_l_05;
inout [47:0]  SP4_h_l_03;
inout [23:0]  SP12_h_l_05;
inout [23:0]  SP12_h_l_06;
inout [47:0]  SP4_h_l_01;
inout [47:0]  SP4_h_l_07;
inout [15:0]  sp4_v_t_08;
inout [23:0]  SP12_h_l_01;
inout [15:0]  sp4_v_b_00_09;
inout [127:0]  vdd_cntl;
inout [127:0]  pgate;
inout [127:0]  wl;
inout [127:0]  reset_b;
inout [23:0]  SP12_h_l_04;

input [7:0]  bnr_op_00_09;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_04;
input [1:1]  last_rsr;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_08;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_02;
input [23:12]  padin;
input [7:0]  rgt_op_07;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net1002;

wire  [0:1]  net1014;

wire  [0:1]  net1013;

wire  [7:0]  glb_netwk_b;

wire  [0:7]  net1016;

wire  [0:15]  net865;

wire  [7:0]  glb_netwk_t;

wire  [0:7]  net1017;

wire  [0:7]  net884;

wire  [0:7]  net1008;

wire  [0:1]  net1000;

wire  [7:0]  colbuf_cntl_b;

wire  [0:15]  net793;

wire  [0:1]  net1005;

wire  [0:15]  net757;

wire  [0:15]  net829;

wire  [0:7]  net1007;

wire  [0:1]  net1012;

wire  [0:1]  net719;

wire  [0:15]  net901;

wire  [0:7]  net704;

wire  [0:15]  net973;

wire  [0:1]  net1009;

wire  [0:15]  net937;

wire  [0:1]  net1010;

wire  [0:1]  net755;

wire  [0:1]  net1001;

wire  [0:1]  net1003;

wire  [7:0]  colbuf_cntl_t;



tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
io_col4_lft_ice8p_v2 I_io_00_08 ( .cbit_colcntl(net704[0:7]),
     .ceb(ceb), .sdo(net743), .sdi(sdi), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(net719[0:1]), .pado(net719[0:1]),
     .padeb(net1000[0:1]), .sp4_v_t(sp4_v_t_08[15:0]),
     .sp4_h_l(SP4_h_l_08[47:0]), .sp12_h_l(SP12_h_l_08[23:0]),
     .prog(prog), .spi_ss_in_b(net1012[0:1]), .tnl_op(tnr_op_08[7:0]),
     .lft_op(rgt_op_08[7:0]), .bnl_op(rgt_op_07[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net757[0:15]), .wl(wl[127:112]), .cf(cf_l[191:168]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_08[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net739));
io_col4_lft_ice8p_v2 I_io_00_07 ( .cbit_colcntl(net1016[0:7]),
     .ceb(ceb), .sdo(net815), .sdi(net743), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(net755[0:1]), .pado(net755[0:1]),
     .padeb(net1001[0:1]), .sp4_v_t(net757[0:15]),
     .sp4_h_l(SP4_h_l_07[47:0]), .sp12_h_l(SP12_h_l_07[23:0]),
     .prog(prog), .spi_ss_in_b(net1013[0:1]), .tnl_op(rgt_op_08[7:0]),
     .lft_op(rgt_op_07[7:0]), .bnl_op(rgt_op_06[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net829[0:15]), .wl(wl[111:96]), .cf(cf_l[167:144]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_07[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net775));
io_col4_lft_ice8p_v2 I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net959), .sdi(net779), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[21:20]), .pado(pado[21:20]),
     .padeb(padeb[21:20]), .sp4_v_t(net793[0:15]),
     .sp4_h_l(SP4_h_l_05[47:0]), .sp12_h_l(SP12_h_l_05[23:0]),
     .prog(prog), .spi_ss_in_b(net1003[0:1]), .tnl_op(rgt_op_06[7:0]),
     .lft_op(rgt_op_05[7:0]), .bnl_op(rgt_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net973[0:15]), .wl(wl[79:64]), .cf(cf_l[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[6]));
io_col4_lft_ice8p_v2 I_io_00_06 ( .cbit_colcntl(net1017[0:7]),
     .ceb(ceb), .sdo(net779), .sdi(net815), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[23:22]), .pado(pado[23:22]),
     .padeb(padeb[23:22]), .sp4_v_t(net829[0:15]),
     .sp4_h_l(SP4_h_l_06[47:0]), .sp12_h_l(SP12_h_l_06[23:0]),
     .prog(prog), .spi_ss_in_b(net1010[0:1]), .tnl_op(rgt_op_07[7:0]),
     .lft_op(rgt_op_06[7:0]), .bnl_op(rgt_op_05[7:0]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net793[0:15]), .wl(wl[95:80]), .cf(cf_l[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[7]));
io_col4_lft_ice8p_v2 I_io_00_02 ( .cbit_colcntl(net1007[0:7]),
     .ceb(ceb), .sdo(net887), .sdi(net851), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[15:14]), .pado(pado[15:14]),
     .padeb(padeb[15:14]), .sp4_v_t(net865[0:15]),
     .sp4_h_l(SP4_h_l_02[47:0]), .sp12_h_l(SP12_h_l_02[23:0]),
     .prog(prog), .spi_ss_in_b(net1014[0:1]), .tnl_op(rgt_op_03[7:0]),
     .lft_op(rgt_op_02[7:0]), .bnl_op(rgt_op_01[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(net901[0:15]), .wl(wl[31:16]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[3]));
io_col4_lft_ice8p_v2 I_io_00_01 ( .cbit_colcntl(net884[0:7]),
     .ceb(ceb), .sdo(sdo), .sdi(net887), .spiout({tiegnd,
     last_rsr[1]}), .cdone_in(jtag_rowtest_mode_rowu1_b),
     .spioeb({tievdd, tiegnd}), .mode(mode), .shift(shift),
     .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[13:12]), .pado(pado[13:12]),
     .padeb(padeb[13:12]), .sp4_v_t(net901[0:15]),
     .sp4_h_l(SP4_h_l_01[47:0]), .sp12_h_l(SP12_h_l_01[23:0]),
     .prog(prog), .spi_ss_in_b(net1005[0:1]), .tnl_op(rgt_op_02[7:0]),
     .lft_op(rgt_op_01[7:0]), .bnl_op(bnr_op_00_09[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_v_b_00_09[15:0]), .wl(wl[15:0]), .cf(cf_l[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_09));
io_col4_lft_ice8p_v2 I_io_00_03 ( .cbit_colcntl(net1008[0:7]),
     .ceb(ceb), .sdo(net851), .sdi(net923), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[17:16]), .pado(pado[17:16]),
     .padeb(padeb[17:16]), .sp4_v_t(net937[0:15]),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b(net1009[0:1]), .tnl_op(rgt_op_04[7:0]),
     .lft_op(rgt_op_03[7:0]), .bnl_op(rgt_op_02[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net865[0:15]), .wl(wl[47:32]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[4]));
io_col4_lft_ice8p_v2 I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net923), .sdi(net959), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[19:18]), .pado(pado[19:18]),
     .padeb(padeb[19:18]), .sp4_v_t(net973[0:15]),
     .sp4_h_l(SP4_h_l_04[47:0]), .sp12_h_l(SP12_h_l_04[23:0]),
     .prog(prog), .spi_ss_in_b(net1002[0:1]), .tnl_op(rgt_op_05[7:0]),
     .lft_op(rgt_op_04[7:0]), .bnl_op(rgt_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net937[0:15]), .wl(wl[63:48]), .cf(cf_l[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[5]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - ice1chip, Cell - io_top_lft_1x6_ice1f, View - schematic
// LAST TIME SAVED: Mar  5 17:03:41 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_top_lft_1x6_ice1f ( bs_en_o, ceb_o, cf_top_l,
     fabric_out_06_17, hiz_b_o, mode_o, padeb_t_l, pado_t_l, r_o, sdo,
     shift_o, slf_op_01_17, slf_op_02_17, slf_op_03_17, slf_op_04_17,
     slf_op_05_17, slf_op_06_17, tclk_o, update_o, bl_01, bl_02, bl_03,
     bl_04, bl_05, bl_06, sp4_h_l_01_17, sp4_h_r_06_17, sp4_v_b_01_17,
     sp4_v_b_02_17, sp4_v_b_03_17, sp4_v_b_04_17, sp4_v_b_05_17,
     sp4_v_b_06_17, sp12_v_b_01_17, sp12_v_b_02_17, sp12_v_b_03_17,
     sp12_v_b_04_17, sp12_v_b_05_17, sp12_v_b_06_17, bnl_op_01_17,
     bnr_op_06_17, bs_en_i, ceb_i, glb_net_01, glb_net_02, glb_net_03,
     glb_net_04, glb_net_05, glb_net_06, hiz_b_i, hold_t_l,
     lft_op_01_17, lft_op_02_17, lft_op_03_17, lft_op_04_17,
     lft_op_05_17, lft_op_06_17, mode_i, padin_t_l, pgate_l, prog, r_i,
     reset_l, sdi, shift_i, tclk_i, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_06_17, hiz_b_o, mode_o, r_o, sdo,
     shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_01_17;
output [3:0]  slf_op_03_17;
output [3:0]  slf_op_04_17;
output [3:0]  slf_op_05_17;
output [11:0]  pado_t_l;
output [11:0]  padeb_t_l;
output [3:0]  slf_op_06_17;
output [3:0]  slf_op_02_17;
output [143:0]  cf_top_l;

inout [23:0]  sp12_v_b_04_17;
inout [23:0]  sp12_v_b_03_17;
inout [47:0]  sp4_v_b_01_17;
inout [23:0]  sp12_v_b_01_17;
inout [23:0]  sp12_v_b_05_17;
inout [15:0]  sp4_h_r_06_17;
inout [53:0]  bl_01;
inout [53:0]  bl_04;
inout [41:0]  bl_03;
inout [15:0]  sp4_h_l_01_17;
inout [53:0]  bl_05;
inout [53:0]  bl_06;
inout [23:0]  sp12_v_b_06_17;
inout [23:0]  sp12_v_b_02_17;
inout [47:0]  sp4_v_b_03_17;
inout [47:0]  sp4_v_b_06_17;
inout [47:0]  sp4_v_b_04_17;
inout [47:0]  sp4_v_b_02_17;
inout [47:0]  sp4_v_b_05_17;
inout [53:0]  bl_02;

input [7:0]  lft_op_03_17;
input [7:0]  glb_net_01;
input [7:0]  glb_net_03;
input [7:0]  bnl_op_01_17;
input [15:0]  wl_l;
input [7:0]  lft_op_01_17;
input [7:0]  glb_net_06;
input [7:0]  lft_op_05_17;
input [7:0]  lft_op_02_17;
input [11:0]  padin_t_l;
input [7:0]  glb_net_02;
input [15:0]  pgate_l;
input [7:0]  bnr_op_06_17;
input [7:0]  lft_op_04_17;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_04;
input [7:0]  lft_op_06_17;
input [7:0]  glb_net_05;
input [15:0]  reset_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net1532;

wire  [0:1]  net1319;

wire  [0:15]  net1427;

wire  [0:1]  net1312;

wire  [0:1]  net1318;

wire  [0:1]  net1361;

wire  [0:15]  net1392;

wire  [0:15]  net1357;

wire  [0:1]  net1501;

wire  [0:1]  net1431;

wire  [0:15]  net1462;



tckbufx32_ice8p I_tck_halfbankcenter ( .in(net0262), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));
scan_buf_ice8p I345 ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net0262), .shift_o(shift_o),
     .sdo(net1482), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_top_ice8p I_IO_02_17 ( .sdo(net1412), .sdi(net1342),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net1427[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_l[3:2]), .pado(pado_t_l[3:2]),
     .padeb(padeb_t_l[3:2]), .sp4_v_b(net1357[0:15]),
     .sp4_h_l(sp4_v_b_02_17[47:0]), .sp12_h_l(sp12_v_b_02_17[23:0]),
     .prog(prog), .spi_ss_in_b(net1361[0:1]),
     .tnl_op(lft_op_01_17[7:0]), .lft_op(lft_op_02_17[7:0]),
     .bnl_op(lft_op_03_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[47:24]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_17[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_t_l), .fabric_out(net1320));
io_col4_top_ice8p I_IO_03_17_bram ( .sdo(net1342), .sdi(net1377),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net1357[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_l[5:4]), .pado(pado_t_l[5:4]),
     .padeb(padeb_t_l[5:4]), .sp4_v_b(net1392[0:15]),
     .sp4_h_l(sp4_v_b_03_17[47:0]), .sp12_h_l(sp12_v_b_03_17[23:0]),
     .prog(prog), .spi_ss_in_b(net1318[0:1]),
     .tnl_op(lft_op_02_17[7:0]), .lft_op(lft_op_03_17[7:0]),
     .bnl_op(lft_op_04_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[71:48]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_17[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_t_l), .fabric_out(net1410));
io_col4_top_ice8p I_IO_01_17 ( .sdo(sdo), .sdi(net1412),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_01_17[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[1:0]),
     .pado(pado_t_l[1:0]), .padeb(padeb_t_l[1:0]),
     .sp4_v_b(net1427[0:15]), .sp4_h_l(sp4_v_b_01_17[47:0]),
     .sp12_h_l(sp12_v_b_01_17[23:0]), .prog(prog),
     .spi_ss_in_b(net1431[0:1]), .tnl_op(bnl_op_01_17[7:0]),
     .lft_op(lft_op_01_17[7:0]), .bnl_op(lft_op_02_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_01[5],
     bl_01[4], bl_01[37], bl_01[36], bl_01[35], bl_01[34], bl_01[33],
     bl_01[32], bl_01[14], bl_01[20], bl_01[19], bl_01[18], bl_01[17],
     bl_01[16], bl_01[27], bl_01[26], bl_01[25], bl_01[23]}),
     .wl(wl_l[15:0]), .cf(cf_top_l[23:0]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_01_17[3:0]),
     .glb_netwk(glb_net_01[7:0]), .hold(hold_t_l),
     .fabric_out(net1445));
io_col4_top_ice8p I_IO_05_17 ( .sdo(net1517), .sdi(net1447),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net1532[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_l[9:8]), .pado(pado_t_l[9:8]),
     .padeb(padeb_t_l[9:8]), .sp4_v_b(net1462[0:15]),
     .sp4_h_l(sp4_v_b_05_17[47:0]), .sp12_h_l(sp12_v_b_05_17[23:0]),
     .prog(prog), .spi_ss_in_b(net1319[0:1]),
     .tnl_op(lft_op_04_17[7:0]), .lft_op(lft_op_05_17[7:0]),
     .bnl_op(lft_op_06_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[119:96]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_17[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_t_l), .fabric_out(net1480));
io_col4_top_ice8p I_IO_06_17 ( .sdo(net1447), .sdi(net1482),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net1462[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_l[11:10]),
     .pado(pado_t_l[11:10]), .padeb(padeb_t_l[11:10]),
     .sp4_v_b(sp4_h_r_06_17[15:0]), .sp4_h_l(sp4_v_b_06_17[47:0]),
     .sp12_h_l(sp12_v_b_06_17[23:0]), .prog(prog),
     .spi_ss_in_b(net1501[0:1]), .tnl_op(lft_op_05_17[7:0]),
     .lft_op(lft_op_06_17[7:0]), .bnl_op(bnr_op_06_17[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_l[15:0]), .cf(cf_top_l[143:120]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_06_17[3:0]),
     .glb_netwk(glb_net_06[7:0]), .hold(hold_t_l),
     .fabric_out(fabric_out_06_17));
io_col4_top_ice8p I_IO_04_17 ( .sdo(net1377), .sdi(net1517),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net1392[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t_l[7:6]), .pado(pado_t_l[7:6]),
     .padeb(padeb_t_l[7:6]), .sp4_v_b(net1532[0:15]),
     .sp4_h_l(sp4_v_b_04_17[47:0]), .sp12_h_l(sp12_v_b_04_17[23:0]),
     .prog(prog), .spi_ss_in_b(net1312[0:1]),
     .tnl_op(lft_op_03_17[7:0]), .lft_op(lft_op_04_17[7:0]),
     .bnl_op(lft_op_05_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[95:72]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_17[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_t_l), .fabric_out(net1313));

endmodule
// Library - ice1chip, Cell - quad_tl_ice1, View - schematic
// LAST TIME SAVED: May 18 11:43:55 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module quad_tl_ice1 ( bm_aa_2bot, bm_ab_2bot, bm_sdo_o, bs_en_o, ceb_o,
     cf_l, cf_t, fabric_out_00_09, fabric_out_06_17, fo_dlyadj,
     hiz_b_o, mode_o, padeb_l_t, padeb_t_l, padin_00_09a, padin_06_17b,
     pado_l_t, pado_t_l, r_o, sdo, shift_o, slf_op_00_09, slf_op_01_09,
     slf_op_02_09, slf_op_03_09, slf_op_04_09, slf_op_05_09,
     slf_op_06_09, slf_op_06_10, slf_op_06_11, slf_op_06_12,
     slf_op_06_13, slf_op_06_14, slf_op_06_15, slf_op_06_16,
     slf_op_06_17, tclk_o, update_o, bl, pgate_l, reset_b_l,
     sp4_h_r_06_09, sp4_h_r_06_10, sp4_h_r_06_11, sp4_h_r_06_12,
     sp4_h_r_06_13, sp4_h_r_06_14, sp4_h_r_06_15, sp4_h_r_06_16,
     sp4_h_r_06_17, sp4_r_v_b_06_09, sp4_r_v_b_06_10, sp4_r_v_b_06_11,
     sp4_r_v_b_06_12, sp4_r_v_b_06_13, sp4_r_v_b_06_14,
     sp4_r_v_b_06_15, sp4_r_v_b_06_16, sp4_v_b_00_09, sp4_v_b_01_09,
     sp4_v_b_02_09, sp4_v_b_03_09, sp4_v_b_04_09, sp4_v_b_05_09,
     sp4_v_b_06_09, sp12_h_r_06_09, sp12_h_r_06_10, sp12_h_r_06_11,
     sp12_h_r_06_12, sp12_h_r_06_13, sp12_h_r_06_14, sp12_h_r_06_15,
     sp12_h_r_06_16, sp12_v_b_01_09, sp12_v_b_02_09, sp12_v_b_03_09,
     sp12_v_b_04_09, sp12_v_b_05_09, sp12_v_b_06_09, vdd_cntl_l, wl_l,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_01_09,
     bnl_op_02_09, bnl_op_03_09, bnl_op_04_09, bnl_op_05_09,
     bnl_op_06_09, bnr_op_00_09, bnr_op_01_09, bnr_op_02_09,
     bnr_op_03_09, bnr_op_04_09, bnr_op_05_09, bnr_op_06_09,
     bot_op_01_09, bot_op_02_09, bot_op_03_09, bot_op_04_09,
     bot_op_05_09, bot_op_06_09, bs_en_i, carry_in_01_09,
     carry_in_02_09, carry_in_04_09, carry_in_05_09, carry_in_06_09,
     ceb_i, glb_in, hiz_b_i, hold_l_t, hold_t_l,
     jtag_rowtest_mode_rowu1_b, last_rsr, lc_bot_01_09, lc_bot_02_09,
     lc_bot_04_09, lc_bot_05_09, lc_bot_06_09, mode_i, padin_l_t,
     padin_t_l, prog, purst, r_i, rgt_op_06_09, rgt_op_06_10,
     rgt_op_06_11, rgt_op_06_12, rgt_op_06_13, rgt_op_06_14,
     rgt_op_06_15, rgt_op_06_16, sdi, shift_i, tclk_i, tnr_op_06_16,
     update_i );
output  bs_en_o, ceb_o, fabric_out_00_09, fabric_out_06_17, hiz_b_o,
     mode_o, padin_00_09a, padin_06_17b, r_o, sdo, shift_o, tclk_o,
     update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, carry_in_01_09, carry_in_02_09,
     carry_in_04_09, carry_in_05_09, carry_in_06_09, ceb_i, hiz_b_i,
     hold_l_t, hold_t_l, jtag_rowtest_mode_rowu1_b, lc_bot_01_09,
     lc_bot_02_09, lc_bot_04_09, lc_bot_05_09, lc_bot_06_09, mode_i,
     prog, purst, r_i, sdi, shift_i, tclk_i, update_i;

output [7:0]  slf_op_04_09;
output [23:12]  pado_l_t;
output [11:0]  padeb_t_l;
output [10:0]  bm_ab_2bot;
output [7:0]  slf_op_06_12;
output [7:0]  slf_op_01_09;
output [3:0]  slf_op_06_17;
output [191:0]  cf_l;
output [7:0]  slf_op_06_13;
output [7:0]  slf_op_06_09;
output [7:0]  slf_op_06_14;
output [23:12]  padeb_l_t;
output [10:0]  bm_aa_2bot;
output [3:0]  slf_op_00_09;
output [143:0]  cf_t;
output [7:0]  slf_op_06_10;
output [11:0]  pado_t_l;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_06_11;
output [7:3]  fo_dlyadj;
output [7:0]  slf_op_06_16;
output [7:0]  slf_op_05_09;
output [7:0]  slf_op_06_15;
output [7:0]  slf_op_02_09;
output [7:0]  slf_op_03_09;

inout [23:0]  sp12_v_b_03_09;
inout [47:0]  sp4_v_b_01_09;
inout [47:0]  sp4_h_r_06_15;
inout [47:0]  sp4_v_b_06_09;
inout [23:0]  sp12_h_r_06_14;
inout [47:0]  sp4_h_r_06_14;
inout [47:0]  sp4_v_b_04_09;
inout [47:0]  sp4_r_v_b_06_11;
inout [47:0]  sp4_r_v_b_06_10;
inout [23:0]  sp12_v_b_04_09;
inout [23:0]  sp12_h_r_06_09;
inout [47:0]  sp4_h_r_06_10;
inout [23:0]  sp12_h_r_06_13;
inout [23:0]  sp12_h_r_06_16;
inout [23:0]  sp12_v_b_06_09;
inout [47:0]  sp4_h_r_06_16;
inout [23:0]  sp12_h_r_06_11;
inout [143:0]  wl_l;
inout [143:0]  reset_b_l;
inout [143:0]  vdd_cntl_l;
inout [23:0]  sp12_v_b_01_09;
inout [23:0]  sp12_h_r_06_12;
inout [47:0]  sp4_h_r_06_11;
inout [47:0]  sp4_r_v_b_06_14;
inout [329:0]  bl;
inout [47:0]  sp4_r_v_b_06_09;
inout [47:0]  sp4_v_b_02_09;
inout [47:0]  sp4_h_r_06_12;
inout [47:0]  sp4_h_r_06_09;
inout [15:0]  sp4_h_r_06_17;
inout [23:0]  sp12_h_r_06_15;
inout [23:0]  sp12_h_r_06_10;
inout [143:0]  pgate_l;
inout [47:0]  sp4_r_v_b_06_15;
inout [23:0]  sp12_v_b_02_09;
inout [15:0]  sp4_v_b_00_09;
inout [47:0]  sp4_v_b_03_09;
inout [47:0]  sp4_r_v_b_06_16;
inout [47:0]  sp4_r_v_b_06_13;
inout [23:0]  sp12_v_b_05_09;
inout [47:0]  sp4_h_r_06_13;
inout [47:0]  sp4_v_b_05_09;
inout [47:0]  sp4_r_v_b_06_12;

input [7:0]  bot_op_06_09;
input [7:0]  rgt_op_06_14;
input [7:0]  rgt_op_06_16;
input [7:0]  bnl_op_02_09;
input [7:0]  bnr_op_06_09;
input [1:0]  bm_sdi_i;
input [7:0]  rgt_op_06_13;
input [7:0]  rgt_op_06_12;
input [7:0]  rgt_op_06_09;
input [1:0]  bm_sweb_i;
input [7:0]  bot_op_01_09;
input [23:12]  padin_l_t;
input [7:0]  bnr_op_00_09;
input [7:0]  bnr_op_03_09;
input [1:0]  bm_sclkrw_i;
input [7:0]  bnl_op_04_09;
input [7:0]  bot_op_04_09;
input [7:0]  bnr_op_02_09;
input [7:0]  bnl_op_01_09;
input [7:0]  glb_in;
input [11:0]  padin_t_l;
input [7:0]  bnr_op_05_09;
input [7:0]  bnr_op_01_09;
input [7:0]  rgt_op_06_11;
input [7:0]  rgt_op_06_10;
input [7:0]  bot_op_05_09;
input [1:1]  last_rsr;
input [7:0]  bnl_op_03_09;
input [7:0]  bot_op_02_09;
input [7:0]  bm_sa_i;
input [7:0]  bnl_op_06_09;
input [7:0]  bnr_op_04_09;
input [7:0]  bot_op_03_09;
input [7:0]  rgt_op_06_15;
input [3:0]  tnr_op_06_16;
input [7:0]  bnl_op_05_09;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  clk_tree_drv_tl;

wire  [3:0]  slf_op_02_17;

wire  [3:0]  slf_op_01_17;

wire  [3:0]  slf_op_05_17;

wire  [3:0]  slf_op_04_17;

wire  [7:0]  clk_center;

wire  [3:0]  slf_op_08_17;

wire  [3:0]  slf_op_00_15;

wire  [0:47]  net795;

wire  [0:23]  net1235;

wire  [0:1]  net1439;

wire  [0:23]  net1141;

wire  [0:47]  net1446;

wire  [0:7]  net1273;

wire  [0:7]  net833;

wire  [0:23]  net950;

wire  [0:47]  net1450;

wire  [0:47]  net1151;

wire  [3:0]  slf_op_00_11;

wire  [1:0]  bm_sdi_b1_o;

wire  [3:0]  slf_op_00_10;

wire  [3:0]  slf_op_00_12;

wire  [0:47]  net1169;

wire  [3:0]  slf_op_00_13;

wire  [3:0]  slf_op_00_14;

wire  [3:0]  slf_op_00_16;

wire  [0:47]  net1291;

wire  [0:47]  net746;

wire  [0:47]  net1445;

wire  [0:47]  net826;

wire  [0:7]  net773;

wire  [0:23]  net951;

wire  [0:23]  net1140;

wire  [0:7]  net939;

wire  [0:47]  net959;

wire  [0:47]  net819;

wire  [0:47]  net765;

wire  [0:47]  net1239;

wire  [0:7]  net929;

wire  [0:7]  net1022;

wire  [0:47]  net732;

wire  [0:47]  net960;

wire  [0:7]  net836;

wire  [0:47]  net1196;

wire  [0:47]  net1003;

wire  [0:47]  net1049;

wire  [0:23]  net1191;

wire  [0:7]  net1214;

wire  [0:23]  net1190;

wire  [0:23]  net998;

wire  [0:7]  net832;

wire  [0:7]  net770;

wire  [0:23]  net749;

wire  [0:23]  net856;

wire  [0:23]  net1284;

wire  [0:7]  net834;

wire  [0:47]  net1018;

wire  [0:47]  net1303;

wire  [0:23]  net1093;

wire  [0:47]  net1050;

wire  [0:7]  net931;

wire  [0:7]  net1026;

wire  [0:47]  net728;

wire  [0:47]  net1055;

wire  [0:47]  net1144;

wire  [0:23]  net716;

wire  [0:47]  net956;

wire  [0:23]  net948;

wire  [0:7]  net769;

wire  [0:23]  net720;

wire  [0:47]  net1267;

wire  [0:23]  net1043;

wire  [0:23]  net1394;

wire  [0:23]  net1096;

wire  [0:23]  net1234;

wire  [0:23]  net851;

wire  [0:7]  net1402;

wire  [0:23]  net721;

wire  [0:47]  net979;

wire  [0:47]  net954;

wire  [0:23]  net1001;

wire  [0:47]  net1288;

wire  [0:7]  net1024;

wire  [0:47]  net1113;

wire  [0:7]  net1460;

wire  [0:23]  net1046;

wire  [0:47]  net1289;

wire  [0:47]  net1290;

wire  [0:47]  net790;

wire  [0:23]  net1094;

wire  [0:47]  net980;

wire  [0:7]  net1452;

wire  [0:23]  net1236;

wire  [0:47]  net794;

wire  [0:23]  net748;

wire  [0:47]  net1243;

wire  [0:47]  net1099;

wire  [0:23]  net949;

wire  [0:47]  net1266;

wire  [0:47]  net982;

wire  [0:47]  net1170;

wire  [0:23]  net850;

wire  [0:7]  net695;

wire  [0:7]  net786;

wire  [0:7]  net987;

wire  [0:47]  net735;

wire  [0:47]  net1193;

wire  [0:7]  net988;

wire  [0:47]  net763;

wire  [0:23]  net1285;

wire  [0:23]  net740;

wire  [0:7]  net1082;

wire  [0:47]  net1100;

wire  [0:47]  net1208;

wire  [0:7]  net1451;

wire  [0:7]  net989;

wire  [0:7]  net1117;

wire  [0:47]  net829;

wire  [0:47]  net1076;

wire  [0:47]  net827;

wire  [0:7]  net1275;

wire  [0:23]  net1299;

wire  [0:7]  net772;

wire  [0:47]  net830;

wire  [0:47]  net1195;

wire  [0:23]  net855;

wire  [0:47]  net825;

wire  [0:47]  net1051;

wire  [0:7]  net1212;

wire  [0:47]  net1146;

wire  [0:47]  net791;

wire  [0:47]  net1240;

wire  [0:47]  net1101;

wire  [0:47]  net793;

wire  [0:7]  net1307;

wire  [0:23]  net756;

wire  [0:47]  net1150;

wire  [0:23]  net718;

wire  [0:47]  net1005;

wire  [0:47]  net1194;

wire  [0:47]  net1172;

wire  [0:23]  net852;

wire  [0:23]  net999;

wire  [0:47]  net764;

wire  [0:1]  net1441;

wire  [0:23]  net1189;

wire  [0:47]  net1074;

wire  [0:47]  net1264;

wire  [0:47]  net1056;

wire  [0:47]  net731;

wire  [0:7]  net1274;

wire  [0:7]  net990;

wire  [0:47]  net961;

wire  [0:23]  net857;

wire  [0:7]  net818;

wire  [0:23]  net1044;

wire  [0:47]  net828;

wire  [0:7]  net768;

wire  [0:23]  net1138;

wire  [0:47]  net1075;

wire  [0:23]  net1204;

wire  [0:47]  net724;

wire  [0:7]  net1453;

wire  [0:23]  net1233;

wire  [0:23]  net1139;

wire  [0:47]  net1245;

wire  [0:47]  net958;

wire  [0:47]  net1145;

wire  [0:7]  net858;

wire  [0:47]  net734;

wire  [0:7]  net1085;

wire  [0:15]  net820;

wire  [0:47]  net955;

wire  [0:23]  net1188;

wire  [0:23]  net1000;

wire  [0:7]  net1083;

wire  [0:47]  net1244;

wire  [0:47]  net1077;

wire  [0:47]  net1098;

wire  [0:23]  net1283;

wire  [0:47]  net1148;

wire  [0:23]  net1109;

wire  [0:23]  net1286;

wire  [0:47]  net1004;

wire  [0:7]  net1084;

wire  [0:47]  net1398;

wire  [0:47]  net1006;

wire  [0:47]  net809;

wire  [0:47]  net1241;

wire  [0:23]  net1014;

wire  [0:7]  net767;

wire  [0:7]  net771;

wire  [0:47]  net981;

wire  [0:23]  net854;

wire  [0:47]  net1053;

wire  [0:7]  net1272;

wire  [0:47]  net1265;

wire  [0:47]  net1449;

wire  [0:47]  net1171;

wire  [0:47]  net1149;

wire  [0:7]  net1118;

wire  [0:7]  net1224;

wire  [0:47]  net792;

wire  [0:23]  net1045;

wire  [0:47]  net1443;

wire  [0:23]  net1095;

wire  [0:23]  net849;

wire  [0:47]  net1448;

wire  [0:47]  net1054;

wire  [0:23]  net704;

wire  [0:47]  net1246;

wire  [0:7]  net831;

wire  [0:7]  net1216;

wire  [0:7]  net1213;

wire  [0:47]  net1444;

wire  [0:7]  net1034;



bram1x4_ice1f I_bram_col_t03 ( .prog(prog),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .reset_b(reset_b_l[127:0]), .bm_wdummymux_en_o(net1440),
     .bm_sreb_o(net1436), .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(net694),
     .bm_sa_o(net695[0:7]), .bm_rcapmux_en_o(net1435),
     .bm_init_o(net697), .lft_op_05(net990[0:7]), .bl(bl[167:126]),
     .sp4_h_l_06(net1076[0:47]), .sp12_h_l_02(net1045[0:23]),
     .lft_op_06(net989[0:7]), .sp12_h_l_03(net1044[0:23]),
     .sp12_h_r_03(net704[0:23]), .sp12_h_l_01(net1046[0:23]),
     .sp4_v_b_04(net1049[0:47]), .sp4_v_b_05(net1098[0:47]),
     .lft_op_07(net988[0:7]), .sp4_v_b_06(net1099[0:47]),
     .sp4_v_b_08(net1101[0:47]), .sp4_v_b_07(net1100[0:47]),
     .lft_op_03(net929[0:7]), .lft_op_01(slf_op_02_09[7:0]),
     .sp4_h_l_02(net1055[0:47]), .sp12_h_l_06(net1094[0:23]),
     .sp12_h_r_07(net716[0:23]), .sp12_h_l_05(net1093[0:23]),
     .sp12_h_r_06(net718[0:23]), .sp12_h_l_04(net1043[0:23]),
     .sp12_h_r_05(net720[0:23]), .sp12_h_r_08(net721[0:23]),
     .sp12_h_l_07(net1095[0:23]), .sp12_h_l_08(net1096[0:23]),
     .sp4_r_v_b_03(net724[0:47]), .vdd_cntl(vdd_cntl_l[127:0]),
     .pgate(pgate_l[127:0]), .bot_op_01(bot_op_03_09[7:0]),
     .sp4_r_v_b_04(net728[0:47]), .sp4_v_b_01(sp4_v_b_03_09[47:0]),
     .sp4_v_b_03(net1050[0:47]), .sp4_h_r_08(net731[0:47]),
     .sp4_r_v_b_05(net732[0:47]), .sp4_v_b_02(net1051[0:47]),
     .sp4_v_t_08(net734[0:47]), .sp4_r_v_b_02(net735[0:47]),
     .bnr_op_01(bnr_op_03_09[7:0]), .bm_sdi_o(bm_sdi_b1_o[1:0]),
     .sp4_h_l_04(net1053[0:47]), .lft_op_08(net987[0:7]),
     .sp12_h_r_01(net740[0:23]), .bm_sdo_i({tiegnd_bram_t,
     bm_sdi_b1_o[0]}), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sweb_o(net1441[0:1]), .sp4_h_l_03(net1054[0:47]),
     .sp4_h_l_01(net1056[0:47]), .sp4_h_r_01(net746[0:47]),
     .tnr_op_08({slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0], slf_op_04_17[3], slf_op_04_17[2],
     slf_op_04_17[1], slf_op_04_17[0]}), .sp12_h_r_02(net748[0:23]),
     .sp12_h_r_04(net749[0:23]), .bm_sclkrw_o(net1439[0:1]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .lft_op_02(net931[0:7]),
     .lft_op_04(net939[0:7]), .bm_sweb_i(bm_sweb_i[1:0]),
     .bnl_op_01(bnl_op_03_09[7:0]), .sp12_v_t_08(net756[0:23]),
     .wl(wl_l[127:0]), .tnl_op_08({slf_op_02_17[3], slf_op_02_17[2],
     slf_op_02_17[1], slf_op_02_17[0], slf_op_02_17[3],
     slf_op_02_17[2], slf_op_02_17[1], slf_op_02_17[0]}),
     .top_op_08({slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0], slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0]}), .bm_ab_2bot(bm_ab_2bot[10:0]),
     .bm_aa_2bot(bm_aa_2bot[10:0]), .sp12_v_b_01(sp12_v_b_03_09[23:0]),
     .sp4_r_v_b_08(net763[0:47]), .sp4_r_v_b_07(net764[0:47]),
     .sp4_r_v_b_06(net765[0:47]), .sp4_r_v_b_01(sp4_v_b_04_09[47:0]),
     .rgt_op_08(net767[0:7]), .rgt_op_07(net768[0:7]),
     .rgt_op_06(net769[0:7]), .rgt_op_05(net770[0:7]),
     .rgt_op_04(net771[0:7]), .rgt_op_03(net772[0:7]),
     .rgt_op_02(net773[0:7]), .rgt_op_01(slf_op_04_09[7:0]),
     .slf_op_02(net1026[0:7]), .slf_op_01(slf_op_03_09[7:0]),
     .slf_op_03(net1024[0:7]), .slf_op_04(net1034[0:7]),
     .slf_op_05(net1085[0:7]), .slf_op_06(net1084[0:7]),
     .slf_op_07(net1083[0:7]), .slf_op_08(net1082[0:7]),
     .bm_ab_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .bm_aa_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .glb_netwk_bot(net1453[0:7]), .glb_netwk_top(net786[0:7]),
     .sp4_h_l_08(net1074[0:47]), .sp4_h_l_07(net1075[0:47]),
     .sp4_h_l_05(net1077[0:47]), .sp4_h_r_02(net790[0:47]),
     .sp4_h_r_03(net791[0:47]), .sp4_h_r_04(net792[0:47]),
     .sp4_h_r_05(net793[0:47]), .sp4_h_r_06(net794[0:47]),
     .sp4_h_r_07(net795[0:47]));
pinlatbuf12p I389 ( .pad_in(padin_t_l[11]), .icegate(hold_t_l),
     .cbit(cf_t[135]), .cout(net675), .prog(prog));
pinlatbuf12p I_pinlatbuf12p_l ( .pad_in(padin_l_t[12]),
     .icegate(hold_l_t), .cbit(cf_l[15]), .cout(net1427), .prog(prog));
io_lft_top_1x8_ice1f I_preio_lt_t00 ( .padin(padin_l_t[23:12]),
     .pado(pado_l_t[23:12]), .padeb(padeb_l_t[23:12]),
     .fo_dlyadj(fo_dlyadj[7:3]), .sp4_v_b_00_09(sp4_v_b_00_09[15:0]),
     .bnr_op_00_09(bnr_op_00_09[7:0]), .tnr_op_08({slf_op_01_17[3],
     slf_op_01_17[2], slf_op_01_17[1], slf_op_01_17[0],
     slf_op_01_17[3], slf_op_01_17[2], slf_op_01_17[1],
     slf_op_01_17[0]}), .shift(shift_o), .bs_en(bs_en_o),
     .mode(mode_o), .sdi(net803), .hiz_b(hiz_b_o), .prog(prog),
     .hold(hold_l_t), .update(update_o), .r(r_o),
     .SP4_h_l_05(net809[0:47]), .slf_op_05(slf_op_00_13[3:0]),
     .slf_op_01(slf_op_00_09[3:0]), .slf_op_06(slf_op_00_14[3:0]),
     .slf_op_02(slf_op_00_10[3:0]), .sdo(sdo), .bl({bl[0], bl[1],
     bl[2], bl[3], bl[4], bl[5], bl[6], bl[7], bl[8], bl[9], bl[10],
     bl[11], bl[12], bl[13], bl[14], bl[15], bl[16], bl[17]}),
     .tclk(net816), .reset_b(reset_b_l[127:0]),
     .rgt_op_02(net818[0:7]), .SP4_h_l_06(net819[0:47]),
     .sp4_v_t_08(net820[0:15]), .slf_op_04(slf_op_00_12[3:0]),
     .slf_op_03(slf_op_00_11[3:0]), .slf_op_07(slf_op_00_15[3:0]),
     .slf_op_08(slf_op_00_16[3:0]), .SP4_h_l_08(net825[0:47]),
     .SP4_h_l_07(net826[0:47]), .SP4_h_l_03(net827[0:47]),
     .SP4_h_l_04(net828[0:47]), .SP4_h_l_02(net829[0:47]),
     .SP4_h_l_01(net830[0:47]), .rgt_op_07(net831[0:7]),
     .rgt_op_06(net832[0:7]), .rgt_op_05(net833[0:7]),
     .rgt_op_03(net834[0:7]), .rgt_op_01(slf_op_01_09[7:0]),
     .rgt_op_08(net836[0:7]), .pgate(pgate_l[127:0]),
     .vdd_cntl(vdd_cntl_l[127:0]), .last_rsr(last_rsr[1]),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .cf_l(cf_l[191:0]), .wl(wl_l[127:0]), .tclk_o(tclk_o),
     .ceb(ceb_o), .fabric_out_09(net1423), .SP12_h_l_02(net849[0:23]),
     .SP12_h_l_04(net850[0:23]), .SP12_h_l_08(net851[0:23]),
     .SP12_h_l_06(net852[0:23]), .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .SP12_h_l_05(net854[0:23]), .SP12_h_l_01(net855[0:23]),
     .SP12_h_l_03(net856[0:23]), .SP12_h_l_07(net857[0:23]),
     .rgt_op_04(net858[0:7]));
io_top_lft_1x6_ice1f I_preio_top_l ( .fabric_out_06_17(net859),
     .cf_top_l(cf_t[143:0]), .wl_l({wl_l[142], wl_l[143], wl_l[141],
     wl_l[140], wl_l[138], wl_l[139], wl_l[137], wl_l[136], wl_l[134],
     wl_l[135], wl_l[133], wl_l[132], wl_l[130], wl_l[131], wl_l[129],
     wl_l[128]}), .lft_op_01_17(net836[0:7]),
     .vdd_cntl_l({vdd_cntl_l[142], vdd_cntl_l[143], vdd_cntl_l[141],
     vdd_cntl_l[140], vdd_cntl_l[138], vdd_cntl_l[139],
     vdd_cntl_l[137], vdd_cntl_l[136], vdd_cntl_l[134],
     vdd_cntl_l[135], vdd_cntl_l[133], vdd_cntl_l[132],
     vdd_cntl_l[130], vdd_cntl_l[131], vdd_cntl_l[129],
     vdd_cntl_l[128]}), .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .reset_l({reset_b_l[142],
     reset_b_l[143], reset_b_l[141], reset_b_l[140], reset_b_l[138],
     reset_b_l[139], reset_b_l[137], reset_b_l[136], reset_b_l[134],
     reset_b_l[135], reset_b_l[133], reset_b_l[132], reset_b_l[130],
     reset_b_l[131], reset_b_l[129], reset_b_l[128]}), .r_i(r_i),
     .prog(prog), .pgate_l({pgate_l[142], pgate_l[143], pgate_l[141],
     pgate_l[140], pgate_l[138], pgate_l[139], pgate_l[137],
     pgate_l[136], pgate_l[134], pgate_l[135], pgate_l[133],
     pgate_l[132], pgate_l[130], pgate_l[131], pgate_l[129],
     pgate_l[128]}), .mode_i(mode_i), .hiz_b_i(hiz_b_i),
     .bs_en_i(bs_en_i), .update_o(net1405), .tclk_o(net1406),
     .shift_o(net1407), .sdo(net1408), .r_o(net1409), .mode_o(net1410),
     .hiz_b_o(net1411), .glb_net_06(net1402[0:7]),
     .glb_net_05(net1212[0:7]), .glb_net_04(net1307[0:7]),
     .glb_net_03(net786[0:7]), .glb_net_02(net1117[0:7]),
     .glb_net_01(net1022[0:7]), .bs_en_o(net1413),
     .sp4_h_r_06_17(sp4_h_r_06_17[15:0]), .bl_06(bl[329:276]),
     .bl_05(bl[275:222]), .bl_04(bl[221:168]), .bl_02(bl[125:72]),
     .bl_01(bl[71:18]), .sp4_h_l_01_17(net820[0:15]),
     .bnl_op_01_17({slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0], slf_op_00_16[3], slf_op_00_16[2],
     slf_op_00_16[1], slf_op_00_16[0]}), .padin_t_l(padin_t_l[11:0]),
     .lft_op_03_17(net1082[0:7]), .sp4_v_b_04_17(net1303[0:47]),
     .lft_op_02_17(net987[0:7]), .lft_op_04_17(net767[0:7]),
     .sp4_v_b_06_17(net1398[0:47]), .sp12_v_b_04_17(net1299[0:23]),
     .sp4_v_b_02_17(net1113[0:47]), .sp12_v_b_05_17(net1204[0:23]),
     .lft_op_06_17(slf_op_06_16[7:0]),
     .slf_op_04_17(slf_op_04_17[3:0]), .sp4_v_b_05_17(net1208[0:47]),
     .sp12_v_b_03_17(net756[0:23]), .slf_op_01_17(slf_op_01_17[3:0]),
     .sp4_v_b_01_17(net1018[0:47]), .sp4_v_b_03_17(net734[0:47]),
     .slf_op_03_17(slf_op_08_17[3:0]), .lft_op_05_17(net1272[0:7]),
     .bnr_op_06_17(rgt_op_06_16[7:0]), .sp12_v_b_01_17(net1014[0:23]),
     .slf_op_06_17(slf_op_06_17[3:0]), .sp12_v_b_06_17(net1394[0:23]),
     .slf_op_02_17(slf_op_02_17[3:0]), .sp12_v_b_02_17(net1109[0:23]),
     .padeb_t_l(padeb_t_l[11:0]), .bl_03(bl[167:126]), .ceb_o(net1412),
     .pado_t_l(pado_t_l[11:0]), .hold_t_l(hold_t_l),
     .slf_op_05_17(slf_op_05_17[3:0]), .ceb_i(ceb_i));
lt_1x8_top_ice1f I_lt_col_t01 ( .glb_netwk_b(net1451[0:7]),
     .rgt_op_03(net929[0:7]), .slf_op_02(net818[0:7]),
     .rgt_op_02(net931[0:7]), .rgt_op_01(slf_op_02_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04({slf_op_00_12[3],
     slf_op_00_12[2], slf_op_00_12[1], slf_op_00_12[0],
     slf_op_00_12[3], slf_op_00_12[2], slf_op_00_12[1],
     slf_op_00_12[0]}), .lft_op_03({slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0], slf_op_00_11[3],
     slf_op_00_11[2], slf_op_00_11[1], slf_op_00_11[0]}),
     .lft_op_02({slf_op_00_10[3], slf_op_00_10[2], slf_op_00_10[1],
     slf_op_00_10[0], slf_op_00_10[3], slf_op_00_10[2],
     slf_op_00_10[1], slf_op_00_10[0]}), .lft_op_01({slf_op_00_09[3],
     slf_op_00_09[2], slf_op_00_09[1], slf_op_00_09[0],
     slf_op_00_09[3], slf_op_00_09[2], slf_op_00_09[1],
     slf_op_00_09[0]}), .rgt_op_04(net939[0:7]),
     .carry_in(carry_in_01_09), .bnl_op_01(bnl_op_01_09[7:0]),
     .slf_op_04(net858[0:7]), .slf_op_03(net834[0:7]),
     .slf_op_01(slf_op_01_09[7:0]), .sp4_h_l_04(net828[0:47]),
     .carry_out(net946), .vdd_cntl(vdd_cntl_l[127:0]),
     .sp12_h_r_04(net948[0:23]), .sp12_h_r_03(net949[0:23]),
     .sp12_h_r_02(net950[0:23]), .sp12_h_r_01(net951[0:23]),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_01_09[47:0]), .sp4_r_v_b_04(net954[0:47]),
     .sp4_r_v_b_03(net955[0:47]), .sp4_r_v_b_02(net956[0:47]),
     .sp4_r_v_b_01(sp4_v_b_02_09[47:0]), .sp4_h_r_04(net958[0:47]),
     .sp4_h_r_03(net959[0:47]), .sp4_h_r_02(net960[0:47]),
     .sp4_h_r_01(net961[0:47]), .sp4_h_l_03(net827[0:47]),
     .sp4_h_l_02(net829[0:47]), .sp4_h_l_01(net830[0:47]),
     .bl(bl[71:18]), .bot_op_01(bot_op_01_09[7:0]),
     .sp12_h_l_01(net855[0:23]), .sp12_h_l_02(net849[0:23]),
     .sp12_h_l_03(net856[0:23]), .sp12_h_l_04(net850[0:23]),
     .sp4_v_b_04(net1449[0:47]), .sp4_v_b_03(net1450[0:47]),
     .sp4_v_b_02(net1448[0:47]), .bnr_op_01(bnr_op_01_09[7:0]),
     .sp4_h_l_05(net809[0:47]), .sp4_h_l_06(net819[0:47]),
     .sp4_h_l_07(net826[0:47]), .sp4_h_l_08(net825[0:47]),
     .sp4_h_r_08(net979[0:47]), .sp4_h_r_07(net980[0:47]),
     .sp4_h_r_06(net981[0:47]), .sp4_h_r_05(net982[0:47]),
     .slf_op_05(net833[0:7]), .slf_op_06(net832[0:7]),
     .slf_op_07(net831[0:7]), .slf_op_08(net836[0:7]),
     .rgt_op_08(net987[0:7]), .rgt_op_07(net988[0:7]),
     .rgt_op_06(net989[0:7]), .rgt_op_05(net990[0:7]),
     .lft_op_08({slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0], slf_op_00_16[3], slf_op_00_16[2],
     slf_op_00_16[1], slf_op_00_16[0]}), .lft_op_07({slf_op_00_15[3],
     slf_op_00_15[2], slf_op_00_15[1], slf_op_00_15[0],
     slf_op_00_15[3], slf_op_00_15[2], slf_op_00_15[1],
     slf_op_00_15[0]}), .lft_op_06({slf_op_00_14[3], slf_op_00_14[2],
     slf_op_00_14[1], slf_op_00_14[0], slf_op_00_14[3],
     slf_op_00_14[2], slf_op_00_14[1], slf_op_00_14[0]}),
     .lft_op_05({slf_op_00_13[3], slf_op_00_13[2], slf_op_00_13[1],
     slf_op_00_13[0], slf_op_00_13[3], slf_op_00_13[2],
     slf_op_00_13[1], slf_op_00_13[0]}), .sp12_h_l_08(net851[0:23]),
     .sp12_h_l_07(net857[0:23]), .sp12_h_l_06(net852[0:23]),
     .sp12_h_r_05(net998[0:23]), .sp12_h_r_06(net999[0:23]),
     .sp12_h_r_07(net1000[0:23]), .sp12_h_r_08(net1001[0:23]),
     .sp12_h_l_05(net854[0:23]), .sp4_r_v_b_05(net1003[0:47]),
     .sp4_r_v_b_06(net1004[0:47]), .sp4_r_v_b_07(net1005[0:47]),
     .sp4_r_v_b_08(net1006[0:47]), .sp4_v_b_08(net1443[0:47]),
     .sp4_v_b_07(net1444[0:47]), .sp4_v_b_06(net1445[0:47]),
     .sp4_v_b_05(net1446[0:47]), .pgate(pgate_l[127:0]),
     .reset_b(reset_b_l[127:0]), .wl(wl_l[127:0]),
     .sp12_v_t_08(net1014[0:23]), .tnr_op_08({slf_op_02_17[3],
     slf_op_02_17[2], slf_op_02_17[1], slf_op_02_17[0],
     slf_op_02_17[3], slf_op_02_17[2], slf_op_02_17[1],
     slf_op_02_17[0]}), .top_op_08({slf_op_01_17[3], slf_op_01_17[2],
     slf_op_01_17[1], slf_op_01_17[0], slf_op_01_17[3],
     slf_op_01_17[2], slf_op_01_17[1], slf_op_01_17[0]}),
     .tnl_op_08({tiegnd_qtl, tiegnd_qtl, tiegnd_qtl, tiegnd_qtl,
     tiegnd_qtl, tiegnd_qtl, tiegnd_qtl, tiegnd_qtl}),
     .sp4_v_t_08(net1018[0:47]), .lc_bot(lc_bot_01_09),
     .op_vic(net1020), .sp12_v_b_01(sp12_v_b_01_09[23:0]),
     .glb_netwk_t(net1022[0:7]));
lt_1x8_top_ice1f I_lt_col_t02 ( .glb_netwk_b(net1452[0:7]),
     .rgt_op_03(net1024[0:7]), .slf_op_02(net931[0:7]),
     .rgt_op_02(net1026[0:7]), .rgt_op_01(slf_op_03_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net858[0:7]),
     .lft_op_03(net834[0:7]), .lft_op_02(net818[0:7]),
     .lft_op_01(slf_op_01_09[7:0]), .rgt_op_04(net1034[0:7]),
     .carry_in(carry_in_02_09), .bnl_op_01(bnl_op_02_09[7:0]),
     .slf_op_04(net939[0:7]), .slf_op_03(net929[0:7]),
     .slf_op_01(slf_op_02_09[7:0]), .sp4_h_l_04(net958[0:47]),
     .carry_out(net1041), .vdd_cntl(vdd_cntl_l[127:0]),
     .sp12_h_r_04(net1043[0:23]), .sp12_h_r_03(net1044[0:23]),
     .sp12_h_r_02(net1045[0:23]), .sp12_h_r_01(net1046[0:23]),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_02_09[47:0]), .sp4_r_v_b_04(net1049[0:47]),
     .sp4_r_v_b_03(net1050[0:47]), .sp4_r_v_b_02(net1051[0:47]),
     .sp4_r_v_b_01(sp4_v_b_03_09[47:0]), .sp4_h_r_04(net1053[0:47]),
     .sp4_h_r_03(net1054[0:47]), .sp4_h_r_02(net1055[0:47]),
     .sp4_h_r_01(net1056[0:47]), .sp4_h_l_03(net959[0:47]),
     .sp4_h_l_02(net960[0:47]), .sp4_h_l_01(net961[0:47]),
     .bl(bl[125:72]), .bot_op_01(bot_op_02_09[7:0]),
     .sp12_h_l_01(net951[0:23]), .sp12_h_l_02(net950[0:23]),
     .sp12_h_l_03(net949[0:23]), .sp12_h_l_04(net948[0:23]),
     .sp4_v_b_04(net954[0:47]), .sp4_v_b_03(net955[0:47]),
     .sp4_v_b_02(net956[0:47]), .bnr_op_01(bnr_op_02_09[7:0]),
     .sp4_h_l_05(net982[0:47]), .sp4_h_l_06(net981[0:47]),
     .sp4_h_l_07(net980[0:47]), .sp4_h_l_08(net979[0:47]),
     .sp4_h_r_08(net1074[0:47]), .sp4_h_r_07(net1075[0:47]),
     .sp4_h_r_06(net1076[0:47]), .sp4_h_r_05(net1077[0:47]),
     .slf_op_05(net990[0:7]), .slf_op_06(net989[0:7]),
     .slf_op_07(net988[0:7]), .slf_op_08(net987[0:7]),
     .rgt_op_08(net1082[0:7]), .rgt_op_07(net1083[0:7]),
     .rgt_op_06(net1084[0:7]), .rgt_op_05(net1085[0:7]),
     .lft_op_08(net836[0:7]), .lft_op_07(net831[0:7]),
     .lft_op_06(net832[0:7]), .lft_op_05(net833[0:7]),
     .sp12_h_l_08(net1001[0:23]), .sp12_h_l_07(net1000[0:23]),
     .sp12_h_l_06(net999[0:23]), .sp12_h_r_05(net1093[0:23]),
     .sp12_h_r_06(net1094[0:23]), .sp12_h_r_07(net1095[0:23]),
     .sp12_h_r_08(net1096[0:23]), .sp12_h_l_05(net998[0:23]),
     .sp4_r_v_b_05(net1098[0:47]), .sp4_r_v_b_06(net1099[0:47]),
     .sp4_r_v_b_07(net1100[0:47]), .sp4_r_v_b_08(net1101[0:47]),
     .sp4_v_b_08(net1006[0:47]), .sp4_v_b_07(net1005[0:47]),
     .sp4_v_b_06(net1004[0:47]), .sp4_v_b_05(net1003[0:47]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .wl(wl_l[127:0]), .sp12_v_t_08(net1109[0:23]),
     .tnr_op_08({slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0], slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0]}), .top_op_08({slf_op_02_17[3],
     slf_op_02_17[2], slf_op_02_17[1], slf_op_02_17[0],
     slf_op_02_17[3], slf_op_02_17[2], slf_op_02_17[1],
     slf_op_02_17[0]}), .tnl_op_08({slf_op_01_17[3], slf_op_01_17[2],
     slf_op_01_17[1], slf_op_01_17[0], slf_op_01_17[3],
     slf_op_01_17[2], slf_op_01_17[1], slf_op_01_17[0]}),
     .sp4_v_t_08(net1113[0:47]), .lc_bot(lc_bot_02_09),
     .op_vic(net1458), .sp12_v_b_01(sp12_v_b_02_09[23:0]),
     .glb_netwk_t(net1117[0:7]));
lt_1x8_top_ice1f I_lt_col_t05 ( .glb_netwk_b(net1118[0:7]),
     .rgt_op_03(slf_op_06_11[7:0]), .slf_op_02(net1216[0:7]),
     .rgt_op_02(slf_op_06_10[7:0]), .rgt_op_01(slf_op_06_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net771[0:7]),
     .lft_op_03(net772[0:7]), .lft_op_02(net773[0:7]),
     .lft_op_01(slf_op_04_09[7:0]), .rgt_op_04(slf_op_06_12[7:0]),
     .carry_in(carry_in_05_09), .bnl_op_01(bnl_op_05_09[7:0]),
     .slf_op_04(net1224[0:7]), .slf_op_03(net1214[0:7]),
     .slf_op_01(slf_op_05_09[7:0]), .sp4_h_l_04(net1243[0:47]),
     .carry_out(net1136), .vdd_cntl(vdd_cntl_l[127:0]),
     .sp12_h_r_04(net1138[0:23]), .sp12_h_r_03(net1139[0:23]),
     .sp12_h_r_02(net1140[0:23]), .sp12_h_r_01(net1141[0:23]),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_05_09[47:0]), .sp4_r_v_b_04(net1144[0:47]),
     .sp4_r_v_b_03(net1145[0:47]), .sp4_r_v_b_02(net1146[0:47]),
     .sp4_r_v_b_01(sp4_v_b_06_09[47:0]), .sp4_h_r_04(net1148[0:47]),
     .sp4_h_r_03(net1149[0:47]), .sp4_h_r_02(net1150[0:47]),
     .sp4_h_r_01(net1151[0:47]), .sp4_h_l_03(net1244[0:47]),
     .sp4_h_l_02(net1245[0:47]), .sp4_h_l_01(net1246[0:47]),
     .bl(bl[275:222]), .bot_op_01(bot_op_05_09[7:0]),
     .sp12_h_l_01(net1236[0:23]), .sp12_h_l_02(net1235[0:23]),
     .sp12_h_l_03(net1234[0:23]), .sp12_h_l_04(net1233[0:23]),
     .sp4_v_b_04(net1239[0:47]), .sp4_v_b_03(net1240[0:47]),
     .sp4_v_b_02(net1241[0:47]), .bnr_op_01(bnr_op_05_09[7:0]),
     .sp4_h_l_05(net1267[0:47]), .sp4_h_l_06(net1266[0:47]),
     .sp4_h_l_07(net1265[0:47]), .sp4_h_l_08(net1264[0:47]),
     .sp4_h_r_08(net1169[0:47]), .sp4_h_r_07(net1170[0:47]),
     .sp4_h_r_06(net1171[0:47]), .sp4_h_r_05(net1172[0:47]),
     .slf_op_05(net1275[0:7]), .slf_op_06(net1274[0:7]),
     .slf_op_07(net1273[0:7]), .slf_op_08(net1272[0:7]),
     .rgt_op_08(slf_op_06_16[7:0]), .rgt_op_07(slf_op_06_15[7:0]),
     .rgt_op_06(slf_op_06_14[7:0]), .rgt_op_05(slf_op_06_13[7:0]),
     .lft_op_08(net767[0:7]), .lft_op_07(net768[0:7]),
     .lft_op_06(net769[0:7]), .lft_op_05(net770[0:7]),
     .sp12_h_l_08(net1286[0:23]), .sp12_h_l_07(net1285[0:23]),
     .sp12_h_l_06(net1284[0:23]), .sp12_h_r_05(net1188[0:23]),
     .sp12_h_r_06(net1189[0:23]), .sp12_h_r_07(net1190[0:23]),
     .sp12_h_r_08(net1191[0:23]), .sp12_h_l_05(net1283[0:23]),
     .sp4_r_v_b_05(net1193[0:47]), .sp4_r_v_b_06(net1194[0:47]),
     .sp4_r_v_b_07(net1195[0:47]), .sp4_r_v_b_08(net1196[0:47]),
     .sp4_v_b_08(net1291[0:47]), .sp4_v_b_07(net1290[0:47]),
     .sp4_v_b_06(net1289[0:47]), .sp4_v_b_05(net1288[0:47]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .wl(wl_l[127:0]), .sp12_v_t_08(net1204[0:23]),
     .tnr_op_08({slf_op_06_17[3], slf_op_06_17[2], slf_op_06_17[1],
     slf_op_06_17[0], slf_op_06_17[3], slf_op_06_17[2],
     slf_op_06_17[1], slf_op_06_17[0]}), .top_op_08({slf_op_05_17[3],
     slf_op_05_17[2], slf_op_05_17[1], slf_op_05_17[0],
     slf_op_05_17[3], slf_op_05_17[2], slf_op_05_17[1],
     slf_op_05_17[0]}), .tnl_op_08({slf_op_04_17[3], slf_op_04_17[2],
     slf_op_04_17[1], slf_op_04_17[0], slf_op_04_17[3],
     slf_op_04_17[2], slf_op_04_17[1], slf_op_04_17[0]}),
     .sp4_v_t_08(net1208[0:47]), .lc_bot(lc_bot_05_09),
     .op_vic(net1462), .sp12_v_b_01(sp12_v_b_05_09[23:0]),
     .glb_netwk_t(net1212[0:7]));
lt_1x8_top_ice1f I_lt_col_t04 ( .glb_netwk_b(net1213[0:7]),
     .rgt_op_03(net1214[0:7]), .slf_op_02(net773[0:7]),
     .rgt_op_02(net1216[0:7]), .rgt_op_01(slf_op_05_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net1034[0:7]),
     .lft_op_03(net1024[0:7]), .lft_op_02(net1026[0:7]),
     .lft_op_01(slf_op_03_09[7:0]), .rgt_op_04(net1224[0:7]),
     .carry_in(carry_in_04_09), .bnl_op_01(bnl_op_04_09[7:0]),
     .slf_op_04(net771[0:7]), .slf_op_03(net772[0:7]),
     .slf_op_01(slf_op_04_09[7:0]), .sp4_h_l_04(net792[0:47]),
     .carry_out(net1231), .vdd_cntl(vdd_cntl_l[127:0]),
     .sp12_h_r_04(net1233[0:23]), .sp12_h_r_03(net1234[0:23]),
     .sp12_h_r_02(net1235[0:23]), .sp12_h_r_01(net1236[0:23]),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_04_09[47:0]), .sp4_r_v_b_04(net1239[0:47]),
     .sp4_r_v_b_03(net1240[0:47]), .sp4_r_v_b_02(net1241[0:47]),
     .sp4_r_v_b_01(sp4_v_b_05_09[47:0]), .sp4_h_r_04(net1243[0:47]),
     .sp4_h_r_03(net1244[0:47]), .sp4_h_r_02(net1245[0:47]),
     .sp4_h_r_01(net1246[0:47]), .sp4_h_l_03(net791[0:47]),
     .sp4_h_l_02(net790[0:47]), .sp4_h_l_01(net746[0:47]),
     .bl(bl[221:168]), .bot_op_01(bot_op_04_09[7:0]),
     .sp12_h_l_01(net740[0:23]), .sp12_h_l_02(net748[0:23]),
     .sp12_h_l_03(net704[0:23]), .sp12_h_l_04(net749[0:23]),
     .sp4_v_b_04(net728[0:47]), .sp4_v_b_03(net724[0:47]),
     .sp4_v_b_02(net735[0:47]), .bnr_op_01(bnr_op_04_09[7:0]),
     .sp4_h_l_05(net793[0:47]), .sp4_h_l_06(net794[0:47]),
     .sp4_h_l_07(net795[0:47]), .sp4_h_l_08(net731[0:47]),
     .sp4_h_r_08(net1264[0:47]), .sp4_h_r_07(net1265[0:47]),
     .sp4_h_r_06(net1266[0:47]), .sp4_h_r_05(net1267[0:47]),
     .slf_op_05(net770[0:7]), .slf_op_06(net769[0:7]),
     .slf_op_07(net768[0:7]), .slf_op_08(net767[0:7]),
     .rgt_op_08(net1272[0:7]), .rgt_op_07(net1273[0:7]),
     .rgt_op_06(net1274[0:7]), .rgt_op_05(net1275[0:7]),
     .lft_op_08(net1082[0:7]), .lft_op_07(net1083[0:7]),
     .lft_op_06(net1084[0:7]), .lft_op_05(net1085[0:7]),
     .sp12_h_l_08(net721[0:23]), .sp12_h_l_07(net716[0:23]),
     .sp12_h_l_06(net718[0:23]), .sp12_h_r_05(net1283[0:23]),
     .sp12_h_r_06(net1284[0:23]), .sp12_h_r_07(net1285[0:23]),
     .sp12_h_r_08(net1286[0:23]), .sp12_h_l_05(net720[0:23]),
     .sp4_r_v_b_05(net1288[0:47]), .sp4_r_v_b_06(net1289[0:47]),
     .sp4_r_v_b_07(net1290[0:47]), .sp4_r_v_b_08(net1291[0:47]),
     .sp4_v_b_08(net763[0:47]), .sp4_v_b_07(net764[0:47]),
     .sp4_v_b_06(net765[0:47]), .sp4_v_b_05(net732[0:47]),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .wl(wl_l[127:0]), .sp12_v_t_08(net1299[0:23]),
     .tnr_op_08({slf_op_05_17[3], slf_op_05_17[2], slf_op_05_17[1],
     slf_op_05_17[0], slf_op_05_17[3], slf_op_05_17[2],
     slf_op_05_17[1], slf_op_05_17[0]}), .top_op_08({slf_op_04_17[3],
     slf_op_04_17[2], slf_op_04_17[1], slf_op_04_17[0],
     slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0]}), .tnl_op_08({slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0], slf_op_08_17[3],
     slf_op_08_17[2], slf_op_08_17[1], slf_op_08_17[0]}),
     .sp4_v_t_08(net1303[0:47]), .lc_bot(lc_bot_04_09),
     .op_vic(net1459), .sp12_v_b_01(sp12_v_b_04_09[23:0]),
     .glb_netwk_t(net1307[0:7]));
lt_1x8_top_ice1f I_lt_col_t06 ( .glb_netwk_b(net1460[0:7]),
     .rgt_op_03(rgt_op_06_11[7:0]), .slf_op_02(slf_op_06_10[7:0]),
     .rgt_op_02(rgt_op_06_10[7:0]), .rgt_op_01(rgt_op_06_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net1224[0:7]),
     .lft_op_03(net1214[0:7]), .lft_op_02(net1216[0:7]),
     .lft_op_01(slf_op_05_09[7:0]), .rgt_op_04(rgt_op_06_12[7:0]),
     .carry_in(carry_in_06_09), .bnl_op_01(bnl_op_06_09[7:0]),
     .slf_op_04(slf_op_06_12[7:0]), .slf_op_03(slf_op_06_11[7:0]),
     .slf_op_01(slf_op_06_09[7:0]), .sp4_h_l_04(net1148[0:47]),
     .carry_out(net1326), .vdd_cntl(vdd_cntl_l[127:0]),
     .sp12_h_r_04(sp12_h_r_06_12[23:0]),
     .sp12_h_r_03(sp12_h_r_06_11[23:0]),
     .sp12_h_r_02(sp12_h_r_06_10[23:0]),
     .sp12_h_r_01(sp12_h_r_06_09[23:0]),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_06_09[47:0]),
     .sp4_r_v_b_04(sp4_r_v_b_06_12[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_06_11[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_06_10[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_06_09[47:0]),
     .sp4_h_r_04(sp4_h_r_06_12[47:0]),
     .sp4_h_r_03(sp4_h_r_06_11[47:0]),
     .sp4_h_r_02(sp4_h_r_06_10[47:0]),
     .sp4_h_r_01(sp4_h_r_06_09[47:0]), .sp4_h_l_03(net1149[0:47]),
     .sp4_h_l_02(net1150[0:47]), .sp4_h_l_01(net1151[0:47]),
     .bl(bl[329:276]), .bot_op_01(bot_op_06_09[7:0]),
     .sp12_h_l_01(net1141[0:23]), .sp12_h_l_02(net1140[0:23]),
     .sp12_h_l_03(net1139[0:23]), .sp12_h_l_04(net1138[0:23]),
     .sp4_v_b_04(net1144[0:47]), .sp4_v_b_03(net1145[0:47]),
     .sp4_v_b_02(net1146[0:47]), .bnr_op_01(bnr_op_06_09[7:0]),
     .sp4_h_l_05(net1172[0:47]), .sp4_h_l_06(net1171[0:47]),
     .sp4_h_l_07(net1170[0:47]), .sp4_h_l_08(net1169[0:47]),
     .sp4_h_r_08(sp4_h_r_06_16[47:0]),
     .sp4_h_r_07(sp4_h_r_06_15[47:0]),
     .sp4_h_r_06(sp4_h_r_06_14[47:0]),
     .sp4_h_r_05(sp4_h_r_06_13[47:0]), .slf_op_05(slf_op_06_13[7:0]),
     .slf_op_06(slf_op_06_14[7:0]), .slf_op_07(slf_op_06_15[7:0]),
     .slf_op_08(slf_op_06_16[7:0]), .rgt_op_08(rgt_op_06_16[7:0]),
     .rgt_op_07(rgt_op_06_15[7:0]), .rgt_op_06(rgt_op_06_14[7:0]),
     .rgt_op_05(rgt_op_06_13[7:0]), .lft_op_08(net1272[0:7]),
     .lft_op_07(net1273[0:7]), .lft_op_06(net1274[0:7]),
     .lft_op_05(net1275[0:7]), .sp12_h_l_08(net1191[0:23]),
     .sp12_h_l_07(net1190[0:23]), .sp12_h_l_06(net1189[0:23]),
     .sp12_h_r_05(sp12_h_r_06_13[23:0]),
     .sp12_h_r_06(sp12_h_r_06_14[23:0]),
     .sp12_h_r_07(sp12_h_r_06_15[23:0]),
     .sp12_h_r_08(sp12_h_r_06_16[23:0]), .sp12_h_l_05(net1188[0:23]),
     .sp4_r_v_b_05(sp4_r_v_b_06_13[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_06_14[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_06_15[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_06_16[47:0]), .sp4_v_b_08(net1196[0:47]),
     .sp4_v_b_07(net1195[0:47]), .sp4_v_b_06(net1194[0:47]),
     .sp4_v_b_05(net1193[0:47]), .pgate(pgate_l[127:0]),
     .reset_b(reset_b_l[127:0]), .wl(wl_l[127:0]),
     .sp12_v_t_08(net1394[0:23]), .tnr_op_08({tnr_op_06_16[3],
     tnr_op_06_16[2], tnr_op_06_16[1], tnr_op_06_16[0],
     tnr_op_06_16[3], tnr_op_06_16[2], tnr_op_06_16[1],
     tnr_op_06_16[0]}), .top_op_08({slf_op_06_17[3], slf_op_06_17[2],
     slf_op_06_17[1], slf_op_06_17[0], slf_op_06_17[3],
     slf_op_06_17[2], slf_op_06_17[1], slf_op_06_17[0]}),
     .tnl_op_08({slf_op_05_17[3], slf_op_05_17[2], slf_op_05_17[1],
     slf_op_05_17[0], slf_op_05_17[3], slf_op_05_17[2],
     slf_op_05_17[1], slf_op_05_17[0]}), .sp4_v_t_08(net1398[0:47]),
     .lc_bot(lc_bot_06_09), .op_vic(net1465),
     .sp12_v_b_01(sp12_v_b_06_09[23:0]), .glb_netwk_t(net1402[0:7]));
tielo I369 ( .tielo(tiegnd_qtl));
tielo I365 ( .tielo(tiegnd_bram_t));
scan_buf_ice8p I_scanbuf_8p_tl ( .update_i(net1405), .tclk_i(net1406),
     .shift_i(net1407), .sdi(net1408), .r_i(net1409), .mode_i(net1410),
     .hiz_b_i(net1411), .ceb_i(net1412), .bs_en_i(net1413),
     .update_o(update_o), .tclk_o(net816), .shift_o(shift_o),
     .sdo(net803), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
fabric_buf_ice8p I385 ( .f_in(net1423), .f_out(fabric_out_00_09));
fabric_buf_ice8p I390 ( .f_in(net675), .f_out(padin_06_17b));
fabric_buf_ice8p I391 ( .f_in(net1427), .f_out(padin_00_09a));
fabric_buf_ice8p I388 ( .f_in(net859), .f_out(fabric_out_06_17));
clk_quad_buf_x8_ice8p I_clk_qtl_center ( .clko(clk_tree_drv_tl[7:0]),
     .clki(clk_center[7:0]));
clk_quad_buf_x8_ice8p I_clktree_quad_drv_tl ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));

endmodule
// Library - leafcell, Cell - pinlatbuf12p_1, View - schematic
// LAST TIME SAVED: Dec 24 09:06:49 2010
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module pinlatbuf12p_1 ( cout, cbit, icegate, pad_in, prog );
output  cout;

input  cbit, icegate, pad_in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I_txgate_lvt_2 ( .in(cout), .out(net13), .pp(net046),
     .nn(net17));
txgate_lvt I_txgate_lvt_1 ( .in(pad_in), .out(net13), .pp(net17),
     .nn(net046));
inv_lvt I6 ( .A(net046), .Y(net17));
inv_lvt I24 ( .A(prog), .Y(net19));
inv_lvt I_inv_lvt ( .A(net044), .Y(cout));
nand2_lvt I_nand2_lvt ( .A(net19), .Y(net044), .B(net13));
nand2_lvt I5 ( .A(icegate), .Y(net046), .B(cbit));

endmodule
// Library - ice1chip, Cell - io_rgt_bot_1x8_ice1f, View - schematic
// LAST TIME SAVED: Mar 10 17:31:55 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_rgt_bot_1x8_ice1f ( cf_r[191:0], fabric_out_01,
     fabric_out_02, fabric_out_08, padeb[12:0], pado[12:0], sdo,
     slf_op_01[3:0], slf_op_02[3:0], slf_op_03[3:0], slf_op_04[3:0],
     slf_op_05[3:0], slf_op_06[3:0], slf_op_07[3:0], slf_op_08[3:0],
     tck_pad, tclk_o, tdi_pad, tms_pad, SP4_h_l_01[47:0],
     SP4_h_l_02[47:0], SP4_h_l_03[47:0], SP4_h_l_04[47:0],
     SP4_h_l_05[47:0], SP4_h_l_06[47:0], SP4_h_l_07[47:0],
     SP4_h_l_08[47:0], SP12_h_l_01[23:0], SP12_h_l_02[23:0],
     SP12_h_l_03[23:0], SP12_h_l_04[23:0], SP12_h_l_05[23:0],
     SP12_h_l_06[23:0], SP12_h_l_07[23:0], SP12_h_l_08[23:0], bl[17:0],
     pgate[127:0], reset_b[127:0], sp4_v_b_13_09[15:0],
     sp4_v_t_08[15:0], vdd_cntl[127:0], wl[127:0], bnl_op_13_09[7:0],
     bs_en, ceb, glb_netwk_col[7:0], hiz_b, hold,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[2],
     last_rsr[3], lft_op_01[7:0], lft_op_02[7:0], lft_op_03[7:0],
     lft_op_04[7:0], lft_op_05[7:0], lft_op_06[7:0], lft_op_07[7:0],
     lft_op_08[7:0], mode, mux_jtag_sel_b, padin[12:0], prog, r, sdi,
     sdo_enable, shift, tclk, tnl_op_08[7:0], totdopad, trstb_pad,
     update );
output  fabric_out_01, fabric_out_02, fabric_out_08, sdo, tck_pad,
     tclk_o, tdi_pad, tms_pad;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, mode, mux_jtag_sel_b, prog, r, sdi,
     sdo_enable, shift, tclk, totdopad, trstb_pad, update;

output [3:0]  slf_op_01;
output [3:0]  slf_op_08;
output [3:0]  slf_op_07;
output [3:0]  slf_op_02;
output [3:0]  slf_op_06;
output [12:0]  pado;
output [3:0]  slf_op_03;
output [191:0]  cf_r;
output [12:0]  padeb;
output [3:0]  slf_op_05;
output [3:0]  slf_op_04;

inout [23:0]  SP12_h_l_02;
inout [23:0]  SP12_h_l_06;
inout [23:0]  SP12_h_l_07;
inout [23:0]  SP12_h_l_03;
inout [47:0]  SP4_h_l_04;
inout [17:0]  bl;
inout [23:0]  SP12_h_l_04;
inout [47:0]  SP4_h_l_05;
inout [15:0]  sp4_v_t_08;
inout [47:0]  SP4_h_l_01;
inout [47:0]  SP4_h_l_06;
inout [47:0]  SP4_h_l_02;
inout [23:0]  SP12_h_l_05;
inout [47:0]  SP4_h_l_08;
inout [47:0]  SP4_h_l_03;
inout [15:0]  sp4_v_b_13_09;
inout [127:0]  reset_b;
inout [127:0]  vdd_cntl;
inout [127:0]  wl;
inout [23:0]  SP12_h_l_01;
inout [127:0]  pgate;
inout [23:0]  SP12_h_l_08;
inout [47:0]  SP4_h_l_07;

input [7:0]  lft_op_01;
input [7:0]  lft_op_06;
input [7:0]  lft_op_04;
input [7:0]  lft_op_03;
input [7:0]  lft_op_05;
input [7:0]  lft_op_07;
input [7:0]  lft_op_02;
input [7:0]  lft_op_08;
input [7:0]  tnl_op_08;
input [2:3]  last_rsr;
input [7:0]  bnl_op_13_09;
input [12:0]  padin;
input [7:0]  glb_netwk_col;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net544;

wire  [0:15]  net400;

wire  [0:1]  net507;

wire  [0:7]  net584;

wire  [7:0]  glb_netwk_t;

wire  [11:36]  cf_rd;

wire  [0:1]  net345;

wire  [0:15]  net472;

wire  [7:0]  colbuf_cntl_t;

wire  [0:15]  net652;

wire  [0:1]  net350;

wire  [0:7]  net548;

wire  [7:0]  colbuf_cntl_b;

wire  [0:1]  net352;

wire  [0:15]  net580;

wire  [0:7]  net346;

wire  [0:1]  net344;

wire  [0:7]  net349;

wire  [0:15]  net616;

wire  [0:7]  net476;

wire  [0:1]  net360;

wire  [7:0]  glb_netwk_b;

wire  [0:1]  net363;

wire  [11:36]  cf_rp;

wire  [0:15]  net508;

wire  [0:1]  net361;

wire  [0:7]  net440;



mux2_hvt I_mux_jtagcf_2_ ( .in1(cf_rp[36]), .in0(vdd_),
     .out(cf_rd[36]), .sel(mux_jtag_sel_b));
mux2_hvt I_mux_jtagcf_1_ ( .in1(cf_rp[12]), .in0(vdd_),
     .out(cf_rd[12]), .sel(mux_jtag_sel_b));
mux2_hvt I_mux_jtagcf_0_ ( .in1(cf_rp[11]), .in0(vdd_),
     .out(cf_rd[11]), .sel(mux_jtag_sel_b));
bram_bufferx4 I_muxedjtagbuf_2_ ( .in(cf_rd[36]), .out(cf_r[36]));
bram_bufferx4 I_muxedjtagbuf_1_ ( .in(cf_rd[12]), .out(cf_r[12]));
bram_bufferx4 I_muxedjtagbuf_0_ ( .in(cf_rd[11]), .out(cf_r[11]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tiegnd));
tckbufx32_ice8p I_tmsbuf ( .in(tms), .out(tms_pad));
tckbufx32_ice8p I_tckbuf ( .in(tck), .out(tck_pad));
tckbufx32_ice8p I_tdibuf ( .in(tdi), .out(tdi_pad));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
io_col4_rgt_ice8p_v2 I_io_00_02 ( .slf_op(slf_op_02[3:0]),
     .cdone_in(trstb_pad), .spioeb({sdo_enable, tievdd}),
     .tnl_op(lft_op_03[7:0]), .spi_ss_in_b({nc_ss, tck}), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_02[23:0]),
     .spiout({totdopad, tiegnd}), .sp4_v_b(net580[0:15]), .prog(prog),
     .cf({cf_r[47:37], cf_rp[36], cf_r[35:24]}),
     .vdd_cntl(vdd_cntl[31:16]), .lft_op(lft_op_02[7:0]),
     .padin(padin[3:2]), .mode(mode), .wl(wl[31:16]), .pado(pado[3:2]),
     .sp4_v_t(net400[0:15]), .padeb(padeb[3:2]),
     .reset(reset_b[31:16]), .bl(bl[17:0]), .cbit_colcntl(net346[0:7]),
     .sdo(net405), .fabric_out(fabric_out_02),
     .glb_netwk(glb_netwk_b[7:0]), .pgate(pgate[31:16]), .sdi(net585),
     .sp4_h_l(SP4_h_l_02[47:0]), .bnl_op(lft_op_01[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_08 ( .slf_op(slf_op_08[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(tnl_op_08[7:0]), .spi_ss_in_b(net361[0:1]), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_08[23:0]),
     .spiout({tiegnd, tiegnd}), .sp4_v_b(net472[0:15]), .prog(prog),
     .cf(cf_r[191:168]), .vdd_cntl(vdd_cntl[127:112]),
     .lft_op(lft_op_08[7:0]), .padin(padin[12:11]), .mode(mode),
     .wl(wl[127:112]), .pado(pado[12:11]), .sp4_v_t(sp4_v_t_08[15:0]),
     .padeb(padeb[12:11]), .reset(reset_b[127:112]), .bl(bl[17:0]),
     .cbit_colcntl(net440[0:7]), .sdo(sdo), .fabric_out(fabric_out_08),
     .glb_netwk(glb_netwk_t[7:0]), .pgate(pgate[127:112]),
     .sdi(net477), .sp4_h_l(SP4_h_l_08[47:0]),
     .bnl_op(lft_op_07[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_07 ( .slf_op(slf_op_07[3:0]),
     .cdone_in(jtag_rowtest_mode_rowu3_b), .spioeb({tievdd, tiegnd}),
     .tnl_op(lft_op_08[7:0]), .spi_ss_in_b(net352[0:1]), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_07[23:0]),
     .spiout({tiegnd, last_rsr[3]}), .sp4_v_b(net544[0:15]),
     .prog(prog), .cf(cf_r[167:144]), .vdd_cntl(vdd_cntl[111:96]),
     .lft_op(lft_op_07[7:0]), .padin(padin[10:9]), .mode(mode),
     .wl(wl[111:96]), .pado(pado[10:9]), .sp4_v_t(net472[0:15]),
     .padeb(padeb[10:9]), .reset(reset_b[111:96]), .bl(bl[17:0]),
     .cbit_colcntl(net476[0:7]), .sdo(net477), .fabric_out(net478),
     .glb_netwk(glb_netwk_t[7:0]), .pgate(pgate[111:96]), .sdi(net549),
     .sp4_h_l(SP4_h_l_07[47:0]), .bnl_op(lft_op_06[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_05 ( .slf_op(slf_op_05[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_06[7:0]), .spi_ss_in_b(net345[0:1]), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_05[23:0]),
     .spiout({tiegnd, tiegnd}), .sp4_v_b(net652[0:15]), .prog(prog),
     .cf(cf_r[119:96]), .vdd_cntl(vdd_cntl[79:64]),
     .lft_op(lft_op_05[7:0]), .padin(net507[0:1]), .mode(mode),
     .wl(wl[79:64]), .pado(net507[0:1]), .sp4_v_t(net508[0:15]),
     .padeb(net363[0:1]), .reset(reset_b[79:64]), .bl(bl[17:0]),
     .cbit_colcntl(colbuf_cntl_t[7:0]), .sdo(net513),
     .fabric_out(net514), .glb_netwk(glb_netwk_t[7:0]),
     .pgate(pgate[79:64]), .sdi(net657), .sp4_h_l(SP4_h_l_05[47:0]),
     .bnl_op(lft_op_04[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_06 ( .slf_op(slf_op_06[3:0]),
     .cdone_in(jtag_rowtest_mode_rowu2_b), .spioeb({tievdd, tiegnd}),
     .tnl_op(lft_op_07[7:0]), .spi_ss_in_b(net360[0:1]), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_06[23:0]),
     .spiout({tiegnd, last_rsr[2]}), .sp4_v_b(net508[0:15]),
     .prog(prog), .cf(cf_r[143:120]), .vdd_cntl(vdd_cntl[95:80]),
     .lft_op(lft_op_06[7:0]), .padin(padin[8:7]), .mode(mode),
     .wl(wl[95:80]), .pado(pado[8:7]), .sp4_v_t(net544[0:15]),
     .padeb(padeb[8:7]), .reset(reset_b[95:80]), .bl(bl[17:0]),
     .cbit_colcntl(net548[0:7]), .sdo(net549), .fabric_out(net550),
     .glb_netwk(glb_netwk_t[7:0]), .pgate(pgate[95:80]), .sdi(net513),
     .sp4_h_l(SP4_h_l_06[47:0]), .bnl_op(lft_op_05[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_01 ( .slf_op(slf_op_01[3:0]),
     .cdone_in(mux_jtag_sel_b), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_02[7:0]), .spi_ss_in_b({tms, tdi}), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_01[23:0]),
     .spiout({tiegnd, tiegnd}), .sp4_v_b(sp4_v_b_13_09[15:0]),
     .prog(prog), .cf({cf_r[23:13], cf_rp[12], cf_rp[11], cf_r[10:0]}),
     .vdd_cntl(vdd_cntl[15:0]), .lft_op(lft_op_01[7:0]),
     .padin(padin[1:0]), .mode(mode), .wl(wl[15:0]), .pado(pado[1:0]),
     .sp4_v_t(net580[0:15]), .padeb(padeb[1:0]), .reset(reset_b[15:0]),
     .bl(bl[17:0]), .cbit_colcntl(net584[0:7]), .sdo(net585),
     .fabric_out(fabric_out_01), .glb_netwk(glb_netwk_b[7:0]),
     .pgate(pgate[15:0]), .sdi(sdi), .sp4_h_l(SP4_h_l_01[47:0]),
     .bnl_op(bnl_op_13_09[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_03 ( .slf_op(slf_op_03[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_04[7:0]), .spi_ss_in_b(net350[0:1]), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_03[23:0]),
     .spiout({tiegnd, tiegnd}), .sp4_v_b(net400[0:15]), .prog(prog),
     .cf(cf_r[71:48]), .vdd_cntl(vdd_cntl[47:32]),
     .lft_op(lft_op_03[7:0]), .padin({padin[4], padin_nc}),
     .mode(mode), .wl(wl[47:32]), .pado({pado[4], pado_nc}),
     .sp4_v_t(net616[0:15]), .padeb({padeb[4], padeb_nc}),
     .reset(reset_b[47:32]), .bl(bl[17:0]), .cbit_colcntl(net349[0:7]),
     .sdo(net621), .fabric_out(net622), .glb_netwk(glb_netwk_b[7:0]),
     .pgate(pgate[47:32]), .sdi(net405), .sp4_h_l(SP4_h_l_03[47:0]),
     .bnl_op(lft_op_02[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_04 ( .slf_op(slf_op_04[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_05[7:0]), .spi_ss_in_b(net344[0:1]), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_04[23:0]),
     .spiout({tiegnd, tiegnd}), .sp4_v_b(net616[0:15]), .prog(prog),
     .cf(cf_r[95:72]), .vdd_cntl(vdd_cntl[63:48]),
     .lft_op(lft_op_04[7:0]), .padin(padin[6:5]), .mode(mode),
     .wl(wl[63:48]), .pado(pado[6:5]), .sp4_v_t(net652[0:15]),
     .padeb(padeb[6:5]), .reset(reset_b[63:48]), .bl(bl[17:0]),
     .cbit_colcntl(colbuf_cntl_b[7:0]), .sdo(net657),
     .fabric_out(net658), .glb_netwk(glb_netwk_b[7:0]),
     .pgate(pgate[63:48]), .sdi(net621), .sp4_h_l(SP4_h_l_04[47:0]),
     .bnl_op(lft_op_03[7:0]));

endmodule
// Library - ice8chip, Cell - io_col4_bot_ice8p, View - schematic
// LAST TIME SAVED: Jan 12 14:58:38 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_col4_bot_ice8p ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [23:0]  cf;
output [1:0]  pado;
output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;

inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;

input [1:0]  padin;
input [1:0]  spiout;
input [15:0]  reset;
input [15:0]  pgate;
input [7:0]  glb_netwk;
input [1:0]  spioeb;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [15:0]  wl;
input [15:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [0:7]  net225;



inv_lvt I_inv1 ( .A(prog), .Y(progb));
inv_lvt I_inv2 ( .A(progb), .Y(progd));
io_gmux_x16bare_v3 I_io_gmux_x16bare_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .cbitb_colcntl(net225[0:7]), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29],
     sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13],
     sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5],
     tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
sbox1_colbdlc_v3 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
rm6w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));

endmodule
// Library - ice1chip, Cell - io_bot_rgt_1x6_ice1f, View - schematic
// LAST TIME SAVED: Jun 22 09:34:02 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_bot_rgt_1x6_ice1f ( cf_b_r[143:0], fabric_out_07_00,
     fabric_out_12_00, padeb_b_r[11], padeb_b_r[23:13], pado_b_r[11],
     pado_b_r[23:13], sdo_pad, slf_op_01_00[3:0], slf_op_02_00[3:0],
     slf_op_03_00[3:0], slf_op_04_00[3:0], slf_op_05_00[3:0],
     slf_op_06_00[3:0], spi_ss_in_bbank[4:0], bl_01[53:0], bl_02[53:0],
     bl_03[53:0], bl_04[41:0], bl_05[53:0], bl_06[53:0],
     sp4_h_l_07_00[15:0], sp4_h_r_12_17[15:0], sp4_v_b_01_00[47:0],
     sp4_v_b_02_00[47:0], sp4_v_b_03_00[47:0], sp4_v_b_04_00[47:0],
     sp4_v_b_05_00[47:0], sp4_v_b_06_00[47:0], sp12_v_b_01_00[23:0],
     sp12_v_b_02_00[23:0], sp12_v_b_03_00[23:0], sp12_v_b_04_00[23:0],
     sp12_v_b_05_00[23:0], sp12_v_b_06_00[23:0], bnl_op_01_00[7:0],
     bs_en_i, ceb_i, end_of_startup, glb_net_01[7:0], glb_net_02[7:0],
     glb_net_03[7:0], glb_net_04[7:0], glb_net_05[7:0],
     glb_net_06[7:0], hiz_b_i, hold_b_r, lft_op_01_00[7:0],
     lft_op_02_00[7:0], lft_op_03_00[7:0], lft_op_04_00[7:0],
     lft_op_05_00[7:0], lft_op_06_00[7:0], md_spi_b, mode_i,
     padin_b_r[11], padin_b_r[23:13], pgate_l[15:0], prog, r_i,
     reset_l[15:0], sdi, shift_i, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk_i, tnr_op_06_00[7:0], update_i, vdd_cntl_l[15:0],
     wl_l[15:0] );
output  fabric_out_07_00, fabric_out_12_00, sdo_pad;


input  bs_en_i, ceb_i, end_of_startup, hiz_b_i, hold_b_r, md_spi_b,
     mode_i, prog, r_i, sdi, shift_i, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk_i, update_i;

output [3:0]  slf_op_06_00;
output [3:0]  slf_op_01_00;
output [3:0]  slf_op_04_00;
output [143:0]  cf_b_r;
output [4:0]  spi_ss_in_bbank;
output [23:11]  pado_b_r;
output [23:11]  padeb_b_r;
output [3:0]  slf_op_02_00;
output [3:0]  slf_op_03_00;
output [3:0]  slf_op_05_00;

inout [47:0]  sp4_v_b_03_00;
inout [23:0]  sp12_v_b_03_00;
inout [47:0]  sp4_v_b_01_00;
inout [15:0]  sp4_h_l_07_00;
inout [53:0]  bl_06;
inout [47:0]  sp4_v_b_05_00;
inout [15:0]  sp4_h_r_12_17;
inout [23:0]  sp12_v_b_06_00;
inout [53:0]  bl_02;
inout [47:0]  sp4_v_b_04_00;
inout [23:0]  sp12_v_b_02_00;
inout [23:0]  sp12_v_b_01_00;
inout [53:0]  bl_01;
inout [53:0]  bl_05;
inout [47:0]  sp4_v_b_02_00;
inout [23:0]  sp12_v_b_05_00;
inout [23:0]  sp12_v_b_04_00;
inout [41:0]  bl_04;
inout [47:0]  sp4_v_b_06_00;
inout [53:0]  bl_03;

input [7:0]  glb_net_06;
input [7:0]  glb_net_04;
input [7:0]  glb_net_01;
input [15:0]  vdd_cntl_l;
input [7:0]  bnl_op_01_00;
input [7:0]  lft_op_06_00;
input [7:0]  lft_op_03_00;
input [15:0]  wl_l;
input [7:0]  lft_op_01_00;
input [7:0]  tnr_op_06_00;
input [15:0]  pgate_l;
input [7:0]  glb_net_03;
input [7:0]  glb_net_05;
input [7:0]  glb_net_02;
input [7:0]  lft_op_04_00;
input [7:0]  lft_op_05_00;
input [7:0]  lft_op_02_00;
input [15:0]  reset_l;
input [23:11]  padin_b_r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net374;

wire  [0:1]  net543;

wire  [0:1]  net545;

wire  [0:15]  net339;

wire  [132:83]  cf_b_r_pd;

wire  [0:1]  net546;

wire  [0:15]  net409;

wire  [132:83]  cf_b_r_p;

wire  [0:15]  net444;

wire  [0:15]  net514;



bram_bufferx4 I_cfbuf_spiss_ck_1_ ( .in(cf_b_r_pd[132]),
     .out(cf_b_r[132]));
bram_bufferx4 I_cfbuf_spiss_ck_0_ ( .in(cf_b_r_pd[131]),
     .out(cf_b_r[131]));
bram_bufferx4 I_buf_spisdi ( .in(cf_b_r_pd[107]), .out(cf_b_r[107]));
bram_bufferx4 I_buf_coldboot_1_ ( .in(cf_b_r_pd[84]),
     .out(cf_b_r[84]));
bram_bufferx4 I_buf_coldboot_0_ ( .in(cf_b_r_pd[83]),
     .out(cf_b_r[83]));
mux2_hvt I_cfmux_spiss_ck_1_ ( .in1(cf_b_r_p[132]),
     .in0(tiegnd_preIO_br), .out(cf_b_r_pd[132]),
     .sel(end_of_startup));
mux2_hvt I_cfmux_spiss_ck_0_ ( .in1(cf_b_r_p[131]),
     .in0(tiegnd_preIO_br), .out(cf_b_r_pd[131]),
     .sel(end_of_startup));
mux2_hvt I_cfmux_spisdi ( .in1(cf_b_r_p[107]), .in0(tiegnd_preIO_br),
     .out(cf_b_r_pd[107]), .sel(end_of_startup));
mux2_hvt I_cfmux_coldboot_1_ ( .in1(cf_b_r_p[84]),
     .in0(tiegnd_preIO_br), .out(cf_b_r_pd[84]), .sel(end_of_startup));
mux2_hvt I_cfmux_coldboot_0_ ( .in1(cf_b_r_p[83]),
     .in0(tiegnd_preIO_br), .out(cf_b_r_pd[83]), .sel(end_of_startup));
bram_bufferx4x6 I_bram_bufferx4x6 ( .in(net463), .out(net301));
lowla_modified I_lowla_modified ( .clk(endtck), .min(net301),
     .lao(sdo_pad));
scan_buf_ice8p I_scanbuf_8p_mb ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net314), .tclk_o(net315), .shift_o(net316),
     .sdo(net317), .r_o(net318), .mode_o(net319), .hiz_b_o(net320),
     .ceb_o(net321), .bs_en_o(net322));
io_col4_bot_ice8p I_IO_08_00 ( .sdo(net323), .sdi(net393),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net409[0:15]), .mode(net319), .shift(net316),
     .hiz_b(net320), .r(net318), .bs_en(net322), .tclk(endtck),
     .update(net314), .padin(padin_b_r[15:14]), .pado(pado_b_r[15:14]),
     .padeb(padeb_b_r[15:14]), .sp4_v_b(net339[0:15]),
     .sp4_h_l(sp4_v_b_02_00[47:0]), .sp12_h_l(sp12_v_b_02_00[23:0]),
     .prog(prog), .spi_ss_in_b(net545[0:1]),
     .tnl_op(lft_op_01_00[7:0]), .lft_op(lft_op_02_00[7:0]),
     .bnl_op(lft_op_03_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_b_r[47:24]), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_00[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_b_r), .fabric_out(net357));
io_col4_bot_ice8p I_IO_10_00_bram ( .sdo(net358), .sdi(net498),
     .spiout({tielow, tielow}), .cdone_in(end_of_startup),
     .spioeb({tievdd, tievdd}), .sp4_v_t(net514[0:15]), .mode(net319),
     .shift(net316), .hiz_b(net320), .r(net318), .bs_en(net322),
     .tclk(endtck), .update(net314), .padin(padin_b_r[19:18]),
     .pado(pado_b_r[19:18]), .padeb(padeb_b_r[19:18]),
     .sp4_v_b(net374[0:15]), .sp4_h_l(sp4_v_b_04_00[47:0]),
     .sp12_h_l(sp12_v_b_04_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_bbank[1:0]), .tnl_op(lft_op_03_00[7:0]),
     .lft_op(lft_op_04_00[7:0]), .bnl_op(lft_op_05_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_04[5],
     bl_04[4], bl_04[37], bl_04[36], bl_04[35], bl_04[34], bl_04[33],
     bl_04[32], bl_04[14], bl_04[20], bl_04[19], bl_04[18], bl_04[17],
     bl_04[16], bl_04[27], bl_04[26], bl_04[25], bl_04[23]}),
     .wl(wl_l[15:0]), .cf({cf_b_r[95:85], cf_b_r_p[84:83],
     cf_b_r[82:72]}), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_00[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_b_r), .fabric_out(net392));
io_col4_bot_ice8p I_IO_07_00 ( .sdo(net393), .sdi(net317),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_07_00[15:0]), .mode(net319),
     .shift(net316), .hiz_b(net320), .r(net318), .bs_en(net322),
     .tclk(endtck), .update(net314), .padin({padin_b_r[13],
     padin_b_r[11]}), .pado({pado_b_r[13], pado_b_r[11]}),
     .padeb({padeb_b_r[13], padeb_b_r[11]}), .sp4_v_b(net409[0:15]),
     .sp4_h_l(sp4_v_b_01_00[47:0]), .sp12_h_l(sp12_v_b_01_00[23:0]),
     .prog(prog), .spi_ss_in_b(net546[0:1]),
     .tnl_op(bnl_op_01_00[7:0]), .lft_op(lft_op_01_00[7:0]),
     .bnl_op(lft_op_02_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_b_r[23:0]), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_00[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_b_r), .fabric_out(fabric_out_07_00));
io_col4_bot_ice8p I_IO_11_00 ( .sdo(net428), .sdi(net358),
     .spiout({tielow, spi_sdo}), .cdone_in(end_of_startup),
     .spioeb({tievdd, spi_sdo_oe_b}), .sp4_v_t(net374[0:15]),
     .mode(net319), .shift(net316), .hiz_b(net320), .r(net318),
     .bs_en(net322), .tclk(endtck), .update(net314),
     .padin(padin_b_r[21:20]), .pado(pado_b_r[21:20]),
     .padeb(padeb_b_r[21:20]), .sp4_v_b(net444[0:15]),
     .sp4_h_l(sp4_v_b_05_00[47:0]), .sp12_h_l(sp12_v_b_05_00[23:0]),
     .prog(prog), .spi_ss_in_b({spi_ss_in_bbank[2], spi_ss_nc}),
     .tnl_op(lft_op_04_00[7:0]), .lft_op(lft_op_05_00[7:0]),
     .bnl_op(lft_op_06_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf({cf_b_r[119:108], cf_b_r_p[107], cf_b_r[106:96]}),
     .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_00[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_b_r), .fabric_out(net462));
io_col4_bot_ice8p I_IO_12_00 ( .sdo(net463), .sdi(net428),
     .spiout({spi_ss_out, spi_clk_out}), .cdone_in(end_of_startup),
     .spioeb({md_spi_b, md_spi_b}), .sp4_v_t(net444[0:15]),
     .mode(net319), .shift(net316), .hiz_b(net320), .r(net318),
     .bs_en(net322), .tclk(endtck), .update(net314),
     .padin(padin_b_r[23:22]), .pado(pado_b_r[23:22]),
     .padeb(padeb_b_r[23:22]), .sp4_v_b(sp4_h_r_12_17[15:0]),
     .sp4_h_l(sp4_v_b_06_00[47:0]), .sp12_h_l(sp12_v_b_06_00[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_bbank[4:3]),
     .tnl_op(lft_op_05_00[7:0]), .lft_op(lft_op_06_00[7:0]),
     .bnl_op(tnr_op_06_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_06[5], bl_06[4], bl_06[37],
     bl_06[36], bl_06[35], bl_06[34], bl_06[33], bl_06[32], bl_06[14],
     bl_06[20], bl_06[19], bl_06[18], bl_06[17], bl_06[16], bl_06[27],
     bl_06[26], bl_06[25], bl_06[23]}), .wl(wl_l[15:0]),
     .cf({cf_b_r[143:133], cf_b_r_p[132:131], cf_b_r[130:120]}),
     .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_00[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_b_r), .fabric_out(fabric_out_12_00));
io_col4_bot_ice8p I_IO_09_00 ( .sdo(net498), .sdi(net323),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net339[0:15]), .mode(net319), .shift(net316),
     .hiz_b(net320), .r(net318), .bs_en(net322), .tclk(endtck),
     .update(net314), .padin(padin_b_r[17:16]), .pado(pado_b_r[17:16]),
     .padeb(padeb_b_r[17:16]), .sp4_v_b(net514[0:15]),
     .sp4_h_l(sp4_v_b_03_00[47:0]), .sp12_h_l(sp12_v_b_03_00[23:0]),
     .prog(prog), .spi_ss_in_b(net543[0:1]),
     .tnl_op(lft_op_02_00[7:0]), .lft_op(lft_op_03_00[7:0]),
     .bnl_op(lft_op_04_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_b_r[71:48]), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_00[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_b_r), .fabric_out(net544));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(net315), .out(endtck));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x tielo4x_t ( .tielo(tiegnd_preIO_br));
tielo4x I483 ( .tielo(tielow));

endmodule
// Library - leafcell, Cell - clkbuffer200u, View - schematic
// LAST TIME SAVED: Jun 30 10:54:26 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module clkbuffer200u ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - ice1chip, Cell - lt_1x8_bot_ice1f, View - schematic
// LAST TIME SAVED: Jun  6 13:25:37 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module lt_1x8_bot_ice1f ( carry_out, glb_netwk_bot, op_vic, slf_op_01,
     slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07,
     slf_op_08, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02, sp4_h_l_03,
     sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07, sp4_h_l_08,
     sp4_h_r_01, sp4_h_r_02, sp4_h_r_03, sp4_h_r_04, sp4_h_r_05,
     sp4_h_r_06, sp4_h_r_07, sp4_h_r_08, sp4_r_v_b_01, sp4_r_v_b_02,
     sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05, sp4_r_v_b_06,
     sp4_r_v_b_07, sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03,
     sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07, sp4_v_b_08,
     sp4_v_t_08, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04,
     sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_r_01,
     sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06,
     sp12_h_r_07, sp12_h_r_08, sp12_v_b_01, sp12_v_t_08, vdd_cntl, wl,
     bnl_op_01, bnr_op_01, bot_op_01, carry_in, glb_netwk_col, lc_bot,
     lft_op_01, lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06,
     lft_op_07, lft_op_08, prog, purst, rgt_op_01, rgt_op_02,
     rgt_op_03, rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08,
     tnl_op_08, tnr_op_08, top_op_08 );
output  carry_out, op_vic;


input  carry_in, lc_bot, prog, purst;

output [7:0]  slf_op_01;
output [7:0]  slf_op_08;
output [7:0]  slf_op_04;
output [7:0]  slf_op_02;
output [7:0]  slf_op_03;
output [7:0]  glb_netwk_bot;
output [7:0]  slf_op_05;
output [7:0]  slf_op_07;
output [7:0]  slf_op_06;

inout [47:0]  sp4_h_l_01;
inout [23:0]  sp12_h_l_06;
inout [23:0]  sp12_v_b_01;
inout [23:0]  sp12_h_l_01;
inout [23:0]  sp12_h_r_05;
inout [23:0]  sp12_h_r_08;
inout [47:0]  sp4_r_v_b_05;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_v_b_03;
inout [47:0]  sp4_h_l_05;
inout [53:0]  bl;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_r_v_b_02;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_v_b_05;
inout [47:0]  sp4_h_l_02;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_01;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_v_b_02;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_v_b_06;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_v_t_08;
inout [47:0]  sp4_h_r_03;
inout [23:0]  sp12_v_t_08;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_v_b_07;
inout [23:0]  sp12_h_l_04;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_h_l_08;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_h_l_07;
inout [23:0]  sp12_h_r_04;
inout [47:0]  sp4_h_r_08;
inout [47:0]  sp4_h_l_06;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_h_l_03;
inout [47:0]  sp4_r_v_b_01;
inout [23:0]  sp12_h_l_05;
inout [127:0]  pgate;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_h_l_04;
inout [127:0]  vdd_cntl;
inout [127:0]  wl;
inout [47:0]  sp4_v_b_04;
inout [127:0]  reset_b;

input [7:0]  rgt_op_06;
input [7:0]  lft_op_08;
input [7:0]  tnl_op_08;
input [7:0]  glb_netwk_col;
input [7:0]  bot_op_01;
input [7:0]  rgt_op_01;
input [7:0]  top_op_08;
input [7:0]  tnr_op_08;
input [7:0]  lft_op_06;
input [7:0]  lft_op_05;
input [7:0]  rgt_op_04;
input [7:0]  lft_op_03;
input [7:0]  bnr_op_01;
input [7:0]  lft_op_01;
input [7:0]  lft_op_02;
input [7:0]  rgt_op_02;
input [7:0]  bnl_op_01;
input [7:0]  rgt_op_08;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_04;
input [7:0]  lft_op_07;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_05;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net0755;

wire  [0:7]  net1056;

wire  [0:23]  net1130;

wire  [7:0]  colbuf_cntl_bot;

wire  [0:7]  net932;

wire  [7:0]  glb_netwk_top;

wire  [0:23]  net1037;

wire  [0:23]  net1068;

wire  [0:23]  net975;

wire  [0:23]  net944;

wire  [0:7]  net1118;

wire  [0:23]  net1099;

wire  [0:7]  net1087;

wire  [0:7]  net963;

wire  [0:23]  net1006;

wire  [7:0]  colbuf_cntl_top;



ltile4_ice1f I_LT06 ( .cntl_cbit(net963[0:7]), .op_bot(net996),
     .op_vic(net965), .prog(prog), .carry_out(net967),
     .lft_op(lft_op_06[7:0]), .sp12_h_l(sp12_h_l_06[23:0]),
     .sp4_h_l(sp4_h_l_06[47:0]), .sp4_v_b(sp4_v_b_06[47:0]),
     .sp12_v_b(net1006[0:23]), .sp12_h_r(sp12_h_r_06[23:0]),
     .sp4_h_r(sp4_h_r_06[47:0]), .sp12_v_t(net975[0:23]),
     .sp4_v_t(sp4_v_b_07[47:0]), .sp4_r_v_b(sp4_r_v_b_06[47:0]),
     .wl(wl[95:80]), .top_op(slf_op_07[7:0]), .rgt_op(rgt_op_06[7:0]),
     .bot_op(slf_op_05[7:0]), .bl(bl[53:0]), .reset_b(reset_b[95:80]),
     .vdd_cntl(vdd_cntl[95:80]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net998), .purst(purst), .slf_op(slf_op_06[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_05[7:0]),
     .bnl_op(lft_op_05[7:0]), .tnr_op(rgt_op_07[7:0]),
     .tnl_op(lft_op_07[7:0]));
ltile4_ice1f I_LT03 ( .cntl_cbit(net1056[0:7]), .op_bot(net1089),
     .op_vic(net1058), .prog(prog), .carry_out(net1060),
     .lft_op(lft_op_03[7:0]), .sp12_h_l(sp12_h_l_03[23:0]),
     .sp4_h_l(sp4_h_l_03[47:0]), .sp4_v_b(sp4_v_b_03[47:0]),
     .sp12_v_b(net1099[0:23]), .sp12_h_r(sp12_h_r_03[23:0]),
     .sp4_h_r(sp4_h_r_03[47:0]), .sp12_v_t(net1068[0:23]),
     .sp4_v_t(sp4_v_b_04[47:0]), .sp4_r_v_b(sp4_r_v_b_03[47:0]),
     .wl(wl[47:32]), .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net1091), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4_ice1f I_LT04 ( .cntl_cbit(colbuf_cntl_bot[7:0]),
     .op_bot(net1058), .op_vic(net1027), .prog(prog),
     .carry_out(net1029), .lft_op(lft_op_04[7:0]),
     .sp12_h_l(sp12_h_l_04[23:0]), .sp4_h_l(sp4_h_l_04[47:0]),
     .sp4_v_b(sp4_v_b_04[47:0]), .sp12_v_b(net1068[0:23]),
     .sp12_h_r(sp12_h_r_04[23:0]), .sp4_h_r(sp4_h_r_04[47:0]),
     .sp12_v_t(net1037[0:23]), .sp4_v_t(sp4_v_b_05[47:0]),
     .sp4_r_v_b(sp4_r_v_b_04[47:0]), .wl(wl[63:48]),
     .top_op(slf_op_05[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net1060), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(rgt_op_05[7:0]),
     .tnl_op(lft_op_05[7:0]));
ltile4_ice1f I_LT05 ( .cntl_cbit(colbuf_cntl_top[7:0]),
     .op_bot(net1027), .op_vic(net996), .prog(prog),
     .carry_out(net998), .lft_op(lft_op_05[7:0]),
     .sp12_h_l(sp12_h_l_05[23:0]), .sp4_h_l(sp4_h_l_05[47:0]),
     .sp4_v_b(sp4_v_b_05[47:0]), .sp12_v_b(net1037[0:23]),
     .sp12_h_r(sp12_h_r_05[23:0]), .sp4_h_r(sp4_h_r_05[47:0]),
     .sp12_v_t(net1006[0:23]), .sp4_v_t(sp4_v_b_06[47:0]),
     .sp4_r_v_b(sp4_r_v_b_05[47:0]), .wl(wl[79:64]),
     .top_op(slf_op_06[7:0]), .rgt_op(rgt_op_05[7:0]),
     .bot_op(slf_op_04[7:0]), .bl(bl[53:0]), .reset_b(reset_b[79:64]),
     .vdd_cntl(vdd_cntl[79:64]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net1029), .purst(purst), .slf_op(slf_op_05[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_04[7:0]),
     .bnl_op(lft_op_04[7:0]), .tnr_op(rgt_op_06[7:0]),
     .tnl_op(lft_op_06[7:0]));
ltile4_ice1f I_LT01 ( .cntl_cbit(net1118[0:7]), .op_bot(lc_bot),
     .op_vic(net1120), .prog(prog), .carry_out(net1122),
     .lft_op(lft_op_01[7:0]), .sp12_h_l(sp12_h_l_01[23:0]),
     .sp4_h_l(sp4_h_l_01[47:0]), .sp4_v_b(sp4_v_b_01[47:0]),
     .sp12_v_b(sp12_v_b_01[23:0]), .sp12_h_r(sp12_h_r_01[23:0]),
     .sp4_h_r(sp4_h_r_01[47:0]), .sp12_v_t(net1130[0:23]),
     .sp4_v_t(sp4_v_b_02[47:0]), .sp4_r_v_b(sp4_r_v_b_01[47:0]),
     .wl(wl[15:0]), .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4_ice1f I_LT02 ( .cntl_cbit(net1087[0:7]), .op_bot(net1120),
     .op_vic(net1089), .prog(prog), .carry_out(net1091),
     .lft_op(lft_op_02[7:0]), .sp12_h_l(sp12_h_l_02[23:0]),
     .sp4_h_l(sp4_h_l_02[47:0]), .sp4_v_b(sp4_v_b_02[47:0]),
     .sp12_v_b(net1130[0:23]), .sp12_h_r(sp12_h_r_02[23:0]),
     .sp4_h_r(sp4_h_r_02[47:0]), .sp12_v_t(net1099[0:23]),
     .sp4_v_t(sp4_v_b_03[47:0]), .sp4_r_v_b(sp4_r_v_b_02[47:0]),
     .wl(wl[31:16]), .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net1122), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));
ltile4_ice1f I_LT08 ( .cntl_cbit(net0755[0:7]), .op_bot(net934),
     .op_vic(op_vic), .prog(prog), .carry_out(carry_out),
     .lft_op(lft_op_08[7:0]), .sp12_h_l(sp12_h_l_08[23:0]),
     .sp4_h_l(sp4_h_l_08[47:0]), .sp4_v_b(sp4_v_b_08[47:0]),
     .sp12_v_b(net944[0:23]), .sp12_h_r(sp12_h_r_08[23:0]),
     .sp4_h_r(sp4_h_r_08[47:0]), .sp12_v_t(sp12_v_t_08[23:0]),
     .sp4_v_t(sp4_v_t_08[47:0]), .sp4_r_v_b(sp4_r_v_b_08[47:0]),
     .wl(wl[127:112]), .top_op(top_op_08[7:0]),
     .rgt_op(rgt_op_08[7:0]), .bot_op(slf_op_07[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[127:112]), .vdd_cntl(vdd_cntl[127:112]),
     .glb_netwk(glb_netwk_top[7:0]), .carry_in(net936), .purst(purst),
     .slf_op(slf_op_08[7:0]), .pgate(pgate[127:112]),
     .bnr_op(rgt_op_07[7:0]), .bnl_op(lft_op_07[7:0]),
     .tnr_op(tnr_op_08[7:0]), .tnl_op(tnl_op_08[7:0]));
ltile4_ice1f I_LT07 ( .cntl_cbit(net932[0:7]), .op_bot(net965),
     .op_vic(net934), .prog(prog), .carry_out(net936),
     .lft_op(lft_op_07[7:0]), .sp12_h_l(sp12_h_l_07[23:0]),
     .sp4_h_l(sp4_h_l_07[47:0]), .sp4_v_b(sp4_v_b_07[47:0]),
     .sp12_v_b(net975[0:23]), .sp12_h_r(sp12_h_r_07[23:0]),
     .sp4_h_r(sp4_h_r_07[47:0]), .sp12_v_t(net944[0:23]),
     .sp4_v_t(sp4_v_b_08[47:0]), .sp4_r_v_b(sp4_r_v_b_07[47:0]),
     .wl(wl[111:96]), .top_op(slf_op_08[7:0]), .rgt_op(rgt_op_07[7:0]),
     .bot_op(slf_op_06[7:0]), .bl(bl[53:0]), .reset_b(reset_b[111:96]),
     .vdd_cntl(vdd_cntl[111:96]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net967), .purst(purst), .slf_op(slf_op_07[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_06[7:0]),
     .bnl_op(lft_op_06[7:0]), .tnr_op(rgt_op_08[7:0]),
     .tnl_op(lft_op_08[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_bot (
     .colbuf_cntl(colbuf_cntl_bot[7:0]), .col_clk(glb_netwk_bot[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_top (
     .colbuf_cntl(colbuf_cntl_top[7:0]), .col_clk(glb_netwk_top[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - ice1chip, Cell - quad_br_ice1, View - schematic
// LAST TIME SAVED: May  3 12:05:59 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module quad_br_ice1 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o[7:0],
     bm_sclk_o, bm_sclkrw_o[1:0], bm_sdi_o[1:0], bm_sdo_o[1:0],
     bm_sreb_o, bm_sweb_o[1:0], bm_wdummymux_en_o, bs_en_o,
     carry_out_07_08, carry_out_08_08, carry_out_09_08,
     carry_out_11_08, carry_out_12_08, ceb_o, cf_b_r[143:0],
     cf_r[191:0], fabric_out_07_00, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fabric_out_13_08, hiz_b_o, mode_o, op_vic_07_08,
     op_vic_08_08, op_vic_09_08, op_vic_11_08, op_vic_12_08,
     padeb_b_r[11], padeb_b_r[23:13], padeb_r[12:0], padin_07_00a,
     padin_13_08b, pado_b_r[11], pado_b_r[23:13], pado_r[12:0], r_o,
     sdo, sdo_pad, shift_o, slf_op_07_00[3:0], slf_op_07_01[7:0],
     slf_op_07_02[7:0], slf_op_07_03[7:0], slf_op_07_04[7:0],
     slf_op_07_05[7:0], slf_op_07_06[7:0], slf_op_07_07[7:0],
     slf_op_07_08[7:0], slf_op_08_08[7:0], slf_op_09_08[7:0],
     slf_op_10_08[7:0], slf_op_11_08[7:0], slf_op_12_08[7:0],
     slf_op_13_08[3:0], spi_ss_in_bbank[4:0], tck_pad, tclk_o, tdi_pad,
     tms_pad, update_o, bl[329:0], pgate_r[143:0], reset_b_r[143:0],
     sp4_h_l_07_00[15:0], sp4_h_l_07_01[47:0], sp4_h_l_07_02[47:0],
     sp4_h_l_07_03[47:0], sp4_h_l_07_04[47:0], sp4_h_l_07_05[47:0],
     sp4_h_l_07_06[47:0], sp4_h_l_07_07[47:0], sp4_h_l_07_08[47:0],
     sp4_v_b_07_01[47:0], sp4_v_b_07_02[47:0], sp4_v_b_07_03[47:0],
     sp4_v_b_07_04[47:0], sp4_v_b_07_05[47:0], sp4_v_b_07_06[47:0],
     sp4_v_b_07_07[47:0], sp4_v_b_07_08[47:0], sp4_v_t_07_08[47:0],
     sp4_v_t_08_08[47:0], sp4_v_t_09_08[47:0], sp4_v_t_10_08[47:0],
     sp4_v_t_11_08[47:0], sp4_v_t_12_08[47:0], sp4_v_t_13_08[15:0],
     sp12_h_l_07_01[23:0], sp12_h_l_07_02[23:0], sp12_h_l_07_03[23:0],
     sp12_h_l_07_04[23:0], sp12_h_l_07_05[23:0], sp12_h_l_07_06[23:0],
     sp12_h_l_07_07[23:0], sp12_h_l_07_08[23:0], sp12_v_t_07_08[23:0],
     sp12_v_t_08_08[23:0], sp12_v_t_09_08[23:0], sp12_v_t_10_08[23:0],
     sp12_v_t_11_08[23:0], sp12_v_t_12_08[23:0], vdd_cntl_r[143:0],
     wl_r[143:0], bm_aa_top[10:0], bm_ab_top[10:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i[1:0],
     bm_sdi_i[1:0], bm_sdo_i[1:0], bm_sreb_i, bm_sweb_i[1:0],
     bm_wdummymux_en_i, bnl_op_07_01[3:0], bs_en_i, bs_en_mi, ceb_i,
     ceb_mi, end_of_startup, glb_in[7:0], hiz_b_i, hiz_b_mi, hold_b_r,
     hold_r_b, jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     last_rsr[2], last_rsr[3], lft_op_07_01[7:0], lft_op_07_02[7:0],
     lft_op_07_03[7:0], lft_op_07_04[7:0], lft_op_07_05[7:0],
     lft_op_07_06[7:0], lft_op_07_07[7:0], lft_op_07_08[7:0], md_spi_b,
     mode_i, mode_mi, mux_jtag_sel_b, padin_b_r[11], padin_b_r[23:13],
     padin_r[12:0], pll_sdo, prog, purst, r_i, r_mi, sdi, sdi_pad,
     sdo_enable, shift_i, shift_mi, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk_i, tclk_mi, tnl_op_07_08[7:0], tnl_op_08_08[7:0],
     tnl_op_09_08[7:0], tnl_op_10_08[7:0], tnl_op_11_08[7:0],
     tnl_op_12_08[7:0], tnl_op_13_08[7:0], tnr_op_07_08[7:0],
     tnr_op_08_08[7:0], tnr_op_09_08[7:0], tnr_op_10_08[7:0],
     tnr_op_11_08[7:0], tnr_op_12_08[7:0], top_op_07_08[7:0],
     top_op_08_08[7:0], top_op_09_08[7:0], top_op_10_08[7:0],
     top_op_11_08[7:0], top_op_12_08[7:0], totdopad, trstb_pad,
     update_i, update_mi );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_07_08, carry_out_08_08,
     carry_out_09_08, carry_out_11_08, carry_out_12_08, ceb_o,
     fabric_out_07_00, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fabric_out_13_08, hiz_b_o, mode_o, op_vic_07_08,
     op_vic_08_08, op_vic_09_08, op_vic_11_08, op_vic_12_08,
     padin_07_00a, padin_13_08b, r_o, sdo, sdo_pad, shift_o, tck_pad,
     tclk_o, tdi_pad, tms_pad, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, bs_en_mi, ceb_i, ceb_mi,
     end_of_startup, hiz_b_i, hiz_b_mi, hold_b_r, hold_r_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode_i, mode_mi, mux_jtag_sel_b, pll_sdo, prog, purst, r_i, r_mi,
     sdi, sdi_pad, sdo_enable, shift_i, shift_mi, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk_i, tclk_mi, totdopad, trstb_pad,
     update_i, update_mi;

output [1:0]  bm_sdo_o;
output [7:0]  slf_op_07_04;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_07_08;
output [7:0]  slf_op_07_05;
output [4:0]  spi_ss_in_bbank;
output [7:0]  slf_op_07_03;
output [7:0]  slf_op_12_08;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_07_07;
output [3:0]  slf_op_13_08;
output [143:0]  cf_b_r;
output [7:0]  slf_op_11_08;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_08_08;
output [7:0]  slf_op_07_01;
output [23:11]  padeb_b_r;
output [191:0]  cf_r;
output [12:0]  padeb_r;
output [23:11]  pado_b_r;
output [3:0]  slf_op_07_00;
output [12:0]  pado_r;
output [7:0]  slf_op_07_02;
output [7:0]  slf_op_07_06;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_10_08;
output [7:0]  slf_op_09_08;

inout [47:0]  sp4_v_b_07_06;
inout [47:0]  sp4_v_t_12_08;
inout [23:0]  sp12_v_t_07_08;
inout [47:0]  sp4_h_l_07_07;
inout [47:0]  sp4_h_l_07_03;
inout [23:0]  sp12_v_t_10_08;
inout [47:0]  sp4_v_b_07_08;
inout [23:0]  sp12_h_l_07_08;
inout [23:0]  sp12_h_l_07_01;
inout [15:0]  sp4_h_l_07_00;
inout [15:0]  sp4_v_t_13_08;
inout [47:0]  sp4_h_l_07_08;
inout [47:0]  sp4_h_l_07_04;
inout [47:0]  sp4_h_l_07_01;
inout [47:0]  sp4_v_b_07_02;
inout [47:0]  sp4_h_l_07_02;
inout [47:0]  sp4_v_t_08_08;
inout [23:0]  sp12_v_t_11_08;
inout [23:0]  sp12_h_l_07_04;
inout [23:0]  sp12_v_t_08_08;
inout [23:0]  sp12_h_l_07_06;
inout [47:0]  sp4_v_t_09_08;
inout [23:0]  sp12_v_t_12_08;
inout [47:0]  sp4_h_l_07_05;
inout [47:0]  sp4_v_b_07_04;
inout [23:0]  sp12_h_l_07_05;
inout [47:0]  sp4_v_b_07_03;
inout [47:0]  sp4_v_t_11_08;
inout [47:0]  sp4_v_t_07_08;
inout [47:0]  sp4_h_l_07_06;
inout [47:0]  sp4_v_b_07_05;
inout [143:0]  wl_r;
inout [143:0]  pgate_r;
inout [23:0]  sp12_h_l_07_07;
inout [47:0]  sp4_v_t_10_08;
inout [47:0]  sp4_v_b_07_07;
inout [143:0]  vdd_cntl_r;
inout [329:0]  bl;
inout [23:0]  sp12_h_l_07_02;
inout [47:0]  sp4_v_b_07_01;
inout [23:0]  sp12_v_t_09_08;
inout [23:0]  sp12_h_l_07_03;
inout [143:0]  reset_b_r;

input [1:0]  bm_sweb_i;
input [7:0]  tnr_op_08_08;
input [7:0]  lft_op_07_03;
input [7:0]  top_op_11_08;
input [7:0]  lft_op_07_07;
input [7:0]  lft_op_07_01;
input [7:0]  glb_in;
input [7:0]  top_op_10_08;
input [23:11]  padin_b_r;
input [7:0]  tnl_op_11_08;
input [7:0]  lft_op_07_08;
input [7:0]  tnr_op_12_08;
input [7:0]  tnl_op_13_08;
input [7:0]  lft_op_07_02;
input [1:0]  bm_sclkrw_i;
input [2:3]  last_rsr;
input [10:0]  bm_aa_top;
input [1:0]  bm_sdi_i;
input [7:0]  tnl_op_08_08;
input [7:0]  tnr_op_09_08;
input [7:0]  tnl_op_07_08;
input [7:0]  top_op_09_08;
input [7:0]  lft_op_07_04;
input [3:0]  bnl_op_07_01;
input [12:0]  padin_r;
input [7:0]  top_op_07_08;
input [7:0]  top_op_08_08;
input [7:0]  lft_op_07_05;
input [7:0]  tnl_op_10_08;
input [1:0]  bm_sdo_i;
input [10:0]  bm_ab_top;
input [7:0]  top_op_12_08;
input [7:0]  tnl_op_12_08;
input [7:0]  tnl_op_09_08;
input [7:0]  tnr_op_07_08;
input [7:0]  lft_op_07_06;
input [7:0]  bm_sa_i;
input [7:0]  tnr_op_11_08;
input [7:0]  tnr_op_10_08;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:47]  net1288;

wire  [0:47]  net1383;

wire  [0:47]  net1484;

wire  [0:23]  net1478;

wire  [0:23]  net1509;

wire  [0:47]  net1192;

wire  [0:7]  net1389;

wire  [0:47]  net907;

wire  [0:23]  net1212;

wire  [0:7]  net784;

wire  [0:7]  net913;

wire  [0:47]  net1119;

wire  [0:23]  net901;

wire  [0:47]  net976;

wire  [0:47]  net1169;

wire  [0:47]  net1264;

wire  [0:23]  net1305;

wire  [0:47]  net1492;

wire  [0:23]  net1464;

wire  [0:23]  net911;

wire  [0:23]  net1210;

wire  [0:7]  net1104;

wire  [0:23]  net1209;

wire  [0:23]  net1480;

wire  [0:47]  net980;

wire  [0:47]  net979;

wire  [0:47]  net1551;

wire  [0:23]  net1500;

wire  [0:47]  net1309;

wire  [0:47]  net1000;

wire  [0:47]  net1310;

wire  [0:23]  net1402;

wire  [0:47]  net1360;

wire  [0:47]  net1550;

wire  [0:7]  net1390;

wire  [0:47]  net1262;

wire  [0:23]  net1020;

wire  [0:7]  net936;

wire  [0:23]  net894;

wire  [0:7]  net1045;

wire  [0:47]  net1261;

wire  [0:47]  net889;

wire  [0:23]  net1022;

wire  [0:23]  net1400;

wire  [0:47]  net1382;

wire  [0:23]  net1114;

wire  [0:47]  net1095;

wire  [0:47]  net1003;

wire  [7:0]  clk_center;

wire  [3:0]  slf_op_13_04;

wire  [3:0]  slf_op_12_00;

wire  [0:47]  net1266;

wire  [0:47]  net1076;

wire  [3:0]  slf_op_13_01;

wire  [3:0]  slf_op_13_03;

wire  [0:7]  net1340;

wire  [0:23]  net1257;

wire  [3:0]  slf_op_13_05;

wire  [3:0]  slf_op_08_00;

wire  [0:23]  net1255;

wire  [0:7]  net934;

wire  [0:7]  net1200;

wire  [3:0]  slf_op_13_06;

wire  [0:23]  net1211;

wire  [0:23]  net1019;

wire  [0:47]  net1495;

wire  [0:23]  net1352;

wire  [0:7]  net910;

wire  [0:47]  net1286;

wire  [0:47]  net1171;

wire  [0:47]  net1071;

wire  [0:10]  net792;

wire  [0:7]  net1105;

wire  [0:7]  net1047;

wire  [0:7]  net01436;

wire  [0:47]  net916;

wire  [0:23]  net1350;

wire  [0:7]  net1199;

wire  [3:0]  slf_op_11_00;

wire  [0:23]  net1306;

wire  [0:47]  net1098;

wire  [0:7]  net1531;

wire  [0:47]  net1191;

wire  [0:47]  net1287;

wire  [0:23]  net1476;

wire  [0:47]  net802;

wire  [0:23]  net1021;

wire  [0:47]  net1096;

wire  [0:7]  net1142;

wire  [0:23]  net1508;

wire  [0:47]  net1193;

wire  [0:47]  net1025;

wire  [0:47]  net805;

wire  [0:23]  net1115;

wire  [0:23]  net1160;

wire  [0:47]  net1122;

wire  [0:47]  net1312;

wire  [0:47]  net977;

wire  [0:47]  net1167;

wire  [0:15]  net948;

wire  [0:47]  net1121;

wire  [0:47]  net1380;

wire  [0:47]  net1120;

wire  [0:47]  net1555;

wire  [3:0]  slf_op_09_00;

wire  [0:23]  net970;

wire  [0:23]  net1162;

wire  [0:23]  net1256;

wire  [0:47]  net1405;

wire  [0:23]  net1399;

wire  [0:47]  net1406;

wire  [0:23]  net903;

wire  [0:7]  net1245;

wire  [0:47]  net1267;

wire  [0:7]  net1529;

wire  [0:23]  net1066;

wire  [0:47]  net1166;

wire  [0:47]  net1072;

wire  [0:7]  net938;

wire  [0:7]  net1106;

wire  [0:23]  net1304;

wire  [0:47]  net1554;

wire  [0:47]  net1214;

wire  [0:47]  net982;

wire  [0:7]  net935;

wire  [0:47]  net1001;

wire  [0:23]  net971;

wire  [0:7]  net1295;

wire  [0:23]  net1067;

wire  [0:47]  net1381;

wire  [0:47]  net1404;

wire  [0:23]  net1064;

wire  [0:7]  net937;

wire  [0:23]  net1117;

wire  [0:47]  net1525;

wire  [0:47]  net1260;

wire  [0:47]  net1172;

wire  [0:7]  net1055;

wire  [0:47]  net1524;

wire  [0:7]  net1391;

wire  [0:47]  net1488;

wire  [0:7]  net1530;

wire  [0:47]  net1027;

wire  [0:7]  net939;

wire  [0:23]  net1254;

wire  [0:47]  net1361;

wire  [0:7]  net1528;

wire  [0:47]  net1362;

wire  [0:47]  net1491;

wire  [0:23]  net1159;

wire  [0:7]  net782;

wire  [0:7]  net1533;

wire  [0:7]  net1532;

wire  [0:10]  net791;

wire  [0:7]  net1237;

wire  [0:47]  net1002;

wire  [0:47]  net1506;

wire  [0:47]  net1215;

wire  [0:47]  net1216;

wire  [0:47]  net1311;

wire  [0:47]  net1285;

wire  [0:47]  net1355;

wire  [7:0]  clk_tree_drv_br;

wire  [0:23]  net1065;

wire  [0:47]  net1190;

wire  [0:23]  net972;

wire  [0:47]  net1407;

wire  [3:0]  slf_op_13_07;

wire  [3:0]  slf_op_10_00;

wire  [0:23]  net1161;

wire  [0:47]  net800;

wire  [0:7]  net1296;

wire  [11:11]  padinlat_b_r;

wire  [0:23]  net899;

wire  [0:23]  net969;

wire  [0:47]  net1359;

wire  [0:7]  net1235;

wire  [0:47]  net1170;

wire  [0:7]  net1150;

wire  [0:7]  net1332;

wire  [0:23]  net898;

wire  [0:23]  net1401;

wire  [0:47]  net1553;

wire  [0:47]  net1077;

wire  [0:47]  net1075;

wire  [0:7]  net1330;

wire  [0:23]  net1351;

wire  [0:47]  net1168;

wire  [0:47]  net799;

wire  [0:23]  net1116;

wire  [0:47]  net1357;

wire  [0:7]  net1294;

wire  [0:47]  net896;

wire  [0:47]  net1070;

wire  [0:47]  net1165;

wire  [0:23]  net1307;

wire  [0:23]  net1349;

wire  [0:47]  net1552;

wire  [0:47]  net1356;

wire  [0:47]  net1265;

wire  [0:47]  net981;

wire  [0:23]  net1481;

wire  [0:7]  net793;

wire  [0:47]  net1523;

wire  [0:47]  net1097;

wire  [0:7]  net1140;

wire  [3:0]  slf_op_13_02;

wire  [0:47]  net1217;

wire  [0:7]  net1201;

wire  [0:47]  net1074;



bram1x4_ice1f I_bram_col_b10 ( .glb_netwk_top(net01436[0:7]),
     .prog(prog), .glb_netwk_col(clk_tree_drv_br[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .reset_b(reset_b_r[143:16]),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sreb_o(bm_sreb_o),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .lft_op_05(net1296[0:7]), .bl(bl[203:162]),
     .sp4_h_l_06(net1097[0:47]), .sp12_h_l_02(net1066[0:23]),
     .lft_op_06(net1295[0:7]), .sp12_h_l_03(net1065[0:23]),
     .sp12_h_r_03(net1464[0:23]), .sp12_h_l_01(net1067[0:23]),
     .sp4_v_b_04(net1070[0:47]), .sp4_v_b_05(net1119[0:47]),
     .lft_op_07(net1294[0:7]), .sp4_v_b_06(net1120[0:47]),
     .sp4_v_b_08(net1122[0:47]), .sp4_v_b_07(net1121[0:47]),
     .lft_op_03(net1235[0:7]), .lft_op_01(net910[0:7]),
     .sp4_h_l_02(net1076[0:47]), .sp12_h_l_06(net1115[0:23]),
     .sp12_h_r_07(net1476[0:23]), .sp12_h_l_05(net1114[0:23]),
     .sp12_h_r_06(net1478[0:23]), .sp12_h_l_04(net1064[0:23]),
     .sp12_h_r_05(net1480[0:23]), .sp12_h_r_08(net1481[0:23]),
     .sp12_h_l_07(net1116[0:23]), .sp12_h_l_08(net1117[0:23]),
     .sp4_r_v_b_03(net1484[0:47]), .vdd_cntl(vdd_cntl_r[143:16]),
     .pgate(pgate_r[143:16]), .bot_op_01({slf_op_10_00[3],
     slf_op_10_00[2], slf_op_10_00[1], slf_op_10_00[0],
     slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0]}), .sp4_r_v_b_04(net1488[0:47]),
     .sp4_v_b_01(net907[0:47]), .sp4_v_b_03(net1071[0:47]),
     .sp4_h_r_08(net1491[0:47]), .sp4_r_v_b_05(net1492[0:47]),
     .sp4_v_b_02(net1072[0:47]), .sp4_v_t_08(sp4_v_t_10_08[47:0]),
     .sp4_r_v_b_02(net1495[0:47]), .bnr_op_01({slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0],
     slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0]}), .bm_sdi_o(bm_sdi_o[1:0]),
     .sp4_h_l_04(net1074[0:47]), .lft_op_08(slf_op_09_08[7:0]),
     .sp12_h_r_01(net1500[0:23]), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .sp4_h_l_03(net1075[0:47]), .sp4_h_l_01(net1077[0:47]),
     .sp4_h_r_01(net1506[0:47]), .tnr_op_08(tnr_op_10_08[7:0]),
     .sp12_h_r_02(net1508[0:23]), .sp12_h_r_04(net1509[0:23]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .lft_op_02(net1237[0:7]), .lft_op_04(net1245[0:7]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bnl_op_01({slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0],
     slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0]}), .sp12_v_t_08(sp12_v_t_10_08[23:0]),
     .wl(wl_r[143:16]), .tnl_op_08(tnl_op_10_08[7:0]),
     .top_op_08(top_op_10_08[7:0]), .bm_ab_2bot(net792[0:10]),
     .bm_aa_2bot(net791[0:10]), .sp12_v_b_01(net899[0:23]),
     .sp4_r_v_b_08(net1523[0:47]), .sp4_r_v_b_07(net1524[0:47]),
     .sp4_r_v_b_06(net1525[0:47]), .sp4_r_v_b_01(net896[0:47]),
     .rgt_op_08(slf_op_11_08[7:0]), .rgt_op_07(net1528[0:7]),
     .rgt_op_06(net1529[0:7]), .rgt_op_05(net1530[0:7]),
     .rgt_op_04(net1531[0:7]), .rgt_op_03(net1532[0:7]),
     .rgt_op_02(net1533[0:7]), .rgt_op_01(net782[0:7]),
     .slf_op_02(net1047[0:7]), .slf_op_01(net784[0:7]),
     .slf_op_03(net1045[0:7]), .slf_op_04(net1055[0:7]),
     .slf_op_05(net1106[0:7]), .slf_op_06(net1105[0:7]),
     .slf_op_07(net1104[0:7]), .slf_op_08(slf_op_10_08[7:0]),
     .bm_ab_top(bm_ab_top[10:0]), .bm_aa_top(bm_aa_top[10:0]),
     .glb_netwk_bot(net936[0:7]), .sp4_h_l_08(net1095[0:47]),
     .sp4_h_l_07(net1096[0:47]), .sp4_h_l_05(net1098[0:47]),
     .sp4_h_r_02(net1550[0:47]), .sp4_h_r_03(net1551[0:47]),
     .sp4_h_r_04(net1552[0:47]), .sp4_h_r_05(net1553[0:47]),
     .sp4_h_r_06(net1554[0:47]), .sp4_h_r_07(net1555[0:47]));
pinlatbuf12p_1 I484 ( .pad_in(padin_r[12]), .icegate(hold_r_b),
     .cbit(cf_r[183]), .cout(net0731), .prog(prog));
pinlatbuf12p_1 I486 ( .pad_in(padin_b_r[11]), .icegate(hold_b_r),
     .cbit(cf_b_r[15]), .cout(padinlat_b_r[11]), .prog(prog));
tielo I369 ( .tielo(tgnd_br_q));
scan_buf_ice8p I_scanbuf_8p_br ( .update_i(update_mi),
     .tclk_i(tclk_mi), .shift_i(shift_mi), .sdi(sdi_pad), .r_i(r_mi),
     .mode_i(mode_mi), .hiz_b_i(hiz_b_mi), .ceb_i(ceb_mi),
     .bs_en_i(bs_en_mi), .update_o(update_o), .tclk_o(net774),
     .shift_o(shift_o), .sdo(net776), .r_o(r_o), .mode_o(mode_o),
     .hiz_b_o(hiz_b_o), .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_rgt_bot_1x8_ice1f I_preio_rgt_b ( cf_r[191:0], net808, net807,
     net809, padeb_r[12:0], pado_r[12:0], sdo, slf_op_13_01[3:0],
     slf_op_13_02[3:0], slf_op_13_03[3:0], slf_op_13_04[3:0],
     slf_op_13_05[3:0], slf_op_13_06[3:0], slf_op_13_07[3:0],
     slf_op_13_08[3:0], tck_pad, tclk_o, tdi_pad, tms_pad,
     net982[0:47], net981[0:47], net980[0:47], net979[0:47],
     net1003[0:47], net1002[0:47], net1001[0:47], net1000[0:47],
     net972[0:23], net971[0:23], net970[0:23], net969[0:23],
     net1019[0:23], net1020[0:23], net1021[0:23], net1022[0:23],
     bl[329:312], pgate_r[143:16], reset_b_r[143:16], net948[0:15],
     sp4_v_t_13_08[15:0], vdd_cntl_r[143:16], wl_r[143:16],
     {slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0], slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0]}, bs_en_o, ceb_o,
     clk_tree_drv_br[7:0], hiz_b_o, hold_r_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[2],
     last_rsr[3], net913[0:7], net1142[0:7], net1140[0:7],
     net1150[0:7], net1201[0:7], net1200[0:7], net1199[0:7],
     slf_op_12_08[7:0], mode_o, mux_jtag_sel_b, padin_r[12:0], prog,
     r_o, net776, sdo_enable, shift_o, net774, tnl_op_13_08[7:0],
     totdopad, trstb_pad, update_o);
io_bot_rgt_1x6_ice1f I_preio_bot_r ( cf_b_r[143:0], net1437, net912,
     padeb_b_r[11], padeb_b_r[23:13], pado_b_r[11], pado_b_r[23:13],
     sdo_pad, slf_op_07_00[3:0], slf_op_08_00[3:0], slf_op_09_00[3:0],
     slf_op_10_00[3:0], slf_op_11_00[3:0], slf_op_12_00[3:0],
     spi_ss_in_bbank[4:0], bl[53:0], bl[107:54], bl[161:108],
     bl[203:162], bl[257:204], bl[311:258], sp4_h_l_07_00[15:0],
     net948[0:15], sp4_v_b_07_01[47:0], net889[0:47], net916[0:47],
     net907[0:47], net896[0:47], net1168[0:47], net903[0:23],
     net901[0:23], net911[0:23], net899[0:23], net894[0:23],
     net898[0:23], lft_op_07_01[7:0], bs_en_i, ceb_i, end_of_startup,
     net939[0:7], net938[0:7], net937[0:7], net936[0:7], net935[0:7],
     net934[0:7], hiz_b_i, hold_b_r, slf_op_07_01[7:0], net793[0:7],
     net910[0:7], net784[0:7], net782[0:7], net913[0:7], md_spi_b,
     mode_i, padin_b_r[11], padin_b_r[23:13], {pgate_r[1], pgate_r[0],
     pgate_r[2], pgate_r[3], pgate_r[5], pgate_r[4], pgate_r[6],
     pgate_r[7], pgate_r[9], pgate_r[8], pgate_r[10], pgate_r[11],
     pgate_r[13], pgate_r[12], pgate_r[14], pgate_r[15]}, prog, r_i,
     {reset_b_r[1], reset_b_r[0], reset_b_r[2], reset_b_r[3],
     reset_b_r[5], reset_b_r[4], reset_b_r[6], reset_b_r[7],
     reset_b_r[9], reset_b_r[8], reset_b_r[10], reset_b_r[11],
     reset_b_r[13], reset_b_r[12], reset_b_r[14], reset_b_r[15]}, sdi,
     shift_i, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out, tclk_i,
     {slf_op_13_01[3], slf_op_13_01[2], slf_op_13_01[1],
     slf_op_13_01[0], slf_op_13_01[3], slf_op_13_01[2],
     slf_op_13_01[1], slf_op_13_01[0]}, update_i, {vdd_cntl_r[1],
     vdd_cntl_r[0], vdd_cntl_r[2], vdd_cntl_r[3], vdd_cntl_r[5],
     vdd_cntl_r[4], vdd_cntl_r[6], vdd_cntl_r[7], vdd_cntl_r[9],
     vdd_cntl_r[8], vdd_cntl_r[10], vdd_cntl_r[11], vdd_cntl_r[13],
     vdd_cntl_r[12], vdd_cntl_r[14], vdd_cntl_r[15]}, {wl_r[1],
     wl_r[0], wl_r[2], wl_r[3], wl_r[5], wl_r[4], wl_r[6], wl_r[7],
     wl_r[9], wl_r[8], wl_r[10], wl_r[11], wl_r[13], wl_r[12],
     wl_r[14], wl_r[15]});
lt_1x8_bot_ice1f I_lt_col_b12 ( .glb_netwk_bot(net934[0:7]),
     .rgt_op_03({slf_op_13_03[3], slf_op_13_03[2], slf_op_13_03[1],
     slf_op_13_03[0], slf_op_13_03[3], slf_op_13_03[2],
     slf_op_13_03[1], slf_op_13_03[0]}), .slf_op_02(net1142[0:7]),
     .rgt_op_02({slf_op_13_02[3], slf_op_13_02[2], slf_op_13_02[1],
     slf_op_13_02[0], slf_op_13_02[3], slf_op_13_02[2],
     slf_op_13_02[1], slf_op_13_02[0]}), .rgt_op_01({slf_op_13_01[3],
     slf_op_13_01[2], slf_op_13_01[1], slf_op_13_01[0],
     slf_op_13_01[3], slf_op_13_01[2], slf_op_13_01[1],
     slf_op_13_01[0]}), .purst(purst), .prog(prog),
     .lft_op_04(net1531[0:7]), .lft_op_03(net1532[0:7]),
     .lft_op_02(net1533[0:7]), .lft_op_01(net782[0:7]),
     .rgt_op_04({slf_op_13_04[3], slf_op_13_04[2], slf_op_13_04[1],
     slf_op_13_04[0], slf_op_13_04[3], slf_op_13_04[2],
     slf_op_13_04[1], slf_op_13_04[0]}), .carry_in(tgnd_br_q),
     .bnl_op_01({slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0], slf_op_11_00[3], slf_op_11_00[2],
     slf_op_11_00[1], slf_op_11_00[0]}), .slf_op_04(net1150[0:7]),
     .slf_op_03(net1140[0:7]), .slf_op_01(net913[0:7]),
     .sp4_h_l_04(net1169[0:47]), .carry_out(carry_out_12_08),
     .vdd_cntl(vdd_cntl_r[143:16]), .sp12_h_r_04(net969[0:23]),
     .sp12_h_r_03(net970[0:23]), .sp12_h_r_02(net971[0:23]),
     .sp12_h_r_01(net972[0:23]), .glb_netwk_col(clk_tree_drv_br[7:0]),
     .sp4_v_b_01(net1168[0:47]), .sp4_r_v_b_04(net799[0:47]),
     .sp4_r_v_b_03(net976[0:47]), .sp4_r_v_b_02(net977[0:47]),
     .sp4_r_v_b_01(net805[0:47]), .sp4_h_r_04(net979[0:47]),
     .sp4_h_r_03(net980[0:47]), .sp4_h_r_02(net981[0:47]),
     .sp4_h_r_01(net982[0:47]), .sp4_h_l_03(net1170[0:47]),
     .sp4_h_l_02(net1171[0:47]), .sp4_h_l_01(net1172[0:47]),
     .bl(bl[311:258]), .bot_op_01({slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0], slf_op_12_00[3],
     slf_op_12_00[2], slf_op_12_00[1], slf_op_12_00[0]}),
     .sp12_h_l_01(net1162[0:23]), .sp12_h_l_02(net1161[0:23]),
     .sp12_h_l_03(net1160[0:23]), .sp12_h_l_04(net1159[0:23]),
     .sp4_v_b_04(net1165[0:47]), .sp4_v_b_03(net1166[0:47]),
     .sp4_v_b_02(net1167[0:47]), .bnr_op_01({pll_sdo, pll_sdo, pll_sdo,
     pll_sdo, pll_sdo, pll_sdo, pll_sdo, pll_sdo}),
     .sp4_h_l_05(net1193[0:47]), .sp4_h_l_06(net1192[0:47]),
     .sp4_h_l_07(net1191[0:47]), .sp4_h_l_08(net1190[0:47]),
     .sp4_h_r_08(net1000[0:47]), .sp4_h_r_07(net1001[0:47]),
     .sp4_h_r_06(net1002[0:47]), .sp4_h_r_05(net1003[0:47]),
     .slf_op_05(net1201[0:7]), .slf_op_06(net1200[0:7]),
     .slf_op_07(net1199[0:7]), .slf_op_08(slf_op_12_08[7:0]),
     .rgt_op_08({slf_op_13_08[3], slf_op_13_08[2], slf_op_13_08[1],
     slf_op_13_08[0], slf_op_13_08[3], slf_op_13_08[2],
     slf_op_13_08[1], slf_op_13_08[0]}), .rgt_op_07({slf_op_13_07[3],
     slf_op_13_07[2], slf_op_13_07[1], slf_op_13_07[0],
     slf_op_13_07[3], slf_op_13_07[2], slf_op_13_07[1],
     slf_op_13_07[0]}), .rgt_op_06({slf_op_13_06[3], slf_op_13_06[2],
     slf_op_13_06[1], slf_op_13_06[0], slf_op_13_06[3],
     slf_op_13_06[2], slf_op_13_06[1], slf_op_13_06[0]}),
     .rgt_op_05({slf_op_13_05[3], slf_op_13_05[2], slf_op_13_05[1],
     slf_op_13_05[0], slf_op_13_05[3], slf_op_13_05[2],
     slf_op_13_05[1], slf_op_13_05[0]}), .lft_op_08(slf_op_11_08[7:0]),
     .lft_op_07(net1528[0:7]), .lft_op_06(net1529[0:7]),
     .lft_op_05(net1530[0:7]), .sp12_h_l_08(net1212[0:23]),
     .sp12_h_l_07(net1211[0:23]), .sp12_h_l_06(net1210[0:23]),
     .sp12_h_r_05(net1019[0:23]), .sp12_h_r_06(net1020[0:23]),
     .sp12_h_r_07(net1021[0:23]), .sp12_h_r_08(net1022[0:23]),
     .sp12_h_l_05(net1209[0:23]), .sp4_r_v_b_05(net802[0:47]),
     .sp4_r_v_b_06(net1025[0:47]), .sp4_r_v_b_07(net800[0:47]),
     .sp4_r_v_b_08(net1027[0:47]), .sp4_v_b_08(net1217[0:47]),
     .sp4_v_b_07(net1216[0:47]), .sp4_v_b_06(net1215[0:47]),
     .sp4_v_b_05(net1214[0:47]), .pgate(pgate_r[143:16]),
     .reset_b(reset_b_r[143:16]), .wl(wl_r[143:16]),
     .sp12_v_t_08(sp12_v_t_12_08[23:0]), .tnr_op_08(tnr_op_12_08[7:0]),
     .top_op_08(top_op_12_08[7:0]), .tnl_op_08(tnl_op_12_08[7:0]),
     .sp4_v_t_08(sp4_v_t_12_08[47:0]), .lc_bot(tgnd_br_q),
     .op_vic(op_vic_12_08), .sp12_v_b_01(net898[0:23]));
lt_1x8_bot_ice1f I_lt_col_b09 ( .glb_netwk_bot(net937[0:7]),
     .rgt_op_03(net1045[0:7]), .slf_op_02(net1237[0:7]),
     .rgt_op_02(net1047[0:7]), .rgt_op_01(net784[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net1340[0:7]), .lft_op_03(net1330[0:7]),
     .lft_op_02(net1332[0:7]), .lft_op_01(net793[0:7]),
     .rgt_op_04(net1055[0:7]), .carry_in(tgnd_br_q),
     .bnl_op_01({slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0], slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0]}), .slf_op_04(net1245[0:7]),
     .slf_op_03(net1235[0:7]), .slf_op_01(net910[0:7]),
     .sp4_h_l_04(net1264[0:47]), .carry_out(carry_out_09_08),
     .vdd_cntl(vdd_cntl_r[143:16]), .sp12_h_r_04(net1064[0:23]),
     .sp12_h_r_03(net1065[0:23]), .sp12_h_r_02(net1066[0:23]),
     .sp12_h_r_01(net1067[0:23]), .glb_netwk_col(clk_tree_drv_br[7:0]),
     .sp4_v_b_01(net916[0:47]), .sp4_r_v_b_04(net1070[0:47]),
     .sp4_r_v_b_03(net1071[0:47]), .sp4_r_v_b_02(net1072[0:47]),
     .sp4_r_v_b_01(net907[0:47]), .sp4_h_r_04(net1074[0:47]),
     .sp4_h_r_03(net1075[0:47]), .sp4_h_r_02(net1076[0:47]),
     .sp4_h_r_01(net1077[0:47]), .sp4_h_l_03(net1265[0:47]),
     .sp4_h_l_02(net1266[0:47]), .sp4_h_l_01(net1267[0:47]),
     .bl(bl[161:108]), .bot_op_01({slf_op_09_00[3], slf_op_09_00[2],
     slf_op_09_00[1], slf_op_09_00[0], slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0]}),
     .sp12_h_l_01(net1257[0:23]), .sp12_h_l_02(net1256[0:23]),
     .sp12_h_l_03(net1255[0:23]), .sp12_h_l_04(net1254[0:23]),
     .sp4_v_b_04(net1260[0:47]), .sp4_v_b_03(net1261[0:47]),
     .sp4_v_b_02(net1262[0:47]), .bnr_op_01({slf_op_10_00[3],
     slf_op_10_00[2], slf_op_10_00[1], slf_op_10_00[0],
     slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0]}), .sp4_h_l_05(net1288[0:47]),
     .sp4_h_l_06(net1287[0:47]), .sp4_h_l_07(net1286[0:47]),
     .sp4_h_l_08(net1285[0:47]), .sp4_h_r_08(net1095[0:47]),
     .sp4_h_r_07(net1096[0:47]), .sp4_h_r_06(net1097[0:47]),
     .sp4_h_r_05(net1098[0:47]), .slf_op_05(net1296[0:7]),
     .slf_op_06(net1295[0:7]), .slf_op_07(net1294[0:7]),
     .slf_op_08(slf_op_09_08[7:0]), .rgt_op_08(slf_op_10_08[7:0]),
     .rgt_op_07(net1104[0:7]), .rgt_op_06(net1105[0:7]),
     .rgt_op_05(net1106[0:7]), .lft_op_08(slf_op_08_08[7:0]),
     .lft_op_07(net1389[0:7]), .lft_op_06(net1390[0:7]),
     .lft_op_05(net1391[0:7]), .sp12_h_l_08(net1307[0:23]),
     .sp12_h_l_07(net1306[0:23]), .sp12_h_l_06(net1305[0:23]),
     .sp12_h_r_05(net1114[0:23]), .sp12_h_r_06(net1115[0:23]),
     .sp12_h_r_07(net1116[0:23]), .sp12_h_r_08(net1117[0:23]),
     .sp12_h_l_05(net1304[0:23]), .sp4_r_v_b_05(net1119[0:47]),
     .sp4_r_v_b_06(net1120[0:47]), .sp4_r_v_b_07(net1121[0:47]),
     .sp4_r_v_b_08(net1122[0:47]), .sp4_v_b_08(net1312[0:47]),
     .sp4_v_b_07(net1311[0:47]), .sp4_v_b_06(net1310[0:47]),
     .sp4_v_b_05(net1309[0:47]), .pgate(pgate_r[143:16]),
     .reset_b(reset_b_r[143:16]), .wl(wl_r[143:16]),
     .sp12_v_t_08(sp12_v_t_09_08[23:0]), .tnr_op_08(tnr_op_09_08[7:0]),
     .top_op_08(top_op_09_08[7:0]), .tnl_op_08(tnl_op_09_08[7:0]),
     .sp4_v_t_08(sp4_v_t_09_08[47:0]), .lc_bot(tgnd_br_q),
     .op_vic(op_vic_09_08), .sp12_v_b_01(net911[0:23]));
lt_1x8_bot_ice1f I_lt_col_b11 ( .glb_netwk_bot(net935[0:7]),
     .rgt_op_03(net1140[0:7]), .slf_op_02(net1533[0:7]),
     .rgt_op_02(net1142[0:7]), .rgt_op_01(net913[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net1055[0:7]), .lft_op_03(net1045[0:7]),
     .lft_op_02(net1047[0:7]), .lft_op_01(net784[0:7]),
     .rgt_op_04(net1150[0:7]), .carry_in(tgnd_br_q),
     .bnl_op_01({slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0], slf_op_10_00[3], slf_op_10_00[2],
     slf_op_10_00[1], slf_op_10_00[0]}), .slf_op_04(net1531[0:7]),
     .slf_op_03(net1532[0:7]), .slf_op_01(net782[0:7]),
     .sp4_h_l_04(net1552[0:47]), .carry_out(carry_out_11_08),
     .vdd_cntl(vdd_cntl_r[143:16]), .sp12_h_r_04(net1159[0:23]),
     .sp12_h_r_03(net1160[0:23]), .sp12_h_r_02(net1161[0:23]),
     .sp12_h_r_01(net1162[0:23]), .glb_netwk_col(clk_tree_drv_br[7:0]),
     .sp4_v_b_01(net896[0:47]), .sp4_r_v_b_04(net1165[0:47]),
     .sp4_r_v_b_03(net1166[0:47]), .sp4_r_v_b_02(net1167[0:47]),
     .sp4_r_v_b_01(net1168[0:47]), .sp4_h_r_04(net1169[0:47]),
     .sp4_h_r_03(net1170[0:47]), .sp4_h_r_02(net1171[0:47]),
     .sp4_h_r_01(net1172[0:47]), .sp4_h_l_03(net1551[0:47]),
     .sp4_h_l_02(net1550[0:47]), .sp4_h_l_01(net1506[0:47]),
     .bl(bl[257:204]), .bot_op_01({slf_op_11_00[3], slf_op_11_00[2],
     slf_op_11_00[1], slf_op_11_00[0], slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0]}),
     .sp12_h_l_01(net1500[0:23]), .sp12_h_l_02(net1508[0:23]),
     .sp12_h_l_03(net1464[0:23]), .sp12_h_l_04(net1509[0:23]),
     .sp4_v_b_04(net1488[0:47]), .sp4_v_b_03(net1484[0:47]),
     .sp4_v_b_02(net1495[0:47]), .bnr_op_01({slf_op_12_00[3],
     slf_op_12_00[2], slf_op_12_00[1], slf_op_12_00[0],
     slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0]}), .sp4_h_l_05(net1553[0:47]),
     .sp4_h_l_06(net1554[0:47]), .sp4_h_l_07(net1555[0:47]),
     .sp4_h_l_08(net1491[0:47]), .sp4_h_r_08(net1190[0:47]),
     .sp4_h_r_07(net1191[0:47]), .sp4_h_r_06(net1192[0:47]),
     .sp4_h_r_05(net1193[0:47]), .slf_op_05(net1530[0:7]),
     .slf_op_06(net1529[0:7]), .slf_op_07(net1528[0:7]),
     .slf_op_08(slf_op_11_08[7:0]), .rgt_op_08(slf_op_12_08[7:0]),
     .rgt_op_07(net1199[0:7]), .rgt_op_06(net1200[0:7]),
     .rgt_op_05(net1201[0:7]), .lft_op_08(slf_op_10_08[7:0]),
     .lft_op_07(net1104[0:7]), .lft_op_06(net1105[0:7]),
     .lft_op_05(net1106[0:7]), .sp12_h_l_08(net1481[0:23]),
     .sp12_h_l_07(net1476[0:23]), .sp12_h_l_06(net1478[0:23]),
     .sp12_h_r_05(net1209[0:23]), .sp12_h_r_06(net1210[0:23]),
     .sp12_h_r_07(net1211[0:23]), .sp12_h_r_08(net1212[0:23]),
     .sp12_h_l_05(net1480[0:23]), .sp4_r_v_b_05(net1214[0:47]),
     .sp4_r_v_b_06(net1215[0:47]), .sp4_r_v_b_07(net1216[0:47]),
     .sp4_r_v_b_08(net1217[0:47]), .sp4_v_b_08(net1523[0:47]),
     .sp4_v_b_07(net1524[0:47]), .sp4_v_b_06(net1525[0:47]),
     .sp4_v_b_05(net1492[0:47]), .pgate(pgate_r[143:16]),
     .reset_b(reset_b_r[143:16]), .wl(wl_r[143:16]),
     .sp12_v_t_08(sp12_v_t_11_08[23:0]), .tnr_op_08(tnr_op_11_08[7:0]),
     .top_op_08(top_op_11_08[7:0]), .tnl_op_08(tnl_op_11_08[7:0]),
     .sp4_v_t_08(sp4_v_t_11_08[47:0]), .lc_bot(tgnd_br_q),
     .op_vic(op_vic_11_08), .sp12_v_b_01(net894[0:23]));
lt_1x8_bot_ice1f I_lt_col_b08 ( .glb_netwk_bot(net938[0:7]),
     .rgt_op_03(net1235[0:7]), .slf_op_02(net1332[0:7]),
     .rgt_op_02(net1237[0:7]), .rgt_op_01(net910[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(slf_op_07_04[7:0]),
     .lft_op_03(slf_op_07_03[7:0]), .lft_op_02(slf_op_07_02[7:0]),
     .lft_op_01(slf_op_07_01[7:0]), .rgt_op_04(net1245[0:7]),
     .carry_in(tgnd_br_q), .bnl_op_01({slf_op_07_00[3],
     slf_op_07_00[2], slf_op_07_00[1], slf_op_07_00[0],
     slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0]}), .slf_op_04(net1340[0:7]),
     .slf_op_03(net1330[0:7]), .slf_op_01(net793[0:7]),
     .sp4_h_l_04(net1359[0:47]), .carry_out(carry_out_08_08),
     .vdd_cntl(vdd_cntl_r[143:16]), .sp12_h_r_04(net1254[0:23]),
     .sp12_h_r_03(net1255[0:23]), .sp12_h_r_02(net1256[0:23]),
     .sp12_h_r_01(net1257[0:23]), .glb_netwk_col(clk_tree_drv_br[7:0]),
     .sp4_v_b_01(net889[0:47]), .sp4_r_v_b_04(net1260[0:47]),
     .sp4_r_v_b_03(net1261[0:47]), .sp4_r_v_b_02(net1262[0:47]),
     .sp4_r_v_b_01(net916[0:47]), .sp4_h_r_04(net1264[0:47]),
     .sp4_h_r_03(net1265[0:47]), .sp4_h_r_02(net1266[0:47]),
     .sp4_h_r_01(net1267[0:47]), .sp4_h_l_03(net1360[0:47]),
     .sp4_h_l_02(net1361[0:47]), .sp4_h_l_01(net1362[0:47]),
     .bl(bl[107:54]), .bot_op_01({slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0], slf_op_08_00[3],
     slf_op_08_00[2], slf_op_08_00[1], slf_op_08_00[0]}),
     .sp12_h_l_01(net1352[0:23]), .sp12_h_l_02(net1351[0:23]),
     .sp12_h_l_03(net1350[0:23]), .sp12_h_l_04(net1349[0:23]),
     .sp4_v_b_04(net1355[0:47]), .sp4_v_b_03(net1356[0:47]),
     .sp4_v_b_02(net1357[0:47]), .bnr_op_01({slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0],
     slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0]}), .sp4_h_l_05(net1383[0:47]),
     .sp4_h_l_06(net1382[0:47]), .sp4_h_l_07(net1381[0:47]),
     .sp4_h_l_08(net1380[0:47]), .sp4_h_r_08(net1285[0:47]),
     .sp4_h_r_07(net1286[0:47]), .sp4_h_r_06(net1287[0:47]),
     .sp4_h_r_05(net1288[0:47]), .slf_op_05(net1391[0:7]),
     .slf_op_06(net1390[0:7]), .slf_op_07(net1389[0:7]),
     .slf_op_08(slf_op_08_08[7:0]), .rgt_op_08(slf_op_09_08[7:0]),
     .rgt_op_07(net1294[0:7]), .rgt_op_06(net1295[0:7]),
     .rgt_op_05(net1296[0:7]), .lft_op_08(slf_op_07_08[7:0]),
     .lft_op_07(slf_op_07_07[7:0]), .lft_op_06(slf_op_07_06[7:0]),
     .lft_op_05(slf_op_07_05[7:0]), .sp12_h_l_08(net1402[0:23]),
     .sp12_h_l_07(net1401[0:23]), .sp12_h_l_06(net1400[0:23]),
     .sp12_h_r_05(net1304[0:23]), .sp12_h_r_06(net1305[0:23]),
     .sp12_h_r_07(net1306[0:23]), .sp12_h_r_08(net1307[0:23]),
     .sp12_h_l_05(net1399[0:23]), .sp4_r_v_b_05(net1309[0:47]),
     .sp4_r_v_b_06(net1310[0:47]), .sp4_r_v_b_07(net1311[0:47]),
     .sp4_r_v_b_08(net1312[0:47]), .sp4_v_b_08(net1407[0:47]),
     .sp4_v_b_07(net1406[0:47]), .sp4_v_b_06(net1405[0:47]),
     .sp4_v_b_05(net1404[0:47]), .pgate(pgate_r[143:16]),
     .reset_b(reset_b_r[143:16]), .wl(wl_r[143:16]),
     .sp12_v_t_08(sp12_v_t_08_08[23:0]), .tnr_op_08(tnr_op_08_08[7:0]),
     .top_op_08(top_op_08_08[7:0]), .tnl_op_08(tnl_op_08_08[7:0]),
     .sp4_v_t_08(sp4_v_t_08_08[47:0]), .lc_bot(tgnd_br_q),
     .op_vic(op_vic_08_08), .sp12_v_b_01(net901[0:23]));
lt_1x8_bot_ice1f I_lt_col_b07 ( .glb_netwk_bot(net939[0:7]),
     .rgt_op_03(net1330[0:7]), .slf_op_02(slf_op_07_02[7:0]),
     .rgt_op_02(net1332[0:7]), .rgt_op_01(net793[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(lft_op_07_04[7:0]),
     .lft_op_03(lft_op_07_03[7:0]), .lft_op_02(lft_op_07_02[7:0]),
     .lft_op_01(lft_op_07_01[7:0]), .rgt_op_04(net1340[0:7]),
     .carry_in(tgnd_br_q), .bnl_op_01({bnl_op_07_01[3],
     bnl_op_07_01[2], bnl_op_07_01[1], bnl_op_07_01[0],
     bnl_op_07_01[3], bnl_op_07_01[2], bnl_op_07_01[1],
     bnl_op_07_01[0]}), .slf_op_04(slf_op_07_04[7:0]),
     .slf_op_03(slf_op_07_03[7:0]), .slf_op_01(slf_op_07_01[7:0]),
     .sp4_h_l_04(sp4_h_l_07_04[47:0]), .carry_out(carry_out_07_08),
     .vdd_cntl(vdd_cntl_r[143:16]), .sp12_h_r_04(net1349[0:23]),
     .sp12_h_r_03(net1350[0:23]), .sp12_h_r_02(net1351[0:23]),
     .sp12_h_r_01(net1352[0:23]), .glb_netwk_col(clk_tree_drv_br[7:0]),
     .sp4_v_b_01(sp4_v_b_07_01[47:0]), .sp4_r_v_b_04(net1355[0:47]),
     .sp4_r_v_b_03(net1356[0:47]), .sp4_r_v_b_02(net1357[0:47]),
     .sp4_r_v_b_01(net889[0:47]), .sp4_h_r_04(net1359[0:47]),
     .sp4_h_r_03(net1360[0:47]), .sp4_h_r_02(net1361[0:47]),
     .sp4_h_r_01(net1362[0:47]), .sp4_h_l_03(sp4_h_l_07_03[47:0]),
     .sp4_h_l_02(sp4_h_l_07_02[47:0]),
     .sp4_h_l_01(sp4_h_l_07_01[47:0]), .bl(bl[53:0]),
     .bot_op_01({slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0], slf_op_07_00[3], slf_op_07_00[2],
     slf_op_07_00[1], slf_op_07_00[0]}),
     .sp12_h_l_01(sp12_h_l_07_01[23:0]),
     .sp12_h_l_02(sp12_h_l_07_02[23:0]),
     .sp12_h_l_03(sp12_h_l_07_03[23:0]),
     .sp12_h_l_04(sp12_h_l_07_04[23:0]),
     .sp4_v_b_04(sp4_v_b_07_04[47:0]),
     .sp4_v_b_03(sp4_v_b_07_03[47:0]),
     .sp4_v_b_02(sp4_v_b_07_02[47:0]), .bnr_op_01({slf_op_08_00[3],
     slf_op_08_00[2], slf_op_08_00[1], slf_op_08_00[0],
     slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0]}), .sp4_h_l_05(sp4_h_l_07_05[47:0]),
     .sp4_h_l_06(sp4_h_l_07_06[47:0]),
     .sp4_h_l_07(sp4_h_l_07_07[47:0]),
     .sp4_h_l_08(sp4_h_l_07_08[47:0]), .sp4_h_r_08(net1380[0:47]),
     .sp4_h_r_07(net1381[0:47]), .sp4_h_r_06(net1382[0:47]),
     .sp4_h_r_05(net1383[0:47]), .slf_op_05(slf_op_07_05[7:0]),
     .slf_op_06(slf_op_07_06[7:0]), .slf_op_07(slf_op_07_07[7:0]),
     .slf_op_08(slf_op_07_08[7:0]), .rgt_op_08(slf_op_08_08[7:0]),
     .rgt_op_07(net1389[0:7]), .rgt_op_06(net1390[0:7]),
     .rgt_op_05(net1391[0:7]), .lft_op_08(lft_op_07_08[7:0]),
     .lft_op_07(lft_op_07_07[7:0]), .lft_op_06(lft_op_07_06[7:0]),
     .lft_op_05(lft_op_07_05[7:0]), .sp12_h_l_08(sp12_h_l_07_08[23:0]),
     .sp12_h_l_07(sp12_h_l_07_07[23:0]),
     .sp12_h_l_06(sp12_h_l_07_06[23:0]), .sp12_h_r_05(net1399[0:23]),
     .sp12_h_r_06(net1400[0:23]), .sp12_h_r_07(net1401[0:23]),
     .sp12_h_r_08(net1402[0:23]), .sp12_h_l_05(sp12_h_l_07_05[23:0]),
     .sp4_r_v_b_05(net1404[0:47]), .sp4_r_v_b_06(net1405[0:47]),
     .sp4_r_v_b_07(net1406[0:47]), .sp4_r_v_b_08(net1407[0:47]),
     .sp4_v_b_08(sp4_v_b_07_08[47:0]),
     .sp4_v_b_07(sp4_v_b_07_07[47:0]),
     .sp4_v_b_06(sp4_v_b_07_06[47:0]),
     .sp4_v_b_05(sp4_v_b_07_05[47:0]), .pgate(pgate_r[143:16]),
     .reset_b(reset_b_r[143:16]), .wl(wl_r[143:16]),
     .sp12_v_t_08(sp12_v_t_07_08[23:0]), .tnr_op_08(tnr_op_07_08[7:0]),
     .top_op_08(top_op_07_08[7:0]), .tnl_op_08(tnl_op_07_08[7:0]),
     .sp4_v_t_08(sp4_v_t_07_08[47:0]), .lc_bot(tgnd_br_q),
     .op_vic(op_vic_07_08), .sp12_v_b_01(net903[0:23]));
fabric_buf_ice8p I485 ( .f_in(net0731), .f_out(padin_13_08b));
fabric_buf_ice8p I481 ( .f_in(net807), .f_out(fabric_out_13_02));
fabric_buf_ice8p I453 ( .f_in(net1437), .f_out(fabric_out_07_00));
fabric_buf_ice8p I482 ( .f_in(net808), .f_out(fabric_out_13_01));
fabric_buf_ice8p I480 ( .f_in(net809), .f_out(fabric_out_13_08));
fabric_buf_ice8p I454 ( .f_in(padinlat_b_r[11]), .f_out(padin_07_00a));
fabric_buf_ice8p I452 ( .f_in(net912), .f_out(fabric_out_12_00));
clk_quad_buf_x8_ice8p I428 ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));
clk_quad_buf_x8_ice8p I427 ( .clko(clk_tree_drv_br[7:0]),
     .clki(clk_center[7:0]));

endmodule
// Library - ice1chip, Cell - io_lft_bot_1x8_ice1f, View - schematic
// LAST TIME SAVED: Apr 11 16:03:08 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_lft_bot_1x8_ice1f ( cf_l, fabric_out_07, fabric_out_08,
     fo_dlyadj, fo_fb, fo_ref, padeb, pado, sdo, slf_op_01, slf_op_02,
     slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07, slf_op_08,
     tclk_o, SP4_h_l_01, SP4_h_l_02, SP4_h_l_03, SP4_h_l_04,
     SP4_h_l_05, SP4_h_l_06, SP4_h_l_07, SP4_h_l_08, SP12_h_l_01,
     SP12_h_l_02, SP12_h_l_03, SP12_h_l_04, SP12_h_l_05, SP12_h_l_06,
     SP12_h_l_07, SP12_h_l_08, bl, pgate, reset_b, sp4_v_b_00_01,
     sp4_v_t_08, vdd_cntl, wl, bnr_op_00_01, bs_en, ceb, glb_netwk_col,
     hiz_b, hold, jtag_rowtest_mode_rowu0_b, last_rsr, mode, padin,
     prog, r, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04, rgt_op_05,
     rgt_op_06, rgt_op_07, rgt_op_08, sdi, shift, tclk, tnr_op_08,
     update );
output  fabric_out_07, fabric_out_08, fo_fb, fo_ref, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu0_b, mode, prog,
     r, sdi, shift, tclk, update;

output [3:0]  slf_op_08;
output [3:0]  slf_op_07;
output [3:0]  slf_op_05;
output [3:0]  slf_op_04;
output [3:0]  slf_op_03;
output [3:0]  slf_op_02;
output [3:0]  slf_op_06;
output [2:0]  fo_dlyadj;
output [11:0]  padeb;
output [3:0]  slf_op_01;
output [11:0]  pado;
output [191:0]  cf_l;

inout [47:0]  SP4_h_l_05;
inout [47:0]  SP4_h_l_02;
inout [47:0]  SP4_h_l_01;
inout [17:0]  bl;
inout [15:0]  sp4_v_t_08;
inout [23:0]  SP12_h_l_04;
inout [23:0]  SP12_h_l_03;
inout [47:0]  SP4_h_l_07;
inout [47:0]  SP4_h_l_03;
inout [23:0]  SP12_h_l_02;
inout [23:0]  SP12_h_l_06;
inout [47:0]  SP4_h_l_06;
inout [47:0]  SP4_h_l_04;
inout [23:0]  SP12_h_l_07;
inout [127:0]  pgate;
inout [127:0]  vdd_cntl;
inout [127:0]  wl;
inout [127:0]  reset_b;
inout [23:0]  SP12_h_l_05;
inout [47:0]  SP4_h_l_08;
inout [23:0]  SP12_h_l_08;
inout [15:0]  sp4_v_b_00_01;
inout [23:0]  SP12_h_l_01;

input [7:0]  bnr_op_00_01;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_02;
input [7:0]  rgt_op_03;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_04;
input [0:0]  last_rsr;
input [11:0]  padin;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_08;
input [7:0]  rgt_op_07;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net1009;

wire  [0:1]  net1014;

wire  [0:1]  net1003;

wire  [7:0]  glb_netwk_t;

wire  [0:1]  net0539;

wire  [0:1]  net1001;

wire  [0:1]  net0540;

wire  [0:1]  net1005;

wire  [0:7]  net884;

wire  [0:1]  net1010;

wire  [0:15]  net937;

wire  [0:1]  net1002;

wire  [0:15]  net901;

wire  [0:7]  net1007;

wire  [0:15]  net829;

wire  [0:1]  net1013;

wire  [0:1]  net1012;

wire  [0:15]  net793;

wire  [0:7]  net704;

wire  [0:7]  net1008;

wire  [0:15]  net757;

wire  [0:1]  net755;

wire  [0:7]  net1017;

wire  [7:0]  colbuf_cntl_b;

wire  [0:7]  net1016;

wire  [0:15]  net973;

wire  [0:1]  net0538;

wire  [7:0]  colbuf_cntl_t;

wire  [0:15]  net865;

wire  [7:0]  glb_netwk_b;



fabric_buf_ice8p I_fabric_buf_8p_0015 ( .f_in(net0546),
     .f_out(fo_ref));
fabric_buf_ice8p I162 ( .f_in(net883), .f_out(fo_fb));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
io_col4_lft_ice8p_v2 I_io_00_08 ( .cbit_colcntl(net704[0:7]),
     .ceb(ceb), .sdo(net743), .sdi(sdi), .spiout({tiegnd,
     last_rsr[0]}), .cdone_in(jtag_rowtest_mode_rowu0_b),
     .spioeb({tievdd, tiegnd}), .mode(mode), .shift(shift),
     .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[11:10]), .pado(pado[11:10]),
     .padeb(padeb[11:10]), .sp4_v_t(sp4_v_t_08[15:0]),
     .sp4_h_l(SP4_h_l_08[47:0]), .sp12_h_l(SP12_h_l_08[23:0]),
     .prog(prog), .spi_ss_in_b(net1012[0:1]), .tnl_op(tnr_op_08[7:0]),
     .lft_op(rgt_op_08[7:0]), .bnl_op(rgt_op_07[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net757[0:15]), .wl(wl[127:112]), .cf(cf_l[191:168]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_08[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_08));
io_col4_lft_ice8p_v2 I_io_00_07 ( .cbit_colcntl(net1016[0:7]),
     .ceb(ceb), .sdo(net815), .sdi(net743), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(net755[0:1]), .pado(net755[0:1]),
     .padeb(net1001[0:1]), .sp4_v_t(net757[0:15]),
     .sp4_h_l(SP4_h_l_07[47:0]), .sp12_h_l(SP12_h_l_07[23:0]),
     .prog(prog), .spi_ss_in_b(net1013[0:1]), .tnl_op(rgt_op_08[7:0]),
     .lft_op(rgt_op_07[7:0]), .bnl_op(rgt_op_06[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net829[0:15]), .wl(wl[111:96]), .cf(cf_l[167:144]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_07[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_07));
io_col4_lft_ice8p_v2 I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net959), .sdi(net779), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[7:6]), .pado(pado[7:6]),
     .padeb(padeb[7:6]), .sp4_v_t(net793[0:15]),
     .sp4_h_l(SP4_h_l_05[47:0]), .sp12_h_l(SP12_h_l_05[23:0]),
     .prog(prog), .spi_ss_in_b(net1003[0:1]), .tnl_op(rgt_op_06[7:0]),
     .lft_op(rgt_op_05[7:0]), .bnl_op(rgt_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net973[0:15]), .wl(wl[79:64]), .cf(cf_l[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[1]));
io_col4_lft_ice8p_v2 I_io_00_06 ( .cbit_colcntl(net1017[0:7]),
     .ceb(ceb), .sdo(net779), .sdi(net815), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[9:8]), .pado(pado[9:8]),
     .padeb(padeb[9:8]), .sp4_v_t(net829[0:15]),
     .sp4_h_l(SP4_h_l_06[47:0]), .sp12_h_l(SP12_h_l_06[23:0]),
     .prog(prog), .spi_ss_in_b(net1010[0:1]), .tnl_op(rgt_op_07[7:0]),
     .lft_op(rgt_op_06[7:0]), .bnl_op(rgt_op_05[7:0]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net793[0:15]), .wl(wl[95:80]), .cf(cf_l[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[2]));
io_col4_lft_ice8p_v2 I_io_00_02 ( .cbit_colcntl(net1007[0:7]),
     .ceb(ceb), .sdo(net887), .sdi(net851), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .sp4_v_t(net865[0:15]),
     .sp4_h_l(SP4_h_l_02[47:0]), .sp12_h_l(SP12_h_l_02[23:0]),
     .prog(prog), .spi_ss_in_b(net1014[0:1]), .tnl_op(rgt_op_03[7:0]),
     .lft_op(rgt_op_02[7:0]), .bnl_op(rgt_op_01[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(net901[0:15]), .wl(wl[31:16]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net883));
io_col4_lft_ice8p_v2 I_io_00_01 ( .cbit_colcntl(net884[0:7]),
     .ceb(ceb), .sdo(sdo), .sdi(net887), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(net0538[0:1]), .pado(net0539[0:1]),
     .padeb(net0540[0:1]), .sp4_v_t(net901[0:15]),
     .sp4_h_l(SP4_h_l_01[47:0]), .sp12_h_l(SP12_h_l_01[23:0]),
     .prog(prog), .spi_ss_in_b(net1005[0:1]), .tnl_op(rgt_op_02[7:0]),
     .lft_op(rgt_op_01[7:0]), .bnl_op(bnr_op_00_01[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_v_b_00_01[15:0]), .wl(wl[15:0]), .cf(cf_l[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold), .fabric_out(net0546));
io_col4_lft_ice8p_v2 I_io_00_03 ( .cbit_colcntl(net1008[0:7]),
     .ceb(ceb), .sdo(net851), .sdi(net923), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[3:2]), .pado(pado[3:2]),
     .padeb(padeb[3:2]), .sp4_v_t(net937[0:15]),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b(net1009[0:1]), .tnl_op(rgt_op_04[7:0]),
     .lft_op(rgt_op_03[7:0]), .bnl_op(rgt_op_02[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net865[0:15]), .wl(wl[47:32]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net955));
io_col4_lft_ice8p_v2 I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net923), .sdi(net959), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[5:4]), .pado(pado[5:4]),
     .padeb(padeb[5:4]), .sp4_v_t(net973[0:15]),
     .sp4_h_l(SP4_h_l_04[47:0]), .sp12_h_l(SP12_h_l_04[23:0]),
     .prog(prog), .spi_ss_in_b(net1002[0:1]), .tnl_op(rgt_op_05[7:0]),
     .lft_op(rgt_op_04[7:0]), .bnl_op(rgt_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net937[0:15]), .wl(wl[63:48]), .cf(cf_l[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - ice1chip, Cell - io_bot_lft_1x6_ice1f, View - schematic
// LAST TIME SAVED: May 19 10:57:01 2011
// NETLIST TIME: Jun 29 10:32:25 2011
`timescale 1ns / 1ns 

module io_bot_lft_1x6_ice1f ( bs_en_o, ceb_o, cf_bot_l[143:0],
     fabric_out_05_00, fabric_out_06_00, fo_bypass, fo_reset, fo_sck,
     fo_sdi, hiz_b_o, mode_o, padeb_b_l[10:0], padeb_b_l[12],
     pado_b_l[10:0], pado_b_l[12], r_o, sdo, shift_o,
     slf_op_01_00[3:0], slf_op_02_00[3:0], slf_op_03_00[3:0],
     slf_op_04_00[3:0], slf_op_05_00[3:0], slf_op_06_00[3:0], tclk_o,
     update_o, bl_01[53:0], bl_02[53:0], bl_03[41:0], bl_04[53:0],
     bl_05[53:0], bl_06[53:0], sp4_h_l_01_00[15:0],
     sp4_h_r_06_00[15:0], sp4_v_b_01_00[47:0], sp4_v_b_02_00[47:0],
     sp4_v_b_03_00[47:0], sp4_v_b_04_00[47:0], sp4_v_b_05_00[47:0],
     sp4_v_b_06_00[47:0], sp12_v_b_01_00[23:0], sp12_v_b_02_00[23:0],
     sp12_v_b_03_00[23:0], sp12_v_b_04_00[23:0], sp12_v_b_05_00[23:0],
     sp12_v_b_06_00[23:0], bnl_op_01_00[7:0], bs_en_i, ceb_i,
     glb_net_01[7:0], glb_net_02[7:0], glb_net_03[7:0],
     glb_net_04[7:0], glb_net_05[7:0], glb_net_06[7:0], hiz_b_i,
     hold_b_l, lft_op_01_00[7:0], lft_op_02_00[7:0], lft_op_03_00[7:0],
     lft_op_04_00[7:0], lft_op_05_00[7:0], lft_op_06_00[7:0], mode_i,
     padin_b_l[10:0], padin_b_l[12], pgate_l[15:0], prog, r_i,
     reset_l[15:0], sdi, shift_i, tclk_i, tnr_op_06_00[7:0], update_i,
     vdd_cntl_l[15:0], wl_l[15:0] );
output  bs_en_o, ceb_o, fabric_out_05_00, fabric_out_06_00, fo_bypass,
     fo_reset, fo_sck, fo_sdi, hiz_b_o, mode_o, r_o, sdo, shift_o,
     tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_01_00;
output [3:0]  slf_op_03_00;
output [3:0]  slf_op_06_00;
output [12:0]  padeb_b_l;
output [143:0]  cf_bot_l;
output [3:0]  slf_op_05_00;
output [12:0]  pado_b_l;
output [3:0]  slf_op_04_00;
output [3:0]  slf_op_02_00;

inout [15:0]  sp4_h_r_06_00;
inout [23:0]  sp12_v_b_04_00;
inout [53:0]  bl_05;
inout [53:0]  bl_02;
inout [53:0]  bl_01;
inout [41:0]  bl_03;
inout [53:0]  bl_04;
inout [23:0]  sp12_v_b_01_00;
inout [47:0]  sp4_v_b_05_00;
inout [23:0]  sp12_v_b_02_00;
inout [15:0]  sp4_h_l_01_00;
inout [47:0]  sp4_v_b_03_00;
inout [23:0]  sp12_v_b_05_00;
inout [47:0]  sp4_v_b_04_00;
inout [53:0]  bl_06;
inout [47:0]  sp4_v_b_01_00;
inout [47:0]  sp4_v_b_02_00;
inout [23:0]  sp12_v_b_06_00;
inout [23:0]  sp12_v_b_03_00;
inout [47:0]  sp4_v_b_06_00;

input [15:0]  pgate_l;
input [7:0]  lft_op_01_00;
input [7:0]  glb_net_01;
input [7:0]  lft_op_03_00;
input [7:0]  lft_op_02_00;
input [15:0]  vdd_cntl_l;
input [7:0]  lft_op_06_00;
input [15:0]  wl_l;
input [12:0]  padin_b_l;
input [7:0]  bnl_op_01_00;
input [7:0]  glb_net_03;
input [15:0]  reset_l;
input [7:0]  glb_net_06;
input [7:0]  tnr_op_06_00;
input [7:0]  lft_op_04_00;
input [7:0]  glb_net_02;
input [7:0]  lft_op_05_00;
input [7:0]  glb_net_05;
input [7:0]  glb_net_04;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net519;

wire  [0:1]  net382;

wire  [0:15]  net483;

wire  [0:1]  net452;

wire  [0:15]  net378;

wire  [0:15]  net413;

wire  [0:15]  net308;

wire  [0:1]  net520;

wire  [0:1]  net487;

wire  [0:1]  net312;

wire  [0:15]  net343;



scan_buf_ice8p I_scanbuf_bl ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net284), .shift_o(shift_o),
     .sdo(net286), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_bot_ice8p I_IO_02_00 ( .sdo(net292), .sdi(net362),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net378[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b_l[3:2]), .pado(pado_b_l[3:2]),
     .padeb(padeb_b_l[3:2]), .sp4_v_b(net308[0:15]),
     .sp4_h_l(sp4_v_b_02_00[47:0]), .sp12_h_l(sp12_v_b_02_00[23:0]),
     .prog(prog), .spi_ss_in_b(net312[0:1]),
     .tnl_op(lft_op_01_00[7:0]), .lft_op(lft_op_02_00[7:0]),
     .bnl_op(lft_op_03_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[47:24]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_00[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_b_l), .fabric_out(fo_reset));
io_col4_bot_ice8p I_IO_03_00_bram ( .sdo(net327), .sdi(net292),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net308[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b_l[5:4]), .pado(pado_b_l[5:4]),
     .padeb(padeb_b_l[5:4]), .sp4_v_b(net343[0:15]),
     .sp4_h_l(sp4_v_b_03_00[47:0]), .sp12_h_l(sp12_v_b_03_00[23:0]),
     .prog(prog), .spi_ss_in_b(net519[0:1]),
     .tnl_op(lft_op_02_00[7:0]), .lft_op(lft_op_03_00[7:0]),
     .bnl_op(lft_op_04_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[71:48]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_00[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_b_l), .fabric_out(fo_sck));
io_col4_bot_ice8p I_IO_01_00 ( .sdo(net362), .sdi(net286),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_01_00[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b_l[1:0]),
     .pado(pado_b_l[1:0]), .padeb(padeb_b_l[1:0]),
     .sp4_v_b(net378[0:15]), .sp4_h_l(sp4_v_b_01_00[47:0]),
     .sp12_h_l(sp12_v_b_01_00[23:0]), .prog(prog),
     .spi_ss_in_b(net382[0:1]), .tnl_op(bnl_op_01_00[7:0]),
     .lft_op(lft_op_01_00[7:0]), .bnl_op(lft_op_02_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_01[5],
     bl_01[4], bl_01[37], bl_01[36], bl_01[35], bl_01[34], bl_01[33],
     bl_01[32], bl_01[14], bl_01[20], bl_01[19], bl_01[18], bl_01[17],
     bl_01[16], bl_01[27], bl_01[26], bl_01[25], bl_01[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[23:0]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_01_00[3:0]),
     .glb_netwk(glb_net_01[7:0]), .hold(hold_b_l),
     .fabric_out(fo_bypass));
io_col4_bot_ice8p I_IO_05_00 ( .sdo(net397), .sdi(net467),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net483[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b_l[9:8]), .pado(pado_b_l[9:8]),
     .padeb(padeb_b_l[9:8]), .sp4_v_b(net413[0:15]),
     .sp4_h_l(sp4_v_b_05_00[47:0]), .sp12_h_l(sp12_v_b_05_00[23:0]),
     .prog(prog), .spi_ss_in_b(net520[0:1]),
     .tnl_op(lft_op_04_00[7:0]), .lft_op(lft_op_05_00[7:0]),
     .bnl_op(lft_op_06_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[119:96]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_00[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_b_l), .fabric_out(fabric_out_05_00));
io_col4_bot_ice8p I_IO_06_00 ( .sdo(sdo), .sdi(net397),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net413[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin({padin_b_l[10], padin_b_l[12]}),
     .pado({pado_b_l[10], pado_b_l[12]}), .padeb({padeb_b_l[10],
     padeb_b_l[12]}), .sp4_v_b(sp4_h_r_06_00[15:0]),
     .sp4_h_l(sp4_v_b_06_00[47:0]), .sp12_h_l(sp12_v_b_06_00[23:0]),
     .prog(prog), .spi_ss_in_b(net452[0:1]),
     .tnl_op(lft_op_05_00[7:0]), .lft_op(lft_op_06_00[7:0]),
     .bnl_op(tnr_op_06_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_06[5], bl_06[4], bl_06[37],
     bl_06[36], bl_06[35], bl_06[34], bl_06[33], bl_06[32], bl_06[14],
     bl_06[20], bl_06[19], bl_06[18], bl_06[17], bl_06[16], bl_06[27],
     bl_06[26], bl_06[25], bl_06[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[143:120]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_00[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_b_l), .fabric_out(fabric_out_06_00));
io_col4_bot_ice8p I_IO_04_00 ( .sdo(net467), .sdi(net327),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(net343[0:15]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b_l[7:6]), .pado(pado_b_l[7:6]),
     .padeb(padeb_b_l[7:6]), .sp4_v_b(net483[0:15]),
     .sp4_h_l(sp4_v_b_04_00[47:0]), .sp12_h_l(sp12_v_b_04_00[23:0]),
     .prog(prog), .spi_ss_in_b(net487[0:1]),
     .tnl_op(lft_op_03_00[7:0]), .lft_op(lft_op_04_00[7:0]),
     .bnl_op(lft_op_05_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[95:72]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_00[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_b_l), .fabric_out(fo_sdi));
tckbufx32_ice8p I354 ( .in(net284), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));

endmodule
// Library - ice1chip, Cell - quad_bl_ice1, View - schematic
// LAST TIME SAVED: May 19 11:18:19 2011
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module quad_bl_ice1 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o[7:0],
     bm_sclk_o, bm_sclkrw_o[1:0], bm_sdi_o[1:0], bm_sdo_o[1:0],
     bm_sreb_o, bm_sweb_o[1:0], bm_wdummymux_en_o, bs_en_o,
     carry_out_01_08, carry_out_02_08, carry_out_04_08,
     carry_out_05_08, carry_out_06_08, ceb_o, cf_b_l[143:0],
     cf_l[191:0], fabric_out_00_07, fabric_out_00_08, fabric_out_05_00,
     fabric_out_06_00, fo_bypass, fo_dlyadj[2:0], fo_fb, fo_ref,
     fo_reset, fo_sck, fo_sdi, hiz_b_o, mode_o, op_vic_01_08,
     op_vic_02_08, op_vic_04_08, op_vic_05_08, op_vic_06_08,
     padeb_b_l[10:0], padeb_b_l[12], padeb_l_b[11:0], padin_00_08,
     padin_06_00, pado_b_l[10:0], pado_b_l[12], pado_l_b[11:0], r_o,
     sdo, shift_o, slf_op_00_08[3:0], slf_op_01_08[7:0],
     slf_op_02_08[7:0], slf_op_03_08[7:0], slf_op_04_08[7:0],
     slf_op_05_08[7:0], slf_op_06_00[3:0], slf_op_06_01[7:0],
     slf_op_06_02[7:0], slf_op_06_03[7:0], slf_op_06_04[7:0],
     slf_op_06_05[7:0], slf_op_06_06[7:0], slf_op_06_07[7:0],
     slf_op_06_08[7:0], tclk_o, update_o, bl[329:0], pgate_l[143:0],
     reset_b_l[143:0], sp4_h_r_06_00[15:0], sp4_h_r_06_01[47:0],
     sp4_h_r_06_02[47:0], sp4_h_r_06_03[47:0], sp4_h_r_06_04[47:0],
     sp4_h_r_06_05[47:0], sp4_h_r_06_06[47:0], sp4_h_r_06_07[47:0],
     sp4_h_r_06_08[47:0], sp4_r_v_b_06_01[47:0], sp4_r_v_b_06_02[47:0],
     sp4_r_v_b_06_03[47:0], sp4_r_v_b_06_04[47:0],
     sp4_r_v_b_06_05[47:0], sp4_r_v_b_06_06[47:0],
     sp4_r_v_b_06_07[47:0], sp4_r_v_b_06_08[47:0], sp4_v_t_00_08[15:0],
     sp4_v_t_01_08[47:0], sp4_v_t_02_08[47:0], sp4_v_t_03_08[47:0],
     sp4_v_t_04_08[47:0], sp4_v_t_05_08[47:0], sp4_v_t_06_08[47:0],
     sp12_h_r_06_01[23:0], sp12_h_r_06_02[23:0], sp12_h_r_06_03[23:0],
     sp12_h_r_06_04[23:0], sp12_h_r_06_05[23:0], sp12_h_r_06_06[23:0],
     sp12_h_r_06_07[23:0], sp12_h_r_06_08[23:0], sp12_v_t_01_08[23:0],
     sp12_v_t_02_08[23:0], sp12_v_t_03_08[23:0], sp12_v_t_04_08[23:0],
     sp12_v_t_05_08[23:0], sp12_v_t_06_08[23:0], vdd_cntl_l[143:0],
     wl_l[143:0], bm_aa_top[10:0], bm_ab_top[10:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i[1:0],
     bm_sdi_i[1:0], bm_sdo_i[1:0], bm_sreb_i, bm_sweb_i[1:0],
     bm_wdummymux_en_i, bnr_op_06_01[3:0], bs_en_i, ceb_i, glb_in[7:0],
     hiz_b_i, hold_b_l, hold_l_b, jtag_rowtest_mode_rowu0_b,
     last_rsr[0], mode_i, padin_b_l[10:0], padin_b_l[12],
     padin_l_b[11:0], pll_lock_out, prog, purst, r_i,
     rgt_op_06_01[7:0], rgt_op_06_02[7:0], rgt_op_06_03[7:0],
     rgt_op_06_04[7:0], rgt_op_06_05[7:0], rgt_op_06_06[7:0],
     rgt_op_06_07[7:0], rgt_op_06_08[7:0], sdi, shift_i, tclk_i,
     tnl_op_01_08[7:0], tnl_op_02_08[7:0], tnl_op_03_08[7:0],
     tnl_op_04_08[7:0], tnl_op_05_08[7:0], tnl_op_06_08[7:0],
     tnr_op_00_08[7:0], tnr_op_01_08[7:0], tnr_op_02_08[7:0],
     tnr_op_03_08[7:0], tnr_op_04_08[7:0], tnr_op_05_08[7:0],
     tnr_op_06_08[7:0], top_op_01_08[7:0], top_op_02_08[7:0],
     top_op_03_08[7:0], top_op_04_08[7:0], top_op_05_08[7:0],
     top_op_06_08[7:0], update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_08, carry_out_02_08,
     carry_out_04_08, carry_out_05_08, carry_out_06_08, ceb_o,
     fabric_out_00_07, fabric_out_00_08, fabric_out_05_00,
     fabric_out_06_00, fo_bypass, fo_fb, fo_ref, fo_reset, fo_sck,
     fo_sdi, hiz_b_o, mode_o, op_vic_01_08, op_vic_02_08, op_vic_04_08,
     op_vic_05_08, op_vic_06_08, padin_00_08, padin_06_00, r_o, sdo,
     shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, ceb_i, hiz_b_i, hold_b_l, hold_l_b,
     jtag_rowtest_mode_rowu0_b, mode_i, pll_lock_out, prog, purst, r_i,
     sdi, shift_i, tclk_i, update_i;

output [7:0]  slf_op_04_08;
output [7:0]  slf_op_06_07;
output [7:0]  slf_op_06_03;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_06_01;
output [7:0]  slf_op_06_02;
output [2:0]  fo_dlyadj;
output [11:0]  pado_l_b;
output [7:0]  slf_op_05_08;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_06_04;
output [7:0]  slf_op_06_06;
output [191:0]  cf_l;
output [11:0]  padeb_l_b;
output [3:0]  slf_op_06_00;
output [12:0]  pado_b_l;
output [143:0]  cf_b_l;
output [12:0]  padeb_b_l;
output [7:0]  slf_op_06_08;
output [3:0]  slf_op_00_08;
output [7:0]  slf_op_02_08;
output [7:0]  slf_op_03_08;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_01_08;
output [7:0]  slf_op_06_05;

inout [47:0]  sp4_r_v_b_06_04;
inout [23:0]  sp12_h_r_06_06;
inout [47:0]  sp4_h_r_06_01;
inout [47:0]  sp4_h_r_06_06;
inout [47:0]  sp4_h_r_06_04;
inout [47:0]  sp4_r_v_b_06_08;
inout [23:0]  sp12_v_t_03_08;
inout [47:0]  sp4_h_r_06_05;
inout [47:0]  sp4_r_v_b_06_06;
inout [15:0]  sp4_h_r_06_00;
inout [47:0]  sp4_v_t_01_08;
inout [23:0]  sp12_v_t_06_08;
inout [23:0]  sp12_v_t_04_08;
inout [47:0]  sp4_v_t_06_08;
inout [47:0]  sp4_h_r_06_07;
inout [23:0]  sp12_h_r_06_07;
inout [47:0]  sp4_v_t_04_08;
inout [47:0]  sp4_h_r_06_08;
inout [47:0]  sp4_h_r_06_03;
inout [23:0]  sp12_h_r_06_01;
inout [47:0]  sp4_r_v_b_06_01;
inout [23:0]  sp12_v_t_02_08;
inout [23:0]  sp12_v_t_01_08;
inout [47:0]  sp4_r_v_b_06_05;
inout [143:0]  pgate_l;
inout [23:0]  sp12_v_t_05_08;
inout [23:0]  sp12_h_r_06_05;
inout [329:0]  bl;
inout [47:0]  sp4_r_v_b_06_07;
inout [143:0]  vdd_cntl_l;
inout [47:0]  sp4_v_t_02_08;
inout [47:0]  sp4_v_t_05_08;
inout [143:0]  reset_b_l;
inout [23:0]  sp12_h_r_06_03;
inout [15:0]  sp4_v_t_00_08;
inout [143:0]  wl_l;
inout [47:0]  sp4_r_v_b_06_02;
inout [23:0]  sp12_h_r_06_02;
inout [47:0]  sp4_r_v_b_06_03;
inout [23:0]  sp12_h_r_06_08;
inout [47:0]  sp4_h_r_06_02;
inout [23:0]  sp12_h_r_06_04;
inout [47:0]  sp4_v_t_03_08;

input [7:0]  tnl_op_01_08;
input [7:0]  tnr_op_00_08;
input [7:0]  rgt_op_06_06;
input [1:0]  bm_sclkrw_i;
input [7:0]  tnl_op_04_08;
input [7:0]  tnr_op_04_08;
input [7:0]  rgt_op_06_08;
input [7:0]  tnr_op_01_08;
input [1:0]  bm_sdi_i;
input [10:0]  bm_aa_top;
input [7:0]  rgt_op_06_04;
input [1:0]  bm_sdo_i;
input [7:0]  tnl_op_02_08;
input [7:0]  tnr_op_02_08;
input [7:0]  rgt_op_06_02;
input [0:0]  last_rsr;
input [7:0]  top_op_05_08;
input [7:0]  top_op_04_08;
input [7:0]  rgt_op_06_07;
input [7:0]  top_op_02_08;
input [7:0]  top_op_01_08;
input [7:0]  tnr_op_03_08;
input [11:0]  padin_l_b;
input [7:0]  tnl_op_05_08;
input [1:0]  bm_sweb_i;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_03_08;
input [7:0]  top_op_06_08;
input [7:0]  rgt_op_06_05;
input [7:0]  tnl_op_06_08;
input [7:0]  top_op_03_08;
input [3:0]  bnr_op_06_01;
input [7:0]  rgt_op_06_03;
input [10:0]  bm_ab_top;
input [7:0]  tnr_op_06_08;
input [7:0]  tnr_op_05_08;
input [7:0]  glb_in;
input [12:0]  padin_b_l;
input [7:0]  rgt_op_06_01;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:47]  net877;

wire  [0:47]  net972;

wire  [0:23]  net940;

wire  [0:47]  net1456;

wire  [0:47]  net792;

wire  [0:23]  net896;

wire  [0:7]  net921;

wire  [0:47]  net1230;

wire  [0:23]  net1363;

wire  [0:7]  net1343;

wire  [0:23]  net744;

wire  [0:47]  net763;

wire  [0:7]  net1168;

wire  [7:0]  clk_center;

wire  [0:7]  net1107;

wire  [0:47]  net791;

wire  [0:7]  net929;

wire  [0:23]  net938;

wire  [0:47]  net820;

wire  [11:11]  padinlat_l_b;

wire  [0:23]  net777;

wire  [0:47]  net1228;

wire  [0:47]  net994;

wire  [0:23]  net989;

wire  [0:47]  net1339;

wire  [0:47]  net1425;

wire  [0:23]  net1357;

wire  [0:47]  net945;

wire  [0:7]  net1438;

wire  [0:10]  net1458;

wire  [0:47]  net1231;

wire  [0:7]  net886;

wire  [0:47]  net899;

wire  [0:47]  net995;

wire  [0:7]  net798;

wire  [0:7]  net814;

wire  [0:47]  net1132;

wire  [0:7]  net1109;

wire  [0:7]  net1329;

wire  [0:47]  net1000;

wire  [0:47]  net1181;

wire  [0:23]  net768;

wire  [0:23]  net1426;

wire  [0:47]  net1184;

wire  [0:23]  net845;

wire  [10:10]  padinlat_b_l;

wire  [0:47]  net819;

wire  [0:47]  net1158;

wire  [0:47]  net962;

wire  [0:47]  net1452;

wire  [0:23]  net941;

wire  [0:47]  net756;

wire  [0:47]  net949;

wire  [0:23]  net1273;

wire  [0:47]  net951;

wire  [7:0]  clk_tree_drv_bl;

wire  [0:47]  net993;

wire  [0:47]  net901;

wire  [0:47]  net774;

wire  [0:47]  net1277;

wire  [0:47]  net944;

wire  [0:47]  net997;

wire  [0:47]  net759;

wire  [0:7]  net1167;

wire  [0:7]  net979;

wire  [0:47]  net1227;

wire  [0:47]  net900;

wire  [0:7]  net980;

wire  [0:7]  net801;

wire  [0:47]  net1319;

wire  [0:47]  net1336;

wire  [0:47]  net1160;

wire  [0:23]  net1445;

wire  [0:23]  net1365;

wire  [0:47]  net1341;

wire  [0:23]  net990;

wire  [0:7]  net1344;

wire  [0:23]  net1127;

wire  [3:0]  slf_op_00_02;

wire  [0:23]  net1392;

wire  [0:7]  net1367;

wire  [0:47]  net1233;

wire  [0:47]  net851;

wire  [0:47]  net971;

wire  [3:0]  slf_op_00_01;

wire  [0:23]  net1178;

wire  [0:47]  net999;

wire  [0:23]  net1271;

wire  [0:7]  net1428;

wire  [0:47]  net948;

wire  [0:7]  net834;

wire  [0:23]  net1272;

wire  [0:7]  net800;

wire  [0:23]  net1360;

wire  [0:7]  net1406;

wire  [0:47]  net946;

wire  [0:47]  net902;

wire  [0:23]  net1128;

wire  [0:7]  net978;

wire  [0:7]  net885;

wire  [0:47]  net1276;

wire  [0:7]  net799;

wire  [0:23]  net1177;

wire  [0:7]  net1404;

wire  [0:7]  net1436;

wire  [0:23]  net1423;

wire  [0:23]  net1179;

wire  [0:23]  net1270;

wire  [0:47]  net1139;

wire  [0:47]  net1138;

wire  [0:23]  net1222;

wire  [0:47]  net1430;

wire  [0:23]  net776;

wire  [0:7]  net826;

wire  [0:23]  net847;

wire  [0:47]  net1133;

wire  [0:23]  net749;

wire  [0:47]  net1254;

wire  [0:47]  net950;

wire  [0:23]  net988;

wire  [0:47]  net1278;

wire  [0:47]  net1136;

wire  [0:47]  net821;

wire  [0:47]  net850;

wire  [0:47]  net1251;

wire  [0:47]  net875;

wire  [0:47]  net852;

wire  [0:47]  net854;

wire  [0:23]  net1126;

wire  [0:47]  net1338;

wire  [0:47]  net1253;

wire  [0:7]  net1427;

wire  [0:47]  net1134;

wire  [0:23]  net846;

wire  [0:23]  net939;

wire  [0:23]  net1356;

wire  [0:23]  net1220;

wire  [0:47]  net1330;

wire  [0:23]  net1358;

wire  [0:15]  net1326;

wire  [3:0]  slf_op_02_00;

wire  [0:47]  net1226;

wire  [0:47]  net855;

wire  [0:47]  net969;

wire  [0:23]  net991;

wire  [3:0]  slf_op_05_00;

wire  [0:23]  net897;

wire  [0:23]  net1223;

wire  [0:23]  net1129;

wire  [0:47]  net1433;

wire  [0:47]  net1454;

wire  [0:7]  net919;

wire  [0:47]  net752;

wire  [0:23]  net1221;

wire  [0:23]  net746;

wire  [0:47]  net1252;

wire  [3:0]  slf_op_00_07;

wire  [0:23]  net894;

wire  [0:7]  net824;

wire  [0:47]  net818;

wire  [0:23]  net844;

wire  [0:23]  net1409;

wire  [3:0]  slf_op_00_05;

wire  [0:47]  net1137;

wire  [0:47]  net760;

wire  [0:47]  net793;

wire  [0:47]  net1182;

wire  [3:0]  slf_op_01_00;

wire  [0:47]  net1183;

wire  [0:47]  net1337;

wire  [0:23]  net1355;

wire  [0:7]  net1166;

wire  [0:23]  net748;

wire  [0:47]  net822;

wire  [0:47]  net996;

wire  [0:47]  net856;

wire  [0:7]  net884;

wire  [0:47]  net998;

wire  [0:47]  net823;

wire  [0:47]  net878;

wire  [0:7]  net1345;

wire  [0:10]  net788;

wire  [0:47]  net1157;

wire  [0:23]  net895;

wire  [3:0]  slf_op_00_06;

wire  [0:7]  net1402;

wire  [0:7]  net1117;

wire  [0:7]  net797;

wire  [0:7]  net1407;

wire  [0:47]  net1421;

wire  [0:47]  net1159;

wire  [0:47]  net1340;

wire  [0:47]  net1431;

wire  [0:47]  net1275;

wire  [0:47]  net1232;

wire  [0:47]  net970;

wire  [0:7]  net1429;

wire  [3:0]  slf_op_00_04;

wire  [3:0]  slf_op_04_00;

wire  [3:0]  slf_op_00_03;

wire  [0:7]  net796;

wire  [0:23]  net1361;

wire  [0:7]  net1342;

wire  [0:47]  net876;

wire  [3:0]  slf_op_03_00;

wire  [0:23]  net1176;

wire  [0:7]  net1403;

wire  [0:23]  net732;

wire  [0:23]  net1432;

wire  [0:7]  net1405;

wire  [0:47]  net857;



bram1x4_ice1f I_bram_col_t03 ( .prog(prog),
     .glb_netwk_col(clk_tree_drv_bl[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .reset_b(reset_b_l[143:16]),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sreb_o(bm_sreb_o),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .lft_op_05(net980[0:7]), .bl(bl[167:126]),
     .sp4_h_l_06(net877[0:47]), .sp12_h_l_02(net846[0:23]),
     .lft_op_06(net979[0:7]), .sp12_h_l_03(net845[0:23]),
     .sp12_h_r_03(net732[0:23]), .sp12_h_l_01(net847[0:23]),
     .sp4_v_b_04(net850[0:47]), .sp4_v_b_05(net899[0:47]),
     .lft_op_07(net978[0:7]), .sp4_v_b_06(net900[0:47]),
     .sp4_v_b_08(net902[0:47]), .sp4_v_b_07(net901[0:47]),
     .lft_op_03(net919[0:7]), .lft_op_01(net1438[0:7]),
     .sp4_h_l_02(net856[0:47]), .sp12_h_l_06(net895[0:23]),
     .sp12_h_r_07(net744[0:23]), .sp12_h_l_05(net894[0:23]),
     .sp12_h_r_06(net746[0:23]), .sp12_h_l_04(net844[0:23]),
     .sp12_h_r_05(net748[0:23]), .sp12_h_r_08(net749[0:23]),
     .sp12_h_l_07(net896[0:23]), .sp12_h_l_08(net897[0:23]),
     .sp4_r_v_b_03(net752[0:47]), .vdd_cntl(vdd_cntl_l[143:16]),
     .pgate(pgate_l[143:16]), .bot_op_01({slf_op_03_00[3],
     slf_op_03_00[2], slf_op_03_00[1], slf_op_03_00[0],
     slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0]}), .sp4_r_v_b_04(net756[0:47]),
     .sp4_v_b_01(net1431[0:47]), .sp4_v_b_03(net851[0:47]),
     .sp4_h_r_08(net759[0:47]), .sp4_r_v_b_05(net760[0:47]),
     .sp4_v_b_02(net852[0:47]), .sp4_v_t_08(sp4_v_t_03_08[47:0]),
     .sp4_r_v_b_02(net763[0:47]), .bnr_op_01({slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0],
     slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0]}), .bm_sdi_o(bm_sdi_o[1:0]),
     .sp4_h_l_04(net854[0:47]), .lft_op_08(slf_op_02_08[7:0]),
     .sp12_h_r_01(net768[0:23]), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .sp4_h_l_03(net855[0:47]), .sp4_h_l_01(net857[0:47]),
     .sp4_h_r_01(net774[0:47]), .tnr_op_08(tnr_op_03_08[7:0]),
     .sp12_h_r_02(net776[0:23]), .sp12_h_r_04(net777[0:23]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .lft_op_02(net921[0:7]), .lft_op_04(net929[0:7]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bnl_op_01({slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0],
     slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0]}), .sp12_v_t_08(sp12_v_t_03_08[23:0]),
     .wl(wl_l[143:16]), .tnl_op_08(tnl_op_03_08[7:0]),
     .top_op_08(top_op_03_08[7:0]), .bm_ab_2bot(net788[0:10]),
     .bm_aa_2bot(net1458[0:10]), .sp12_v_b_01(net1432[0:23]),
     .sp4_r_v_b_08(net791[0:47]), .sp4_r_v_b_07(net792[0:47]),
     .sp4_r_v_b_06(net793[0:47]), .sp4_r_v_b_01(net1433[0:47]),
     .rgt_op_08(slf_op_04_08[7:0]), .rgt_op_07(net796[0:7]),
     .rgt_op_06(net797[0:7]), .rgt_op_05(net798[0:7]),
     .rgt_op_04(net799[0:7]), .rgt_op_03(net800[0:7]),
     .rgt_op_02(net801[0:7]), .rgt_op_01(net1427[0:7]),
     .slf_op_02(net826[0:7]), .slf_op_01(net1429[0:7]),
     .slf_op_03(net824[0:7]), .slf_op_04(net834[0:7]),
     .slf_op_05(net886[0:7]), .slf_op_06(net885[0:7]),
     .slf_op_07(net884[0:7]), .slf_op_08(slf_op_03_08[7:0]),
     .bm_ab_top(bm_ab_top[10:0]), .bm_aa_top(bm_aa_top[10:0]),
     .glb_netwk_bot(net1405[0:7]), .glb_netwk_top(net814[0:7]),
     .sp4_h_l_08(net875[0:47]), .sp4_h_l_07(net876[0:47]),
     .sp4_h_l_05(net878[0:47]), .sp4_h_r_02(net818[0:47]),
     .sp4_h_r_03(net819[0:47]), .sp4_h_r_04(net820[0:47]),
     .sp4_h_r_05(net821[0:47]), .sp4_h_r_06(net822[0:47]),
     .sp4_h_r_07(net823[0:47]));
lt_1x8_bot_ice1f I_lt_col_t02 ( .rgt_op_03(net824[0:7]),
     .slf_op_02(net921[0:7]), .rgt_op_02(net826[0:7]),
     .rgt_op_01(net1429[0:7]), .purst(purst), .prog(prog),
     .lft_op_04(net1367[0:7]), .lft_op_03(net1345[0:7]),
     .lft_op_02(net1329[0:7]), .lft_op_01(net1436[0:7]),
     .rgt_op_04(net834[0:7]), .glb_netwk_bot(net1406[0:7]),
     .carry_in(tiegnd_bl), .bnl_op_01({slf_op_01_00[3],
     slf_op_01_00[2], slf_op_01_00[1], slf_op_01_00[0],
     slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0]}), .slf_op_04(net929[0:7]),
     .slf_op_03(net919[0:7]), .slf_op_01(net1438[0:7]),
     .sp4_h_l_04(net948[0:47]), .carry_out(carry_out_02_08),
     .vdd_cntl(vdd_cntl_l[143:16]), .sp12_h_r_04(net844[0:23]),
     .sp12_h_r_03(net845[0:23]), .sp12_h_r_02(net846[0:23]),
     .sp12_h_r_01(net847[0:23]), .glb_netwk_col(clk_tree_drv_bl[7:0]),
     .sp4_v_b_01(net1430[0:47]), .sp4_r_v_b_04(net850[0:47]),
     .sp4_r_v_b_03(net851[0:47]), .sp4_r_v_b_02(net852[0:47]),
     .sp4_r_v_b_01(net1431[0:47]), .sp4_h_r_04(net854[0:47]),
     .sp4_h_r_03(net855[0:47]), .sp4_h_r_02(net856[0:47]),
     .sp4_h_r_01(net857[0:47]), .sp4_h_l_03(net949[0:47]),
     .sp4_h_l_02(net950[0:47]), .sp4_h_l_01(net951[0:47]),
     .bl(bl[125:72]), .bot_op_01({slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0], slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0]}),
     .sp12_h_l_01(net941[0:23]), .sp12_h_l_02(net940[0:23]),
     .sp12_h_l_03(net939[0:23]), .sp12_h_l_04(net938[0:23]),
     .sp4_v_b_04(net944[0:47]), .sp4_v_b_03(net945[0:47]),
     .sp4_v_b_02(net946[0:47]), .bnr_op_01({slf_op_03_00[3],
     slf_op_03_00[2], slf_op_03_00[1], slf_op_03_00[0],
     slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0]}), .sp4_h_l_05(net972[0:47]),
     .sp4_h_l_06(net971[0:47]), .sp4_h_l_07(net970[0:47]),
     .sp4_h_l_08(net969[0:47]), .sp4_h_r_08(net875[0:47]),
     .sp4_h_r_07(net876[0:47]), .sp4_h_r_06(net877[0:47]),
     .sp4_h_r_05(net878[0:47]), .slf_op_05(net980[0:7]),
     .slf_op_06(net979[0:7]), .slf_op_07(net978[0:7]),
     .slf_op_08(slf_op_02_08[7:0]), .rgt_op_08(slf_op_03_08[7:0]),
     .rgt_op_07(net884[0:7]), .rgt_op_06(net885[0:7]),
     .rgt_op_05(net886[0:7]), .lft_op_08(slf_op_01_08[7:0]),
     .lft_op_07(net1342[0:7]), .lft_op_06(net1343[0:7]),
     .lft_op_05(net1344[0:7]), .sp12_h_l_08(net991[0:23]),
     .sp12_h_l_07(net990[0:23]), .sp12_h_l_06(net989[0:23]),
     .sp12_h_r_05(net894[0:23]), .sp12_h_r_06(net895[0:23]),
     .sp12_h_r_07(net896[0:23]), .sp12_h_r_08(net897[0:23]),
     .sp12_h_l_05(net988[0:23]), .sp4_r_v_b_05(net899[0:47]),
     .sp4_r_v_b_06(net900[0:47]), .sp4_r_v_b_07(net901[0:47]),
     .sp4_r_v_b_08(net902[0:47]), .sp4_v_b_08(net996[0:47]),
     .sp4_v_b_07(net995[0:47]), .sp4_v_b_06(net994[0:47]),
     .sp4_v_b_05(net993[0:47]), .pgate(pgate_l[143:16]),
     .reset_b(reset_b_l[143:16]), .wl(wl_l[143:16]),
     .top_op_08(top_op_02_08[7:0]), .tnr_op_08(tnr_op_02_08[7:0]),
     .tnl_op_08(tnl_op_02_08[7:0]), .sp12_v_t_08(sp12_v_t_02_08[23:0]),
     .sp4_v_t_08(sp4_v_t_02_08[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_02_08), .sp12_v_b_01(net1409[0:23]));
lt_1x8_bot_ice1f I_lt_col_t01 ( .glb_netwk_bot(net1407[0:7]),
     .rgt_op_03(net919[0:7]), .slf_op_02(net1329[0:7]),
     .rgt_op_02(net921[0:7]), .rgt_op_01(net1438[0:7]), .purst(purst),
     .prog(prog), .lft_op_04({slf_op_00_04[3], slf_op_00_04[2],
     slf_op_00_04[1], slf_op_00_04[0], slf_op_00_04[3],
     slf_op_00_04[2], slf_op_00_04[1], slf_op_00_04[0]}),
     .lft_op_03({slf_op_00_03[3], slf_op_00_03[2], slf_op_00_03[1],
     slf_op_00_03[0], slf_op_00_03[3], slf_op_00_03[2],
     slf_op_00_03[1], slf_op_00_03[0]}), .lft_op_02({slf_op_00_02[3],
     slf_op_00_02[2], slf_op_00_02[1], slf_op_00_02[0],
     slf_op_00_02[3], slf_op_00_02[2], slf_op_00_02[1],
     slf_op_00_02[0]}), .lft_op_01({slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0], slf_op_00_01[3],
     slf_op_00_01[2], slf_op_00_01[1], slf_op_00_01[0]}),
     .rgt_op_04(net929[0:7]), .carry_in(tiegnd_bl),
     .bnl_op_01({pll_lock_out, pll_lock_out, pll_lock_out,
     pll_lock_out, pll_lock_out, pll_lock_out, pll_lock_out,
     pll_lock_out}), .slf_op_04(net1367[0:7]),
     .slf_op_03(net1345[0:7]), .slf_op_01(net1436[0:7]),
     .sp4_h_l_04(net1339[0:47]), .carry_out(carry_out_01_08),
     .vdd_cntl(vdd_cntl_l[143:16]), .sp12_h_r_04(net938[0:23]),
     .sp12_h_r_03(net939[0:23]), .sp12_h_r_02(net940[0:23]),
     .sp12_h_r_01(net941[0:23]), .glb_netwk_col(clk_tree_drv_bl[7:0]),
     .sp4_v_b_01(net1456[0:47]), .sp4_r_v_b_04(net944[0:47]),
     .sp4_r_v_b_03(net945[0:47]), .sp4_r_v_b_02(net946[0:47]),
     .sp4_r_v_b_01(net1430[0:47]), .sp4_h_r_04(net948[0:47]),
     .sp4_h_r_03(net949[0:47]), .sp4_h_r_02(net950[0:47]),
     .sp4_h_r_01(net951[0:47]), .sp4_h_l_03(net1338[0:47]),
     .sp4_h_l_02(net1340[0:47]), .sp4_h_l_01(net1341[0:47]),
     .bl(bl[71:18]), .bot_op_01({slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0], slf_op_01_00[3],
     slf_op_01_00[2], slf_op_01_00[1], slf_op_01_00[0]}),
     .sp12_h_l_01(net1361[0:23]), .sp12_h_l_02(net1355[0:23]),
     .sp12_h_l_03(net1363[0:23]), .sp12_h_l_04(net1356[0:23]),
     .sp4_v_b_04(net1452[0:47]), .sp4_v_b_03(net962[0:47]),
     .sp4_v_b_02(net1454[0:47]), .bnr_op_01({slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0],
     slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0]}), .sp4_h_l_05(net1319[0:47]),
     .sp4_h_l_06(net1330[0:47]), .sp4_h_l_07(net1337[0:47]),
     .sp4_h_l_08(net1336[0:47]), .sp4_h_r_08(net969[0:47]),
     .sp4_h_r_07(net970[0:47]), .sp4_h_r_06(net971[0:47]),
     .sp4_h_r_05(net972[0:47]), .slf_op_05(net1344[0:7]),
     .slf_op_06(net1343[0:7]), .slf_op_07(net1342[0:7]),
     .slf_op_08(slf_op_01_08[7:0]), .rgt_op_08(slf_op_02_08[7:0]),
     .rgt_op_07(net978[0:7]), .rgt_op_06(net979[0:7]),
     .rgt_op_05(net980[0:7]), .lft_op_08({slf_op_00_08[3],
     slf_op_00_08[2], slf_op_00_08[1], slf_op_00_08[0],
     slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0]}), .lft_op_07({slf_op_00_07[3], slf_op_00_07[2],
     slf_op_00_07[1], slf_op_00_07[0], slf_op_00_07[3],
     slf_op_00_07[2], slf_op_00_07[1], slf_op_00_07[0]}),
     .lft_op_06({slf_op_00_06[3], slf_op_00_06[2], slf_op_00_06[1],
     slf_op_00_06[0], slf_op_00_06[3], slf_op_00_06[2],
     slf_op_00_06[1], slf_op_00_06[0]}), .lft_op_05({slf_op_00_05[3],
     slf_op_00_05[2], slf_op_00_05[1], slf_op_00_05[0],
     slf_op_00_05[3], slf_op_00_05[2], slf_op_00_05[1],
     slf_op_00_05[0]}), .sp12_h_l_08(net1357[0:23]),
     .sp12_h_l_07(net1365[0:23]), .sp12_h_l_06(net1358[0:23]),
     .sp12_h_r_05(net988[0:23]), .sp12_h_r_06(net989[0:23]),
     .sp12_h_r_07(net990[0:23]), .sp12_h_r_08(net991[0:23]),
     .sp12_h_l_05(net1360[0:23]), .sp4_r_v_b_05(net993[0:47]),
     .sp4_r_v_b_06(net994[0:47]), .sp4_r_v_b_07(net995[0:47]),
     .sp4_r_v_b_08(net996[0:47]), .sp4_v_b_08(net997[0:47]),
     .sp4_v_b_07(net998[0:47]), .sp4_v_b_06(net999[0:47]),
     .sp4_v_b_05(net1000[0:47]), .pgate(pgate_l[143:16]),
     .reset_b(reset_b_l[143:16]), .wl(wl_l[143:16]),
     .sp12_v_t_08(sp12_v_t_01_08[23:0]), .tnr_op_08(tnr_op_01_08[7:0]),
     .top_op_08(top_op_01_08[7:0]), .tnl_op_08(tnl_op_01_08[7:0]),
     .sp4_v_t_08(sp4_v_t_01_08[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_01_08), .sp12_v_b_01(net1392[0:23]));
lt_1x8_bot_ice1f I_lt_col_t06 ( .glb_netwk_bot(net1402[0:7]),
     .rgt_op_03(rgt_op_06_03[7:0]), .slf_op_02(slf_op_06_02[7:0]),
     .rgt_op_02(rgt_op_06_02[7:0]), .rgt_op_01(rgt_op_06_01[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net1117[0:7]),
     .lft_op_03(net1107[0:7]), .lft_op_02(net1109[0:7]),
     .lft_op_01(net1428[0:7]), .rgt_op_04(rgt_op_06_04[7:0]),
     .carry_in(tiegnd_bl), .bnl_op_01({slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0],
     slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0]}), .slf_op_04(slf_op_06_04[7:0]),
     .slf_op_03(slf_op_06_03[7:0]), .slf_op_01(slf_op_06_01[7:0]),
     .sp4_h_l_04(net1230[0:47]), .carry_out(carry_out_06_08),
     .vdd_cntl(vdd_cntl_l[143:16]), .sp12_h_r_04(sp12_h_r_06_04[23:0]),
     .sp12_h_r_03(sp12_h_r_06_03[23:0]),
     .sp12_h_r_02(sp12_h_r_06_02[23:0]),
     .sp12_h_r_01(sp12_h_r_06_01[23:0]),
     .glb_netwk_col(clk_tree_drv_bl[7:0]), .sp4_v_b_01(net1425[0:47]),
     .sp4_r_v_b_04(sp4_r_v_b_06_04[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_06_03[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_06_02[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_06_01[47:0]),
     .sp4_h_r_04(sp4_h_r_06_04[47:0]),
     .sp4_h_r_03(sp4_h_r_06_03[47:0]),
     .sp4_h_r_02(sp4_h_r_06_02[47:0]),
     .sp4_h_r_01(sp4_h_r_06_01[47:0]), .sp4_h_l_03(net1231[0:47]),
     .sp4_h_l_02(net1232[0:47]), .sp4_h_l_01(net1233[0:47]),
     .bl(bl[329:276]), .bot_op_01({slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0], slf_op_06_00[3],
     slf_op_06_00[2], slf_op_06_00[1], slf_op_06_00[0]}),
     .sp12_h_l_01(net1223[0:23]), .sp12_h_l_02(net1222[0:23]),
     .sp12_h_l_03(net1221[0:23]), .sp12_h_l_04(net1220[0:23]),
     .sp4_v_b_04(net1226[0:47]), .sp4_v_b_03(net1227[0:47]),
     .sp4_v_b_02(net1228[0:47]), .bnr_op_01({bnr_op_06_01[3],
     bnr_op_06_01[2], bnr_op_06_01[1], bnr_op_06_01[0],
     bnr_op_06_01[3], bnr_op_06_01[2], bnr_op_06_01[1],
     bnr_op_06_01[0]}), .sp4_h_l_05(net1254[0:47]),
     .sp4_h_l_06(net1253[0:47]), .sp4_h_l_07(net1252[0:47]),
     .sp4_h_l_08(net1251[0:47]), .sp4_h_r_08(sp4_h_r_06_08[47:0]),
     .sp4_h_r_07(sp4_h_r_06_07[47:0]),
     .sp4_h_r_06(sp4_h_r_06_06[47:0]),
     .sp4_h_r_05(sp4_h_r_06_05[47:0]), .slf_op_05(slf_op_06_05[7:0]),
     .slf_op_06(slf_op_06_06[7:0]), .slf_op_07(slf_op_06_07[7:0]),
     .slf_op_08(slf_op_06_08[7:0]), .rgt_op_08(rgt_op_06_08[7:0]),
     .rgt_op_07(rgt_op_06_07[7:0]), .rgt_op_06(rgt_op_06_06[7:0]),
     .rgt_op_05(rgt_op_06_05[7:0]), .lft_op_08(slf_op_05_08[7:0]),
     .lft_op_07(net1166[0:7]), .lft_op_06(net1167[0:7]),
     .lft_op_05(net1168[0:7]), .sp12_h_l_08(net1273[0:23]),
     .sp12_h_l_07(net1272[0:23]), .sp12_h_l_06(net1271[0:23]),
     .sp12_h_r_05(sp12_h_r_06_05[23:0]),
     .sp12_h_r_06(sp12_h_r_06_06[23:0]),
     .sp12_h_r_07(sp12_h_r_06_07[23:0]),
     .sp12_h_r_08(sp12_h_r_06_08[23:0]), .sp12_h_l_05(net1270[0:23]),
     .sp4_r_v_b_05(sp4_r_v_b_06_05[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_06_06[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_06_07[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_06_08[47:0]), .sp4_v_b_08(net1278[0:47]),
     .sp4_v_b_07(net1277[0:47]), .sp4_v_b_06(net1276[0:47]),
     .sp4_v_b_05(net1275[0:47]), .pgate(pgate_l[143:16]),
     .reset_b(reset_b_l[143:16]), .wl(wl_l[143:16]),
     .sp12_v_t_08(sp12_v_t_06_08[23:0]), .tnr_op_08(tnr_op_06_08[7:0]),
     .top_op_08(top_op_06_08[7:0]), .tnl_op_08(tnl_op_06_08[7:0]),
     .sp4_v_t_08(sp4_v_t_06_08[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_06_08), .sp12_v_b_01(net1426[0:23]));
lt_1x8_bot_ice1f I_lt_col_t04 ( .glb_netwk_bot(net1404[0:7]),
     .rgt_op_03(net1107[0:7]), .slf_op_02(net801[0:7]),
     .rgt_op_02(net1109[0:7]), .rgt_op_01(net1428[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net834[0:7]), .lft_op_03(net824[0:7]),
     .lft_op_02(net826[0:7]), .lft_op_01(net1429[0:7]),
     .rgt_op_04(net1117[0:7]), .carry_in(tiegnd_bl),
     .bnl_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .slf_op_04(net799[0:7]),
     .slf_op_03(net800[0:7]), .slf_op_01(net1427[0:7]),
     .sp4_h_l_04(net820[0:47]), .carry_out(carry_out_04_08),
     .vdd_cntl(vdd_cntl_l[143:16]), .sp12_h_r_04(net1126[0:23]),
     .sp12_h_r_03(net1127[0:23]), .sp12_h_r_02(net1128[0:23]),
     .sp12_h_r_01(net1129[0:23]), .glb_netwk_col(clk_tree_drv_bl[7:0]),
     .sp4_v_b_01(net1433[0:47]), .sp4_r_v_b_04(net1132[0:47]),
     .sp4_r_v_b_03(net1133[0:47]), .sp4_r_v_b_02(net1134[0:47]),
     .sp4_r_v_b_01(net1421[0:47]), .sp4_h_r_04(net1136[0:47]),
     .sp4_h_r_03(net1137[0:47]), .sp4_h_r_02(net1138[0:47]),
     .sp4_h_r_01(net1139[0:47]), .sp4_h_l_03(net819[0:47]),
     .sp4_h_l_02(net818[0:47]), .sp4_h_l_01(net774[0:47]),
     .bl(bl[221:168]), .bot_op_01({slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0], slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0]}),
     .sp12_h_l_01(net768[0:23]), .sp12_h_l_02(net776[0:23]),
     .sp12_h_l_03(net732[0:23]), .sp12_h_l_04(net777[0:23]),
     .sp4_v_b_04(net756[0:47]), .sp4_v_b_03(net752[0:47]),
     .sp4_v_b_02(net763[0:47]), .bnr_op_01({slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0],
     slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0]}), .sp4_h_l_05(net821[0:47]),
     .sp4_h_l_06(net822[0:47]), .sp4_h_l_07(net823[0:47]),
     .sp4_h_l_08(net759[0:47]), .sp4_h_r_08(net1157[0:47]),
     .sp4_h_r_07(net1158[0:47]), .sp4_h_r_06(net1159[0:47]),
     .sp4_h_r_05(net1160[0:47]), .slf_op_05(net798[0:7]),
     .slf_op_06(net797[0:7]), .slf_op_07(net796[0:7]),
     .slf_op_08(slf_op_04_08[7:0]), .rgt_op_08(slf_op_05_08[7:0]),
     .rgt_op_07(net1166[0:7]), .rgt_op_06(net1167[0:7]),
     .rgt_op_05(net1168[0:7]), .lft_op_08(slf_op_03_08[7:0]),
     .lft_op_07(net884[0:7]), .lft_op_06(net885[0:7]),
     .lft_op_05(net886[0:7]), .sp12_h_l_08(net749[0:23]),
     .sp12_h_l_07(net744[0:23]), .sp12_h_l_06(net746[0:23]),
     .sp12_h_r_05(net1176[0:23]), .sp12_h_r_06(net1177[0:23]),
     .sp12_h_r_07(net1178[0:23]), .sp12_h_r_08(net1179[0:23]),
     .sp12_h_l_05(net748[0:23]), .sp4_r_v_b_05(net1181[0:47]),
     .sp4_r_v_b_06(net1182[0:47]), .sp4_r_v_b_07(net1183[0:47]),
     .sp4_r_v_b_08(net1184[0:47]), .sp4_v_b_08(net791[0:47]),
     .sp4_v_b_07(net792[0:47]), .sp4_v_b_06(net793[0:47]),
     .sp4_v_b_05(net760[0:47]), .pgate(pgate_l[143:16]),
     .reset_b(reset_b_l[143:16]), .wl(wl_l[143:16]),
     .sp12_v_t_08(sp12_v_t_04_08[23:0]), .tnr_op_08(tnr_op_04_08[7:0]),
     .top_op_08(top_op_04_08[7:0]), .tnl_op_08(tnl_op_04_08[7:0]),
     .sp4_v_t_08(sp4_v_t_04_08[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_04_08), .sp12_v_b_01(net1423[0:23]));
lt_1x8_bot_ice1f I_lt_col_t05 ( .glb_netwk_bot(net1403[0:7]),
     .rgt_op_03(slf_op_06_03[7:0]), .slf_op_02(net1109[0:7]),
     .rgt_op_02(slf_op_06_02[7:0]), .rgt_op_01(slf_op_06_01[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net799[0:7]),
     .lft_op_03(net800[0:7]), .lft_op_02(net801[0:7]),
     .lft_op_01(net1427[0:7]), .rgt_op_04(slf_op_06_04[7:0]),
     .carry_in(tiegnd_bl), .bnl_op_01({slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0],
     slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0]}), .slf_op_04(net1117[0:7]),
     .slf_op_03(net1107[0:7]), .slf_op_01(net1428[0:7]),
     .sp4_h_l_04(net1136[0:47]), .carry_out(carry_out_05_08),
     .vdd_cntl(vdd_cntl_l[143:16]), .sp12_h_r_04(net1220[0:23]),
     .sp12_h_r_03(net1221[0:23]), .sp12_h_r_02(net1222[0:23]),
     .sp12_h_r_01(net1223[0:23]), .glb_netwk_col(clk_tree_drv_bl[7:0]),
     .sp4_v_b_01(net1421[0:47]), .sp4_r_v_b_04(net1226[0:47]),
     .sp4_r_v_b_03(net1227[0:47]), .sp4_r_v_b_02(net1228[0:47]),
     .sp4_r_v_b_01(net1425[0:47]), .sp4_h_r_04(net1230[0:47]),
     .sp4_h_r_03(net1231[0:47]), .sp4_h_r_02(net1232[0:47]),
     .sp4_h_r_01(net1233[0:47]), .sp4_h_l_03(net1137[0:47]),
     .sp4_h_l_02(net1138[0:47]), .sp4_h_l_01(net1139[0:47]),
     .bl(bl[275:222]), .bot_op_01({slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0], slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0]}),
     .sp12_h_l_01(net1129[0:23]), .sp12_h_l_02(net1128[0:23]),
     .sp12_h_l_03(net1127[0:23]), .sp12_h_l_04(net1126[0:23]),
     .sp4_v_b_04(net1132[0:47]), .sp4_v_b_03(net1133[0:47]),
     .sp4_v_b_02(net1134[0:47]), .bnr_op_01({slf_op_06_00[3],
     slf_op_06_00[2], slf_op_06_00[1], slf_op_06_00[0],
     slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0]}), .sp4_h_l_05(net1160[0:47]),
     .sp4_h_l_06(net1159[0:47]), .sp4_h_l_07(net1158[0:47]),
     .sp4_h_l_08(net1157[0:47]), .sp4_h_r_08(net1251[0:47]),
     .sp4_h_r_07(net1252[0:47]), .sp4_h_r_06(net1253[0:47]),
     .sp4_h_r_05(net1254[0:47]), .slf_op_05(net1168[0:7]),
     .slf_op_06(net1167[0:7]), .slf_op_07(net1166[0:7]),
     .slf_op_08(slf_op_05_08[7:0]), .rgt_op_08(slf_op_06_08[7:0]),
     .rgt_op_07(slf_op_06_07[7:0]), .rgt_op_06(slf_op_06_06[7:0]),
     .rgt_op_05(slf_op_06_05[7:0]), .lft_op_08(slf_op_04_08[7:0]),
     .lft_op_07(net796[0:7]), .lft_op_06(net797[0:7]),
     .lft_op_05(net798[0:7]), .sp12_h_l_08(net1179[0:23]),
     .sp12_h_l_07(net1178[0:23]), .sp12_h_l_06(net1177[0:23]),
     .sp12_h_r_05(net1270[0:23]), .sp12_h_r_06(net1271[0:23]),
     .sp12_h_r_07(net1272[0:23]), .sp12_h_r_08(net1273[0:23]),
     .sp12_h_l_05(net1176[0:23]), .sp4_r_v_b_05(net1275[0:47]),
     .sp4_r_v_b_06(net1276[0:47]), .sp4_r_v_b_07(net1277[0:47]),
     .sp4_r_v_b_08(net1278[0:47]), .sp4_v_b_08(net1184[0:47]),
     .sp4_v_b_07(net1183[0:47]), .sp4_v_b_06(net1182[0:47]),
     .sp4_v_b_05(net1181[0:47]), .pgate(pgate_l[143:16]),
     .reset_b(reset_b_l[143:16]), .wl(wl_l[143:16]),
     .sp12_v_t_08(sp12_v_t_05_08[23:0]), .tnr_op_08(tnr_op_05_08[7:0]),
     .top_op_08(top_op_05_08[7:0]), .tnl_op_08(tnl_op_05_08[7:0]),
     .sp4_v_t_08(sp4_v_t_05_08[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_05_08), .sp12_v_b_01(net1445[0:23]));
clk_quad_buf_x8_ice8p I_clktree_quad_drv_tl ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));
clk_quad_buf_x8_ice8p I_clk_qtl_center ( .clko(clk_tree_drv_bl[7:0]),
     .clki(clk_center[7:0]));
tielo I450 ( .tielo(tiegnd_bl));
pinlatbuf12p I_pinlatbuf12p_b ( .pad_in(padin_b_l[10]),
     .icegate(hold_l_b), .cbit(cf_b_l[135]), .cout(padinlat_b_l[10]),
     .prog(prog));
io_lft_bot_1x8_ice1f I_io_bot_00 ( .padeb(padeb_l_b[11:0]),
     .pado(pado_l_b[11:0]), .padin(padin_l_b[11:0]), .fo_fb(fo_fb),
     .fo_dlyadj(fo_dlyadj[2:0]), .fo_ref(fo_ref), .shift(net1310),
     .bs_en(net1311), .mode(net1312), .sdi(net1313), .hiz_b(net1314),
     .prog(prog), .hold(hold_l_b), .update(net1317), .r(net1318),
     .SP4_h_l_05(net1319[0:47]), .slf_op_05(slf_op_00_05[3:0]),
     .slf_op_01(slf_op_00_01[3:0]), .slf_op_06(slf_op_00_06[3:0]),
     .slf_op_02(slf_op_00_02[3:0]), .sdo(net1324), .bl({bl[0], bl[1],
     bl[2], bl[3], bl[4], bl[5], bl[6], bl[7], bl[8], bl[9], bl[10],
     bl[11], bl[12], bl[13], bl[14], bl[15], bl[16], bl[17]}),
     .sp4_v_b_00_01(net1326[0:15]), .tclk(net1327),
     .reset_b(reset_b_l[143:16]), .rgt_op_02(net1329[0:7]),
     .SP4_h_l_06(net1330[0:47]), .sp4_v_t_08(sp4_v_t_00_08[15:0]),
     .slf_op_04(slf_op_00_04[3:0]), .slf_op_03(slf_op_00_03[3:0]),
     .slf_op_07(slf_op_00_07[3:0]), .slf_op_08(slf_op_00_08[3:0]),
     .SP4_h_l_08(net1336[0:47]), .SP4_h_l_07(net1337[0:47]),
     .SP4_h_l_03(net1338[0:47]), .SP4_h_l_04(net1339[0:47]),
     .SP4_h_l_02(net1340[0:47]), .SP4_h_l_01(net1341[0:47]),
     .rgt_op_07(net1342[0:7]), .rgt_op_06(net1343[0:7]),
     .rgt_op_05(net1344[0:7]), .rgt_op_03(net1345[0:7]),
     .rgt_op_01(net1436[0:7]), .rgt_op_08(slf_op_01_08[7:0]),
     .pgate(pgate_l[143:16]), .vdd_cntl(vdd_cntl_l[143:16]),
     .cf_l(cf_l[191:0]), .wl(wl_l[143:16]),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .tclk_o(net1353), .ceb(net1354), .SP12_h_l_02(net1355[0:23]),
     .SP12_h_l_04(net1356[0:23]), .SP12_h_l_08(net1357[0:23]),
     .SP12_h_l_06(net1358[0:23]), .glb_netwk_col(clk_tree_drv_bl[7:0]),
     .SP12_h_l_05(net1360[0:23]), .SP12_h_l_01(net1361[0:23]),
     .fabric_out_07(fo_00_07), .SP12_h_l_03(net1363[0:23]),
     .fabric_out_08(fo_00_08), .SP12_h_l_07(net1365[0:23]),
     .last_rsr(last_rsr[0]), .rgt_op_04(net1367[0:7]),
     .bnr_op_00_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}),
     .tnr_op_08(tnr_op_00_08[7:0]));
io_bot_lft_1x6_ice1f I_preio_bot_l ( bs_en_o, ceb_o, cf_b_l[143:0],
     net1480, net1478, fo_bypass, fo_reset, fo_sck, fo_sdi, hiz_b_o,
     mode_o, padeb_b_l[10:0], padeb_b_l[12], pado_b_l[10:0],
     pado_b_l[12], r_o, sdo, shift_o, slf_op_01_00[3:0],
     slf_op_02_00[3:0], slf_op_03_00[3:0], slf_op_04_00[3:0],
     slf_op_05_00[3:0], slf_op_06_00[3:0], tclk_o, update_o, bl[71:18],
     bl[125:72], bl[167:126], bl[221:168], bl[275:222], bl[329:276],
     net1326[0:15], sp4_h_r_06_00[15:0], net1456[0:47], net1430[0:47],
     net1431[0:47], net1433[0:47], net1421[0:47], net1425[0:47],
     net1392[0:23], net1409[0:23], net1432[0:23], net1423[0:23],
     net1445[0:23], net1426[0:23], {slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0], slf_op_00_01[3],
     slf_op_00_01[2], slf_op_00_01[1], slf_op_00_01[0]}, net1311,
     net1354, net1407[0:7], net1406[0:7], net1405[0:7], net1404[0:7],
     net1403[0:7], net1402[0:7], net1314, hold_b_l, net1436[0:7],
     net1438[0:7], net1429[0:7], net1427[0:7], net1428[0:7],
     slf_op_06_01[7:0], net1312, padin_b_l[10:0], padin_b_l[12],
     {pgate_l[1], pgate_l[0], pgate_l[2], pgate_l[3], pgate_l[5],
     pgate_l[4], pgate_l[6], pgate_l[7], pgate_l[9], pgate_l[8],
     pgate_l[10], pgate_l[11], pgate_l[13], pgate_l[12], pgate_l[14],
     pgate_l[15]}, prog, net1318, {reset_b_l[1], reset_b_l[0],
     reset_b_l[2], reset_b_l[3], reset_b_l[5], reset_b_l[4],
     reset_b_l[6], reset_b_l[7], reset_b_l[9], reset_b_l[8],
     reset_b_l[10], reset_b_l[11], reset_b_l[13], reset_b_l[12],
     reset_b_l[14], reset_b_l[15]}, net1324, net1310, net1353,
     rgt_op_06_01[7:0], net1317, {vdd_cntl_l[1], vdd_cntl_l[0],
     vdd_cntl_l[2], vdd_cntl_l[3], vdd_cntl_l[5], vdd_cntl_l[4],
     vdd_cntl_l[6], vdd_cntl_l[7], vdd_cntl_l[9], vdd_cntl_l[8],
     vdd_cntl_l[10], vdd_cntl_l[11], vdd_cntl_l[13], vdd_cntl_l[12],
     vdd_cntl_l[14], vdd_cntl_l[15]}, {wl_l[1], wl_l[0], wl_l[2],
     wl_l[3], wl_l[5], wl_l[4], wl_l[6], wl_l[7], wl_l[9], wl_l[8],
     wl_l[10], wl_l[11], wl_l[13], wl_l[12], wl_l[14], wl_l[15]});
scan_buf_ice8p I_scanbuf_8p_ml ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net1317), .tclk_o(net1327), .shift_o(net1310),
     .sdo(net1313), .r_o(net1318), .mode_o(net1312), .hiz_b_o(net1314),
     .ceb_o(net1354), .bs_en_o(net1311));
fabric_buf_ice8p I785 ( .f_in(net1478), .f_out(fabric_out_06_00));
fabric_buf_ice8p I786 ( .f_in(net1480), .f_out(fabric_out_05_00));
fabric_buf_ice8p I_fabric_buf_8p_0016 ( .f_in(fo_00_08),
     .f_out(fabric_out_00_08));
fabric_buf_ice8p I_fabric_buf_8p_0015 ( .f_in(fo_00_07),
     .f_out(fabric_out_00_07));
fabric_buf_ice8p I_fabric_buf8p_25 ( .f_in(padinlat_l_b[11]),
     .f_out(padin_00_08));
fabric_buf_ice8p I784 ( .f_in(padinlat_b_l[10]), .f_out(padin_06_00));
pinlatbuf12p_1 I_pinlatbuf12p ( .pad_in(padin_l_b[11]),
     .icegate(hold_l_b), .cbit(cf_l[183]), .cout(padinlat_l_b[11]),
     .prog(prog));

endmodule
// Library - leafcell, Cell - bram_bufferx2e, View - schematic
// LAST TIME SAVED: May 13 10:18:51 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module bram_bufferx2e ( out, en, in );
output  out;

input  en, in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I391 ( .A(net7), .Y(out));
nand2 I193 ( .A(en), .Y(net7), .B(in));

endmodule
// Library - leafcell, Cell - bram_bank_logic_bot, View - schematic
// LAST TIME SAVED: Jul  8 10:16:10 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module bram_bank_logic_bot ( bm_sclkrw_o, bm_sdo_o, bm_sweb_o,
     bm_banksel_i, bm_sclk_i, bm_sclkrw_i, bm_sdo_i, bm_sweb_i );

input  bm_sclk_i, bm_sclkrw_i, bm_sweb_i;

output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sclkrw_o;

input [1:0]  bm_banksel_i;
input [1:0]  bm_sdo_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net26;

wire  [0:1]  net25;



ml_dff I52_1_ ( .R(net020), .D(bm_sdo_i[1]), .CLK(bm_sclk_i),
     .QN(net25[0]), .Q(net26[1]));
ml_dff I52_0_ ( .R(net020), .D(bm_sdo_i[0]), .CLK(bm_sclk_i),
     .QN(net25[1]), .Q(net26[0]));
bram_bufferx16_2inv I51_1_ ( .in(net26[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I51_0_ ( .in(net26[0]), .out(bm_sdo_o[0]));
bram_bufferx2e I54_1_ ( .in(bm_sweb_i), .en(bm_banksel_i[1]),
     .out(bm_sweb_o[1]));
bram_bufferx2e I54_0_ ( .in(bm_sweb_i), .en(bm_banksel_i[0]),
     .out(bm_sweb_o[0]));
bram_bufferx2e I48_1_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[1]),
     .out(bm_sclkrw_o[1]));
bram_bufferx2e I48_0_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[0]),
     .out(bm_sclkrw_o[0]));
tielo I55 ( .tielo(net020));

endmodule
// Library - leafcell, Cell - bram_icg, View - schematic
// LAST TIME SAVED: Oct 22 11:07:43 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module bram_icg ( clkout, clk, en );
output  clkout;

input  clk, en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I391 ( .A(net014), .Y(clkout));
inv I6 ( .A(net023), .Y(net027));
inv I4 ( .A(cn), .Y(c));
inv I3 ( .A(clk), .Y(cn));
nand2 I193 ( .A(net027), .Y(net014), .B(c));
inv_tri_2 I7 ( .Tb(cn), .T(c), .A(net027), .Y(net023));
inv_tri_2 I5 ( .Tb(c), .T(cn), .A(en), .Y(net023));

endmodule
// Library - leafcell, Cell - bram_hbuffer_dff_2xbank, View - schematic
// LAST TIME SAVED: Oct 22 09:16:56 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module bram_hbuffer_dff_2xbank ( bm_banksel_o, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclkrw_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [3:0]  bm_sdi_o;
output [3:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [3:0]  bm_banksel_o;
output [1:0]  bm_sclk_o;

input [3:0]  bm_sdi_i;
input [7:0]  bm_sa_i;
input [3:0]  bm_sdo_i;
input [3:0]  bm_banksel_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net103;

wire  [0:3]  net102;



ml_dff I48_3_ ( .R(net057), .D(bm_sdo_i[3]), .CLK(bm_sclk_i),
     .QN(net102[0]), .Q(net103[0]));
ml_dff I48_2_ ( .R(net057), .D(bm_sdo_i[2]), .CLK(bm_sclk_i),
     .QN(net102[1]), .Q(net103[1]));
ml_dff I48_1_ ( .R(net057), .D(bm_sdo_i[1]), .CLK(bm_sclk_i),
     .QN(net102[2]), .Q(net103[2]));
ml_dff I48_0_ ( .R(net057), .D(bm_sdo_i[0]), .CLK(bm_sclk_i),
     .QN(net102[3]), .Q(net103[3]));
nor2 I20 ( .A(bm_banksel_i[2]), .B(bm_banksel_i[3]), .Y(net67));
nor2 I49 ( .A(bm_banksel_i[0]), .B(bm_banksel_i[1]), .Y(net70));
inv I21 ( .A(net67), .Y(net72));
inv I17 ( .A(net70), .Y(net74));
tielo I23 ( .tielo(net057));
bram_icg I47 ( .en(net74), .clk(bm_sclk_i), .clkout(net61));
bram_icg I19 ( .en(net72), .clk(bm_sclk_i), .clkout(net64));
bram_bufferx16_2inv I16_3_ ( .in(net103[0]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I16_2_ ( .in(net103[1]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I16_1_ ( .in(net103[2]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I16_0_ ( .in(net103[3]), .out(bm_sdo_o[0]));
bram_bufferx4 I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx4 I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx4 I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx4 I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx4 I22 ( .in(net64), .out(bm_sclk_o[1]));
bram_bufferx4 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx4 I13_3_ ( .in(bm_banksel_i[3]), .out(bm_banksel_o[3]));
bram_bufferx4 I13_2_ ( .in(bm_banksel_i[2]), .out(bm_banksel_o[2]));
bram_bufferx4 I13_1_ ( .in(bm_banksel_i[1]), .out(bm_banksel_o[1]));
bram_bufferx4 I13_0_ ( .in(bm_banksel_i[0]), .out(bm_banksel_o[0]));
bram_bufferx4 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx4 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx4 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx4 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx4 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx4 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx4 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx4 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx4 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx4 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx4 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx4 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx4 I18 ( .in(net61), .out(bm_sclk_o[0]));
bram_bufferx4 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_hbuffer_1xbank, View - schematic
// LAST TIME SAVED: Jun 11 17:38:23 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module bram_hbuffer_1xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [1:0]  bm_banksel_o;
output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;

input [1:0]  bm_sdi_i;
input [1:0]  bm_sdo_i;
input [1:0]  bm_banksel_i;
input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - clkmux4to1, View - schematic
// LAST TIME SAVED: Jun 30 10:55:11 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module clkmux4to1 ( mout, cbit, .cdsNet0(min[0]), .cdsNet0(min[1]),
     .cdsNet0(min[2]), .cdsNet0(min[3]) );
output  mout;


input [3:0]  min;
input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cbit_b;



txgate_hvt I4 ( .in(net_2_0), .out(net52), .pp(cbit[1]),
     .nn(cbit_b[1]));
txgate_hvt I3 ( .in(net_2_1), .out(net52), .pp(cbit_b[1]),
     .nn(cbit[1]));
txgate_hvt I6 ( .in(min[2]), .out(net_2_1), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I5 ( .in(min[3]), .out(net_2_1), .pp(cbit_b[0]),
     .nn(cbit[0]));
txgate_hvt Itg20 ( .in(min[0]), .out(net_2_0), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I7 ( .in(min[1]), .out(net_2_0), .pp(cbit_b[0]),
     .nn(cbit[0]));
inv_hvt I2 ( .A(net046), .Y(mout));
inv_hvt I1_1_ ( .A(cbit[1]), .Y(cbit_b[1]));
inv_hvt I1_0_ ( .A(cbit[0]), .Y(cbit_b[0]));
inv_hvt I0 ( .A(net52), .Y(net046));

endmodule
// Library - ice1chip, Cell - quad_x4_ice1, View - schematic
// LAST TIME SAVED: May  3 11:40:33 2011
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module quad_x4_ice1 ( bm_sdo_o[3:0], cf_b[287:0], cf_l[383:0],
     cf_r[383:0], cf_t[287:0], fabric_out_05_00_bicegate,
     fabric_out_06_00, fabric_out_07_00, fabric_out_12_00_wb,
     fabric_out_13_01, fabric_out_13_02, fo_bypass, fo_dlyadj[7:0],
     fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, padeb_b[23:0],
     padeb_l[23:0], padeb_r[24:0], padeb_t[23:0], pado_b[23:0],
     pado_l[23:0], pado_r[24:0], pado_t[23:0], sdo_pad,
     spi_ss_in_bbank[4:0], tck_pad, tdi_pad, tms_pad, bl_bot[663:0],
     bl_top[663:0], bm_banksel_i[3:0], bm_init_i, bm_rcapmux_en_i,
     bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i, bm_sdi_i[3:0], bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb, end_of_startup,
     gclk_l2clktv[1:0], gclk_r2clktv[1:0], hiz_b,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[0],
     last_rsr[1], last_rsr[2], last_rsr[3], md_spi_b, mode,
     mux_jtag_sel_b, padin_b[23:0], padin_l[23:0], padin_r[24:0],
     padin_t[23:0], pgate_l[287:0], pgate_r[287:0], pll_lock_out,
     pll_sdo, prog, purst, r, reset_b_l[287:0], reset_b_r[287:0],
     sdi_pad, sdo_enable, shift, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk, totdopad, trstb_pad, update, vdd_cntl_l[287:0],
     vdd_cntl_r[287:0], wl_l[287:0], wl_r[287:0] );
output  fabric_out_05_00_bicegate, fabric_out_06_00, fabric_out_07_00,
     fabric_out_12_00_wb, fabric_out_13_01, fabric_out_13_02,
     fo_bypass, fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, sdo_pad,
     tck_pad, tdi_pad, tms_pad;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb, end_of_startup, hiz_b,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode, mux_jtag_sel_b, pll_lock_out, pll_sdo, prog, purst, r,
     sdi_pad, sdo_enable, shift, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk, totdopad, trstb_pad, update;

output [4:0]  spi_ss_in_bbank;
output [3:0]  bm_sdo_o;
output [23:0]  pado_l;
output [23:0]  padeb_l;
output [383:0]  cf_l;
output [23:0]  pado_t;
output [383:0]  cf_r;
output [24:0]  padeb_r;
output [23:0]  padeb_b;
output [23:0]  padeb_t;
output [287:0]  cf_t;
output [287:0]  cf_b;
output [7:0]  fo_dlyadj;
output [23:0]  pado_b;
output [24:0]  pado_r;

inout [663:0]  bl_bot;
inout [663:0]  bl_top;

input [3:0]  bm_sdi_i;
input [7:0]  bm_sa_i;
input [1:0]  gclk_r2clktv;
input [3:0]  bm_banksel_i;
input [287:0]  pgate_l;
input [23:0]  padin_l;
input [287:0]  pgate_r;
input [287:0]  vdd_cntl_r;
input [287:0]  reset_b_r;
input [287:0]  wl_r;
input [1:0]  gclk_l2clktv;
input [23:0]  padin_b;
input [0:3]  last_rsr;
input [287:0]  reset_b_l;
input [23:0]  padin_t;
input [24:0]  padin_r;
input [287:0]  wl_l;
input [287:0]  vdd_cntl_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  slf_op_07_13;

wire  [7:0]  slf_op_07_14;

wire  [0:23]  net1208;

wire  [0:23]  net983;

wire  [0:47]  net816;

wire  [3:0]  slf_op_06_17;

wire  [0:23]  net984;

wire  [0:23]  net1171;

wire  [0:23]  net1209;

wire  [0:7]  net995;

wire  [0:15]  net818;

wire  [0:23]  net1103;

wire  [7:0]  slf_op_07_11;

wire  [0:23]  net777;

wire  [7:0]  slf_op_01_09;

wire  [0:47]  net1225;

wire  [0:23]  net772;

wire  [0:47]  net1220;

wire  [0:23]  net771;

wire  [0:23]  net1198;

wire  [7:0]  slf_op_12_09;

wire  [0:10]  net1046;

wire  [0:1]  net1147;

wire  [7:0]  slf_op_08_09;

wire  [0:47]  net811;

wire  [0:47]  net1165;

wire  [0:47]  net1213;

wire  [0:47]  net849;

wire  [7:0]  slf_op_09_09;

wire  [7:0]  slf_op_07_08;

wire  [0:47]  net1218;

wire  [0:47]  net1001;

wire  [0:7]  net1190;

wire  [7:0]  slf_op_07_05;

wire  [0:47]  net1215;

wire  [0:23]  net985;

wire  [0:47]  net1224;

wire  [7:0]  slf_op_06_08;

wire  [0:23]  net1231;

wire  [0:47]  net1219;

wire  [0:23]  net986;

wire  [7:0]  slf_op_06_05;

wire  [0:47]  net1227;

wire  [0:23]  net1205;

wire  [7:0]  slf_op_06_06;

wire  [0:47]  net1115;

wire  [7:0]  slf_op_07_16;

wire  [0:7]  net1149;

wire  [0:47]  net1223;

wire  [7:0]  slf_op_04_08;

wire  [7:0]  slf_op_01_08;

wire  [0:47]  net921;

wire  [0:47]  net1212;

wire  [0:23]  net1222;

wire  [1:0]  bm_sweb_b2_o;

wire  [0:47]  net1242;

wire  [0:47]  net1228;

wire  [3:0]  slf_op_07_00;

wire  [0:47]  net998;

wire  [0:47]  net812;

wire  [0:1]  net1275;

wire  [1:0]  bm_sdo_b1_o;

wire  [0:23]  net773;

wire  [0:23]  net1206;

wire  [0:47]  net819;

wire  [7:0]  slf_op_07_15;

wire  [0:23]  net1170;

wire  [7:0]  slf_op_08_08;

wire  [7:0]  slf_op_07_12;

wire  [7:0]  slf_op_02_08;

wire  [0:23]  net1207;

wire  [7:0]  slf_op_06_11;

wire  [7:0]  slf_op_07_06;

wire  [0:47]  net820;

wire  [7:0]  slf_op_07_07;

wire  [7:0]  slf_op_04_09;

wire  [0:23]  net776;

wire  [0:47]  net1200;

wire  [7:0]  slf_op_02_09;

wire  [7:0]  slf_op_06_07;

wire  [7:0]  slf_op_06_03;

wire  [7:0]  slf_op_06_02;

wire  [7:0]  slf_op_07_01;

wire  [0:1]  net1146;

wire  [7:0]  slf_op_11_08;

wire  [7:0]  slf_op_07_03;

wire  [1:0]  bm_bank10_banksel_o;

wire  [7:0]  bm_bank30_sa_o;

wire  [7:0]  slf_op_03_09;

wire  [0:47]  net824;

wire  [0:47]  net1000;

wire  [0:23]  net774;

wire  [0:10]  net1232;

wire  [0:1]  net952;

wire  [7:0]  slf_op_05_08;

wire  [3:0]  slf_op_07_17;

wire  [0:47]  net814;

wire  [0:10]  net1071;

wire  [0:47]  net1221;

wire  [0:23]  net1195;

wire  [0:47]  net1241;

wire  [0:47]  net815;

wire  [7:0]  slf_op_06_14;

wire  [7:0]  slf_op_06_01;

wire  [7:0]  slf_op_05_09;

wire  [0:47]  net1217;

wire  [0:47]  net822;

wire  [7:0]  slf_op_06_16;

wire  [7:0]  slf_op_06_10;

wire  [7:0]  slf_op_03_08;

wire  [7:0]  slf_op_10_09;

wire  [0:47]  net848;

wire  [1:0]  bm_sdo_b0_o;

wire  [0:15]  net1250;

wire  [3:0]  slf_op_13_09;

wire  [0:47]  net810;

wire  [7:0]  gclk;

wire  [7:0]  slf_op_06_12;

wire  [1:0]  bm_sdo_b3_o;

wire  [0:47]  net813;

wire  [3:0]  slf_op_06_00;

wire  [1:0]  bm_sclkrw_b0_o;

wire  [1:0]  bm_bank30_sclk_o;

wire  [7:0]  slf_op_07_10;

wire  [0:47]  net1216;

wire  [1:0]  bm_sweb_b0_o;

wire  [3:0]  slf_op_00_08;

wire  [0:23]  net1197;

wire  [7:0]  slf_op_09_08;

wire  [1:0]  bm_sdi_b0_o;

wire  [7:0]  slf_op_12_08;

wire  [0:47]  net967;

wire  [7:0]  slf_op_06_15;

wire  [0:47]  net1214;

wire  [0:23]  net982;

wire  [7:0]  slf_op_06_04;

wire  [0:47]  net823;

wire  [0:23]  net775;

wire  [1:0]  bm_sclkrw_b2_o;

wire  [0:23]  net770;

wire  [0:47]  net1226;

wire  [1:0]  bm_sdi_b2_o;

wire  [0:47]  net999;

wire  [7:0]  slf_op_07_04;

wire  [3:0]  bm_bank30_sdi_o;

wire  [0:23]  net1196;

wire  [7:0]  slf_op_11_09;

wire  [7:0]  slf_op_07_02;

wire  [7:0]  slf_op_06_13;

wire  [0:47]  net821;

wire  [0:47]  net1199;

wire  [7:0]  slf_op_07_09;

wire  [3:0]  bm_bank30_sdo_i;

wire  [0:23]  net981;

wire  [0:15]  net911;

wire  [7:0]  slf_op_06_09;

wire  [0:1]  net1143;

wire  [3:0]  slf_op_00_09;

wire  [0:1]  net948;

wire  [0:10]  net1138;

wire  [7:0]  slf_op_10_08;

wire  [3:0]  bm_bank30_banksel_o;

wire  [0:15]  net1154;

wire  [3:0]  slf_op_13_08;

wire  [1:0]  bm_sdo_b2_o;



ice1f_cram_row142col4 I64 ( .vdd_cntl_l(vdd_cntl_l[287:146]),
     .bl(bl_top[333:330]), .vdd_cntl_r(vdd_cntl_r[287:146]),
     .reset_r(reset_b_r[287:146]), .pgate_r(pgate_r[287:146]),
     .reset_l(reset_b_l[287:146]), .pgate_l(pgate_l[287:146]),
     .wl_r(wl_r[287:146]), .wl_l(wl_l[287:146]));
ice1f_cram_row142col4 I65 ( .vdd_cntl_l(vdd_cntl_l[141:0]),
     .bl(bl_bot[333:330]), .vdd_cntl_r(vdd_cntl_r[141:0]),
     .reset_r(reset_b_r[141:0]), .pgate_r(pgate_r[141:0]),
     .reset_l(reset_b_l[141:0]), .pgate_l(pgate_l[141:0]),
     .wl_r(wl_r[141:0]), .wl_l(wl_l[141:0]));
bram_sdo_reg I_bm_sdo_reg_b0 ( .do(bm_sdo_b0_o_0), .di(bm_sdo_b0_o[0]),
     .clk(bm_sck_b0_i), .tielo(net1262));
bram_sdo_reg I_bm_sdo_reg_b2 ( .do(bm_sdo_b2_o_0), .di(bm_sdo_b2_o[0]),
     .clk(bm_bank30_sclk_o[1]), .tielo(net1256));
bram_sdo_reg I_bm_sdo_reg_b3 ( .do(bm_sdo_b3_o_0), .di(bm_sdo_b3_o[0]),
     .clk(bm_sck_b2_o), .tielo(tielo_4bram3));
bram_sdo_reg I_bm_sdo_reg_b1 ( .do(bm_sdo_b1_o_0), .di(bm_sdo_b1_o[0]),
     .clk(bm_sck_b0_o), .tielo(tielo_4bram1));
clk_mux2to1_ice8p I_glb_ck_tree_top5432 ( .bl(bl_top[333:330]),
     .gnet(gclk[5:2]), .reset_r(reset_b_r[145:144]),
     .min0({padin_0717a_ck, fabric_out_13_09}), .min1({gclk_r2clktv[0],
     fabric_out_00_09}), .min2({padin_0009a_ck, fabric_out_06_17}),
     .min3({padin_1309a_ck, gclk_l2clktv[1]}),
     .pgate_l(pgate_l[145:144]), .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[145:144]), .reset_l(reset_b_l[145:144]),
     .wl_l(wl_l[145:144]), .wl_r(wl_r[145:144]),
     .pgate_r(pgate_r[145:144]), .vdd_cntl_r(vdd_cntl_r[145:144]));
clk_mux2to1_ice8p I_glb_ck_tree_bot7610 ( .bl(bl_bot[333:330]),
     .gnet({gclk[7], gclk[6], gclk[1], gclk[0]}),
     .reset_r(reset_b_r[143:142]), .min0({padin_1308b_ck,
     gclk_r2clktv[1]}), .min1({padin_0008b_ck, fabric_out_07_17}),
     .min2({gclk_l2clktv[0], fabric_out_00_08}), .min3({padin_0617b_ck,
     fabric_out_13_08}), .pgate_l(pgate_l[143:142]), .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[143:142]), .reset_l(reset_b_l[143:142]),
     .wl_l(wl_l[143:142]), .wl_r(wl_r[143:142]),
     .pgate_r(pgate_r[143:142]), .vdd_cntl_r(vdd_cntl_r[143:142]));
quad_tr_ice1 i_tr_quad ( .update_i(net957),
     .sp4_h_l_07_17(net818[0:15]), .lc_bot_07_09(n_inter_07),
     .bm_sdi_i({tielo_4bram3, bm_sdi_b2_o[1]}),
     .lc_bot_09_09(n_inter_09), .tclk_i(tclkio_mr), .shift_i(net969),
     .sdi(sdio_mr), .r_i(net971), .purst(purst), .prog(prog),
     .mode_i(net974), .slf_op_07_16(slf_op_07_16[7:0]),
     .slf_op_07_15(slf_op_07_15[7:0]),
     .slf_op_07_14(slf_op_07_14[7:0]),
     .slf_op_07_13(slf_op_07_13[7:0]),
     .slf_op_07_12(slf_op_07_12[7:0]),
     .slf_op_07_11(slf_op_07_11[7:0]),
     .slf_op_07_10(slf_op_07_10[7:0]),
     .slf_op_07_09(slf_op_07_09[7:0]),
     .hold_t_r(fabric_out_08_17_ticegate),
     .hold_r_t(fabric_out_13_10_ricegate), .hiz_b_i(net975),
     .glb_in(gclk[7:0]), .ceb_i(net980),
     .carry_in_12_09(carry_io_12_0809),
     .carry_in_11_09(carry_io_11_0809),
     .carry_in_09_09(carry_io_09_0809),
     .carry_in_08_09(carry_io_08_0809), .bs_en_i(net987),
     .sp4_v_b_12_09(net999[0:47]), .sp4_v_b_11_09(net1000[0:47]),
     .sp4_v_b_10_09(net1001[0:47]), .sp4_v_b_09_09(net998[0:47]),
     .sp4_v_b_08_09(net967[0:47]), .bnl_op_12_09(slf_op_11_08[7:0]),
     .bnl_op_11_09(slf_op_10_08[7:0]),
     .bnl_op_10_09(slf_op_09_08[7:0]),
     .bnl_op_09_09(slf_op_08_08[7:0]),
     .slf_op_08_09(slf_op_08_09[7:0]),
     .bot_op_12_09(slf_op_12_08[7:0]),
     .bot_op_11_09(slf_op_11_08[7:0]),
     .bot_op_10_09(slf_op_10_08[7:0]),
     .bot_op_09_09(slf_op_09_08[7:0]),
     .bot_op_08_09(slf_op_08_08[7:0]),
     .bot_op_07_09(slf_op_07_08[7:0]), .update_o(net863),
     .tclk_o(tclkio_mt), .bm_wdummymux_en_i(net988),
     .lft_op_07_09(slf_op_06_09[7:0]),
     .carry_in_07_09(carry_io_07_0809),
     .lft_op_07_16(slf_op_06_16[7:0]),
     .slf_op_13_09(slf_op_13_09[3:0]),
     .fabric_out_13_10(fabric_out_13_10_ricegate),
     .slf_op_12_09(slf_op_12_09[7:0]),
     .slf_op_11_09(slf_op_11_09[7:0]),
     .slf_op_10_09(slf_op_10_09[7:0]),
     .slf_op_09_09(slf_op_09_09[7:0]),
     .slf_op_07_17(slf_op_07_17[3:0]), .sp12_h_l_07_16(net770[0:23]),
     .sp12_h_l_07_15(net771[0:23]), .sp12_h_l_07_14(net772[0:23]),
     .sp12_h_l_07_13(net773[0:23]), .sp12_h_l_07_12(net774[0:23]),
     .sp12_h_l_07_11(net775[0:23]), .sp12_h_l_07_10(net776[0:23]),
     .sp12_v_b_07_09(net986[0:23]), .shift_o(net866), .sdo(sdio_mt),
     .r_o(net876), .padin_13_09a(padin_1309a_ck),
     .fabric_out_07_17(fabric_out_07_17),
     .padin_07_17a(padin_0717a_ck), .mode_o(net880), .hiz_b_o(net883),
     .cf_r(cf_r[383:192]), .ceb_o(net858), .bs_en_o(net888),
     .bnr_op_12_09({slf_op_13_08[3], slf_op_13_08[2], slf_op_13_08[1],
     slf_op_13_08[0], slf_op_13_08[3], slf_op_13_08[2],
     slf_op_13_08[1], slf_op_13_08[0]}),
     .bnr_op_11_09(slf_op_12_08[7:0]),
     .bnr_op_10_09(slf_op_11_08[7:0]),
     .bnr_op_09_09(slf_op_10_08[7:0]),
     .bnr_op_08_09(slf_op_09_08[7:0]),
     .bnr_op_07_09(slf_op_08_08[7:0]), .sp4_v_b_07_16(net810[0:47]),
     .sp4_v_b_07_15(net811[0:47]), .sp4_v_b_07_14(net812[0:47]),
     .sp4_v_b_07_13(net813[0:47]), .sp4_v_b_07_12(net814[0:47]),
     .sp4_v_b_07_11(net815[0:47]), .sp4_v_b_07_10(net816[0:47]),
     .sp4_v_b_07_09(net921[0:47]), .sp12_v_b_12_09(net981[0:23]),
     .sp12_v_b_11_09(net982[0:23]), .sp12_v_b_10_09(net983[0:23]),
     .sp12_v_b_09_09(net984[0:23]), .sp12_v_b_08_09(net985[0:23]),
     .fabric_out_13_09(fabric_out_13_09), .pado_t_r(pado_t[23:12]),
     .sp4_h_l_07_16(net819[0:47]), .sp4_h_l_07_15(net820[0:47]),
     .sp4_h_l_07_14(net821[0:47]), .sp4_h_l_07_13(net822[0:47]),
     .sp4_h_l_07_12(net823[0:47]), .sp4_h_l_07_11(net824[0:47]),
     .sp4_h_l_07_10(net849[0:47]), .bnl_op_08_09(slf_op_07_08[7:0]),
     .bnl_op_13_09(slf_op_12_08[7:0]),
     .lft_op_07_15(slf_op_06_15[7:0]),
     .lft_op_07_14(slf_op_06_14[7:0]),
     .lft_op_07_13(slf_op_06_13[7:0]),
     .lft_op_07_12(slf_op_06_12[7:0]),
     .lft_op_07_11(slf_op_06_11[7:0]),
     .lft_op_07_10(slf_op_06_10[7:0]),
     .vdd_cntl_r(vdd_cntl_r[287:144]), .wl_r(wl_r[287:144]),
     .reset_b_r(reset_b_r[287:144]), .pado_r(pado_r[24:13]),
     .padeb_r(padeb_r[24:13]), .padin_r(padin_r[24:13]),
     .bnl_op_07_09(slf_op_06_08[7:0]), .sp4_h_l_07_09(net848[0:47]),
     .sp12_h_l_07_09(net777[0:23]), .lc_bot_11_09(n_inter_11),
     .lc_bot_12_09(n_inter_12), .sp4_h_r_13_09(net911[0:15]),
     .bl(bl_top[663:334]), .pgate_r(pgate_r[287:144]),
     .cf_t(cf_t[287:144]), .lc_bot_08_09(n_inter_08),
     .bm_aa_2bot(net1071[0:10]), .bm_ab_2bot(net1046[0:10]),
     .bm_init_i(net997), .bm_rcapmux_en_i(net996),
     .bm_sa_i(net995[0:7]), .bm_sclk_i(bm_sck_b2_o),
     .bm_sclkrw_i({tielo_4bram3, bm_sclkrw_b2_o[1]}),
     .bm_sdo_o(bm_sdo_b3_o[1:0]), .padin_t_r(padin_t[23:12]),
     .bm_sreb_i(net990), .bm_sweb_i({tielo_4bram3, bm_sweb_b2_o[1]}),
     .padeb_t_r(padeb_t[23:12]),
     .fabric_out_08_17(fabric_out_08_17_ticegate),
     .tnl_op_07_16(slf_op_06_17[3:0]));
quad_tl_ice1 i_tl_quad ( .padin_l_t(padin_l[23:12]),
     .pado_l_t(pado_l[23:12]), .padeb_l_t(padeb_l[23:12]),
     .fo_dlyadj(fo_dlyadj[7:3]), .padin_06_17b(padin_0617b_ck),
     .padin_00_09a(padin_0009a_ck), .padeb_t_l(padeb_t[11:0]),
     .mode_o(net1135), .hiz_b_o(net1136),
     .fabric_out_06_17(fabric_out_06_17),
     .fabric_out_00_09(fabric_out_00_09), .cf_t(cf_t[143:0]),
     .cf_l(cf_l[383:192]), .ceb_o(net1139), .bs_en_o(net1140),
     .bm_sdi_i({tielo_4bram1, bm_sdi_b0_o[1]}),
     .bm_sdo_o(bm_sdo_b1_o[1:0]), .sp12_v_b_02_09(net1171[0:23]),
     .sp12_v_b_01_09(net1103[0:23]), .sp12_h_r_06_16(net770[0:23]),
     .sp12_h_r_06_15(net771[0:23]), .sp12_h_r_06_14(net772[0:23]),
     .sp12_h_r_06_13(net773[0:23]), .sp12_h_r_06_12(net774[0:23]),
     .sp12_h_r_06_11(net775[0:23]), .sp12_h_r_06_10(net776[0:23]),
     .sp12_h_r_06_09(net777[0:23]), .vdd_cntl_l(vdd_cntl_l[287:144]),
     .sp12_v_b_05_09(net1170[0:23]), .slf_op_06_17(slf_op_06_17[3:0]),
     .tclk_o(tclkio_ml), .update_o(net1102), .wl_l(wl_l[287:144]),
     .slf_op_06_16(slf_op_06_16[7:0]),
     .slf_op_06_15(slf_op_06_15[7:0]),
     .slf_op_06_14(slf_op_06_14[7:0]),
     .slf_op_06_13(slf_op_06_13[7:0]),
     .slf_op_06_12(slf_op_06_12[7:0]),
     .slf_op_06_11(slf_op_06_11[7:0]), .bm_wdummymux_en_i(net1183),
     .bm_sreb_i(net1185), .bm_sweb_i({tielo_4bram1, bm_sweb_b0_o[1]}),
     .sp12_v_b_03_09(net1231[0:23]), .shift_o(net1124), .sdo(sdio_ml),
     .r_o(net1132), .pado_t_l(pado_t[11:0]),
     .sp12_v_b_04_09(net1196[0:23]), .sp12_v_b_06_09(net1195[0:23]),
     .sp4_v_b_06_09(net1212[0:47]), .slf_op_06_10(slf_op_06_10[7:0]),
     .sp4_v_b_05_09(net1213[0:47]), .sp4_v_b_04_09(net1214[0:47]),
     .bnl_op_04_09(slf_op_03_08[7:0]),
     .bnl_op_05_09(slf_op_04_08[7:0]), .lc_bot_05_09(n_inter_05),
     .sp4_v_b_02_09(net1216[0:47]), .sp4_v_b_01_09(net1115[0:47]),
     .sp4_v_b_00_09(net1250[0:15]), .sp4_r_v_b_06_16(net810[0:47]),
     .sp4_r_v_b_06_15(net811[0:47]), .sp4_r_v_b_06_14(net812[0:47]),
     .sp4_r_v_b_06_13(net813[0:47]), .sp4_r_v_b_06_12(net814[0:47]),
     .sp4_r_v_b_06_11(net815[0:47]), .sp4_r_v_b_06_10(net816[0:47]),
     .sp4_r_v_b_06_09(net921[0:47]), .sp4_h_r_06_17(net818[0:15]),
     .sp4_h_r_06_16(net819[0:47]), .sp4_h_r_06_15(net820[0:47]),
     .sp4_h_r_06_14(net821[0:47]), .sp4_h_r_06_13(net822[0:47]),
     .sp4_h_r_06_12(net823[0:47]), .sp4_h_r_06_11(net824[0:47]),
     .bnl_op_03_09(slf_op_02_08[7:0]),
     .bnl_op_02_09(slf_op_01_08[7:0]), .bnl_op_01_09({slf_op_00_08[3],
     slf_op_00_08[2], slf_op_00_08[1], slf_op_00_08[0],
     slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0]}), .slf_op_00_09(slf_op_00_09[3:0]),
     .slf_op_06_09(slf_op_06_09[7:0]),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .lc_bot_01_09(n_inter_01), .lc_bot_02_09(n_inter_02),
     .lc_bot_04_09(n_inter_04), .bnl_op_06_09(slf_op_05_08[7:0]),
     .bnr_op_00_09(slf_op_01_08[7:0]),
     .bnr_op_01_09(slf_op_02_08[7:0]),
     .bnr_op_02_09(slf_op_03_08[7:0]),
     .bnr_op_03_09(slf_op_04_08[7:0]), .last_rsr(last_rsr[1]),
     .slf_op_05_09(slf_op_05_09[7:0]),
     .slf_op_04_09(slf_op_04_09[7:0]),
     .slf_op_03_09(slf_op_03_09[7:0]),
     .slf_op_02_09(slf_op_02_09[7:0]),
     .slf_op_01_09(slf_op_01_09[7:0]), .bl(bl_top[329:0]),
     .pgate_l(pgate_l[287:144]), .reset_b_l(reset_b_l[287:144]),
     .sp4_h_r_06_09(net848[0:47]), .sp4_h_r_06_10(net849[0:47]),
     .bnr_op_04_09(slf_op_05_08[7:0]),
     .bnr_op_05_09(slf_op_06_08[7:0]),
     .bnr_op_06_09(slf_op_07_08[7:0]),
     .bot_op_01_09(slf_op_01_08[7:0]),
     .carry_in_05_09(carry_io_05_0809),
     .carry_in_02_09(carry_io_02_0809),
     .carry_in_04_09(carry_io_04_0809),
     .carry_in_06_09(carry_io_06_0809), .ceb_i(net858),
     .bot_op_05_09(slf_op_05_08[7:0]),
     .bot_op_02_09(slf_op_02_08[7:0]),
     .bot_op_03_09(slf_op_03_08[7:0]),
     .bot_op_04_09(slf_op_04_08[7:0]), .update_i(net863),
     .tnr_op_06_16(slf_op_07_17[3:0]), .tclk_i(tclkio_mt),
     .shift_i(net866), .sdi(sdio_mt), .rgt_op_06_16(slf_op_07_16[7:0]),
     .rgt_op_06_15(slf_op_07_15[7:0]),
     .rgt_op_06_14(slf_op_07_14[7:0]),
     .rgt_op_06_13(slf_op_07_13[7:0]),
     .rgt_op_06_12(slf_op_07_12[7:0]),
     .rgt_op_06_11(slf_op_07_11[7:0]),
     .rgt_op_06_10(slf_op_07_10[7:0]),
     .rgt_op_06_09(slf_op_07_09[7:0]), .r_i(net876), .purst(purst),
     .prog(prog), .padin_t_l(padin_t[11:0]), .mode_i(net880),
     .hold_t_l(fabric_out_08_17_ticegate),
     .hold_l_t(fabric_out_00_07_licegate), .hiz_b_i(net883),
     .glb_in(gclk[7:0]), .lc_bot_06_09(n_inter_06),
     .sp4_v_b_03_09(net1215[0:47]), .carry_in_01_09(carry_io_01_0809),
     .bs_en_i(net888), .bot_op_06_09(slf_op_06_08[7:0]),
     .bm_ab_2bot(net1232[0:10]), .bm_aa_2bot(net1138[0:10]),
     .bm_init_i(net1192), .bm_rcapmux_en_i(net1191),
     .bm_sa_i(net1190[0:7]), .bm_sclk_i(bm_sck_b0_o),
     .bm_sclkrw_i({tielo_4bram1, bm_sclkrw_b0_o[1]}));
quad_br_ice1 i_br_quad ( net997, net996, net995[0:7], bm_sck_b2_o,
     bm_sclkrw_b2_o[1:0], bm_sdi_b2_o[1:0], bm_sdo_b2_o[1:0], net990,
     bm_sweb_b2_o[1:0], net988, net987, carry_io_07_0809,
     carry_io_08_0809, carry_io_09_0809, carry_io_11_0809,
     carry_io_12_0809, net980, cf_b[287:144], cf_r[191:0],
     fabric_out_07_00, fabric_out_12_00_wb, fabric_out_13_01,
     fabric_out_13_02, fabric_out_13_08, net975, net974, n_inter_07,
     n_inter_08, n_inter_09, n_inter_11, n_inter_12, padeb_b[11],
     padeb_b[23:13], padeb_r[12:0], padin_0700a_ck, padin_1308b_ck,
     pado_b[11], pado_b[23:13], pado_r[12:0], net971, sdio_mr, sdo_pad,
     net969, slf_op_07_00[3:0], slf_op_07_01[7:0], slf_op_07_02[7:0],
     slf_op_07_03[7:0], slf_op_07_04[7:0], slf_op_07_05[7:0],
     slf_op_07_06[7:0], slf_op_07_07[7:0], slf_op_07_08[7:0],
     slf_op_08_08[7:0], slf_op_09_08[7:0], slf_op_10_08[7:0],
     slf_op_11_08[7:0], slf_op_12_08[7:0], slf_op_13_08[3:0],
     spi_ss_in_bbank[4:0], tck_pad, tclkio_mr, tdi_pad, tms_pad,
     net957, bl_bot[663:334], pgate_r[143:0], reset_b_r[143:0],
     net1154[0:15], net1227[0:47], net1226[0:47], net1225[0:47],
     net1224[0:47], net1223[0:47], net1228[0:47], net1242[0:47],
     net1241[0:47], net1221[0:47], net1220[0:47], net1219[0:47],
     net1218[0:47], net1217[0:47], net1199[0:47], net1200[0:47],
     net1165[0:47], net921[0:47], net967[0:47], net998[0:47],
     net1001[0:47], net1000[0:47], net999[0:47], net911[0:15],
     net1209[0:23], net1208[0:23], net1207[0:23], net1206[0:23],
     net1205[0:23], net1198[0:23], net1197[0:23], net1222[0:23],
     net986[0:23], net985[0:23], net984[0:23], net983[0:23],
     net982[0:23], net981[0:23], vdd_cntl_r[143:0], wl_r[143:0],
     net1071[0:10], net1046[0:10], bm_bank30_init_o,
     bm_bank30_rcapmux_en_o, bm_bank30_sa_o[7:0], bm_bank30_sclk_o[1],
     net952[0:1], bm_bank30_sdi_o[3:2], {bm_sdo_b3_o_0,
     bm_sdi_b2_o[0]}, bm_bank30_sreb_o, net948[0:1], bm_wdummymux_en_o,
     slf_op_06_00[3:0], net1182, bs_en, net1176, ceb, end_of_startup,
     gclk[7:0], net1167, hiz_b, fabric_out_05_00_bicegate,
     fabric_out_13_10_ricegate, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr[2], last_rsr[3],
     slf_op_06_01[7:0], slf_op_06_02[7:0], slf_op_06_03[7:0],
     slf_op_06_04[7:0], slf_op_06_05[7:0], slf_op_06_06[7:0],
     slf_op_06_07[7:0], slf_op_06_08[7:0], md_spi_b, net1166, mode,
     mux_jtag_sel_b, padin_b[11], padin_b[23:13], padin_r[12:0],
     pll_sdo, prog, purst, net1164, r, sdio_mb, sdi_pad, sdo_enable,
     net1162, shift, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out,
     tclkio_mb, tclk, slf_op_06_09[7:0], slf_op_07_09[7:0],
     slf_op_08_09[7:0], slf_op_09_09[7:0], slf_op_10_09[7:0],
     slf_op_11_09[7:0], slf_op_12_09[7:0], slf_op_08_09[7:0],
     slf_op_09_09[7:0], slf_op_10_09[7:0], slf_op_11_09[7:0],
     slf_op_12_09[7:0], {slf_op_13_09[3], slf_op_13_09[2],
     slf_op_13_09[1], slf_op_13_09[0], slf_op_13_09[3],
     slf_op_13_09[2], slf_op_13_09[1], slf_op_13_09[0]},
     slf_op_07_09[7:0], slf_op_08_09[7:0], slf_op_09_09[7:0],
     slf_op_10_09[7:0], slf_op_11_09[7:0], slf_op_12_09[7:0], totdopad,
     trstb_pad, net1152, update);
quad_bl_ice1 i_bl_quad ( net1192, net1191, net1190[0:7], bm_sck_b0_o,
     bm_sclkrw_b0_o[1:0], bm_sdi_b0_o[1:0], bm_sdo_b0_o[1:0], net1185,
     bm_sweb_b0_o[1:0], net1183, net1182, carry_io_01_0809,
     carry_io_02_0809, carry_io_04_0809, carry_io_05_0809,
     carry_io_06_0809, net1176, cf_b[143:0], cf_l[191:0],
     fabric_out_00_07_licegate, fabric_out_00_08,
     fabric_out_05_00_bicegate, fabric_out_06_00, fo_bypass,
     fo_dlyadj[2:0], fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, net1167,
     net1166, n_inter_01, n_inter_02, n_inter_04, n_inter_05,
     n_inter_06, padeb_b[10:0], padeb_b[12], padeb_l[11:0],
     padin_0008b_ck, padin_0600b_ck, pado_b[10:0], pado_b[12],
     pado_l[11:0], net1164, sdio_mb, net1162, slf_op_00_08[3:0],
     slf_op_01_08[7:0], slf_op_02_08[7:0], slf_op_03_08[7:0],
     slf_op_04_08[7:0], slf_op_05_08[7:0], slf_op_06_00[3:0],
     slf_op_06_01[7:0], slf_op_06_02[7:0], slf_op_06_03[7:0],
     slf_op_06_04[7:0], slf_op_06_05[7:0], slf_op_06_06[7:0],
     slf_op_06_07[7:0], slf_op_06_08[7:0], tclkio_mb, net1152,
     bl_bot[329:0], pgate_l[143:0], reset_b_l[143:0], net1154[0:15],
     net1227[0:47], net1226[0:47], net1225[0:47], net1224[0:47],
     net1223[0:47], net1228[0:47], net1242[0:47], net1241[0:47],
     net1221[0:47], net1220[0:47], net1219[0:47], net1218[0:47],
     net1217[0:47], net1199[0:47], net1200[0:47], net1165[0:47],
     net1250[0:15], net1115[0:47], net1216[0:47], net1215[0:47],
     net1214[0:47], net1213[0:47], net1212[0:47], net1209[0:23],
     net1208[0:23], net1207[0:23], net1206[0:23], net1205[0:23],
     net1198[0:23], net1197[0:23], net1222[0:23], net1103[0:23],
     net1171[0:23], net1231[0:23], net1196[0:23], net1170[0:23],
     net1195[0:23], vdd_cntl_l[143:0], wl_l[143:0], net1138[0:10],
     net1232[0:10], net1151, net1150, net1149[0:7], bm_sck_b0_i,
     net1147[0:1], net1146[0:1], {bm_sdo_b1_o_0, bm_sdi_b0_o[0]},
     net1144, net1143[0:1], net1142, slf_op_07_00[3:0], net1140,
     net1139, gclk[7:0], net1136, fabric_out_05_00_bicegate,
     fabric_out_00_07_licegate, jtag_rowtest_mode_rowu0_b, last_rsr[0],
     net1135, padin_b[10:0], padin_b[12], padin_l[11:0], pll_lock_out,
     prog, purst, net1132, slf_op_07_01[7:0], slf_op_07_02[7:0],
     slf_op_07_03[7:0], slf_op_07_04[7:0], slf_op_07_05[7:0],
     slf_op_07_06[7:0], slf_op_07_07[7:0], slf_op_07_08[7:0], sdio_ml,
     net1124, tclkio_ml, {slf_op_00_09[3], slf_op_00_09[2],
     slf_op_00_09[1], slf_op_00_09[0], slf_op_00_09[3],
     slf_op_00_09[2], slf_op_00_09[1], slf_op_00_09[0]},
     slf_op_01_09[7:0], slf_op_02_09[7:0], slf_op_03_09[7:0],
     slf_op_04_09[7:0], slf_op_05_09[7:0], slf_op_01_09[7:0],
     slf_op_02_09[7:0], slf_op_03_09[7:0], slf_op_04_09[7:0],
     slf_op_05_09[7:0], slf_op_06_09[7:0], slf_op_07_09[7:0],
     slf_op_01_09[7:0], slf_op_02_09[7:0], slf_op_03_09[7:0],
     slf_op_04_09[7:0], slf_op_05_09[7:0], slf_op_06_09[7:0], net1102);
bram_bank_logic_bot I21 ( .bm_sdo_i({bm_sdo_b2_o[1], bm_sdo_b2_o_0}),
     .bm_sclk_i(bm_bank30_sclk_o[1]), .bm_sclkrw_i(bm_bank30_sclkrw_o),
     .bm_sweb_i(bm_bank30_sweb_o), .bm_sdo_o(bm_bank30_sdo_i[3:2]),
     .bm_sweb_o(net948[0:1]), .bm_sclkrw_o(net952[0:1]),
     .bm_banksel_i(bm_bank30_banksel_o[3:2]));
bram_bank_logic_bot I63 ( .bm_sdo_i({bm_sdo_b0_o[1], bm_sdo_b0_o_0}),
     .bm_sclk_i(bm_sck_b0_i), .bm_sclkrw_i(net1273),
     .bm_sweb_i(net1274), .bm_sdo_o(net1275[0:1]),
     .bm_sweb_o(net1143[0:1]), .bm_sclkrw_o(net1147[0:1]),
     .bm_banksel_i(bm_bank10_banksel_o[1:0]));
bram_hbuffer_dff_2xbank I_bram_buf1 ( .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_banksel_o(bm_bank30_banksel_o[3:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sweb_o(bm_bank30_sweb_o), .bm_sreb_o(bm_bank30_sreb_o),
     .bm_sclk_o(bm_bank30_sclk_o[1:0]), .bm_sa_o(bm_bank30_sa_o[7:0]),
     .bm_init_o(bm_bank30_init_o), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclkrw_o(bm_bank30_sclkrw_o), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sdo_o(bm_sdo_o[3:0]), .bm_sdi_o(bm_bank30_sdi_o[3:0]),
     .bm_rcapmux_en_o(bm_bank30_rcapmux_en_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_banksel_i(bm_banksel_i[3:0]),
     .bm_sdo_i(bm_bank30_sdo_i[3:0]));
bram_hbuffer_1xbank I2 ( .bm_sa_o(net1149[0:7]),
     .bm_wdummymux_en_o(net1142), .bm_sweb_i(bm_bank30_sweb_o),
     .bm_sreb_i(bm_bank30_sreb_o), .bm_sdi_i(bm_bank30_sdi_o[1:0]),
     .bm_sclk_i(bm_bank30_sclk_o[0]), .bm_init_i(bm_bank30_init_o),
     .bm_banksel_o(bm_bank10_banksel_o[1:0]),
     .bm_rcapmux_en_i(bm_bank30_rcapmux_en_o),
     .bm_wdummymux_en_i(bm_wdummymux_en_o), .bm_sweb_o(net1274),
     .bm_sreb_o(net1144), .bm_sdi_o(net1146[0:1]),
     .bm_sclk_o(bm_sck_b0_i), .bm_init_o(net1151),
     .bm_sa_i(bm_bank30_sa_o[7:0]), .bm_rcapmux_en_o(net1150),
     .bm_sclkrw_i(bm_bank30_sclkrw_o), .bm_sclkrw_o(net1273),
     .bm_sdo_i(net1275[0:1]), .bm_banksel_i(bm_bank30_banksel_o[1:0]),
     .bm_sdo_o(bm_bank30_sdo_i[1:0]));

endmodule
// Library - misc, Cell - nvcm_top_ice8p, View - schematic
// LAST TIME SAVED: Nov 17 16:51:37 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_top_ice8p ( bp0, fsm_blkadd, fsm_blkadd_b, fsm_coladd,
     fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_redrow,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_recall,
     fsm_rowadd, fsm_sample, fsm_tm_allbank_sel, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_bgr_dis,
     fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_ref,
     fsm_tm_rprd, fsm_tm_tcol, fsm_tm_testdec, fsm_tm_testdec_wr,
     fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvpp, fsm_tm_xvpxa_int, fsm_trim_ipp,
     fsm_trim_multibl_read, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_trim_vbg, fsm_trim_vpgmwl, fsm_trim_vrdwl, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b, status_wip, clk,
     nv_dataout, nvcm_ce_b, nvcm_max_coladd, nvcm_max_rowadd, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_redrow, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_recall, fsm_sample, fsm_tm_allbank_sel,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_bgr_dis, fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_tcol, fsm_tm_testdec, fsm_tm_testdec_wr,
     fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvpp, fsm_tm_xvpxa_int, fsm_trim_multibl_read, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b, status_wip;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

output [3:0]  fsm_blkadd_b;
output [8:0]  fsm_rowadd;
output [1:0]  fsm_tm_ref;
output [11:0]  fsm_coladd;
output [2:0]  fsm_trim_vrdwl;
output [3:0]  fsm_trim_vbg;
output [3:0]  fsm_blkadd;
output [3:0]  fsm_trim_ipp;
output [2:0]  fsm_trim_vpgmwl;
output [2:0]  fsm_trim_rrefrd;
output [2:0]  fsm_trim_rrefpgm;

input [11:0]  nvcm_max_coladd;
input [8:0]  nvcm_max_rowadd;
input [8:0]  nv_dataout;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - sbtlibn65lp, Cell - vddp_tiehigh, View - schematic
// LAST TIME SAVED: Jun 21 10:52:52 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module vddp_tiehigh ( vddp_tieh );
inout  vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M8 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net9), .S(vddp_));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_rows, View - schematic
// LAST TIME SAVED: Jul 27 16:24:09 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_testdec_rows ( dec_bias, dec_det, vddp_tieh, wp, wr );
inout  dec_bias, dec_det;

input  vddp_tieh, wp, wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M8 ( .D(dec_det), .B(GND_), .G(wr), .S(gnd_));
nch  M6 ( .D(dec_det), .B(GND_), .G(net20), .S(gnd_));
nch  M5 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(net20));
nch  M7 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(wr));
nch_25  M12 ( .D(net20), .B(gnd_), .G(vddp_tieh), .S(wp));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_rowsx108_1f, View - schematic
// LAST TIME SAVED: Dec 23 16:24:55 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_testdec_rowsx108_1f ( dec_det_buf, dec_bias, dec_det, wp, wr
     );
output  dec_det_buf;

inout  dec_bias, dec_det;


input [107:0]  wr;
input [107:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(dec_det), .Y(net25));
inv_hvt I27 ( .A(net25), .Y(dec_det_buf));
vddp_tiehigh I25 ( .vddp_tieh(vddp_tiel));
ml_testdec_rows Itestdec_rows_107_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[107]), .wp(wp[107]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_106_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[106]), .wp(wp[106]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_105_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[105]), .wp(wp[105]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_104_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[104]), .wp(wp[104]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_103_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[103]), .wp(wp[103]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_102_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[102]), .wp(wp[102]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_101_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[101]), .wp(wp[101]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_100_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[100]), .wp(wp[100]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_99_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[99]), .wp(wp[99]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_98_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[98]), .wp(wp[98]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_97_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[97]), .wp(wp[97]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_96_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[96]), .wp(wp[96]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_95_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[95]), .wp(wp[95]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_94_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[94]), .wp(wp[94]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_93_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[93]), .wp(wp[93]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_92_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[92]), .wp(wp[92]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_91_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[91]), .wp(wp[91]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_90_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[90]), .wp(wp[90]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_89_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[89]), .wp(wp[89]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_88_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[88]), .wp(wp[88]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_87_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[87]), .wp(wp[87]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_86_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[86]), .wp(wp[86]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_85_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[85]), .wp(wp[85]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_84_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[84]), .wp(wp[84]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_83_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[83]), .wp(wp[83]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_82_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[82]), .wp(wp[82]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_81_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[81]), .wp(wp[81]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_80_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[80]), .wp(wp[80]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_79_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[79]), .wp(wp[79]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_78_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[78]), .wp(wp[78]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_77_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[77]), .wp(wp[77]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_76_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[76]), .wp(wp[76]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_75_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[75]), .wp(wp[75]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_74_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[74]), .wp(wp[74]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_73_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[73]), .wp(wp[73]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_72_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[72]), .wp(wp[72]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_71_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[71]), .wp(wp[71]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_70_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[70]), .wp(wp[70]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_69_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[69]), .wp(wp[69]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_68_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[68]), .wp(wp[68]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_67_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[67]), .wp(wp[67]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_66_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[66]), .wp(wp[66]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_65_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[65]), .wp(wp[65]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_64_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[64]), .wp(wp[64]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_63_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[63]), .wp(wp[63]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_62_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[62]), .wp(wp[62]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_61_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[61]), .wp(wp[61]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_60_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[60]), .wp(wp[60]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_59_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[59]), .wp(wp[59]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_58_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[58]), .wp(wp[58]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_57_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[57]), .wp(wp[57]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_56_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[56]), .wp(wp[56]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_55_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[55]), .wp(wp[55]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_54_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[54]), .wp(wp[54]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_53_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[53]), .wp(wp[53]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_52_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[52]), .wp(wp[52]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_51_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[51]), .wp(wp[51]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_50_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[50]), .wp(wp[50]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_49_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[49]), .wp(wp[49]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_48_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[48]), .wp(wp[48]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_47_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[47]), .wp(wp[47]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_46_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[46]), .wp(wp[46]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_45_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[45]), .wp(wp[45]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_44_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[44]), .wp(wp[44]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_43_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[43]), .wp(wp[43]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_42_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[42]), .wp(wp[42]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_41_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[41]), .wp(wp[41]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_40_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[40]), .wp(wp[40]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_39_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[39]), .wp(wp[39]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_38_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[38]), .wp(wp[38]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_37_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[37]), .wp(wp[37]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_36_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[36]), .wp(wp[36]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_35_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[35]), .wp(wp[35]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_34_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[34]), .wp(wp[34]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_33_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[33]), .wp(wp[33]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_32_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[32]), .wp(wp[32]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_31_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[31]), .wp(wp[31]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_30_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[30]), .wp(wp[30]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_29_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[29]), .wp(wp[29]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_28_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[28]), .wp(wp[28]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_27_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[27]), .wp(wp[27]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_26_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[26]), .wp(wp[26]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_25_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[25]), .wp(wp[25]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_24_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[24]), .wp(wp[24]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_23_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[23]), .wp(wp[23]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_22_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[22]), .wp(wp[22]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_21_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[21]), .wp(wp[21]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_20_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[20]), .wp(wp[20]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_19_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[19]), .wp(wp[19]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_18_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[18]), .wp(wp[18]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_17_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[17]), .wp(wp[17]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_16_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[16]), .wp(wp[16]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_15_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[15]), .wp(wp[15]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_14_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[14]), .wp(wp[14]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_13_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[13]), .wp(wp[13]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_12_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[12]), .wp(wp[12]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_11_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[11]), .wp(wp[11]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_10_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[10]), .wp(wp[10]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_9_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[9]), .wp(wp[9]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_8_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[8]), .wp(wp[8]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_7_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[7]), .wp(wp[7]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_6_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[6]), .wp(wp[6]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_5_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[5]), .wp(wp[5]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_4_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[4]), .wp(wp[4]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_3_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[3]), .wp(wp[3]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_2_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[2]), .wp(wp[2]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_1_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[1]), .wp(wp[1]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_0_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[0]), .wp(wp[0]),
     .dec_bias(dec_bias));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd2vdd25, View - schematic
// LAST TIME SAVED: Jun 11 16:25:15 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
nch_25  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));
pch_25  M0 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
pch_25  M1 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
pch_25  M2 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
pch_25  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));

endmodule
// Library - tsmcN40, Cell - nor2_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:25 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nor2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  M2 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  M1 ( .D(net15), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(net15));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_columns, View - schematic
// LAST TIME SAVED: Jun 24 12:15:49 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_testdec_columns ( bl, vdd_drv, dec_det_even_25,
     dec_det_odd_25 );
inout  vdd_drv;

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(vdd_drv), .B(gnd_), .G(dec_det_even_25), .S(bl[0]));
nch_25  M4 ( .D(vdd_drv), .B(gnd_), .G(dec_det_odd_25), .S(bl[1]));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_columnsx330_1f, View -
//schematic
// LAST TIME SAVED: Dec 28 17:38:01 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_testdec_columnsx330_1f ( bl, bl_dummyl, bl_dummyr, bl_test,
     dec_det_buf, testdec_even_b_25, testdec_odd_b_25 );

input  dec_det_buf, testdec_even_b_25, testdec_odd_b_25;

inout [327:0]  bl;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I134 ( .A(dec_det_buf), .Y(net40));
inv_hvt I55 ( .A(net40), .Y(net36));
ml_ls_vdd2vdd25 I144 ( .in(net36), .sup(vddp_), .out_vddio_b(net38),
     .out_vddio(dec_det_25), .in_b(net40));
nor2_25 I26 ( .A(testdec_odd_b_25), .Y(dec_det_odd_25), .Gb(GND_),
     .G(GND_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
nor2_25 I59 ( .A(testdec_even_b_25), .Y(dec_det_even_25), .Gb(GND_),
     .G(GND_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
rppolywo  R1 ( .MINUS(vdd_drv), .PLUS(vdd_));
rppolywo  R2 ( .MINUS(vdd_drv), .PLUS(vdd_));
rppolywo  R3 ( .MINUS(vdd_drv), .PLUS(vdd_));
rppolywo  R0 ( .MINUS(vdd_drv), .PLUS(vdd_));
ml_testdec_columns Itestdec_columns_dml ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyl[1:0]));
ml_testdec_columns Itestdec_columns_163_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[327:326]));
ml_testdec_columns Itestdec_columns_162_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[325:324]));
ml_testdec_columns Itestdec_columns_161_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[323:322]));
ml_testdec_columns Itestdec_columns_160_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[321:320]));
ml_testdec_columns Itestdec_columns_159_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[319:318]));
ml_testdec_columns Itestdec_columns_158_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[317:316]));
ml_testdec_columns Itestdec_columns_157_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[315:314]));
ml_testdec_columns Itestdec_columns_156_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[313:312]));
ml_testdec_columns Itestdec_columns_155_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[311:310]));
ml_testdec_columns Itestdec_columns_154_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[309:308]));
ml_testdec_columns Itestdec_columns_153_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[307:306]));
ml_testdec_columns Itestdec_columns_152_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[305:304]));
ml_testdec_columns Itestdec_columns_151_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[303:302]));
ml_testdec_columns Itestdec_columns_150_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[301:300]));
ml_testdec_columns Itestdec_columns_149_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[299:298]));
ml_testdec_columns Itestdec_columns_148_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[297:296]));
ml_testdec_columns Itestdec_columns_147_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[295:294]));
ml_testdec_columns Itestdec_columns_146_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[293:292]));
ml_testdec_columns Itestdec_columns_145_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[291:290]));
ml_testdec_columns Itestdec_columns_144_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[289:288]));
ml_testdec_columns Itestdec_columns_143_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[287:286]));
ml_testdec_columns Itestdec_columns_142_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[285:284]));
ml_testdec_columns Itestdec_columns_141_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[283:282]));
ml_testdec_columns Itestdec_columns_140_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[281:280]));
ml_testdec_columns Itestdec_columns_139_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[279:278]));
ml_testdec_columns Itestdec_columns_138_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[277:276]));
ml_testdec_columns Itestdec_columns_137_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[275:274]));
ml_testdec_columns Itestdec_columns_136_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[273:272]));
ml_testdec_columns Itestdec_columns_135_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[271:270]));
ml_testdec_columns Itestdec_columns_134_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[269:268]));
ml_testdec_columns Itestdec_columns_133_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[267:266]));
ml_testdec_columns Itestdec_columns_132_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[265:264]));
ml_testdec_columns Itestdec_columns_131_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[263:262]));
ml_testdec_columns Itestdec_columns_130_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[261:260]));
ml_testdec_columns Itestdec_columns_129_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[259:258]));
ml_testdec_columns Itestdec_columns_128_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[257:256]));
ml_testdec_columns Itestdec_columns_127_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[255:254]));
ml_testdec_columns Itestdec_columns_126_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[253:252]));
ml_testdec_columns Itestdec_columns_125_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[251:250]));
ml_testdec_columns Itestdec_columns_124_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[249:248]));
ml_testdec_columns Itestdec_columns_123_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[247:246]));
ml_testdec_columns Itestdec_columns_122_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[245:244]));
ml_testdec_columns Itestdec_columns_121_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[243:242]));
ml_testdec_columns Itestdec_columns_120_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[241:240]));
ml_testdec_columns Itestdec_columns_119_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[239:238]));
ml_testdec_columns Itestdec_columns_118_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[237:236]));
ml_testdec_columns Itestdec_columns_117_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[235:234]));
ml_testdec_columns Itestdec_columns_116_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[233:232]));
ml_testdec_columns Itestdec_columns_115_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[231:230]));
ml_testdec_columns Itestdec_columns_114_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[229:228]));
ml_testdec_columns Itestdec_columns_113_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[227:226]));
ml_testdec_columns Itestdec_columns_112_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[225:224]));
ml_testdec_columns Itestdec_columns_111_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[223:222]));
ml_testdec_columns Itestdec_columns_110_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[221:220]));
ml_testdec_columns Itestdec_columns_109_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[219:218]));
ml_testdec_columns Itestdec_columns_108_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[217:216]));
ml_testdec_columns Itestdec_columns_107_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[215:214]));
ml_testdec_columns Itestdec_columns_106_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[213:212]));
ml_testdec_columns Itestdec_columns_105_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[211:210]));
ml_testdec_columns Itestdec_columns_104_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[209:208]));
ml_testdec_columns Itestdec_columns_103_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[207:206]));
ml_testdec_columns Itestdec_columns_102_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[205:204]));
ml_testdec_columns Itestdec_columns_101_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[203:202]));
ml_testdec_columns Itestdec_columns_100_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[201:200]));
ml_testdec_columns Itestdec_columns_99_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[199:198]));
ml_testdec_columns Itestdec_columns_98_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[197:196]));
ml_testdec_columns Itestdec_columns_97_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[195:194]));
ml_testdec_columns Itestdec_columns_96_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[193:192]));
ml_testdec_columns Itestdec_columns_95_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[191:190]));
ml_testdec_columns Itestdec_columns_94_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[189:188]));
ml_testdec_columns Itestdec_columns_93_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[187:186]));
ml_testdec_columns Itestdec_columns_92_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[185:184]));
ml_testdec_columns Itestdec_columns_91_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[183:182]));
ml_testdec_columns Itestdec_columns_90_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[181:180]));
ml_testdec_columns Itestdec_columns_89_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[179:178]));
ml_testdec_columns Itestdec_columns_88_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[177:176]));
ml_testdec_columns Itestdec_columns_87_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[175:174]));
ml_testdec_columns Itestdec_columns_86_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[173:172]));
ml_testdec_columns Itestdec_columns_85_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[171:170]));
ml_testdec_columns Itestdec_columns_84_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[169:168]));
ml_testdec_columns Itestdec_columns_83_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[167:166]));
ml_testdec_columns Itestdec_columns_82_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[165:164]));
ml_testdec_columns Itestdec_columns_81_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[163:162]));
ml_testdec_columns Itestdec_columns_80_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[161:160]));
ml_testdec_columns Itestdec_columns_79_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[159:158]));
ml_testdec_columns Itestdec_columns_78_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[157:156]));
ml_testdec_columns Itestdec_columns_77_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[155:154]));
ml_testdec_columns Itestdec_columns_76_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[153:152]));
ml_testdec_columns Itestdec_columns_75_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[151:150]));
ml_testdec_columns Itestdec_columns_74_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[149:148]));
ml_testdec_columns Itestdec_columns_73_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[147:146]));
ml_testdec_columns Itestdec_columns_72_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[145:144]));
ml_testdec_columns Itestdec_columns_71_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[143:142]));
ml_testdec_columns Itestdec_columns_70_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[141:140]));
ml_testdec_columns Itestdec_columns_69_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[139:138]));
ml_testdec_columns Itestdec_columns_68_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[137:136]));
ml_testdec_columns Itestdec_columns_67_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[135:134]));
ml_testdec_columns Itestdec_columns_66_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[133:132]));
ml_testdec_columns Itestdec_columns_65_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[131:130]));
ml_testdec_columns Itestdec_columns_64_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[129:128]));
ml_testdec_columns Itestdec_columns_63_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[127:126]));
ml_testdec_columns Itestdec_columns_62_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[125:124]));
ml_testdec_columns Itestdec_columns_61_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[123:122]));
ml_testdec_columns Itestdec_columns_60_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[121:120]));
ml_testdec_columns Itestdec_columns_59_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[119:118]));
ml_testdec_columns Itestdec_columns_58_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[117:116]));
ml_testdec_columns Itestdec_columns_57_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[115:114]));
ml_testdec_columns Itestdec_columns_56_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[113:112]));
ml_testdec_columns Itestdec_columns_55_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[111:110]));
ml_testdec_columns Itestdec_columns_54_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[109:108]));
ml_testdec_columns Itestdec_columns_53_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[107:106]));
ml_testdec_columns Itestdec_columns_52_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[105:104]));
ml_testdec_columns Itestdec_columns_51_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[103:102]));
ml_testdec_columns Itestdec_columns_50_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[101:100]));
ml_testdec_columns Itestdec_columns_49_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[99:98]));
ml_testdec_columns Itestdec_columns_48_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[97:96]));
ml_testdec_columns Itestdec_columns_47_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[95:94]));
ml_testdec_columns Itestdec_columns_46_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[93:92]));
ml_testdec_columns Itestdec_columns_45_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[91:90]));
ml_testdec_columns Itestdec_columns_44_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[89:88]));
ml_testdec_columns Itestdec_columns_43_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[87:86]));
ml_testdec_columns Itestdec_columns_42_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[85:84]));
ml_testdec_columns Itestdec_columns_41_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[83:82]));
ml_testdec_columns Itestdec_columns_40_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[81:80]));
ml_testdec_columns Itestdec_columns_39_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[79:78]));
ml_testdec_columns Itestdec_columns_38_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[77:76]));
ml_testdec_columns Itestdec_columns_37_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[75:74]));
ml_testdec_columns Itestdec_columns_36_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[73:72]));
ml_testdec_columns Itestdec_columns_35_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[71:70]));
ml_testdec_columns Itestdec_columns_34_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[69:68]));
ml_testdec_columns Itestdec_columns_33_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[67:66]));
ml_testdec_columns Itestdec_columns_32_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[65:64]));
ml_testdec_columns Itestdec_columns_31_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[63:62]));
ml_testdec_columns Itestdec_columns_30_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[61:60]));
ml_testdec_columns Itestdec_columns_29_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[59:58]));
ml_testdec_columns Itestdec_columns_28_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[57:56]));
ml_testdec_columns Itestdec_columns_27_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[55:54]));
ml_testdec_columns Itestdec_columns_26_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[53:52]));
ml_testdec_columns Itestdec_columns_25_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[51:50]));
ml_testdec_columns Itestdec_columns_24_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[49:48]));
ml_testdec_columns Itestdec_columns_23_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[47:46]));
ml_testdec_columns Itestdec_columns_22_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[45:44]));
ml_testdec_columns Itestdec_columns_21_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[43:42]));
ml_testdec_columns Itestdec_columns_20_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[41:40]));
ml_testdec_columns Itestdec_columns_19_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[39:38]));
ml_testdec_columns Itestdec_columns_18_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[37:36]));
ml_testdec_columns Itestdec_columns_17_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[35:34]));
ml_testdec_columns Itestdec_columns_16_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[33:32]));
ml_testdec_columns Itestdec_columns_15_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[31:30]));
ml_testdec_columns Itestdec_columns_14_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[29:28]));
ml_testdec_columns Itestdec_columns_13_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[27:26]));
ml_testdec_columns Itestdec_columns_12_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[25:24]));
ml_testdec_columns Itestdec_columns_11_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[23:22]));
ml_testdec_columns Itestdec_columns_10_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[21:20]));
ml_testdec_columns Itestdec_columns_9_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[19:18]));
ml_testdec_columns Itestdec_columns_8_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[17:16]));
ml_testdec_columns Itestdec_columns_7_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[15:14]));
ml_testdec_columns Itestdec_columns_6_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[13:12]));
ml_testdec_columns Itestdec_columns_5_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[11:10]));
ml_testdec_columns Itestdec_columns_4_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[9:8]));
ml_testdec_columns Itestdec_columns_3_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[7:6]));
ml_testdec_columns Itestdec_columns_2_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[5:4]));
ml_testdec_columns Itestdec_columns_1_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[3:2]));
ml_testdec_columns Itestdec_columns_0_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[1:0]));
ml_testdec_columns Itestdec_columns_dmr ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyr[1:0]));
ml_testdec_columns Itestdec_columns_tst ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_test[1:0]));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tielow, View - schematic
// LAST TIME SAVED: Jul 20 11:25:32 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module vdd_tielow ( gnd_tiel );
inout  gnd_tiel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(gnd_tiel), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(net9), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - leafcell, Cell - buffer500um, View - schematic
// LAST TIME SAVED: May 13 11:02:42 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module buffer500um ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - NVCM_40nm, Cell - cell_1x1, View - schematic
// LAST TIME SAVED: Oct 15 17:03:11 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module cell_1x1 ( bl, wp, wr );
inout  bl;

input  wp, wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nchx  WR_CELL ( .D(net08), .G(wr), .S(bl));
nchx  WP_CELL ( .D(net011), .G(wp), .S(net08));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x1, View - schematic
// LAST TIME SAVED: Jul 12 16:56:42 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_cell_2x1 ( bl, wp, wr );

input  wp, wr;

inout [1:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cell_1x1 I11 ( .wp(wp), .wr(wr), .bl(bl[0]));
cell_1x1 I12 ( .wp(wp), .wr(wr), .bl(bl[1]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x8, View - schematic
// LAST TIME SAVED: Feb 26 14:36:29 2008
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_cell_2x8 ( bl, wp, wr );


inout [1:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m7 ( .bl(bl[1:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_2x1 m6 ( .bl(bl[1:0]), .wr(wr[6]), .wp(wp[6]));
nvcm_cell_2x1 m5 ( .bl(bl[1:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_2x1 m4 ( .bl(bl[1:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_2x1 m3 ( .bl(bl[1:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_2x1 m2 ( .bl(bl[1:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_1x8, View - schematic
// LAST TIME SAVED: Jul  8 17:57:53 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_cell_1x8 ( bl, wp, wr );

input  wp, wr;

inout [7:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cell_1x1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
cell_1x1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));
cell_1x1 m2 ( .wp(wp), .wr(wr), .bl(bl[2]));
cell_1x1 m3 ( .wp(wp), .wr(wr), .bl(bl[3]));
cell_1x1 m4 ( .wp(wp), .wr(wr), .bl(bl[4]));
cell_1x1 m5 ( .wp(wp), .wr(wr), .bl(bl[5]));
cell_1x1 m6 ( .wp(wp), .wr(wr), .bl(bl[6]));
cell_1x1 m7 ( .wp(wp), .wr(wr), .bl(bl[7]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_8x8, View - schematic
// LAST TIME SAVED: Jun 24 17:57:01 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_cell_8x8 ( bl, wp, wr );


inout [7:0]  bl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 m0 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 m1 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 m2 ( .bl(bl[7:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_1x8 m3 ( .bl(bl[7:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_1x8 m7 ( .bl(bl[7:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_1x8 m4 ( .bl(bl[7:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_1x8 m5 ( .bl(bl[7:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_1x8 m6 ( .bl(bl[7:0]), .wr(wr[6]), .wp(wp[6]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_16x8, View - schematic
// LAST TIME SAVED: Jun 24 17:57:26 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_cell_16x8 ( bl, wp, wr );


inout [15:0]  bl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_8x8 m0 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[7:0]));
nvcm_cell_8x8 m1 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[15:8]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_336x8, View - schematic
// LAST TIME SAVED: Dec 30 14:06:16 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_cell_336x8 ( bl, bl_dummyl, bl_dummyr, bl_test, wp, wr );


inout [5:0]  bl_dummyr;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [327:0]  bl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x8 Invcm_cell_2x8 ( .wp(wp[7:0]), .wr(wr[7:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_16x8 Invcm_cell_16x8_19_ ( .wp(wp[7:0]), .bl(bl[319:304]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_18_ ( .wp(wp[7:0]), .bl(bl[303:288]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_17_ ( .wp(wp[7:0]), .bl(bl[287:272]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_16_ ( .wp(wp[7:0]), .bl(bl[271:256]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_15_ ( .wp(wp[7:0]), .bl(bl[255:240]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_14_ ( .wp(wp[7:0]), .bl(bl[239:224]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_13_ ( .wp(wp[7:0]), .bl(bl[223:208]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_12_ ( .wp(wp[7:0]), .bl(bl[207:192]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_11_ ( .wp(wp[7:0]), .bl(bl[191:176]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_10_ ( .wp(wp[7:0]), .bl(bl[175:160]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_9_ ( .wp(wp[7:0]), .bl(bl[159:144]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_8_ ( .wp(wp[7:0]), .bl(bl[143:128]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_7_ ( .wp(wp[7:0]), .bl(bl[127:112]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_6_ ( .wp(wp[7:0]), .bl(bl[111:96]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_5_ ( .wp(wp[7:0]), .bl(bl[95:80]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_4_ ( .wp(wp[7:0]), .bl(bl[79:64]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_3_ ( .wp(wp[7:0]), .bl(bl[63:48]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_2_ ( .wp(wp[7:0]), .bl(bl[47:32]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_1_ ( .wp(wp[7:0]), .bl(bl[31:16]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_0_ ( .wp(wp[7:0]), .bl(bl[15:0]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_20_ ( .wp(wp[7:0]), .bl({bl_dummyr[5:0],
     bl_test[1:0], bl[327:320]}), .wr(wr[7:0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_338x112_1f, View - schematic
// LAST TIME SAVED: Dec 28 17:18:26 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nvcm_cell_338x112_1f ( bl, bl_dummyl, bl_dummyr, bl_test, wp,
     wp_dummyb, wp_dummyt, wr, wr_dummyb, wr_dummyt );


inout [1:0]  bl_dummyr;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [327:0]  bl;

input [1:0]  wp_dummyb;
input [1:0]  wr_dummyb;
input [1:0]  wr_dummyt;
input [107:0]  wp;
input [1:0]  wp_dummyt;
input [107:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_336x8 Invcm_cell_336x8_11_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[101:94]), .wp(wp[101:94]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_10_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[93:86]), .wp(wp[93:86]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_9_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[85:78]), .wp(wp[85:78]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_8_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[77:70]), .wp(wp[77:70]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_7_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[69:62]), .wp(wp[69:62]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_6_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[61:54]), .wp(wp[61:54]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_5_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[53:46]), .wp(wp[53:46]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_4_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[45:38]), .wp(wp[45:38]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_3_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[37:30]), .wp(wp[37:30]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_2_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[29:22]), .wp(wp[29:22]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_1_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[21:14]), .wp(wp[21:14]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_0_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[13:6]), .wp(wp[13:6]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_t ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr({wr[5:0], wr_dummyt[1:0]}), .wp({wp[5:0], wp_dummyt[1:0]}),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_b ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr({wr_dummyb[1:0], wr[107:102]}), .wp({wp_dummyb[1:0],
     wp[107:102]}), .bl_dummyl(bl_dummyl[1:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_bgen, View - schematic
// LAST TIME SAVED: Jul 15 18:50:47 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_testdec_bgen ( dec_ok, dec_bias, dec_det, testdec_en_b,
     testdec_prec_b );
output  dec_ok;

inout  dec_bias, dec_det;

input  testdec_en_b, testdec_prec_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M4 ( .D(dec_det), .B(GND_), .G(testdec_en_b), .S(gnd_));
pch_hvt  M0 ( .D(dec_det), .B(vdd_), .G(testdec_prec_b), .S(vdd_));
inv_hvt I134 ( .A(dec_det), .Y(dec_ok));
nch  M13 ( .D(dec_bias), .B(GND_), .G(testdec_en_b), .S(gnd_));
nch  M6 ( .D(dec_bias), .B(GND_), .G(dec_bias), .S(gnd_));
nch  M7 ( .D(dec_bias_p), .B(GND_), .G(dec_bias), .S(gnd_));
nch  M14 ( .D(ngate), .B(GND_), .G(dec_bias), .S(gnd_));
nch  M15 ( .D(ngate), .B(GND_), .G(testdec_en_b), .S(gnd_));
nch  M10 ( .D(dec_bias_sup), .B(GND_), .G(ngate), .S(dec_bias));
pch  M19 ( .D(ngate), .B(vdd_), .G(testdec_en_b), .S(net76));
pch  M16 ( .D(net76), .B(vdd_), .G(testdec_en_b), .S(vdd_));
pch  M18_1_ ( .D(dec_bias_sup), .B(vdd_), .G(testdec_en_b), .S(vdd_));
pch  M18_0_ ( .D(dec_bias_sup), .B(vdd_), .G(testdec_en_b), .S(vdd_));
pch  M9_2_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));
pch  M9_1_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));
pch  M9_0_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));
pch  M8 ( .D(dec_bias_p), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_yp3_x8, View - schematic
// LAST TIME SAVED: Jul 13 16:32:00 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_yp3_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M17 ( .D(bl[5]), .B(GND_), .G(yp3_25[5]), .S(bl_out));
nch_25  M16 ( .D(bl[6]), .B(GND_), .G(yp3_25[6]), .S(bl_out));
nch_25  M18 ( .D(bl[4]), .B(GND_), .G(yp3_25[4]), .S(bl_out));
nch_25  M19 ( .D(bl[3]), .B(GND_), .G(yp3_25[3]), .S(bl_out));
nch_25  M26 ( .D(bl[0]), .B(GND_), .G(yp3_b_25[0]), .S(vblinhi_rde));
nch_25  M0 ( .D(bl[1]), .B(GND_), .G(yp3_b_25[1]), .S(vblinhi_rdo));
nch_25  M3 ( .D(bl[3]), .B(GND_), .G(yp3_b_25[3]), .S(vblinhi_rdo));
nch_25  M2 ( .D(bl[2]), .B(GND_), .G(yp3_b_25[2]), .S(vblinhi_rde));
nch_25  M4 ( .D(bl[4]), .B(GND_), .G(yp3_b_25[4]), .S(vblinhi_rde));
nch_25  M6 ( .D(bl[5]), .B(GND_), .G(yp3_b_25[5]), .S(vblinhi_rdo));
nch_25  M22 ( .D(bl[0]), .B(GND_), .G(yp3_25[0]), .S(bl_out));
nch_25  M20 ( .D(bl[2]), .B(GND_), .G(yp3_25[2]), .S(bl_out));
nch_25  M21 ( .D(bl[1]), .B(GND_), .G(yp3_25[1]), .S(bl_out));
nch_25  M8 ( .D(bl[7]), .B(GND_), .G(yp3_b_25[7]), .S(vblinhi_rdo));
nch_25  M15 ( .D(bl[7]), .B(GND_), .G(yp3_25[7]), .S(bl_out));
nch_25  M7 ( .D(bl[6]), .B(GND_), .G(yp3_b_25[6]), .S(vblinhi_rde));
pch_25  M5_7_ ( .D(bl[7]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_6_ ( .D(bl[6]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_5_ ( .D(bl[5]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_4_ ( .D(bl[4]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_3_ ( .D(bl[3]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_2_ ( .D(bl[2]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_1_ ( .D(bl[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_0_ ( .D(bl[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));

endmodule
// Library - leafcell, Cell - cfg4pllreset, View - schematic
// LAST TIME SAVED: Jul  7 08:09:12 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module cfg4pllreset ( out, in, prog );
output  out;

input  in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2 I1 ( .A(net012), .B(prog), .Y(net8));
inv I2 ( .A(in), .Y(net012));
inv I3 ( .A(net8), .Y(out));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x8, View - schematic
// LAST TIME SAVED: May  4 13:03:21 2008
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_dummy, View - schematic
// LAST TIME SAVED: Jun 23 14:12:41 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_dummy ( bl_dummyr, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, pgminhi_dmmy_b_25, vdd_tieh );
inout  vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo;

input  pgminhi_dmmy_b_25, vdd_tieh;

inout [1:0]  bl_dummyr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(bl_dummyr[1]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rdo));
nch_25  M2 ( .D(bl_dummyr[0]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rde));
pch_25  M8 ( .D(bl_dummyr[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M0 ( .D(bl_dummyr[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_yp2_8, View - schematic
// LAST TIME SAVED: Jun 23 14:36:38 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_yp2_8 ( bl, bl_out, vblinhi_rde, vblinhi_rdo, yp2,
     yp2_b_25 );
inout  bl_out, vblinhi_rde, vblinhi_rdo;


inout [7:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M6 ( .D(bl[6]), .B(GND_), .G(yp2[6]), .S(bl_out));
nch_hvt  M7 ( .D(bl[7]), .B(GND_), .G(yp2[7]), .S(bl_out));
nch_hvt  M0 ( .D(bl[1]), .B(GND_), .G(yp2[1]), .S(bl_out));
nch_hvt  M5 ( .D(bl[5]), .B(GND_), .G(yp2[5]), .S(bl_out));
nch_hvt  M4 ( .D(bl[4]), .B(GND_), .G(yp2[4]), .S(bl_out));
nch_hvt  M3 ( .D(bl[3]), .B(GND_), .G(yp2[3]), .S(bl_out));
nch_hvt  M2 ( .D(bl[0]), .B(GND_), .G(yp2[0]), .S(bl_out));
nch_hvt  M1 ( .D(bl[2]), .B(GND_), .G(yp2[2]), .S(bl_out));
nch_25  M14 ( .D(bl[7]), .B(GND_), .G(yp2_b_25[7]), .S(vblinhi_rdo));
nch_25  M13 ( .D(bl[6]), .B(GND_), .G(yp2_b_25[6]), .S(vblinhi_rde));
nch_25  M8 ( .D(bl[1]), .B(GND_), .G(yp2_b_25[1]), .S(vblinhi_rdo));
nch_25  M20 ( .D(bl[0]), .B(GND_), .G(yp2_b_25[0]), .S(vblinhi_rde));
nch_25  M12 ( .D(bl[5]), .B(GND_), .G(yp2_b_25[5]), .S(vblinhi_rdo));
nch_25  M11 ( .D(bl[4]), .B(GND_), .G(yp2_b_25[4]), .S(vblinhi_rde));
nch_25  M10 ( .D(bl[3]), .B(GND_), .G(yp2_b_25[3]), .S(vblinhi_rdo));
nch_25  M9 ( .D(bl[2]), .B(GND_), .G(yp2_b_25[2]), .S(vblinhi_rde));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x64, View - schematic
// LAST TIME SAVED: Feb 26 14:34:16 2008
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_x64 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp2, yp2_b_25, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [63:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
input [7:0]  yp3_25;
input [7:0]  yp3_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  bl_med;



ml_ymux_yp2_8 Iml_ymux_yp2_x8 ( .bl(bl_med[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[0]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_2 ( .vdd_tieh(vdd_tieh), .bl(bl[23:16]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[2]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_3 ( .vdd_tieh(vdd_tieh), .bl(bl[31:24]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[3]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_6 ( .vdd_tieh(vdd_tieh), .bl(bl[55:48]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[6]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_7 ( .vdd_tieh(vdd_tieh), .bl(bl[63:56]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[7]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_5 ( .vdd_tieh(vdd_tieh), .bl(bl[47:40]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[5]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_4 ( .vdd_tieh(vdd_tieh), .bl(bl[39:32]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[4]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_1 ( .vdd_tieh(vdd_tieh), .bl(bl[15:8]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[1]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x328_1f, View - schematic
// LAST TIME SAVED: Jan 17 11:59:56 2011
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_x328_1f ( bl, bl_dummyl, bl_dummyr, bl_out, bl_test,
     vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh,
     pgminhi_dmmy_b_25, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test, yp_test_25, yp_test_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25;

inout [327:0]  bl;
inout [1:0]  bl_test;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;

input [7:0]  yp2;
input [7:0]  yp3_b_25;
input [5:0]  yp1_b_25;
input [1:0]  yp_test_b_25;
input [1:0]  yp_test;
input [7:0]  yp2_b_25;
input [1:0]  yp_test_25;
input [5:0]  yp1;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:5]  blx8_out;

wire  [0:4]  blx64_out;



nch_hvt  M21 ( .D(net224), .B(GND_), .G(yp_test[1]), .S(bl_out));
nch_hvt  M19 ( .D(net228), .B(GND_), .G(yp_test[1]), .S(net224));
nch_hvt  M23 ( .D(net232), .B(GND_), .G(yp_test[0]), .S(bl_out));
nch_hvt  M28 ( .D(net236), .B(GND_), .G(yp1[5]), .S(bl_out));
nch_hvt  M0 ( .D(blx64_out[2]), .B(GND_), .G(yp1[2]), .S(bl_out));
nch_hvt  M22 ( .D(net244), .B(GND_), .G(yp_test[0]), .S(net232));
nch_hvt  M24 ( .D(blx64_out[0]), .B(GND_), .G(yp1[0]), .S(bl_out));
nch_hvt  M30 ( .D(blx8_out[5]), .B(GND_), .G(yp1[5]), .S(net236));
nch_hvt  M3 ( .D(blx64_out[4]), .B(GND_), .G(yp1[4]), .S(bl_out));
nch_hvt  M4 ( .D(blx64_out[3]), .B(GND_), .G(yp1[3]), .S(bl_out));
nch_hvt  M2 ( .D(blx64_out[1]), .B(GND_), .G(yp1[1]), .S(bl_out));
pch_25  M7 ( .D(bl_test[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M8 ( .D(bl_test[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
nch_25  M1 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[0]),
     .S(blx64_out[0]));
nch_25  M26 ( .D(vblinhi_rdo), .B(GND_), .G(yp_test_b_25[1]),
     .S(bl_test[1]));
nch_25  M25 ( .D(bl_test[1]), .B(GND_), .G(yp_test_25[1]), .S(net228));
nch_25  M18 ( .D(vblinhi_rde), .B(GND_), .G(yp_test_b_25[0]),
     .S(bl_test[0]));
nch_25  M11 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[5]),
     .S(blx8_out[5]));
nch_25  M17 ( .D(bl_test[0]), .B(GND_), .G(yp_test_25[0]), .S(net244));
nch_25  M6 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[2]),
     .S(blx64_out[2]));
nch_25  M5 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[1]),
     .S(blx64_out[1]));
nch_25  M10 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[4]),
     .S(blx64_out[4]));
nch_25  M9 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[3]),
     .S(blx64_out[3]));
ml_ymux_bls_x8 Iml_ymux_bls_x8 ( .bl_out(blx8_out[5]),
     .bl(bl[327:320]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_r ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyr[1:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_l ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyl[1:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_0 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[0]), .bl(bl[63:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_2 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[2]), .bl(bl[191:128]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_4 ( .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]), .bl(bl[319:256]),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .bl_out(blx64_out[4]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo));
ml_ymux_bls_x64 Iml_ymux_bls_x64_1 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[1]), .bl(bl[127:64]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_3 ( .yp2(yp2[7:0]), .bl_out(blx64_out[3]),
     .bl(bl[255:192]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .yp2_b_25(yp2_b_25[7:0]), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));

endmodule
// Library - tsmcN40, Cell - inv_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:17 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module inv_25 ( OUT, G, Gb, IN, P, Pb );
output  OUT;

input  G, Gb, IN, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(OUT), .B(Gb), .G(IN), .S(G));
pch_25  M1 ( .D(OUT), .B(Pb), .G(IN), .S(P));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_sup_25, View - schematic
// LAST TIME SAVED: Jul 23 11:45:41 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module oai21x2_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
nch_25  M4 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
nch_25  M7 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));
pch_25  M2 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
pch_25  M0 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));
pch_25  M3 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd25_nor2, View - schematic
// LAST TIME SAVED: Sep 14 15:26:13 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ls_vdd25_nor2 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_25 I79 ( .A(in), .Y(out_vddio_b), .Gb(gnd_), .G(gnd_), .Pb(sup),
     .P(sup), .B(out_vddio));
nor2_25 I151 ( .A(out_vddio_b), .Y(out_vddio), .Gb(gnd_), .G(gnd_),
     .Pb(sup), .P(sup), .B(in_b));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yptest, View - schematic
// LAST TIME SAVED: Jul 21 11:48:14 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yptest ( yp_test_25, yp_test_b_25, yp_test,
     yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25, ysup_25 );
output  yp_test_25, yp_test_b_25;

input  yp_test, yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25,
     ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I181 ( .A(yp_test), .Y(net40));
inv_25 I182 ( .IN(net028), .OUT(yp_test_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));
oai21x2_sup_25 I180 ( .A1(yp_test_b_low_ysup_25), .Y(yp_test_b_25),
     .A0(net37), .B0(yp_test_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(yp_test), .sup(ysup_25),
     .out_vddio_b(net028), .out_vddio(net37), .in_b(net40));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_yp3_sup_25, View - schematic
// LAST TIME SAVED: Jul 23 14:26:50 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module oai21x2_yp3_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M12 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
nch_25  M1 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
nch_25  M0 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));
pch_25  M4 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
pch_25  M6 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));
pch_25  M5 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));

endmodule
// Library - leafcell, Cell - delay150to600ps, View - schematic
// LAST TIME SAVED: Apr 24 15:51:58 2009
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module delay150to600ps ( dly600psout, dlyout, cbit, dlyin );
output  dly600psout, dlyout;

input  dlyin;

input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  min;



delay150ps I0 ( .in(dlyin), .out(min[0]));
delay150ps I4 ( .in(min[2]), .out(dly600psout));
delay150ps I3 ( .in(min[1]), .out(min[2]));
delay150ps I2 ( .in(min[0]), .out(min[1]));
mux4plldly I1 ( .min({dly600psout, min[2:0]}), .cbit(cbit[1:0]),
     .mout(dlyout));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yp3, View - schematic
// LAST TIME SAVED: Jul 23 14:27:58 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp3 ( yp3_25, yp3_b_25, yp3_b_high_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, ysup_25 );
output  yp3_25, yp3_b_25;

input  yp3_b_high_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



oai21x2_yp3_sup_25 I209 ( .A1(yp3_b_low_ysup_25), .Y(yp3_b_25),
     .A0(net069), .B0(yp3_b_high_b_ysup_25), .ysup_25(ysup_25));
inv_hvt I201 ( .A(yp3_sel), .Y(net075));
inv_hvt I101 ( .A(net075), .Y(net070));
inv_25 I204 ( .IN(yp3_25_b), .OUT(yp3_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd25_nor2 I192 ( .in(net070), .sup(ysup_25),
     .out_vddio_b(yp3_25_b), .out_vddio(net069), .in_b(net075));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yp21, View - schematic
// LAST TIME SAVED: Jul 21 11:47:41 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp21 ( yp21, yp21_b_25, yp21_b_low_b, yp21_sel,
     ysup_25 );
output  yp21, yp21_b_25;

input  yp21_b_low_b, yp21_sel, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I213 ( .IN(yp21_b_25_b), .OUT(yp21_b_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
nand2_hvt I206 ( .A(yp21_sel_b), .Y(net50), .B(yp21_b_low_b));
inv_hvt I207 ( .A(net50), .Y(net68));
inv_hvt I208 ( .A(yp21_sel), .Y(yp21_sel_b));
inv_hvt I209 ( .A(yp21_sel_b), .Y(yp21));
ml_ls_vdd25_nor2 I194 ( .in(net68), .sup(ysup_25),
     .out_vddio_b(yp21_b_25_b), .out_vddio(net72), .in_b(net50));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_vblinhi_pgm_drv, View -
//schematic
// LAST TIME SAVED: Jul 29 15:49:55 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_vblinhi_pgm_drv ( vblinhi_pgm_25, ysup_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25 );
inout  vblinhi_pgm_25, ysup_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd_), .B(GND_), .G(en_blinhi_pgm_b_ysup_25),
     .S(vblinhi_pgm_25));
pch_25  M5 ( .D(net10), .B(ysup_25), .G(en_blinhi_pgm_b_ysup_25),
     .S(ysup_25));
pch_25  M0 ( .D(net10), .B(vblinhi_pgm_25), .G(en_blinhi_pgm_b),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_1f, View - schematic
// LAST TIME SAVED: Dec 28 15:35:42 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_1f ( yp1, yp1_b_25, yp2, yp2_b_25, yp3_25,
     yp3_b_25, yp_test_25, yp_test_b_25, vblinhi_pgm_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b, yp1_sel,
     yp2_b_low_b, yp2_sel, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, yp_test,
     ysup_25 );

inout  vblinhi_pgm_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b,
     yp2_b_low_b, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, ysup_25;

output [7:0]  yp3_b_25;
output [7:0]  yp3_25;
output [7:0]  yp2;
output [5:0]  yp1;
output [1:0]  yp_test_25;
output [1:0]  yp_test_b_25;
output [7:0]  yp2_b_25;
output [5:0]  yp1_b_25;

input [7:0]  yp3_sel;
input [5:0]  yp1_sel;
input [7:0]  yp2_sel;
input [1:0]  yp_test;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_1_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1]), .yp_test(yp_test[1]),
     .yp_test_25(yp_test_25[1]));
ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_0_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[0]), .yp_test(yp_test[0]),
     .yp_test_25(yp_test_25[0]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_7_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[7]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[7]), .yp3_25(yp3_25[7]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_6_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[6]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[6]), .yp3_25(yp3_25[6]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_5_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[5]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[5]), .yp3_25(yp3_25[5]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_4_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[4]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[4]), .yp3_25(yp3_25[4]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_3_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[3]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[3]), .yp3_25(yp3_25[3]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_2_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[2]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[2]), .yp3_25(yp3_25[2]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_1_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[1]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[1]), .yp3_25(yp3_25[1]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_0_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[0]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[0]), .yp3_25(yp3_25[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_7_ ( .yp21_sel(yp2_sel[7]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[7]), .yp21(yp2[7]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_6_ ( .yp21_sel(yp2_sel[6]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[6]), .yp21(yp2[6]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_5_ ( .yp21_sel(yp2_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[5]), .yp21(yp2[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_4_ ( .yp21_sel(yp2_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[4]), .yp21(yp2[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_3_ ( .yp21_sel(yp2_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[3]), .yp21(yp2[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_2_ ( .yp21_sel(yp2_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[2]), .yp21(yp2[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_1_ ( .yp21_sel(yp2_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[1]), .yp21(yp2[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_0_ ( .yp21_sel(yp2_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[0]), .yp21(yp2[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_5_ ( .yp21_sel(yp1_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[5]), .yp21(yp1[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_4_ ( .yp21_sel(yp1_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[4]), .yp21(yp1[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_3_ ( .yp21_sel(yp1_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[3]), .yp21(yp1[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_2_ ( .yp21_sel(yp1_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[2]), .yp21(yp1[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_1_ ( .yp21_sel(yp1_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[1]), .yp21(yp1[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_0_ ( .yp21_sel(yp1_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[0]), .yp21(yp1[0]));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_1_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_0_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_a_clkdly, View - schematic
// LAST TIME SAVED: Jul 15 18:44:33 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_pump_a_clkdly ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I206 ( .A(in), .Y(net66));
inv_hvt I205 ( .A(net66), .Y(net70));
inv_hvt I207 ( .A(net70), .Y(out));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(net66), .S(vdd_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_logic_8f_sbb, View -
//schematic
// LAST TIME SAVED: Jul 15 18:44:43 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_8f_sbb ( out_hv_winv, out_hv_woinv, in );
output  out_hv_winv, out_hv_woinv;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_pump_a_clkdly I141 ( .in(net262), .out(net270));
ml_pump_a_clkdly I219 ( .in(net266), .out(net268));
ml_ls_vdd2vdd25 I144 ( .in(net266), .sup(vddp_),
     .out_vddio_b(out_hv_winv), .out_vddio(net279), .in_b(net258));
ml_ls_vdd2vdd25 I148 ( .in(net262), .sup(vddp_),
     .out_vddio_b(out_hv_woinv), .out_vddio(net274), .in_b(net255));
nor2_hvt I140 ( .A(net268), .B(in), .Y(net255));
nor2_hvt I227 ( .A(net264), .B(net270), .Y(net258));
inv_hvt I225 ( .A(net258), .Y(net266));
inv_hvt I134 ( .A(in), .Y(net264));
inv_hvt I226 ( .A(net255), .Y(net262));

endmodule
// Library - sbtlibn65lp, Cell - oai2211x2_hvt, View - schematic
// LAST TIME SAVED: Jul 23 15:48:12 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module oai2211x2_hvt ( Y, A0, A1, B0, B1, C0, D0 );
output  Y;

input  A0, A1, B0, B1, C0, D0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M10 ( .D(net040), .B(GND_), .G(A1), .S(net024));
nch_hvt  M13 ( .D(net040), .B(GND_), .G(A0), .S(net024));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
nch_hvt  M11 ( .D(Y), .B(GND_), .G(C0), .S(net044));
nch_hvt  M0 ( .D(net044), .B(GND_), .G(D0), .S(net040));
nch_hvt  M1 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
pch_hvt  M12 ( .D(Y), .B(VDD_), .G(D0), .S(vdd_));
pch_hvt  M2 ( .D(Y), .B(VDD_), .G(C0), .S(vdd_));
pch_hvt  M18 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M8 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M19 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M7 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - sbtlibn65lp, Cell - anor31_hvt, View - schematic
// LAST TIME SAVED: Jul 23 15:32:42 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module anor31_hvt ( Y, A, B, C, D );
output  Y;

input  A, B, C, D;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(Y), .B(gnd_), .G(A), .S(net23));
nch_hvt  M6 ( .D(net030), .B(gnd_), .G(C), .S(gnd_));
nch_hvt  M5 ( .D(net23), .B(gnd_), .G(B), .S(net030));
nch_hvt  M7 ( .D(Y), .B(gnd_), .G(D), .S(gnd_));
pch_hvt  M3 ( .D(Y), .B(vdd_), .G(D), .S(net35));
pch_hvt  M4 ( .D(net35), .B(vdd_), .G(A), .S(vdd_));
pch_hvt  M0 ( .D(net35), .B(vdd_), .G(B), .S(vdd_));
pch_hvt  M2 ( .D(net35), .B(vdd_), .G(C), .S(vdd_));

endmodule
// Library - sbtlibn65lp, Cell - oai22x2_hvt, View - schematic
// LAST TIME SAVED: Jul 23 15:55:46 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module oai22x2_hvt ( Y, A0, A1, B0, B1 );
output  Y;

input  A0, A1, B0, B1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(Y), .B(GND_), .G(A0), .S(net024));
nch_hvt  M4 ( .D(Y), .B(GND_), .G(A1), .S(net024));
nch_hvt  M1 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M0 ( .D(Y), .B(VDD_), .G(A0), .S(net017));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_logic_1f, View - schematic
// LAST TIME SAVED: Dec 30 13:06:02 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_1f ( dec_trim, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, s_rd, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25, yp1_sel,
     yp2_sel, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, yp21_b_low_b, yp_test, vdd_tieh,
     fsm_blkadd, fsm_coladd, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     tm_allbank_sel, tm_tcol, ysup_25 );
output  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp21_b_low_b;

inout  vdd_tieh;

input  fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h,
     fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec,
     fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis, tm_allbank_sel,
     tm_tcol, ysup_25;

output [3:0]  sb25_high_25;
output [3:0]  sb25_gnd_25;
output [7:0]  yp3_sel;
output [3:0]  sbhv_high_25;
output [7:5]  dec_trim;
output [7:0]  yp2_sel;
output [5:0]  yp1_sel;
output [3:0]  s_rd;
output [3:0]  sbhv_gnd_25;
output [1:0]  yp_test;

input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefpgm;
input [9:0]  fsm_coladd;
input [1:0]  fsm_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp2_sel_b;

wire  [7:0]  yp3_sel_b;

wire  [7:5]  dec_trim_b;

wire  [3:0]  sb25low_b;

wire  [5:0]  yp1_sel_b;

wire  [1:0]  yp_test_b;

wire  [3:0]  s_rd_b;

wire  [2:0]  tdec;

wire  [3:0]  sbhvlow_b;

wire  [1:0]  xadd_b;

wire  [1:0]  xadd;

wire  [0:9]  yadd;

wire  [0:9]  yadd_b;

wire  [0:3]  net561;

wire  [2:0]  tdec_b;



inv_25 I104 ( .IN(net302), .OUT(en_blinhi_pgm_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I285 ( .IN(net311), .OUT(yp3_b_low_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I284 ( .IN(net306), .OUT(yp3_b_high_odd_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I283 ( .IN(net316), .OUT(yp3_b_high_even_b_ysup_25),
     .P(ysup_25), .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
ml_core_ctrl_logic_8f_sbb Isb25_3_ ( .in(sb25low_b[3]),
     .out_hv_woinv(sb25_gnd_25[3]), .out_hv_winv(sb25_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isb25_2_ ( .in(sb25low_b[2]),
     .out_hv_woinv(sb25_gnd_25[2]), .out_hv_winv(sb25_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isb25_1_ ( .in(sb25low_b[1]),
     .out_hv_woinv(sb25_gnd_25[1]), .out_hv_winv(sb25_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isb25_0_ ( .in(sb25low_b[0]),
     .out_hv_woinv(sb25_gnd_25[0]), .out_hv_winv(sb25_high_25[0]));
ml_core_ctrl_logic_8f_sbb Isbhv_3_ ( .in(sbhvlow_b[3]),
     .out_hv_woinv(sbhv_gnd_25[3]), .out_hv_winv(sbhv_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isbhv_2_ ( .in(sbhvlow_b[2]),
     .out_hv_woinv(sbhv_gnd_25[2]), .out_hv_winv(sbhv_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isbhv_1_ ( .in(sbhvlow_b[1]),
     .out_hv_woinv(sbhv_gnd_25[1]), .out_hv_winv(sbhv_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isbhv_0_ ( .in(sbhvlow_b[0]),
     .out_hv_woinv(sbhv_gnd_25[0]), .out_hv_winv(sbhv_high_25[0]));
ml_ls_vdd25_nor2 I106 ( .in(net343), .sup(ysup_25),
     .out_vddio_b(net301), .out_vddio(net302), .in_b(en_blinhi_pgm_b));
ml_ls_vdd25_nor2 I68 ( .in(net576), .sup(ysup_25),
     .out_vddio_b(net306), .out_vddio(net307), .in_b(net308));
ml_ls_vdd25_nor2 I192 ( .in(net396), .sup(ysup_25),
     .out_vddio_b(net311), .out_vddio(net312), .in_b(net544));
ml_ls_vdd25_nor2 I65 ( .in(net571), .sup(ysup_25),
     .out_vddio_b(net316), .out_vddio(net317), .in_b(net318));
exor2_hvt I151_3_ ( .A(net561[0]), .Y(sb25low_b[3]), .B(pgm_hvact_b));
exor2_hvt I151_2_ ( .A(net561[1]), .Y(sb25low_b[2]), .B(pgm_hvact_b));
exor2_hvt I151_1_ ( .A(net561[2]), .Y(sb25low_b[1]), .B(pgm_hvact_b));
exor2_hvt I151_0_ ( .A(net561[3]), .Y(sb25low_b[0]), .B(pgm_hvact_b));
mux2_hvt I152 ( .in1(net504), .in0(net514), .out(ensb25_dec),
     .sel(pgm_hvact));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(tdec[2]), .sel(ref_pgm));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(tdec[1]), .sel(ref_pgm));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(tdec[0]), .sel(ref_pgm));
oai21x2_hvt I55 ( .A1(sa_bl_to_blsa), .Y(net331), .A0(blk_dec),
     .B0(ymux_dis_b));
nor3_hvt I324 ( .B(fsm_tm_testdec), .Y(net335), .A(fsm_tm_allbl_l),
     .C(fsm_tm_allbl_h));
nor3_hvt I321 ( .B(fsm_tm_allbl_h), .Y(net339), .A(nvcmen_buf_b),
     .C(yp3_b_high_b));
nor4_hvt I326 ( .B(fsm_tm_allbl_l), .Y(net343), .D(nvcmen_buf_b),
     .A(net384), .C(fsm_tm_allbl_l));
nor4_hvt I327 ( .B(fsm_tm_allbl_h), .Y(ymux_dis_b), .D(net405),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_h));
nand3_hvt I227 ( .Y(net352), .B(pgm_hvact), .C(fsm_tm_allwl_h),
     .A(fsm_lshven));
nand3_hvt I236_3_ ( .Y(s_rd_b[3]), .B(xadd[0]), .C(en_rdp),
     .A(xadd[1]));
nand3_hvt I236_2_ ( .Y(s_rd_b[2]), .B(xadd_b[0]), .C(en_rdp),
     .A(xadd[1]));
nand3_hvt I236_1_ ( .Y(s_rd_b[1]), .B(xadd[0]), .C(en_rdp),
     .A(xadd_b[1]));
nand3_hvt I236_0_ ( .Y(s_rd_b[0]), .B(xadd_b[0]), .C(en_rdp),
     .A(xadd_b[1]));
nand3_hvt I230 ( .Y(pgm_hvact_b), .B(fsm_pgm), .C(net502),
     .A(fsm_lshven));
nand3_hvt I232 ( .Y(net364), .B(sa_bl_to_blsa), .C(tm_allwl_l_b),
     .A(fsm_vpxaset));
nand3_hvt I233 ( .Y(net368), .B(net492), .C(nvcmen_buf), .A(net387));
nand3_hvt I234_7_ ( .Y(dec_trim_b[7]), .B(tdec[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I234_6_ ( .Y(dec_trim_b[6]), .B(tdec[1]), .C(tdec_b[0]),
     .A(tdec[2]));
nand3_hvt I234_5_ ( .Y(dec_trim_b[5]), .B(tdec_b[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I231_7_ ( .Y(yp2_sel_b[7]), .B(yadd[4]), .C(yadd[3]),
     .A(yadd[5]));
nand3_hvt I231_6_ ( .Y(yp2_sel_b[6]), .B(yadd[4]), .C(yadd_b[3]),
     .A(yadd[5]));
nand3_hvt I231_5_ ( .Y(yp2_sel_b[5]), .B(yadd_b[4]), .C(yadd[3]),
     .A(yadd[5]));
nand3_hvt I231_4_ ( .Y(yp2_sel_b[4]), .B(yadd_b[4]), .C(yadd_b[3]),
     .A(yadd[5]));
nand3_hvt I231_3_ ( .Y(yp2_sel_b[3]), .B(yadd[4]), .C(yadd[3]),
     .A(yadd_b[5]));
nand3_hvt I231_2_ ( .Y(yp2_sel_b[2]), .B(yadd[4]), .C(yadd_b[3]),
     .A(yadd_b[5]));
nand3_hvt I231_1_ ( .Y(yp2_sel_b[1]), .B(yadd_b[4]), .C(yadd[3]),
     .A(yadd_b[5]));
nand3_hvt I231_0_ ( .Y(yp2_sel_b[0]), .B(yadd_b[4]), .C(yadd_b[3]),
     .A(yadd_b[5]));
nand2_hvt I299 ( .A(fsm_tm_rd_mode), .Y(one_blk_sel_b), .B(blk_dec));
nand2_hvt I301 ( .A(pgm_hvact), .Y(net384), .B(pgm_hvact));
nand2_hvt I293 ( .A(fsm_lshven), .Y(net387), .B(pgm_hvact));
nand2_hvt I297 ( .A(blk_dec_b), .Y(blk_dec), .B(tm_pgm_rd_allblk_n));
nand2_hvt I296 ( .A(blk_dec), .Y(net393), .B(fsm_pgmien));
nand2_hvt I294 ( .A(net387), .Y(net396), .B(net335));
nand2_hvt I298 ( .A(all_blk_sel_b), .Y(sa_bl_to_blsa),
     .B(one_blk_sel_b));
nand2_hvt I300 ( .A(tm_allwl_l_b), .Y(net503), .B(blk_dec));
nand2_hvt I295 ( .A(fsm_nvcmen), .Y(net405), .B(fsm_lshven));
nand2_hvt I291_1_ ( .A(yadd[0]), .Y(yp_test_b[1]), .B(ymux_test_en));
nand2_hvt I291_0_ ( .A(yadd_b[0]), .Y(yp_test_b[0]), .B(ymux_test_en));
nand2_hvt I245 ( .A(rd_and_vfy), .Y(all_blk_sel_b), .B(net536));
nand4_hvt I306 ( .D(fsm_blkadd[0]), .A(fsm_blkadd[3]),
     .C(fsm_blkadd[1]), .Y(blk_dec_b), .B(fsm_blkadd[2]));
nand4_hvt I307_5_ ( .D(yadd[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[5]), .B(yadd[8]));
nand4_hvt I307_4_ ( .D(yadd_b[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[4]), .B(yadd[8]));
nand4_hvt I304_7_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[7]), .B(yadd[2]));
nand4_hvt I304_6_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[6]), .B(yadd[2]));
nand4_hvt I304_5_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[5]), .B(yadd[2]));
nand4_hvt I304_4_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[4]), .B(yadd[2]));
nand4_hvt I304_3_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[3]), .B(yadd_b[2]));
nand4_hvt I304_2_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[2]), .B(yadd_b[2]));
nand4_hvt I304_1_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[1]), .B(yadd_b[2]));
nand4_hvt I304_0_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[0]), .B(yadd_b[2]));
nand4_hvt I239 ( .D(fsm_tm_rprd), .Y(net429), .B(fsm_lshven),
     .C(nvcmen_buf), .A(rd_and_vfy));
nand4_hvt I308 ( .D(fsm_lshven), .A(tm_allwl_l_b), .C(pgm_hvact),
     .Y(net436), .B(blk_dec));
nor2_hvt I316_5_ ( .A(yp1_sel_b[5]), .B(tm_tcol), .Y(yp1_sel[5]));
nor2_hvt I316_4_ ( .A(yp1_sel_b[4]), .B(tm_tcol), .Y(yp1_sel[4]));
nor2_hvt I310 ( .A(fsm_pgmvfy), .B(fsm_pgm), .Y(net443));
nor2_hvt I315 ( .A(net331), .B(net530), .Y(ymux_test_en));
nor2_hvt I312 ( .A(net579), .B(net532), .Y(net449));
nor2_hvt I319 ( .A(fsm_rd), .B(fsm_pgmvfy), .Y(net452));
nor2_hvt I328 ( .A(net331), .B(tm_tcol), .Y(ymux_en_core));
nor2_hvt I317_3_ ( .A(yp1_sel_b[3]), .B(tm_tcol), .Y(yp1_sel[3]));
nor2_hvt I317_2_ ( .A(yp1_sel_b[2]), .B(tm_tcol), .Y(yp1_sel[2]));
nor2_hvt I317_1_ ( .A(yp1_sel_b[1]), .B(tm_tcol), .Y(yp1_sel[1]));
nor2_hvt I317_0_ ( .A(yp1_sel_b[0]), .B(tm_tcol), .Y(yp1_sel[0]));
nor2_hvt I313 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I318 ( .A(fsm_tm_rd_mode), .B(fsm_pgmvfy), .Y(net464));
anor21_hvt I119_1_ ( .A(fsm_rowadd[1]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I119_0_ ( .A(fsm_rowadd[0]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
anor21_hvt I109 ( .A(pgm_hvact), .B(fsm_tm_allwl_h), .Y(net505),
     .C(nvcmen_buf_b));
inv_hvt I271_9_ ( .A(yadd[9]), .Y(yadd_b[9]));
inv_hvt I272_9_ ( .A(vdd_tieh), .Y(yadd[9]));
inv_hvt I247 ( .A(net452), .Y(rd_and_vfy));
inv_hvt I265 ( .A(net464), .Y(net484));
inv_hvt I323 ( .A(fsm_tm_allbl_l), .Y(yp3_b_high_b));
inv_hvt I237_3_ ( .A(s_rd_b[3]), .Y(s_rd[3]));
inv_hvt I237_2_ ( .A(s_rd_b[2]), .Y(s_rd[2]));
inv_hvt I237_1_ ( .A(s_rd_b[1]), .Y(s_rd[1]));
inv_hvt I237_0_ ( .A(s_rd_b[0]), .Y(s_rd[0]));
inv_hvt I252_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I252_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I200 ( .A(fsm_tm_testdec), .Y(net492));
inv_hvt I261 ( .A(net393), .Y(sa_bl_to_pgm_glb));
inv_hvt I271_8_ ( .A(yadd_b[8]), .Y(yadd[8]));
inv_hvt I271_7_ ( .A(yadd_b[7]), .Y(yadd[7]));
inv_hvt I271_6_ ( .A(yadd_b[6]), .Y(yadd[6]));
inv_hvt I271_5_ ( .A(yadd_b[5]), .Y(yadd[5]));
inv_hvt I271_4_ ( .A(yadd_b[4]), .Y(yadd[4]));
inv_hvt I271_3_ ( .A(yadd_b[3]), .Y(yadd[3]));
inv_hvt I271_2_ ( .A(yadd_b[2]), .Y(yadd[2]));
inv_hvt I271_1_ ( .A(yadd_b[1]), .Y(yadd[1]));
inv_hvt I271_0_ ( .A(yadd_b[0]), .Y(yadd[0]));
inv_hvt I268 ( .A(net579), .Y(vddp_rd_overw));
inv_hvt I260 ( .A(nvcmen_buf_b), .Y(nvcmen_buf));
inv_hvt I254 ( .A(net576), .Y(net308));
inv_hvt I278 ( .A(fsm_pgmvfy), .Y(net502));
inv_hvt I281 ( .A(net503), .Y(net504));
inv_hvt I279 ( .A(net505), .Y(net506));
inv_hvt I251 ( .A(net352), .Y(net508));
inv_hvt I258 ( .A(net368), .Y(yp21_b_low_b));
inv_hvt I263 ( .A(fsm_nvcmen), .Y(nvcmen_buf_b));
inv_hvt I280 ( .A(net364), .Y(net514));
inv_hvt I264 ( .A(tm_allbank_sel), .Y(tm_pgm_rd_allblk_n));
inv_hvt I250 ( .A(net436), .Y(net518));
inv_hvt I241 ( .A(net429), .Y(en_rdp));
inv_hvt I255 ( .A(net343), .Y(en_blinhi_pgm_b));
inv_hvt I249 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I277 ( .A(pgm_hvact_b), .Y(pgm_hvact));
inv_hvt I266 ( .A(net443), .Y(ref_pgm));
inv_hvt I259 ( .A(tm_tcol), .Y(net530));
inv_hvt I267 ( .A(fsm_multibl_read), .Y(net532));
inv_hvt I262 ( .A(all_blk_sel_b), .Y(net534));
inv_hvt I272_8_ ( .A(fsm_coladd[8]), .Y(yadd_b[8]));
inv_hvt I272_7_ ( .A(fsm_coladd[7]), .Y(yadd_b[7]));
inv_hvt I272_6_ ( .A(fsm_coladd[6]), .Y(yadd_b[6]));
inv_hvt I272_5_ ( .A(fsm_coladd[5]), .Y(yadd_b[5]));
inv_hvt I272_4_ ( .A(fsm_coladd[4]), .Y(yadd_b[4]));
inv_hvt I272_3_ ( .A(fsm_coladd[3]), .Y(yadd_b[3]));
inv_hvt I272_2_ ( .A(fsm_coladd[2]), .Y(yadd_b[2]));
inv_hvt I272_1_ ( .A(fsm_coladd[1]), .Y(yadd_b[1]));
inv_hvt I272_0_ ( .A(fsm_coladd[0]), .Y(yadd_b[0]));
inv_hvt I201 ( .A(fsm_tm_rd_mode), .Y(net536));
inv_hvt I270_2_ ( .A(tdec[2]), .Y(tdec_b[2]));
inv_hvt I270_1_ ( .A(tdec[1]), .Y(tdec_b[1]));
inv_hvt I270_0_ ( .A(tdec[0]), .Y(tdec_b[0]));
inv_hvt I273_7_ ( .A(yp2_sel_b[7]), .Y(yp2_sel[7]));
inv_hvt I273_6_ ( .A(yp2_sel_b[6]), .Y(yp2_sel[6]));
inv_hvt I273_5_ ( .A(yp2_sel_b[5]), .Y(yp2_sel[5]));
inv_hvt I273_4_ ( .A(yp2_sel_b[4]), .Y(yp2_sel[4]));
inv_hvt I273_3_ ( .A(yp2_sel_b[3]), .Y(yp2_sel[3]));
inv_hvt I273_2_ ( .A(yp2_sel_b[2]), .Y(yp2_sel[2]));
inv_hvt I273_1_ ( .A(yp2_sel_b[1]), .Y(yp2_sel[1]));
inv_hvt I273_0_ ( .A(yp2_sel_b[0]), .Y(yp2_sel[0]));
inv_hvt I256_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I256_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I256_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I257 ( .A(net396), .Y(net544));
inv_hvt I274_7_ ( .A(yp3_sel_b[7]), .Y(yp3_sel[7]));
inv_hvt I274_6_ ( .A(yp3_sel_b[6]), .Y(yp3_sel[6]));
inv_hvt I274_5_ ( .A(yp3_sel_b[5]), .Y(yp3_sel[5]));
inv_hvt I274_4_ ( .A(yp3_sel_b[4]), .Y(yp3_sel[4]));
inv_hvt I274_3_ ( .A(yp3_sel_b[3]), .Y(yp3_sel[3]));
inv_hvt I274_2_ ( .A(yp3_sel_b[2]), .Y(yp3_sel[2]));
inv_hvt I274_1_ ( .A(yp3_sel_b[1]), .Y(yp3_sel[1]));
inv_hvt I274_0_ ( .A(yp3_sel_b[0]), .Y(yp3_sel[0]));
inv_hvt I253 ( .A(net571), .Y(net318));
inv_hvt I275_1_ ( .A(yp_test_b[1]), .Y(yp_test[1]));
inv_hvt I275_0_ ( .A(yp_test_b[0]), .Y(yp_test[0]));
oai2211x2_hvt I86_3_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[3]), .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai2211x2_hvt I86_2_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[2]), .A0(yadd[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
oai2211x2_hvt I86_1_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[1]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd[6]));
oai2211x2_hvt I86_0_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[0]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
anor31_hvt I155_3_ ( .A(ensb25_dec), .D(net506), .B(xadd[1]),
     .Y(net561[0]), .C(xadd[0]));
anor31_hvt I155_2_ ( .A(ensb25_dec), .D(net506), .B(xadd[1]),
     .Y(net561[1]), .C(xadd_b[0]));
anor31_hvt I155_1_ ( .A(ensb25_dec), .D(net506), .B(xadd_b[1]),
     .Y(net561[2]), .C(xadd[0]));
anor31_hvt I155_0_ ( .A(ensb25_dec), .D(net506), .B(xadd_b[1]),
     .Y(net561[3]), .C(xadd_b[0]));
anor31_hvt I121_3_ ( .A(net518), .D(net508), .B(xadd[1]),
     .Y(sbhvlow_b[3]), .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net518), .D(net508), .B(xadd[1]),
     .Y(sbhvlow_b[2]), .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net518), .D(net508), .B(xadd_b[1]),
     .Y(sbhvlow_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net518), .D(net508), .B(xadd_b[1]),
     .Y(sbhvlow_b[0]), .C(xadd_b[0]));
anor31_hvt I107 ( .A(fsm_tm_testdec), .D(net339), .B(nvcmen_buf),
     .Y(net571), .C(yadd[0]));
anor31_hvt I108 ( .A(fsm_tm_testdec), .D(net339), .B(nvcmen_buf),
     .Y(net576), .C(yadd_b[0]));
oai22x2_hvt I93 ( .A1(net534), .Y(net579), .A0(net484),
     .B0(fsm_nv_rri_trim), .B1(fsm_nv_sisi_ui));

endmodule
// Library - leafcell, Cell - pll_finedly, View - schematic
// LAST TIME SAVED: May 11 17:26:27 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pll_finedly ( pll_fbout, cbit, pll_fbin );
output  pll_fbout;

input  pll_fbin;

input [3:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  min;



delay150to600ps I6 ( .dly600psout(net40), .cbit(cbit[1:0]),
     .dlyin(net44), .dlyout(min[2]));
delay150to600ps I5 ( .dly600psout(net44), .cbit(cbit[1:0]),
     .dlyin(net52), .dlyout(min[1]));
delay150to600ps I4 ( .dly600psout(net48), .cbit(cbit[1:0]),
     .dlyin(net40), .dlyout(min[3]));
delay150to600ps I0 ( .dly600psout(net52), .cbit(cbit[1:0]),
     .dlyin(pll_fbin), .dlyout(min[0]));
mux4plldly I1 ( .min(min[3:0]), .cbit(cbit[3:2]), .mout(pll_fbout));

endmodule
// Library - ice1chip, Cell - pll_bufwrap_ice1f, View - schematic
// LAST TIME SAVED: Apr  8 12:23:22 2011
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pll_bufwrap_ice1f ( f_out, f_in );
output  f_out;

input  f_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



fabric_buf_ice8p I6 ( .f_in(f_in), .f_out(f_out));

endmodule
// Library - NVCM_40nm, Cell - ml_dff_nvcm, View - schematic
// LAST TIME SAVED: Jun 21 11:02:43 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_dff_nvcm ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I132 ( .A(clk_b), .Y(clk_buf));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I146 ( .A(net57), .Y(Q));
inv_hvt I147 ( .A(net60), .Y(QN));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net64), .Y(net57));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net64), .Y(net53));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net60), .Y(net57));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net53));
nor2_hvt I129 ( .A(net57), .B(R), .Y(net60));
nor2_hvt I125 ( .A(net53), .B(R), .Y(net64));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_resref_40nm, View - schematic
// LAST TIME SAVED: Sep 11 14:49:31 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_sa_resref_40nm ( bl_in, bl_out, ref );
inout  bl_in, bl_out;

inout [3:0]  ref;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R9 ( .MINUS(ref[3]), .PLUS(ref[2]), .BULK(gnd_));
rppolywo_m  R11 ( .MINUS(ref[1]), .PLUS(ref[0]), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(net41), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(ref[2]), .PLUS(ref[1]), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(ref[0]), .PLUS(net41), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(ref[3]), .BULK(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_restop_40nm, View - schematic
// LAST TIME SAVED: Sep 16 19:06:55 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_sa_restop_40nm ( bl_bot, bl_top );
inout  bl_bot, bl_top;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R24 ( .MINUS(bl_top), .PLUS(net66), .BULK(gnd_));
rppolywo_m  R23 ( .MINUS(net66), .PLUS(bl_bot), .BULK(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_resbot_40nm, View - schematic
// LAST TIME SAVED: Sep 16 11:24:37 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_sa_resbot_40nm ( bl_in, bl_out, in_dec, sa_ngate );
inout  bl_in, bl_out, in_dec;


input [4:1]  sa_ngate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M9 ( .D(net026), .B(GND_), .G(sa_ngate[2]), .S(gnd_));
nch_hvt  M20 ( .D(in_dec), .B(GND_), .G(sa_ngate[1]), .S(gnd_));
nch_hvt  M10 ( .D(net072), .B(GND_), .G(sa_ngate[3]), .S(gnd_));
nch_hvt  M11 ( .D(net132), .B(GND_), .G(sa_ngate[4]), .S(gnd_));
rppolywo_m  R15 ( .MINUS(bl_in), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(bl_in), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(net026), .PLUS(in_dec), .BULK(gnd_));
rppolywo_m  R12 ( .MINUS(bl_in), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(in_dec), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R9 ( .MINUS(bl_out), .PLUS(net132), .BULK(gnd_));
rppolywo_m  R8 ( .MINUS(net072), .PLUS(net026), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(net132), .PLUS(net072), .BULK(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_gwlgnd_nor2, View - schematic
// LAST TIME SAVED: Jul 10 13:02:38 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_gwlgnd_nor2 ( gwl_gnd_25, gwl_b_sup_25, gwl_b_25,
     gwl_b_gnden_25 );
output  gwl_gnd_25;

inout  gwl_b_sup_25;

input  gwl_b_25, gwl_b_gnden_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(net14), .B(GND_), .G(gwl_b_gnden_25), .S(GND_));
nch_25  M0 ( .D(gwl_gnd_25), .B(GND_), .G(gwl_b_25), .S(net14));
pch_25  M2 ( .D(gwl_gnd_25), .B(gwl_b_sup_25), .G(gwl_b_25),
     .S(gwl_b_sup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp, View - schematic
// LAST TIME SAVED: Nov 30 17:03:56 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp ( wp, gwl_gnd_rp_25, ngate_25, gwl_b_25,
     gwl_gnd_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv );
output  wp;

inout  gwl_gnd_rp_25, ngate_25;

input  gwl_b_25, gwl_gnd_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M11 ( .D(net18), .B(GND_), .G(s_b_25), .S(gwl_gnd_25));
nch_25  M12 ( .D(wp), .B(GND_), .G(ngate_25), .S(net18));
nch_25  M10 ( .D(net18), .B(GND_), .G(gwl_b_25), .S(gwl_gnd_25));
pch_25  M0 ( .D(gwl_gnd_rp_25), .B(gwp_hv), .G(s_rd_b_hv), .S(wp));
pch_25  M6 ( .D(wp), .B(gwp_hv), .G(s_b_hv), .S(gwp_hv));

endmodule
// Library - tsmcN40, Cell - nand2_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:22 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nand2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(Y), .B(Gb), .G(A), .S(net16));
nch_25  M3 ( .D(net16), .B(Gb), .G(B), .S(G));
pch_25  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M2 ( .D(Y), .B(Pb), .G(B), .S(P));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp, View - schematic
// LAST TIME SAVED: Aug 27 14:09:22 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_b_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(out_ref), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M2 ( .D(out_div), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M8 ( .D(out_ref), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M5 ( .D(out_div), .B(GND_), .G(saen_b_25), .S(gnd_));
pch_25  M4_1_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M3 ( .D(out_ref), .B(vddp_), .G(in_ref), .S(net65));
pch_25  M6 ( .D(out_div), .B(vddp_), .G(in_div), .S(net65));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_top, View - schematic
// LAST TIME SAVED: Sep 15 18:21:46 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp_top ( sa_out, vdd_tieh, in_div, in_ref, saen_25
     );
output  sa_out;

inout  vdd_tieh;

input  in_div, in_ref, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M6 ( .D(sa_out_b_25), .B(gnd_), .G(saen_b_25), .S(gnd_));
nch_25  M0 ( .D(net053), .B(gnd_), .G(saen_25), .S(gnd_));
nch_25  M5 ( .D(sa_out_b_25), .B(gnd_), .G(out_div2), .S(gnd_));
nch_25  M1 ( .D(sa_bias), .B(gnd_), .G(vdd_tieh), .S(net45));
rppolywo_m  R0 ( .MINUS(net039), .PLUS(net45), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net053), .PLUS(net039), .BULK(gnd_));
pch_25  M43 ( .D(sa_bias), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M4_1_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M7 ( .D(sa_out_b_25), .B(vddp_), .G(out_div2), .S(net089));
pch_25  M3 ( .D(net089), .B(vddp_), .G(sa_bias), .S(vddp_));
nand2_25 I80 ( .G(gnd_), .Pb(vdd_), .A(net051), .Y(net038), .P(vdd_),
     .B(saen_25), .Gb(gnd_));
inv_25 I89 ( .IN(sa_out_b_25), .OUT(net051), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I91 ( .IN(saen_25), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net038), .OUT(sa_out), .P(vdd_), .Pb(vdd_), .G(gnd_),
     .Gb(gnd_));
ml_core_sa_comp Icore_sa_comp0 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp Icore_sa_comp1 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref2), .in_div(in_div2),
     .out_ref(out_ref), .out_div(out_div2));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa, View - schematic
// LAST TIME SAVED: Jun 17 16:48:48 2011
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_sa ( nv_dataout, blsa, vdd_tieh, vddp_tieh, vpxa,
     dec_ok, dec_trim, fsm_rst_b, fsm_sample, fsm_tm_ref,
     fsm_tm_testdec, sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, tm_testdec_wr );
output  nv_dataout;

inout  blsa, vdd_tieh, vddp_tieh, vpxa;

input  dec_ok, fsm_rst_b, fsm_sample, fsm_tm_testdec, saen_25,
     saen_b_vpxa, saprd_b_vpxa, testdec_en_b, tm_testdec_wr;

input [7:5]  dec_trim;
input [1:0]  fsm_tm_ref;
input [4:1]  sa_ngate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  ref;



nmoscap_25  C0 ( .MINUS(GND_), .PLUS(in_ref));
ml_dff_nvcm I132 ( .R(net273), .D(net274), .CLK(fsm_sample),
     .QN(net276), .Q(nv_dataout));
nch  WR_CELL ( .D(net0159), .B(GND_), .G(testdec_b), .S(net167));
rppolywo_m  R6 ( .MINUS(net0150), .PLUS(blsa), .BULK(GND_));
rppolywo_m  R9 ( .MINUS(net171), .PLUS(net175), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(net0160), .PLUS(net0210), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net0137), .PLUS(net171), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net220), .PLUS(net0137), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(blsa), .PLUS(blsa), .BULK(GND_));
rppolywo_m  R11 ( .MINUS(net0210), .PLUS(net0131), .BULK(GND_));
rppolywo_m  R7 ( .MINUS(net0117), .PLUS(net0150), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net0131), .PLUS(net0134), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net0134), .PLUS(net0117), .BULK(GND_));
rppolywo_m  R13 ( .MINUS(gnd_), .PLUS(net0160), .BULK(GND_));
ml_core_sa_resref_40nm Irref_bot ( .bl_in(net142), .bl_out(net236),
     .ref(ref[3:0]));
ml_core_sa_restop_40nm Irref_top ( .bl_top(net0221), .bl_bot(net0159));
ml_core_sa_resbot_40nm Irsen_bot ( .bl_in(net0141), .bl_out(net175),
     .sa_ngate(sa_ngate[4:1]), .in_dec(net0247));
pch  M0 ( .D(net167), .B(vdd_), .G(testdec_en_b), .S(vdd_));
nor2_hvt I214 ( .B(high_res_b), .Y(net214), .A(fsm_tm_testdec));
nor3_hvt I102 ( .B(dec_trim[6]), .Y(high_res_b), .A(dec_trim[5]),
     .C(dec_trim[7]));
mux2_hvt I206 ( .in1(blsa), .in0(net0150), .out(in_div),
     .sel(testdec_b));
mux2_hvt I270 ( .in1(ref[1]), .in0(ref[0]), .out(net185),
     .sel(fsm_tm_ref[0]));
mux2_hvt I271 ( .in1(ref[3]), .in0(ref[2]), .out(net184),
     .sel(fsm_tm_ref[0]));
mux2_hvt I279 ( .in1(net0195), .in0(ref[2]), .out(in_ref),
     .sel(testdec_b));
mux2_hvt I234 ( .in1(dec_ok), .in0(sa_out), .out(net274),
     .sel(tm_testdec_wr));
mux2_hvt I272 ( .in1(net184), .in0(net185), .out(net0195),
     .sel(fsm_tm_ref[1]));
inv_hvt I247 ( .A(fsm_rst_b), .Y(net273));
inv_hvt I208 ( .A(fsm_tm_testdec), .Y(testdec_b));
inv_hvt I248 ( .A(net214), .Y(net226));
nch_hvt  M24 ( .D(gnd_), .B(GND_), .G(sa_ngate[1]), .S(net0150));
nch_hvt  M23 ( .D(net220), .B(GND_), .G(dec_trim[7]), .S(gnd_));
nch_hvt  M31 ( .D(gnd_), .B(GND_), .G(net226), .S(net0131));
nch_hvt  M16 ( .D(net175), .B(GND_), .G(net226), .S(gnd_));
nch_hvt  M13 ( .D(net228), .B(GND_), .G(vdd_tieh), .S(net240));
nch_hvt  M18 ( .D(net151), .B(GND_), .G(vdd_tieh), .S(net142));
nch_hvt  M25 ( .D(gnd_), .B(GND_), .G(sa_ngate[2]), .S(net0117));
nch_hvt  M29 ( .D(gnd_), .B(GND_), .G(dec_trim[6]), .S(net0160));
nch_hvt  M21 ( .D(net0137), .B(GND_), .G(dec_trim[6]), .S(gnd_));
nch_hvt  M28 ( .D(gnd_), .B(GND_), .G(dec_trim[5]), .S(net0210));
nch_hvt  M19 ( .D(net236), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M26 ( .D(gnd_), .B(GND_), .G(sa_ngate[3]), .S(net0134));
nch_hvt  M20 ( .D(net171), .B(GND_), .G(dec_trim[5]), .S(gnd_));
nch_hvt  M30 ( .D(gnd_), .B(GND_), .G(dec_trim[7]), .S(gnd_));
nch_hvt  M27 ( .D(gnd_), .B(GND_), .G(sa_ngate[4]), .S(net0131));
nch_hvt  M12 ( .D(net240), .B(GND_), .G(vdd_tieh), .S(net151));
nch_25  M22 ( .D(net167), .B(GND_), .G(vddp_tieh), .S(net228));
vdd_tielow I204 ( .gnd_tiel(gnd_tlow));
ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 ( .gwl_b_gnden_25(vddp_tieh),
     .gwl_b_sup_25(vpxa), .gwl_b_25(saen_b_vpxa),
     .gwl_gnd_25(gwl_gnd_25_ref));
ml_rock_lwldrv_wp Irock_lwldrv_wp ( .gwl_gnd_rp_25(gwl_gnd_25_ref),
     .s_rd_b_hv(saprd_b_vpxa), .gwl_gnd_25(gwl_gnd_25_ref),
     .s_b_hv(gwl_gnd_25_ref), .gwp_hv(gwl_gnd_25_ref),
     .gwl_b_25(gnd_tlow), .ngate_25(vpxa), .s_b_25(saprd_b_vpxa),
     .wp(net0221));
ml_core_sa_comp_top Icore_sa_comp_top ( .vdd_tieh(vdd_tieh),
     .saen_25(saen_25), .in_ref(in_ref), .in_div(in_div),
     .sa_out(sa_out));

endmodule
// Library - leafcell, Cell - pllmate_40lp, View - schematic
// LAST TIME SAVED: Nov  3 07:32:44 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pllmate_40lp ( pll_bypass, pll_cbit, pll_fb, pll_fse, pll_out1,
     pll_out2, pll_ref, pll_reset, pll_sdo, cbit, fo_dlyadj,
     fo_pll_bypass, fo_pll_sck, fo_pll_sdi, fo_pllfb, fo_pllref,
     fo_pllreset, pad_pllref, pllout_in, prog );
output  pll_bypass, pll_fb, pll_fse, pll_out1, pll_out2, pll_ref,
     pll_reset, pll_sdo;

input  fo_pll_bypass, fo_pll_sck, fo_pll_sdi, fo_pllfb, fo_pllref,
     fo_pllreset, pad_pllref, pllout_in, prog;

output [16:0]  pll_cbit;

input [7:0]  fo_dlyadj;
input [36:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [25:0]  q;

wire  [0:25]  net137;

wire  [24:17]  obit;

wire  [0:1]  net165;

wire  [0:3]  net114;

wire  [0:3]  net119;

wire  [0:1]  net157;



pllcfg_sr26_40lp I_pllcfg_sr ( .q(q[25:0]), .reset(prog),
     .pll_sdi(fo_pll_sdi), .pll_sck(fo_pll_sck));
fabric_buf_ice8p I_BUF4PLL_SDO ( .f_in(net176), .f_out(pll_sdo));
tiehi I_tiehi ( .tiehi(net100));
tielo I_tielo ( .tielo(pll_tielo));
mux4plldly I14 ( .min({pll_tielo, pll_tielo, pll_tielo, pllout2_d1}),
     .cbit({pll_tielo, pll_tielo}), .mout(pllout2_d2));
mux4plldly I15 ( .min({pll_tielo, pll_tielo, pll_tielo, pllout2_d2}),
     .cbit({pll_tielo, pll_tielo}), .mout(net107));
delay150ps I12 ( .in(net108), .out(pllout2_d1));
oa4plldly_40lp I_oa4plldly_fb_3_ ( .cbit(cbit[29]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[3]), .out(net114[0]));
oa4plldly_40lp I_oa4plldly_fb_2_ ( .cbit(cbit[28]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[2]), .out(net114[1]));
oa4plldly_40lp I_oa4plldly_fb_1_ ( .cbit(cbit[27]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[1]), .out(net114[2]));
oa4plldly_40lp I_oa4plldly_fb_0_ ( .cbit(cbit[26]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[0]), .out(net114[3]));
oa4plldly_40lp I_oa4plldly_out_3_ ( .cbit(cbit[34]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[7]), .out(net119[0]));
oa4plldly_40lp I_oa4plldly_out_2_ ( .cbit(cbit[33]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[6]), .out(net119[1]));
oa4plldly_40lp I_oa4plldly_out_1_ ( .cbit(cbit[32]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[5]), .out(net119[2]));
oa4plldly_40lp I_oa4plldly_out_0_ ( .cbit(cbit[31]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[4]), .out(net119[3]));
nand2_hvt I9_1_ ( .A(obit[24]), .Y(net157[0]), .B(net140));
nand2_hvt I9_0_ ( .A(obit[23]), .Y(net157[1]), .B(net140));
nand2_hvt I2_1_ ( .A(obit[20]), .B(net140), .Y(net165[0]));
nand2_hvt I2_0_ ( .A(obit[19]), .B(net140), .Y(net165[1]));
pllphase_sr_40lp I_pllphase_sr ( .tielo(pll_tielo), .tiehi(net100),
     .f_out(f_out), .cbit(obit[21]), .f_dvd2(f_dvd2),
     .f_dvd4_p0(f_dvd4_p0), .f_dvd4_p90(f_dvd4_p90), .sr(pll_reset),
     .CLK(pllout_in));
mux2_hvt I_MUX4ShftCbit_25_ ( .in1(q[25]), .in0(cbit[36]),
     .out(net137[0]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_24_ ( .in1(q[24]), .in0(cbit[24]),
     .out(net137[1]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_23_ ( .in1(q[23]), .in0(cbit[23]),
     .out(net137[2]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_22_ ( .in1(q[22]), .in0(cbit[22]),
     .out(net137[3]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_21_ ( .in1(q[21]), .in0(cbit[21]),
     .out(net137[4]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_20_ ( .in1(q[20]), .in0(cbit[20]),
     .out(net137[5]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_19_ ( .in1(q[19]), .in0(cbit[19]),
     .out(net137[6]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_18_ ( .in1(q[18]), .in0(cbit[18]),
     .out(net137[7]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_17_ ( .in1(q[17]), .in0(cbit[17]),
     .out(net137[8]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_16_ ( .in1(q[16]), .in0(cbit[16]),
     .out(net137[9]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_15_ ( .in1(q[15]), .in0(cbit[15]),
     .out(net137[10]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_14_ ( .in1(q[14]), .in0(cbit[14]),
     .out(net137[11]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_13_ ( .in1(q[13]), .in0(cbit[13]),
     .out(net137[12]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_12_ ( .in1(q[12]), .in0(cbit[12]),
     .out(net137[13]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_11_ ( .in1(q[11]), .in0(cbit[11]),
     .out(net137[14]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_10_ ( .in1(q[10]), .in0(cbit[10]),
     .out(net137[15]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_9_ ( .in1(q[9]), .in0(cbit[9]),
     .out(net137[16]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_8_ ( .in1(q[8]), .in0(cbit[8]),
     .out(net137[17]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_7_ ( .in1(q[7]), .in0(cbit[7]),
     .out(net137[18]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_6_ ( .in1(q[6]), .in0(cbit[6]),
     .out(net137[19]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_5_ ( .in1(q[5]), .in0(cbit[5]),
     .out(net137[20]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_4_ ( .in1(q[4]), .in0(cbit[4]),
     .out(net137[21]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_3_ ( .in1(q[3]), .in0(cbit[3]),
     .out(net137[22]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_2_ ( .in1(q[2]), .in0(cbit[2]),
     .out(net137[23]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_1_ ( .in1(q[1]), .in0(cbit[1]),
     .out(net137[24]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_0_ ( .in1(q[0]), .in0(cbit[0]),
     .out(net137[25]), .sel(net178));
inv_hvt I0 ( .A(pll_bypass), .Y(net140));
clkmux2buffer I_MUX4PLLRef ( .in1(fo_pllref_buf), .in0(pad_pllref),
     .out(pll_ref), .sel(obit[22]));
clkbuffer500um BUF_PLL_OUT1 ( .in(net189), .out(pll_out1));
clkbuffer500um BUF_PLL_OUT2 ( .in(net107), .out(pll_out2));
clkbuffer500um I_BUF4PLL_FB ( .in(net186), .out(pll_fb));
clkbuffer200u Ifo_pllfb_buf ( .in(fo_pllfb), .out(fo_pllfb_buf));
clkbuffer200u Ifo_pllref_buf ( .in(fo_pllref), .out(fo_pllref_buf));
clkmux4to1 I7 ( net158, net157[0:1], f_dvd4_p0, f_dvd4_p90, f_dvd2,
     f_out);
clkmux4to1 I_mux4PhaseOut ( net108, net165[0:1], f_dvd4_p0, f_dvd4_p90,
     f_dvd2, f_out);
clkmux4to1 I_clkmux4finedly ( net172, obit[18:17], pllout_in,
     f_dvd4_p0, f_dvd4_p0, fo_pllfb_buf);
buffer500um I_BUF4PLL_BYPASS ( .in(fo_pll_bypass), .out(pll_bypass));
bram_bufferx4 I3 ( .in(q[25]), .out(net176));
bram_bufferx4 I_cbit23_buffer ( .in(cbit[25]), .out(net178));
bram_bufferx4 I_cbit_buffer_25_ ( .in(net137[0]), .out(pll_fse));
bram_bufferx4 I_cbit_buffer_24_ ( .in(net137[1]), .out(obit[24]));
bram_bufferx4 I_cbit_buffer_23_ ( .in(net137[2]), .out(obit[23]));
bram_bufferx4 I_cbit_buffer_22_ ( .in(net137[3]), .out(obit[22]));
bram_bufferx4 I_cbit_buffer_21_ ( .in(net137[4]), .out(obit[21]));
bram_bufferx4 I_cbit_buffer_20_ ( .in(net137[5]), .out(obit[20]));
bram_bufferx4 I_cbit_buffer_19_ ( .in(net137[6]), .out(obit[19]));
bram_bufferx4 I_cbit_buffer_18_ ( .in(net137[7]), .out(obit[18]));
bram_bufferx4 I_cbit_buffer_17_ ( .in(net137[8]), .out(obit[17]));
bram_bufferx4 I_cbit_buffer_16_ ( .in(net137[9]), .out(pll_cbit[16]));
bram_bufferx4 I_cbit_buffer_15_ ( .in(net137[10]), .out(pll_cbit[15]));
bram_bufferx4 I_cbit_buffer_14_ ( .in(net137[11]), .out(pll_cbit[14]));
bram_bufferx4 I_cbit_buffer_13_ ( .in(net137[12]), .out(pll_cbit[13]));
bram_bufferx4 I_cbit_buffer_12_ ( .in(net137[13]), .out(pll_cbit[12]));
bram_bufferx4 I_cbit_buffer_11_ ( .in(net137[14]), .out(pll_cbit[11]));
bram_bufferx4 I_cbit_buffer_10_ ( .in(net137[15]), .out(pll_cbit[10]));
bram_bufferx4 I_cbit_buffer_9_ ( .in(net137[16]), .out(pll_cbit[9]));
bram_bufferx4 I_cbit_buffer_8_ ( .in(net137[17]), .out(pll_cbit[8]));
bram_bufferx4 I_cbit_buffer_7_ ( .in(net137[18]), .out(pll_cbit[7]));
bram_bufferx4 I_cbit_buffer_6_ ( .in(net137[19]), .out(pll_cbit[6]));
bram_bufferx4 I_cbit_buffer_5_ ( .in(net137[20]), .out(pll_cbit[5]));
bram_bufferx4 I_cbit_buffer_4_ ( .in(net137[21]), .out(pll_cbit[4]));
bram_bufferx4 I_cbit_buffer_3_ ( .in(net137[22]), .out(pll_cbit[3]));
bram_bufferx4 I_cbit_buffer_2_ ( .in(net137[23]), .out(pll_cbit[2]));
bram_bufferx4 I_cbit_buffer_1_ ( .in(net137[24]), .out(pll_cbit[1]));
bram_bufferx4 I_cbit_buffer_0_ ( .in(net137[25]), .out(pll_cbit[0]));
cfg4pllreset I_cfg4pllreset ( .prog(prog), .in(fo_pllreset),
     .out(pll_reset));
pll_finedly I11 ( .cbit(net114[0:3]), .pll_fbin(net172),
     .pll_fbout(net186));
pll_finedly I_pll_finedly ( .cbit(net119[0:3]), .pll_fbin(net158),
     .pll_fbout(net189));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_top, View - schematic
// LAST TIME SAVED: Sep 11 13:36:38 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_sa_top ( nv_dataout, bl_out, bl_pgm_glb, vdd_tieh,
     vddp_tieh, vpxa, dec_ok, dec_trim, fsm_rst_b, fsm_sample,
     fsm_tm_ref, fsm_tm_testdec, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     tm_dma, tm_testdec_wr );
output  nv_dataout;

inout  bl_out, bl_pgm_glb, vdd_tieh, vddp_tieh, vpxa;

input  dec_ok, fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, tm_dma, tm_testdec_wr;

input [1:0]  fsm_tm_ref;
input [4:1]  sa_ngate;
input [7:5]  dec_trim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(net073), .Y(net048));
inv_hvt I45 ( .A(net048), .Y(nv_dataout));
nch_hvt  M2 ( .D(bl_out), .B(GND_), .G(sa_bl_to_blsa), .S(net71));
nch_hvt  M1 ( .D(bl_out), .B(GND_), .G(sa_bl_to_pgm_glb),
     .S(bl_pgm_glb));
nch_hvt  M4 ( .D(net71), .B(GND_), .G(tm_dma), .S(gnd_));
ml_core_sa Iml_core_sa ( .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .vddp_tieh(vddp_tieh),
     .vdd_tieh(vdd_tieh), .sa_ngate(sa_ngate[4:1]), .dec_ok(dec_ok),
     .testdec_en_b(testdec_en_b), .tm_testdec_wr(tm_testdec_wr),
     .fsm_tm_testdec(fsm_tm_testdec), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .dec_trim(dec_trim[7:5]), .nv_dataout(net073), .vpxa(vpxa),
     .blsa(net71));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_core_40nm, View - schematic
// LAST TIME SAVED: Jul 15 18:30:49 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_hv_ls_inv_core_40nm ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net26), .G(sel_25), .S(net26));
pch_25  M5 ( .D(net19), .B(net22), .G(sel_b_25), .S(net22));
pch_25  M7 ( .D(net26), .B(in_hv), .G(net19), .S(in_hv));
pch_25  M6 ( .D(net22), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(net19), .B(GND_), .G(vddp_tieh), .S(net37));
nch_25  M15 ( .D(net37), .B(GND_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(GND_), .G(vddp_tieh), .S(net29));
nch_25  M14 ( .D(net29), .B(GND_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_s_b_hv_sw, View - schematic
// LAST TIME SAVED: Sep  7 10:32:39 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_s_b_hv_sw ( sbout_hv, ssup_hv, sbout_gnd_25, sbout_high_25,
     vddp_tieh );
inout  sbout_hv, ssup_hv;

input  sbout_gnd_25, sbout_high_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_core_40nm Iml_hv_ls_inv_core_40nm ( .sel_b_25(net62),
     .sel_25(sbout_high_25), .out_b_hv(sbout_hv_b), .in_hv(ssup_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M23 ( .D(sbout_hv), .B(GND_), .G(vddp_tieh), .S(net34));
nch_25  M7 ( .D(net34), .B(GND_), .G(sbout_gnd_25), .S(gnd_));
inv_25 I114 ( .IN(sbout_high_25), .OUT(net62), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M0 ( .D(net46), .B(ssup_hv), .G(sbout_hv_b), .S(ssup_hv));
pch_25  M2 ( .D(sbout_hv), .B(net46), .G(sbout_gnd_25), .S(net46));

endmodule
// Library - NVCM_40nm, Cell - ml_wp_ctrl, View - schematic
// LAST TIME SAVED: Jul 27 15:30:44 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_wp_ctrl ( s_b_25, s_b_hv, sb25sup_25, sbhvsup_hv, vddp_tieh,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25 );
inout  sb25sup_25, sbhvsup_hv, vddp_tieh;


inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [3:0]  sbhv_gnd_25;
input [3:0]  sb25_high_25;
input [3:0]  sb25_gnd_25;
input [3:0]  sbhv_high_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_s_b_hv_sw Iml_s_b_25_sw_3_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[3]),
     .sbout_hv(s_b_25[3]), .sbout_high_25(sb25_high_25[3]));
ml_s_b_hv_sw Iml_s_b_25_sw_2_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[2]),
     .sbout_hv(s_b_25[2]), .sbout_high_25(sb25_high_25[2]));
ml_s_b_hv_sw Iml_s_b_25_sw_1_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[1]),
     .sbout_hv(s_b_25[1]), .sbout_high_25(sb25_high_25[1]));
ml_s_b_hv_sw Iml_s_b_25_sw_0_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[0]),
     .sbout_hv(s_b_25[0]), .sbout_high_25(sb25_high_25[0]));
ml_s_b_hv_sw Iml_s_b_hv_sw_3_ ( .sbout_high_25(sbhv_high_25[3]),
     .sbout_hv(s_b_hv[3]), .sbout_gnd_25(sbhv_gnd_25[3]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_2_ ( .sbout_high_25(sbhv_high_25[2]),
     .sbout_hv(s_b_hv[2]), .sbout_gnd_25(sbhv_gnd_25[2]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_1_ ( .sbout_high_25(sbhv_high_25[1]),
     .sbout_hv(s_b_hv[1]), .sbout_gnd_25(sbhv_gnd_25[1]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_0_ ( .sbout_high_25(sbhv_high_25[0]),
     .sbout_hv(s_b_hv[0]), .sbout_gnd_25(sbhv_gnd_25[0]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_top_1f, View - schematic
// LAST TIME SAVED: Dec 29 14:16:08 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_ctrl_top_1f ( gwl_b_gnden_25, nv_dataout, s_rd, yp1,
     yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25, yp_test, yp_test_25,
     yp_test_b_25, bl_out, bl_pgm_glb, s_b_25, s_b_hv, sb25sup_25,
     sbhvsup_hv, vblinhi_pgm_25, vdd_tieh, vpxa, ysup_25, dec_ok,
     fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, testdec_en_b, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );
output  gwl_b_gnden_25, nv_dataout;

inout  bl_out, bl_pgm_glb, sb25sup_25, sbhvsup_hv, vblinhi_pgm_25,
     vdd_tieh, vpxa, ysup_25;

input  dec_ok, fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [7:0]  yp2;
output [5:0]  yp1_b_25;
output [1:0]  yp_test_25;
output [7:0]  yp3_b_25;
output [1:0]  yp_test_b_25;
output [7:0]  yp2_b_25;
output [1:0]  yp_test;
output [5:0]  yp1;
output [7:0]  yp3_25;
output [3:0]  s_rd;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [2:0]  fsm_trim_rrefrd;
input [9:0]  fsm_coladd;
input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefpgm;
input [1:0]  fsm_tm_ref;
input [3:0]  fsm_blkadd;
input [4:1]  sa_ngate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp2_sel;

wire  [3:0]  sb25_gnd_25;

wire  [3:0]  sbhv_gnd_25;

wire  [3:0]  sbhv_high_25;

wire  [5:0]  yp1_sel;

wire  [3:0]  sb25_high_25;

wire  [7:5]  dec_trim;

wire  [7:0]  yp3_sel;



ml_ymux_ctrl_1f Iml_ymux_ctrl_1f ( .yp1_b_25(yp1_b_25[5:0]),
     .yp1(yp1[5:0]), .yp1_sel(yp1_sel[5:0]), .yp2(yp2[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2_sel(yp2_sel[7:0]),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_sel(yp3_sel[7:0]), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test(yp_test[1:0]),
     .yp2_b_low_b(yp21_b_low_b), .yp1_b_low_b(yp21_b_low_b),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .yp_test_25(yp_test_25[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_core_ctrl_logic_1f Icore_ctrl_logic_1f (
     .fsm_coladd(fsm_coladd[9:0]), .yp1_sel(yp1_sel[5:0]),
     .vdd_tieh(vdd_tieh), .fsm_tm_rprd(fsm_tm_rprd), .s_rd(s_rd[3:0]),
     .tm_allbank_sel(tm_allbank_sel), .yp2_sel(yp2_sel[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_tm_allwl_l(tm_allwl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25), .tm_tcol(tm_tcol),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_allbl_l(tm_allbl_l), .fsm_pgm(fsm_pgm),
     .fsm_tm_allbl_h(tm_allbl_h), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_nvcmen(fsm_nvcmen), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_blkadd(fsm_blkadd[3:0]),
     .yp_test(yp_test[1:0]), .yp21_b_low_b(yp21_b_low_b),
     .yp3_sel(yp3_sel[7:0]), .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .sbhv_high_25(sbhv_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sb25_gnd_25(sb25_gnd_25[3:0]),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .dec_trim(dec_trim[7:5]));
pch_hvt  M0 ( .D(vdd_tieh), .B(vdd_), .G(net223), .S(vdd_));
pch_25  M4 ( .D(vddp_tieh), .B(vddp_), .G(net223), .S(vddp_));
nch_hvt  M3 ( .D(net223), .B(GND_), .G(net223), .S(gnd_));
inv_25 I38 ( .IN(net240), .OUT(gwl_b_gnden_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I30 ( .IN(fsm_gwlbdis_b_25), .OUT(net240), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_core_sa_top Icore_sa_top ( .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .vddp_tieh(vddp_tieh),
     .vdd_tieh(vdd_tieh), .sa_ngate(sa_ngate[4:1]), .dec_ok(dec_ok),
     .testdec_en_b(testdec_en_b), .tm_dma(tm_dma),
     .fsm_tm_testdec(fsm_tm_testdec), .tm_testdec_wr(tm_testdec_wr),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .dec_trim(dec_trim[7:5]), .nv_dataout(nv_dataout), .vpxa(vpxa),
     .bl_pgm_glb(bl_pgm_glb), .bl_out(bl_out));
ml_wp_ctrl Iml_wp_ctrl ( .vddp_tieh(vddp_tieh),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .sbhv_high_25(sbhv_high_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_gnd_25(sb25_gnd_25[3:0]), .s_b_25(s_b_25[3:0]),
     .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp_x4, View - schematic
// LAST TIME SAVED: Nov 30 17:14:06 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x4 ( wp, gwl_b_sup_25, ngate_25, gwl_b_25,
     gwl_b_gnden_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_25, gwl_b_gnden_25, gwp_hv;

output [3:0]  wp;

input [3:0]  s_b_25;
input [3:0]  s_rd_b_hv;
input [3:0]  s_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwl_b_25(gwl_b_25), .gwl_gnd_25(gwl_gnd_25));
ml_rock_lwldrv_wp Iml_lwldrv_1 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[1]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[1]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[1]), .wp(wp[1]));
ml_rock_lwldrv_wp Iml_lwldrv_2 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[2]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[2]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[2]), .wp(wp[2]));
ml_rock_lwldrv_wp Iml_lwldrv_3 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[3]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[3]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3]), .wp(wp[3]));
ml_rock_lwldrv_wp Iml_lwldrv_0 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[0]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[0]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp_x108_1f, View -
//schematic
// LAST TIME SAVED: Dec 29 14:15:11 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x108_1f ( wp, gwl_b_sup_25, ngate_25, s_b_25,
     s_b_hv, gwl_b_25, gwl_b_gnden_25, gwp_hv, s_rd_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_gnden_25;

output [107:0]  wp;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [26:0]  gwp_hv;
input [26:0]  gwl_b_25;
input [3:0]  s_rd_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_26_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[26]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[107:104]),
     .gwl_b_25(gwl_b_25[26]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_25_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[25]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[103:100]),
     .gwl_b_25(gwl_b_25[25]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_24_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[24]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[99:96]),
     .gwl_b_25(gwl_b_25[24]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_23_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[23]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[95:92]),
     .gwl_b_25(gwl_b_25[23]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_22_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[22]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[91:88]),
     .gwl_b_25(gwl_b_25[22]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_21_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[21]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[87:84]),
     .gwl_b_25(gwl_b_25[21]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_20_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[20]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[83:80]),
     .gwl_b_25(gwl_b_25[20]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_19_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[19]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[79:76]),
     .gwl_b_25(gwl_b_25[19]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_18_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[18]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[75:72]),
     .gwl_b_25(gwl_b_25[18]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_17_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[17]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[71:68]),
     .gwl_b_25(gwl_b_25[17]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_16_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[16]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[67:64]),
     .gwl_b_25(gwl_b_25[16]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_15_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[15]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[63:60]),
     .gwl_b_25(gwl_b_25[15]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_14_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[14]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[59:56]),
     .gwl_b_25(gwl_b_25[14]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_13_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[13]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[55:52]),
     .gwl_b_25(gwl_b_25[13]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_12_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[12]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[51:48]),
     .gwl_b_25(gwl_b_25[12]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_11_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[11]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[47:44]),
     .gwl_b_25(gwl_b_25[11]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_10_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[10]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[43:40]),
     .gwl_b_25(gwl_b_25[10]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_9_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[9]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[39:36]),
     .gwl_b_25(gwl_b_25[9]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_8_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[8]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[35:32]),
     .gwl_b_25(gwl_b_25[8]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_7_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[7]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[31:28]),
     .gwl_b_25(gwl_b_25[7]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_6_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[6]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[27:24]),
     .gwl_b_25(gwl_b_25[6]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_5_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[5]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[23:20]),
     .gwl_b_25(gwl_b_25[5]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_4_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[4]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[19:16]),
     .gwl_b_25(gwl_b_25[4]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_3_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[3]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[15:12]),
     .gwl_b_25(gwl_b_25[3]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_2_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[2]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[11:8]),
     .gwl_b_25(gwl_b_25[2]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_1_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[1]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[7:4]),
     .gwl_b_25(gwl_b_25[1]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_0_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[0]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[3:0]),
     .gwl_b_25(gwl_b_25[0]), .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_338x112_top_1f, View - schematic
// LAST TIME SAVED: Dec 29 14:19:40 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_338x112_top_1f ( nv_dataout, s_rd, bl_pgm_glb,
     gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde,
     vblinhi_rdo, vpxa, ysup_25, fsm_blkadd, fsm_coladd,
     fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25,
     s_rd_b_hv, sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );
output  nv_dataout;

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  s_rd;

input [1:0]  fsm_rowadd;
input [107:0]  wr;
input [9:0]  fsm_coladd;
input [26:0]  gwl_b_25;
input [2:0]  fsm_trim_rrefrd;
input [26:0]  gwp_hv;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [4:1]  sa_ngate;
input [1:0]  fsm_tm_ref;
input [3:0]  s_rd_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp3_b_25;

wire  [1:0]  bl_dummyl;

wire  [5:0]  yp1;

wire  [107:0]  wp;

wire  [7:0]  yp2_b_25;

wire  [1:0]  bl_dummyr;

wire  [327:0]  bl;

wire  [7:0]  yp3;

wire  [5:0]  yp1_b_25;

wire  [1:0]  yp_test_25;

wire  [1:0]  bl_test;

wire  [3:0]  s_b_hv;

wire  [1:0]  yp_test_b_25;

wire  [1:0]  yp_test;

wire  [7:0]  yp2;

wire  [3:0]  s_b_25;



ml_testdec_rowsx108_1f Iml_testdec_rowsx108_1f (
     .dec_det_buf(dec_det_buf), .dec_bias(dec_bias), .dec_det(dec_det),
     .wr(wr[107:0]), .wp(wp[107:0]));
ml_testdec_columnsx330_1f Iml_testdec_columnsx330_1f ( .bl(bl[327:0]),
     .dec_det_buf(dec_det_buf), .bl_test(bl_test[1:0]),
     .bl_dummyl(bl_dummyl[1:0]), .bl_dummyr(bl_dummyr[1:0]),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25));
vdd_tielow I47 ( .gnd_tiel(net148));
nvcm_cell_338x112_1f Invcm_cell_338x112_1f ( .wr_dummyt({net148,
     net148}), .wr_dummyb({net148, net148}), .wp_dummyt({net148,
     net148}), .wp_dummyb({net148, net148}), .bl_test(bl_test[1:0]),
     .bl_dummyr(bl_dummyr[1:0]), .bl_dummyl(bl_dummyl[1:0]),
     .bl(bl[327:0]), .wp(wp[107:0]), .wr(wr[107:0]));
ml_testdec_bgen Itestdec_bgen ( .dec_ok(dec_ok_l),
     .testdec_en_b(testdec_en_b), .testdec_prec_b(testdec_prec_b),
     .dec_bias(dec_bias), .dec_det(dec_det));
ml_ymux_bls_x328_1f Iml_ymux_bls_x328_1f (
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_25(yp_test_25[1:0]),
     .yp_test(yp_test[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .yp2_b_25(yp2_b_25[7:0]),
     .vblinhi_rdo(vblinhi_rdo), .bl_dummyr(bl_dummyr[1:0]),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyl(bl_dummyl[1:0]), .bl_test(bl_test[1:0]),
     .bl_out(bl_out), .bl(bl[327:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vdd_tieh(vdd_tieh),
     .yp1(yp1[5:0]), .yp2(yp2[7:0]), .yp1_b_25(yp1_b_25[5:0]));
ml_core_ctrl_top_1f Icore_ctrl_top_1f ( .yp1(yp1[5:0]),
     .yp1_b_25(yp1_b_25[5:0]), .dec_ok(dec_ok_l),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .s_rd(s_rd[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .sa_ngate(sa_ngate[4:1]), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .fsm_coladd(fsm_coladd[9:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .gwl_b_gnden_25(gwl_b_gnden_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .vdd_tieh(vdd_tieh), .tm_testdec_wr(tm_testdec_wr),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_blkadd(fsm_blkadd[3:0]), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .nv_dataout(nv_dataout), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_pgm_25(vblinhi_pgm_25),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .bl_out(bl_out),
     .yp_test(yp_test[1:0]));
ml_rock_lwldrv_wp_x108_1f Iml_rock_lwldrv_wp_x108_1f (
     .gwp_hv(gwp_hv[26:0]), .gwl_b_25(gwl_b_25[26:0]),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .ngate_25(ngate_25),
     .gwl_b_sup_25(gwl_b_sup_25), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .gwl_b_gnden_25(gwl_b_gnden_25), .wp(wp[107:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_bank_1_1f, View - schematic
// LAST TIME SAVED: Dec 30 15:03:13 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_bank_1_1f ( nv_dataout, s_rd, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  s_rd;
output [8:4]  nv_dataout;

input [2:0]  fsm_trim_rrefrd;
input [26:0]  gwl_b_25;
input [1:0]  fsm_tm_ref;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [7:0]  fsm_rowadd;
input [26:0]  gwp_hv;
input [4:1]  sa_ngate;
input [3:0]  s_rd_b_hv;
input [107:0]  wr;
input [9:0]  fsm_coladd;
input [3:0]  fsm_blkadd_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net530;

wire  [0:3]  net524;

wire  [0:3]  net297;

wire  [0:3]  net355;

wire  [0:3]  net523;

wire  [0:3]  net529;



ml_core_338x112_top_1f Iblk_4 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net523[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[4]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f Iblk_7 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net530[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd[1], fsm_blkadd[0]}), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .ysup_25(ysup_25), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .testdec_odd_b_25(testdec_odd_b_25),
     .vpxa(vpxa), .testdec_even_b_25(testdec_even_b_25),
     .saen_b_vpxa(saen_b_vpxa), .vblinhi_rdo(vblinhi_rdo),
     .saen_25(saen_25), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[7]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f blk_6 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net355[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[6]),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_tm_trow(fsm_tm_trow),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_rd(fsm_rd),
     .bl_pgm_glb(bl_pgm_glb), .fsm_rowadd(fsm_rowadd[1:0]),
     .gwl_b_sup_25(gwl_b_sup_25), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .ngate_25(ngate_25), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .saen_25(saen_25), .vblinhi_rdo(vblinhi_rdo),
     .saen_b_vpxa(saen_b_vpxa), .testdec_even_b_25(testdec_even_b_25),
     .vpxa(vpxa), .testdec_odd_b_25(testdec_odd_b_25),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ysup_25(ysup_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd[2], fsm_blkadd[1],
     fsm_blkadd_b[0]}), .tm_testdec_wr(tm_testdec_wr),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_338x112_top_1f Iblk_5 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net297[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[5]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f Iblk_8 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net529[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[8]),
     .fsm_coladd(fsm_coladd[9:0]));
inv_hvt I66_3_ ( .A(net523[0]), .Y(net524[0]));
inv_hvt I66_2_ ( .A(net523[1]), .Y(net524[1]));
inv_hvt I66_1_ ( .A(net523[2]), .Y(net524[2]));
inv_hvt I66_0_ ( .A(net523[3]), .Y(net524[3]));
inv_hvt I6_3_ ( .A(net524[0]), .Y(s_rd[3]));
inv_hvt I6_2_ ( .A(net524[1]), .Y(s_rd[2]));
inv_hvt I6_1_ ( .A(net524[2]), .Y(s_rd[1]));
inv_hvt I6_0_ ( .A(net524[3]), .Y(s_rd[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_bank_0_1f, View - schematic
// LAST TIME SAVED: Dec 30 14:58:14 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_core_bank_0_1f ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  nv_dataout;

input [9:0]  fsm_coladd;
input [1:0]  fsm_tm_ref;
input [3:0]  s_rd_b_hv;
input [2:0]  fsm_trim_rrefrd;
input [107:0]  wr;
input [26:0]  gwp_hv;
input [7:0]  fsm_rowadd;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefpgm;
input [26:0]  gwl_b_25;
input [4:1]  sa_ngate;
input [3:0]  fsm_blkadd_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net378;

wire  [0:3]  net320;

wire  [0:3]  net431;

wire  [0:3]  net432;



ml_core_338x112_top_1f Iblk_2 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net320[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[2]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f blk_1 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net431[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[1]),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_tm_trow(fsm_tm_trow),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_rd(fsm_rd),
     .bl_pgm_glb(bl_pgm_glb), .fsm_rowadd(fsm_rowadd[1:0]),
     .gwl_b_sup_25(gwl_b_sup_25), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .ngate_25(ngate_25), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .saen_25(saen_25), .vblinhi_rdo(vblinhi_rdo),
     .saen_b_vpxa(saen_b_vpxa), .testdec_even_b_25(testdec_even_b_25),
     .vpxa(vpxa), .testdec_odd_b_25(testdec_odd_b_25),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ysup_25(ysup_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd[0]}), .tm_testdec_wr(tm_testdec_wr),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_338x112_top_1f Iblk_0 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net432[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[0]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f Iblk_3 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd(net378[0:3]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd[1], fsm_blkadd[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[3]),
     .fsm_coladd(fsm_coladd[9:0]));

endmodule
// Library - leafcell, Cell - pinlatbuf12p, View - schematic
// LAST TIME SAVED: Dec 24 09:07:59 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pinlatbuf12p ( cout, cbit, icegate, pad_in, prog );
output  cout;

input  cbit, icegate, pad_in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I_txgate_lvt_2 ( .in(cout), .out(net13), .pp(net046),
     .nn(net17));
txgate_lvt I_txgate_lvt_1 ( .in(pad_in), .out(net13), .pp(net17),
     .nn(net046));
nand2_lvt I_nand2_lvt ( .A(net19), .Y(net044), .B(net13));
nand2_lvt I5 ( .A(icegate), .Y(net046), .B(cbit));
inv_lvt I6 ( .A(net046), .Y(net17));
inv_lvt I24 ( .A(prog), .Y(net19));
inv_lvt I_inv_lvt ( .A(net044), .Y(cout));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr, View - schematic
// LAST TIME SAVED: Jul 28 11:15:51 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr ( wr, gwl_wr_25, s_25, wr_sup_25 );
output  wr;

input  gwl_wr_25, s_25, wr_sup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I59 ( .A(gwl_wr_25), .Y(net27), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(s_25));
inv_25 I38 ( .IN(net27), .OUT(wr), .P(wr_sup_25), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr_x4, View - schematic
// LAST TIME SAVED: Jan 21 18:09:38 2008
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x4 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  gwl_wr_25, wr_sup_25;

output [3:0]  wr;

input [3:0]  s_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr Iml_lwldrv_2 ( .gwl_wr_25(gwl_wr_25), .wr(wr[2]),
     .s_25(s_25[2]), .wr_sup_25(wr_sup_25));
ml_rock_lwldrv_wr Iml_lwldrv_1 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[1]), .wr(wr[1]));
ml_rock_lwldrv_wr Iml_lwldrv_3 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3]), .wr(wr[3]));
ml_rock_lwldrv_wr Iml_lwldrv_0 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[0]), .wr(wr[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr_x108_1f, View -
//schematic
// LAST TIME SAVED: Dec 29 14:33:23 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x108_1f ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  wr_sup_25;

output [107:0]  wr;

input [26:0]  gwl_wr_25;
input [3:0]  s_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_26_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[107:104]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[26]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_25_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[103:100]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[25]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_24_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[99:96]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[24]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_23_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[95:92]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[23]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_22_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[91:88]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[22]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_21_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[87:84]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[21]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_20_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[83:80]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[20]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_19_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[79:76]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[19]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_18_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[75:72]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[18]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_17_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[71:68]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[17]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_16_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[67:64]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[16]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_15_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[63:60]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[15]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_14_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[59:56]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[14]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_13_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[55:52]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[13]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_12_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[51:48]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[12]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_11_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[47:44]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[11]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_10_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[43:40]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[10]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_9_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[39:36]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[9]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_8_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[35:32]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[8]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_7_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[31:28]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[7]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_6_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[27:24]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[6]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_5_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[23:20]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[5]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_4_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[19:16]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[4]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_3_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[15:12]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[3]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_2_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[11:8]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[2]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_1_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[7:4]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[1]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_0_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[3:0]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[0]));

endmodule
// Library - tsmcN40, Cell - nor3_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:26 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nor3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(Y), .B(Gb), .G(B), .S(G));
nch_25  M5 ( .D(Y), .B(Gb), .G(C), .S(G));
nch_25  M4 ( .D(Y), .B(Gb), .G(A), .S(G));
pch_25  M0 ( .D(net16), .B(Pb), .G(B), .S(net12));
pch_25  M1 ( .D(net12), .B(Pb), .G(A), .S(P));
pch_25  M2 ( .D(Y), .B(Pb), .G(C), .S(net16));

endmodule
// Library - tsmcN40, Cell - nand3_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:23 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module nand3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(net21), .B(Gb), .G(C), .S(G));
nch_25  M3 ( .D(Y), .B(Gb), .G(A), .S(net25));
nch_25  M4 ( .D(net25), .B(Gb), .G(B), .S(net21));
pch_25  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(P));
pch_25  M2 ( .D(Y), .B(Pb), .G(C), .S(P));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vddp2vpxa, View - schematic
// LAST TIME SAVED: Jul 28 11:31:26 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_ls_vddp2vpxa ( out_33, out_b_33, sup, in_25, in_b_25 );
output  out_33, out_b_33;

inout  sup;

input  in_25, in_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(out_33), .B(gnd_), .G(in_b_25), .S(gnd_));
nch_25  M7 ( .D(out_b_33), .B(gnd_), .G(in_25), .S(gnd_));
pch_25  M1 ( .D(out_b_33), .B(sup), .G(in_25), .S(net60));
pch_25  M2 ( .D(out_33), .B(sup), .G(in_b_25), .S(net56));
pch_25  M3 ( .D(net56), .B(sup), .G(out_b_33), .S(sup));
pch_25  M5 ( .D(net60), .B(sup), .G(out_33), .S(sup));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_gwhv, View - schematic
// LAST TIME SAVED: Jul 13 15:44:38 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_gwhv ( gwp_hv, gwp_sup_hv, gwl_25, gwl_25_b,
     vddp_tieh );
output  gwp_hv;

inout  gwp_sup_hv;

input  gwl_25, gwl_25_b, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M10 ( .D(net0129), .B(gnd_), .G(vddp_tieh), .S(net050));
nch_25  M12 ( .D(gwp_hv), .B(gnd_), .G(vddp_tieh), .S(net034));
nch_25  M11 ( .D(net034), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M13 ( .D(net050), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M14 ( .D(net054), .B(gnd_), .G(vddp_tieh), .S(net058));
nch_25  M15 ( .D(net058), .B(gnd_), .G(gwl_25), .S(gnd_));
pch_25  M6 ( .D(net067), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M16 ( .D(gwp_hv), .B(net067), .G(gwl_25_b), .S(net067));
pch_25  M5 ( .D(net054), .B(net087), .G(gwl_25), .S(net087));
pch_25  M8 ( .D(net087), .B(gwp_sup_hv), .G(net0129), .S(gwp_sup_hv));
pch_25  M9 ( .D(net091), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M7 ( .D(net0129), .B(net091), .G(gwl_25_b), .S(net091));

endmodule
// Library - NVCM_40nm, Cell - ml_gwl_drv, View - schematic
// LAST TIME SAVED: Aug  2 17:23:15 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_gwl_drv ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25,
     radd_1_25, radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );
output  gwl_b_25, gwl_wr_25, gwp_hv;

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25, radd_1_25,
     radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I133 ( .IN(gwl_wp_25), .OUT(gwl_wp_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I100 ( .IN(out_33), .OUT(gwl_b_25), .P(gwl_b_sup_25),
     .Pb(gwl_b_sup_25), .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(gwlb_25), .OUT(gwlb_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nor3_25 I123 ( .B(net76), .A(net68), .C(net84), .Y(dec_sel_25),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nand3_25 I44 ( .B(radd_4_25), .A(radd_5_25), .Y(net76), .C(radd_3_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I122 ( .B(radd_1_25), .A(radd_2_25), .Y(net84), .C(radd_0_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I121 ( .B(gwlgrpsel_25), .A(gwlgrpsel_25), .Y(net68),
     .C(radd_6_25), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nor2_25 I128 ( .A(wr_frcen_25), .Y(net056), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(dec_sel_25));
nor2_25 I127 ( .A(wr_dis_25), .Y(gwl_wr_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(net056));
nor2_25 I129 ( .A(dec_sel_25), .Y(net096), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_en_25));
nor2_25 I130 ( .A(net096), .Y(gwlb_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_dis_25));
nor2_25 I131 ( .A(dec_sel_25), .Y(net058), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_frcen_25));
nor2_25 I132 ( .A(net058), .Y(gwl_wp_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_dis_25));
ml_ls_vddp2vpxa I99 ( .in_25(gwlb_25), .sup(gwl_b_sup_25),
     .in_b_25(gwlb_b_25), .out_33(out_33), .out_b_33(net053));
ml_rock_lwldrv_gwhv Iml_rock_lwldrv_gwhv ( .gwp_sup_hv(gwp_sup_hv),
     .vddp_tieh(vddp_tieh), .gwp_hv(gwp_hv), .gwl_25(gwl_wp_25),
     .gwl_25_b(gwl_wp_b_25));

endmodule
// Library - NVCM_40nm, Cell - ml_gwl_drv_x27_1f, View - schematic
// LAST TIME SAVED: Dec 29 15:02:09 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_gwl_drv_x27_1f ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25,
     gnv2_b_25, gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25,
     gnv5_b_25, gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1,
     gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25, gnv2_b_25,
     gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25, gnv5_b_25,
     gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1, gwl_misc_25,
     gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

output [26:0]  gwp_hv;
output [26:0]  gwl_b_25;
output [26:0]  gwl_wr_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_gwl_drv Igwl_drv_25_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[25]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[25]), .gwl_wr_25(gwl_wr_25[25]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_24_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[24]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[24]), .gwl_wr_25(gwl_wr_25[24]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_23_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[23]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[23]), .gwl_wr_25(gwl_wr_25[23]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_22_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[22]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[22]), .gwl_wr_25(gwl_wr_25[22]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_21_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[21]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[21]), .gwl_wr_25(gwl_wr_25[21]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_20_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[20]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[20]), .gwl_wr_25(gwl_wr_25[20]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_19_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[19]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[19]), .gwl_wr_25(gwl_wr_25[19]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_18_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[18]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[18]), .gwl_wr_25(gwl_wr_25[18]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_17_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[17]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[17]), .gwl_wr_25(gwl_wr_25[17]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_16_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[16]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[16]), .gwl_wr_25(gwl_wr_25[16]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_misc_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[26]),
     .radd_0_25(vddp_tieh), .radd_1_25(vddp_tieh),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_misc_25),
     .gwp_hv(gwp_hv[26]), .gwl_wr_25(gwl_wr_25[26]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_15_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[15]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[15]), .gwl_wr_25(gwl_wr_25[15]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_14_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[14]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[14]), .gwl_wr_25(gwl_wr_25[14]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_13_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[13]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[13]), .gwl_wr_25(gwl_wr_25[13]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_12_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[12]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[12]), .gwl_wr_25(gwl_wr_25[12]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_11_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[11]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[11]), .gwl_wr_25(gwl_wr_25[11]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_10_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[10]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[10]), .gwl_wr_25(gwl_wr_25[10]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_9_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[9]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[9]), .gwl_wr_25(gwl_wr_25[9]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_8_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[8]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[8]),
     .gwl_wr_25(gwl_wr_25[8]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_7_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[7]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[7]),
     .gwl_wr_25(gwl_wr_25[7]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_6_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[6]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[6]),
     .gwl_wr_25(gwl_wr_25[6]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_5_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[5]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[5]),
     .gwl_wr_25(gwl_wr_25[5]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_4_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[4]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[4]),
     .gwl_wr_25(gwl_wr_25[4]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[3]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[3]),
     .gwl_wr_25(gwl_wr_25[3]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[2]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[2]),
     .gwl_wr_25(gwl_wr_25[2]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[1]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[1]),
     .gwl_wr_25(gwl_wr_25[1]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[0]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25),
     .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[0]), .gwl_wr_25(gwl_wr_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_1f, View - schematic
// LAST TIME SAVED: Dec 30 14:56:08 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_gwlwr_1f ( gwl_b_25, gwp_hv, wr, gwl_b_sup_25, gwp_sup_hv,
     gnv_25, gnv_b_25, gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25,
     gwl_red_25, gwlb_dis_25, gwlb_en_25, s_25, vddp_tieh, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, wr_sup_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wr_sup_25;

output [26:0]  gwl_b_25;
output [107:0]  wr;
output [26:0]  gwp_hv;

input [3:0]  s_25;
input [1:0]  gred_25;
input [1:0]  gred_b_25;
input [5:0]  gnv_b_25;
input [5:0]  gnv_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [26:0]  gwl_wr_25;



ml_rock_lwldrv_wr_x108_1f Iml_rock_lwldrv_wr_x108_1f (
     .gwl_wr_25(gwl_wr_25[26:0]), .wr(wr[107:0]),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3:0]));
ml_gwl_drv_x27_1f Igwl_drv_x27 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_wr_25(gwl_wr_25[26:0]), .gwl_b_25(gwl_b_25[26:0]),
     .gwlb_en_25(gwlb_en_25), .gwlb_dis_25(gwlb_dis_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25_1(gred_b_25[1]), .gred_b_25_0(gred_b_25[0]),
     .gred_25_1(gred_25[1]), .gred_25_0(gred_25[0]),
     .gnv5_b_25(gnv_b_25[5]), .gnv5_25(gnv_25[5]),
     .gnv4_b_25(gnv_b_25[4]), .gnv4_25(gnv_25[4]),
     .gnv3_b_25(gnv_b_25[3]), .gnv3_25(gnv_25[3]),
     .gnv2_b_25(gnv_b_25[2]), .gnv2_25(gnv_25[2]),
     .gnv1_b_25(gnv_b_25[1]), .gnv1_25(gnv_25[1]),
     .gnv0_b_25(gnv_b_25[0]), .gnv0_25(gnv_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));

endmodule
// Library - ice8chip, Cell - pllclkbuf_n40, View - schematic
// LAST TIME SAVED: Nov  2 13:03:26 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pllclkbuf_n40 ( gclk_l2clktv, gclk_r2clktv, padin_clkl_out,
     padin_clkr_out, pll_bypass, pll_cbit, pll_fb, pll_fse,
     pll_lock_out, pll_ref, pll_reset, pll_sdo, cbit, fabric_clkl_in,
     fabric_clkr_in, fo_bypass, fo_dlyadj, fo_fb, fo_ref, fo_reset,
     fo_sck, fo_sdi, icegate, padin_clkl_in, padin_clkr_in,
     pll_lock_in, pll_out, prog );
output  padin_clkl_out, padin_clkr_out, pll_bypass, pll_fb, pll_fse,
     pll_lock_out, pll_ref, pll_reset, pll_sdo;

input  fabric_clkl_in, fabric_clkr_in, fo_bypass, fo_fb, fo_ref,
     fo_reset, fo_sck, fo_sdi, icegate, padin_clkl_in, padin_clkr_in,
     pll_lock_in, pll_out, prog;

output [1:0]  gclk_l2clktv;
output [16:0]  pll_cbit;
output [1:0]  gclk_r2clktv;

input [7:0]  fo_dlyadj;
input [40:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



fabric_buf_ice8p I_GBUF_R_1_ ( .f_in(fabric_clkr_in),
     .f_out(gclk_r2clktv[1]));
fabric_buf_ice8p I_GBUF_R_0_ ( .f_in(padin_clkr_gate),
     .f_out(gclk_r2clktv[0]));
fabric_buf_ice8p I_GBUF_L_1_ ( .f_in(fabric_clkl_in),
     .f_out(gclk_l2clktv[1]));
fabric_buf_ice8p I_GBUF_L_0_ ( .f_in(padin_clkl_gate),
     .f_out(gclk_l2clktv[0]));
fabric_buf_ice8p I_buf4pll_lock ( .f_in(pll_lock_in),
     .f_out(pll_lock_out));
pllmate_40lp I_pllmate ( .pll_cbit(pll_cbit[16:0]), .cbit({cbit[40],
     cbit[35], cbit[34], cbit[33], cbit[32], cbit[31], cbit[30],
     cbit[29], cbit[28], cbit[27], cbit[26], cbit[25], cbit[24],
     cbit[23], cbit[22], cbit[21], cbit[20], cbit[19], cbit[18],
     cbit[17], cbit[16], cbit[15], cbit[14], cbit[13], cbit[12],
     cbit[11], cbit[10], cbit[9], cbit[8], cbit[7], cbit[6], cbit[5],
     cbit[4], cbit[3], cbit[2], cbit[1], cbit[0]}),
     .fo_dlyadj(fo_dlyadj[7:0]), .pll_out2(superpll_out2),
     .pll_out1(superpll_out1), .prog(prog), .pllout_in(pll_out),
     .pad_pllref(padin_clkl_in), .pll_bypass(pll_bypass),
     .fo_pllreset(fo_reset), .fo_pllref(fo_ref), .fo_pllfb(fo_fb),
     .pll_sdo(pll_sdo), .pll_reset(pll_reset), .pll_ref(pll_ref),
     .pll_fse(pll_fse), .pll_fb(pll_fb), .fo_pll_sck(fo_sck),
     .fo_pll_sdi(fo_sdi), .fo_pll_bypass(fo_bypass));
clkmux2buffer I_PadPLLMux_R ( .in1(superpll_out2), .in0(padin_clkr_in),
     .out(padin_clkr_out), .sel(cbit[38]));
clkmux2buffer I_PadPLLMux_L ( .in1(superpll_out1), .in0(padin_clkl_in),
     .out(padin_clkl_out), .sel(cbit[36]));
pinlatbuf12p I_GBUF_CLKGAT_L ( .pad_in(padin_clkl_out),
     .icegate(icegate), .cbit(cbit[37]), .cout(padin_clkl_gate),
     .prog(prog));
pinlatbuf12p I_GBUF_CLKGAT_R ( .pad_in(padin_clkr_out),
     .icegate(icegate), .cbit(cbit[39]), .cout(padin_clkr_gate),
     .prog(prog));

endmodule
// Library - NVCM_40nm, Cell - ml_rdhv_inv, View - schematic
// LAST TIME SAVED: Jul 27 12:11:18 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_rdhv_inv ( s_rd_b_hv, srdsup_hv, s_rdin_hv, vddp_tieh );
output  s_rd_b_hv;

inout  srdsup_hv;

input  s_rdin_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M1 ( .D(rd_in_25), .B(GND_), .G(vddp_tieh), .S(s_rdin_hv));
pch_25  M0 ( .D(net12), .B(srdsup_hv), .G(s_rdin_hv), .S(srdsup_hv));
pch_25  M3 ( .D(s_rd_b_hv), .B(net12), .G(rd_in_25), .S(net12));
nch_25  M21 ( .D(s_rd_b_hv), .B(GND_), .G(vddp_tieh), .S(net19));
nch_25  M29 ( .D(net19), .B(GND_), .G(rd_in_25), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_invx3_enhance, View - schematic
// LAST TIME SAVED: Oct  1 12:05:13 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_hv_invx3_enhance ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh
     );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));
pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_lshv_6v_switch_enhance, View -
//schematic
// LAST TIME SAVED: Oct  1 12:06:46 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_lshv_6v_switch_enhance ( out_b_hv, out_hv, in_hv, sel_25,
     sel_b_25, vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M0 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
pch_25  M1 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_hotsw_enhance, View -
//schematic
// LAST TIME SAVED: Jun 30 18:50:37 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw_enhance ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3_enhance Ihv_invx3 ( .vddp_tieh(vddp_tieh),
     .out_b_hv(out_b_hv), .sel_25(sel_25), .in_hv(in_hv),
     .sel_hv(sel_hv));
ml_lshv_6v_switch_enhance Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_hotswitch_enhance, View -
//schematic
// LAST TIME SAVED: Sep  8 10:25:27 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_hv_hotswitch_enhance ( hv_in_hv, hv_out_hv, selhv_25,
     vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net042));
nch_25  M2 ( .D(net031), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
nch_25  M4 ( .D(net031), .B(GND_), .G(selhv_25), .S(net042));
inv_25 I112 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M6 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_hotswitch_enhance, View -
//schematic
// LAST TIME SAVED: Apr 30 11:28:27 2008
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch_enhance ( hvin_a_hv, hvin_b_hv, out_hv,
     sel_hv_a_25, sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch_enhance Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tiehigh, View - schematic
// LAST TIME SAVED: May 13 15:28:20 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module vdd_tiehigh ( vdd_tieh );
inout  vdd_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(vdd_tieh), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_logic, View - schematic
// LAST TIME SAVED: Sep 14 11:51:05 2010
// NETLIST TIME: Jun 29 10:32:26 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_logic ( gnv, gred, gwl_misc, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, s, sa_trim, saen, testdec_en_b, testdec_even_b,
     testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd, fsm_coladd, fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rprd, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr );
output  gwl_misc, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, saen, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [3:0]  s;
output [2:0]  sa_trim;
output [5:0]  gnv;
output [1:0]  gred;

input [2:0]  fsm_trim_rrefpgm;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [0:0]  fsm_coladd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  net390;

wire  [3:0]  s_b;

wire  [5:0]  gnv_b;

wire  [2:0]  sa_trim_b;

wire  [1:0]  xadd_b;

wire  [1:0]  gred_b;

wire  [1:0]  xadd;

wire  [0:1]  net386;



anor21_hvt I109_1_ ( .A(net386[0]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I109_0_ ( .A(net386[1]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
nor4_hvt I287 ( .B(fsm_nvcmen_b), .Y(net216), .D(testdec_wp),
     .A(fsm_wren_b), .C(net331));
nor4_hvt I286 ( .B(fsm_pgmvfy), .Y(net211), .D(fsm_tm_allwl_h),
     .A(fsm_pgmvfy), .C(fsm_rd));
nor4_hvt I282 ( .B(fsm_tm_allbl_l), .Y(net0258), .D(net282),
     .A(fsm_tm_allbl_l), .C(fsm_nvcmen_b));
nor4_hvt I284 ( .B(pgm_hvpulse), .Y(wrsup_2vdd), .D(fsm_nvcmen_b),
     .A(pgm_hvpulse), .C(testdec_wr));
nor4_hvt I285 ( .B(fsm_nvcmen_b), .Y(net226), .D(fsm_wpen_b),
     .A(testdec_wr), .C(fsm_tm_allwl_l));
nand2_hvt I302 ( .A(net0341), .Y(net307), .B(tm_testdec));
nand2_hvt I297 ( .A(tm_testdec_wr), .Y(testwr_wpgnd_b),
     .B(tm_testdec));
nand2_hvt I269 ( .A(net355), .Y(testdec_even_b), .B(testdec_en));
nand2_hvt I268 ( .A(testdec_en), .Y(testdec_odd_b), .B(fsm_coladd[0]));
nand2_hvt I267 ( .A(fsm_rd), .Y(net0266), .B(tm_testdec));
nand3_hvt I298 ( .Y(net282), .B(net341), .C(fsm_lshven), .A(fsm_pgm));
nand3_hvt I299 ( .Y(net0278), .B(fsm_rd), .C(fsm_ymuxdis),
     .A(tm_testdec));
nand3_hvt I293 ( .Y(net286), .B(fsm_pgm), .C(fsm_tm_allwl_h),
     .A(fsm_wren));
nand3_hvt I288 ( .Y(net274), .B(fsm_tm_allwl_h), .C(fsm_tm_allwl_h),
     .A(stress2));
nand3_hvt I292 ( .Y(net292), .B(tm_allwl_l_b), .C(net307),
     .A(fsm_nvcmen));
nand3_hvt I303 ( .Y(gwlb_dis), .B(fsm_nvcmen), .C(testwr_wpgnd_b),
     .A(net0332));
inv_hvt I307_5_ ( .A(fsm_rowadd[7]), .Y(gnv_b[5]));
inv_hvt I307_4_ ( .A(fsm_rowadd[6]), .Y(gnv_b[4]));
inv_hvt I307_3_ ( .A(fsm_rowadd[5]), .Y(gnv_b[3]));
inv_hvt I307_2_ ( .A(fsm_rowadd[4]), .Y(gnv_b[2]));
inv_hvt I307_1_ ( .A(fsm_rowadd[3]), .Y(gnv_b[1]));
inv_hvt I307_0_ ( .A(fsm_rowadd[2]), .Y(gnv_b[0]));
inv_hvt I238 ( .A(net0274), .Y(gwl_misc));
inv_hvt I234 ( .A(testdec_en), .Y(testdec_en_b));
inv_hvt I240 ( .A(gwlbsup_vddp), .Y(net202));
inv_hvt I236 ( .A(net0300), .Y(testdec_prec_b));
inv_hvt I305_1_ ( .A(gred_b[1]), .Y(gred[1]));
inv_hvt I305_0_ ( .A(gred_b[0]), .Y(gred[0]));
inv_hvt I314_2_ ( .A(sa_trim_b[2]), .Y(sa_trim[2]));
inv_hvt I314_1_ ( .A(sa_trim_b[1]), .Y(sa_trim[1]));
inv_hvt I314_0_ ( .A(sa_trim_b[0]), .Y(sa_trim[0]));
inv_hvt I315_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I315_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I306_5_ ( .A(gnv_b[5]), .Y(gnv[5]));
inv_hvt I306_4_ ( .A(gnv_b[4]), .Y(gnv[4]));
inv_hvt I306_3_ ( .A(gnv_b[3]), .Y(gnv[3]));
inv_hvt I306_2_ ( .A(gnv_b[2]), .Y(gnv[2]));
inv_hvt I306_1_ ( .A(gnv_b[1]), .Y(gnv[1]));
inv_hvt I306_0_ ( .A(gnv_b[0]), .Y(gnv[0]));
inv_hvt I261 ( .A(pgm_hvpulse), .Y(net0390));
inv_hvt I291 ( .A(net0428), .Y(net331));
inv_hvt I263 ( .A(net282), .Y(pgm_hvpulse));
inv_hvt I250 ( .A(fsm_coladd[0]), .Y(net355));
inv_hvt I255 ( .A(net307), .Y(testdec_wp));
inv_hvt I248 ( .A(net246), .Y(net359));
inv_hvt I252 ( .A(fsm_wren), .Y(fsm_wren_b));
inv_hvt I241 ( .A(gwlbsup_vpxa), .Y(net204));
inv_hvt I244 ( .A(net0278), .Y(net0300));
inv_hvt I264 ( .A(fsm_pgmvfy), .Y(net341));
inv_hvt I246_2_ ( .A(net390[0]), .Y(sa_trim_b[2]));
inv_hvt I246_1_ ( .A(net390[1]), .Y(sa_trim_b[1]));
inv_hvt I246_0_ ( .A(net390[2]), .Y(sa_trim_b[0]));
inv_hvt I254 ( .A(net292), .Y(net365));
inv_hvt I242 ( .A(gwphv_vddp), .Y(net206));
inv_hvt I249 ( .A(net0266), .Y(testdec_en));
inv_hvt I266 ( .A(net0388), .Y(net0327));
inv_hvt I243 ( .A(gwphv_vppint), .Y(net200));
inv_hvt I256 ( .A(net286), .Y(net0343));
inv_hvt I258 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I257 ( .A(tm_testdec_wr), .Y(net0341));
inv_hvt I259 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I304_1_ ( .A(fsm_rowadd[3]), .Y(gred_b[1]));
inv_hvt I304_0_ ( .A(fsm_rowadd[2]), .Y(gred_b[0]));
inv_hvt I253 ( .A(net196), .Y(net351));
inv_hvt I251 ( .A(fsm_wpen), .Y(fsm_wpen_b));
inv_hvt I262 ( .A(fsm_pgm), .Y(fsm_pgm_b));
inv_hvt I309 ( .A(net211), .Y(wp_frcen));
inv_hvt I310 ( .A(net216), .Y(wr_dis));
inv_hvt I308 ( .A(net226), .Y(wp_dis));
inv_hvt I311 ( .A(net274), .Y(wr_frcen));
inv_hvt I312 ( .A(testwr_wpgnd_b), .Y(testdec_wr));
inv_hvt I147_3_ ( .A(s_b[3]), .Y(s[3]));
inv_hvt I147_2_ ( .A(s_b[2]), .Y(s[2]));
inv_hvt I147_1_ ( .A(s_b[1]), .Y(s[1]));
inv_hvt I147_0_ ( .A(s_b[0]), .Y(s[0]));
nor2_hvt I272 ( .A(net0258), .B(tm_testdec), .Y(pgminhi_dmmy_b));
nor2_hvt I279 ( .A(fsm_pgm), .B(fsm_pgmvfy), .Y(net0388));
nor2_hvt I313 ( .A(net0288), .B(net0390), .Y(gwlb_en));
nor2_hvt I274 ( .A(net359), .B(net201), .Y(gwphv_vddp));
nor2_hvt I273 ( .A(fsm_nvcmen_b), .B(tm_dma), .Y(saen));
nor2_hvt I278 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I300 ( .A(fsm_pgmdisc), .B(fsm_pgmhv), .Y(net0231));
nor2_hvt I316 ( .A(net207), .B(net246), .Y(gwphv_vppint));
nor2_hvt I275 ( .A(net0232), .B(fsm_nvcmen_b), .Y(net246));
nor2_hvt I276 ( .A(net203), .B(net351), .Y(gwlbsup_vpxa));
nor2_hvt I296 ( .A(fsm_pgmvfy), .B(fsm_pgm_b), .Y(stress2));
nor2_hvt I277 ( .A(net196), .B(net205), .Y(gwlbsup_vddp));
nor3_hvt I290 ( .B(fsm_tm_allwl_l), .Y(net0428), .A(fsm_tm_allwl_l),
     .C(fsm_tm_allwl_l));
nor3_hvt I324 ( .B(fsm_tm_allwl_h), .Y(net0288), .A(fsm_tm_allwl_h),
     .C(fsm_tm_allwl_h));
nor3_hvt I295 ( .B(fsm_tm_trow), .Y(net0274), .A(fsm_nv_rri_trim),
     .C(fsm_nv_sisi_ui));
nor3_hvt I294 ( .B(fsm_tm_rprd), .Y(net196), .A(fsm_tm_rprd),
     .C(fsm_tm_rprd));
mux2_hvt I180_1_ ( .in1(fsm_rowadd[1]), .in0(fsm_rowadd[1]),
     .out(net386[0]), .sel(fsm_nv_rrow));
mux2_hvt I180_0_ ( .in1(fsm_rowadd[0]), .in0(fsm_rowadd[0]),
     .out(net386[1]), .sel(fsm_nv_rrow));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net390[0]), .sel(net0327));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net390[1]), .sel(net0327));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net390[2]), .sel(net0327));
mux2_hvt I221 ( .in1(fsm_wpen), .in0(fsm_wgnden), .out(net0332),
     .sel(pgm_hvpulse));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_pump_a_clkdly I230 ( .in(net0231), .out(net0232));
ml_pump_a_clkdly I208 ( .in(net200), .out(net201));
ml_pump_a_clkdly I202 ( .in(net202), .out(net203));
ml_pump_a_clkdly I198 ( .in(net204), .out(net205));
ml_pump_a_clkdly I207 ( .in(net206), .out(net207));
anor31_hvt I121_3_ ( .A(net365), .D(net0343), .B(xadd[1]), .Y(s_b[3]),
     .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net365), .D(net0343), .B(xadd[1]), .Y(s_b[2]),
     .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net365), .D(net0343), .B(xadd_b[1]),
     .Y(s_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net365), .D(net0343), .B(xadd_b[1]),
     .Y(s_b[0]), .C(xadd_b[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_invx3, View - schematic
// LAST TIME SAVED: Jul 29 12:21:23 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hv_invx3 ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));
pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_lshv_6v_switch, View - schematic
// LAST TIME SAVED: Jul 29 12:23:54 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_lshv_6v_switch ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M3 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M0 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));

endmodule
// Library - ice1chip, Cell - pll_wrapbuf_ice1f, View - schematic
// LAST TIME SAVED: May  3 11:46:09 2011
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pll_wrapbuf_ice1f ( gclk_l2clktv[1:0], gclk_r2clktv[1:0],
     padin_clkl_out, padin_clkr_out, pll_bypass, pll_cbit[16:0],
     pll_fb, pll_fse, pll_lock_out, pll_ref, pll_reset, pll_sdo,
     cf_bbank[159], cf_bbank[135], cf_lbank[9:1], cf_lbank[33:25],
     cf_lbank[57:49], cf_lbank[81:73], cf_lbank[97], cf_lbank[99],
     cf_lbank[101], fabric_clkl_in, fabric_clkr_in, fo_bypass,
     fo_dlyadj[7:0], fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, icegate,
     padin_clkl_in, padin_clkr_in, pll_lock_in, pll_out, prog );
output  padin_clkl_out, padin_clkr_out, pll_bypass, pll_fb, pll_fse,
     pll_lock_out, pll_ref, pll_reset, pll_sdo;

input  fabric_clkl_in, fabric_clkr_in, fo_bypass, fo_fb, fo_ref,
     fo_reset, fo_sck, fo_sdi, icegate, padin_clkl_in, padin_clkr_in,
     pll_lock_in, pll_out, prog;

output [1:0]  gclk_r2clktv;
output [16:0]  pll_cbit;
output [1:0]  gclk_l2clktv;

input [7:0]  fo_dlyadj;
input [101:1]  cf_lbank;
input [135:159]  cf_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [40:0]  cbit;

wire  [0:1]  net129;

wire  [0:1]  net88;

wire  [0:1]  net82;

wire  [0:1]  net130;



pll_bufwrap_ice1f I8_1_ ( .f_in(net130[0]), .f_out(net82[0]));
pll_bufwrap_ice1f I8_0_ ( .f_in(net130[1]), .f_out(net82[1]));
pll_bufwrap_ice1f I15 ( .f_in(net145), .f_out(padin_clkr_out));
pll_bufwrap_ice1f I12_1_ ( .f_in(net88[0]), .f_out(gclk_l2clktv[1]));
pll_bufwrap_ice1f I12_0_ ( .f_in(net88[1]), .f_out(gclk_l2clktv[0]));
pll_bufwrap_ice1f I9_1_ ( .f_in(net129[0]), .f_out(net88[0]));
pll_bufwrap_ice1f I9_0_ ( .f_in(net129[1]), .f_out(net88[1]));
pll_bufwrap_ice1f I10 ( .f_in(fabric_clkl_in), .f_out(net142));
pll_bufwrap_ice1f I14 ( .f_in(net144), .f_out(padin_clkl_out));
pll_bufwrap_ice1f I11 ( .f_in(fabric_clkr_in), .f_out(net143));
pll_bufwrap_ice1f I13_1_ ( .f_in(net82[0]), .f_out(gclk_r2clktv[1]));
pll_bufwrap_ice1f I13_0_ ( .f_in(net82[1]), .f_out(gclk_r2clktv[0]));
pll_bufwrap_ice1f I16 ( .f_in(padin_clkl_in), .f_out(net124));
pll_bufwrap_ice1f I17 ( .f_in(padin_clkr_in), .f_out(net125));
bram_bufferx4 I25_39_ ( .in(cf_bbank[159]), .out(cbit[39]));
bram_bufferx4 I4_40_ ( .in(cf_lbank[101]), .out(cbit[40]));
bram_bufferx4 I4_26_ ( .in(cf_lbank[57]), .out(cbit[26]));
bram_bufferx4 I4_25_ ( .in(cf_lbank[56]), .out(cbit[25]));
bram_bufferx4 I4_24_ ( .in(cf_lbank[55]), .out(cbit[24]));
bram_bufferx4 I4_23_ ( .in(cf_lbank[54]), .out(cbit[23]));
bram_bufferx4 I4_22_ ( .in(cf_lbank[53]), .out(cbit[22]));
bram_bufferx4 I4_21_ ( .in(cf_lbank[52]), .out(cbit[21]));
bram_bufferx4 I4_20_ ( .in(cf_lbank[51]), .out(cbit[20]));
bram_bufferx4 I4_19_ ( .in(cf_lbank[50]), .out(cbit[19]));
bram_bufferx4 I4_18_ ( .in(cf_lbank[49]), .out(cbit[18]));
bram_bufferx4 I4_8_ ( .in(cf_lbank[9]), .out(cbit[8]));
bram_bufferx4 I4_7_ ( .in(cf_lbank[8]), .out(cbit[7]));
bram_bufferx4 I4_6_ ( .in(cf_lbank[7]), .out(cbit[6]));
bram_bufferx4 I4_5_ ( .in(cf_lbank[6]), .out(cbit[5]));
bram_bufferx4 I4_4_ ( .in(cf_lbank[5]), .out(cbit[4]));
bram_bufferx4 I4_3_ ( .in(cf_lbank[4]), .out(cbit[3]));
bram_bufferx4 I4_2_ ( .in(cf_lbank[3]), .out(cbit[2]));
bram_bufferx4 I4_1_ ( .in(cf_lbank[2]), .out(cbit[1]));
bram_bufferx4 I4_0_ ( .in(cf_lbank[1]), .out(cbit[0]));
bram_bufferx4 I4_36_ ( .in(cf_lbank[97]), .out(cbit[36]));
bram_bufferx4 I4_35_ ( .in(cf_lbank[81]), .out(cbit[35]));
bram_bufferx4 I4_34_ ( .in(cf_lbank[80]), .out(cbit[34]));
bram_bufferx4 I4_33_ ( .in(cf_lbank[79]), .out(cbit[33]));
bram_bufferx4 I4_32_ ( .in(cf_lbank[78]), .out(cbit[32]));
bram_bufferx4 I4_31_ ( .in(cf_lbank[77]), .out(cbit[31]));
bram_bufferx4 I4_30_ ( .in(cf_lbank[76]), .out(cbit[30]));
bram_bufferx4 I4_29_ ( .in(cf_lbank[75]), .out(cbit[29]));
bram_bufferx4 I4_28_ ( .in(cf_lbank[74]), .out(cbit[28]));
bram_bufferx4 I4_27_ ( .in(cf_lbank[73]), .out(cbit[27]));
bram_bufferx4 I4_38_ ( .in(cf_lbank[99]), .out(cbit[38]));
bram_bufferx4 I4_37_ ( .in(cf_bbank[135]), .out(cbit[37]));
bram_bufferx4 I4_17_ ( .in(cf_lbank[33]), .out(cbit[17]));
bram_bufferx4 I4_16_ ( .in(cf_lbank[32]), .out(cbit[16]));
bram_bufferx4 I4_15_ ( .in(cf_lbank[31]), .out(cbit[15]));
bram_bufferx4 I4_14_ ( .in(cf_lbank[30]), .out(cbit[14]));
bram_bufferx4 I4_13_ ( .in(cf_lbank[29]), .out(cbit[13]));
bram_bufferx4 I4_12_ ( .in(cf_lbank[28]), .out(cbit[12]));
bram_bufferx4 I4_11_ ( .in(cf_lbank[27]), .out(cbit[11]));
bram_bufferx4 I4_10_ ( .in(cf_lbank[26]), .out(cbit[10]));
bram_bufferx4 I4_9_ ( .in(cf_lbank[25]), .out(cbit[9]));
pllclkbuf_n40 I_pllclkbuf_cbuf_bot8p ( .fo_ref(fo_ref),
     .fo_sck(fo_sck), .fo_sdi(fo_sdi), .padin_clkl_in(net124),
     .padin_clkr_in(net125), .pll_lock_in(pll_lock_in),
     .pll_out(pll_out), .prog(prog), .gclk_l2clktv(net129[0:1]),
     .gclk_r2clktv(net130[0:1]), .pll_bypass(pll_bypass),
     .pll_cbit(pll_cbit[16:0]), .pll_fb(pll_fb), .pll_fse(pll_fse),
     .pll_lock_out(pll_lock_out), .pll_ref(pll_ref),
     .pll_reset(pll_reset), .pll_sdo(pll_sdo), .fo_bypass(fo_bypass),
     .fo_dlyadj(fo_dlyadj[7:0]), .fo_fb(fo_fb),
     .fabric_clkl_in(net142), .fabric_clkr_in(net143),
     .padin_clkl_out(net144), .padin_clkr_out(net145),
     .icegate(icegate), .fo_reset(fo_reset), .cbit(cbit[40:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_hotsw, View - schematic
// LAST TIME SAVED: Jul  1 14:28:58 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3 Ihv_invx3 ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));
ml_lshv_6v_switch Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_hotswitch, View - schematic
// LAST TIME SAVED: Sep 10 14:28:35 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hv_hotswitch ( hv_in_hv, hv_out_hv, selhv_25, vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M3 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
nch_25  M4 ( .D(net15), .B(GND_), .G(selhv_25), .S(net12));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_hotswitch, View - schematic
// LAST TIME SAVED: Jan 26 19:35:53 2008
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch ( hvin_a_hv, hvin_b_hv, out_hv, sel_hv_a_25,
     sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_bldrv, View - schematic
// LAST TIME SAVED: Nov 17 19:02:34 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_gwlwr_bldrv ( bgr, bl_pgm_glb, bl_frc_gnd, fsm_din, fsm_pgm,
     fsm_pgmien, fsm_trim_ipp, tm_dma );
inout  bgr, bl_pgm_glb;

input  bl_frc_gnd, fsm_din, fsm_pgm, fsm_pgmien, tm_dma;

input [3:0]  fsm_trim_ipp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net0115;

wire  [0:7]  net0152;

wire  [0:1]  net0160;

wire  [0:1]  net0180;

wire  [0:3]  net0172;

wire  [0:3]  net0156;



rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(gnd_), .PLUS(net0141), .BULK(GND_));
nch_25  M20 ( .D(net0173), .B(GND_), .G(pgm_inhi_bias),
     .S(bl_pgm_glb));
nch_25  M21 ( .D(pgm_inhi_bias), .B(GND_), .G(pgm_inhi_bias),
     .S(gnd_));
nch_25  M12_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[0]));
nch_25  M12_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[1]));
nch_25  M13_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[0]));
nch_25  M13_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[1]));
nch_25  M13_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[2]));
nch_25  M13_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[3]));
nch_25  M6 ( .D(net0164), .B(GND_), .G(net0164), .S(gnd_));
nch_25  M3 ( .D(dec_bias_p), .B(GND_), .G(bgr), .S(net0141));
nch_25  M10 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net089));
nch_25  M18_7_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[0]));
nch_25  M18_6_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[1]));
nch_25  M18_5_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[2]));
nch_25  M18_4_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[3]));
nch_25  M18_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[4]));
nch_25  M18_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[5]));
nch_25  M18_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[6]));
nch_25  M18_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[7]));
nch_25  M9 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net0135));
nch_25  M8 ( .D(net0164), .B(GND_), .G(pgmen_b_25), .S(gnd_));
nch_hvt  M36 ( .D(net0173), .B(GND_), .G(pgm_trim0_en), .S(net0107));
nch_hvt  M37 ( .D(net0107), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M31_7_ ( .D(net0115[0]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[0]));
nch_hvt  M31_6_ ( .D(net0115[1]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[1]));
nch_hvt  M31_5_ ( .D(net0115[2]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[2]));
nch_hvt  M31_4_ ( .D(net0115[3]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[3]));
nch_hvt  M31_3_ ( .D(net0115[4]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[4]));
nch_hvt  M31_2_ ( .D(net0115[5]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[5]));
nch_hvt  M31_1_ ( .D(net0115[6]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[6]));
nch_hvt  M31_0_ ( .D(net0115[7]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[7]));
nch_hvt  M19 ( .D(net0135), .B(GND_), .G(fsm_trim_ipp[0]),
     .S(net0131));
nch_hvt  M38_7_ ( .D(net0152[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_6_ ( .D(net0152[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_5_ ( .D(net0152[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_4_ ( .D(net0152[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_3_ ( .D(net0152[4]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_2_ ( .D(net0152[5]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_1_ ( .D(net0152[6]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_0_ ( .D(net0152[7]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_3_ ( .D(net0156[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_2_ ( .D(net0156[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_1_ ( .D(net0156[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_0_ ( .D(net0156[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_1_ ( .D(net0160[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_0_ ( .D(net0160[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M26 ( .D(net0131), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M33 ( .D(bl_pgm_glb), .B(GND_), .G(net0187), .S(gnd_));
nch_hvt  M30_3_ ( .D(net0172[0]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[0]));
nch_hvt  M30_2_ ( .D(net0172[1]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[1]));
nch_hvt  M30_1_ ( .D(net0172[2]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[2]));
nch_hvt  M30_0_ ( .D(net0172[3]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[3]));
nch_hvt  M34 ( .D(net089), .B(GND_), .G(pgm_trim0_en), .S(gnd_));
nch_hvt  M27_1_ ( .D(net0180[0]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[0]));
nch_hvt  M27_0_ ( .D(net0180[1]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[1]));
pch_25  M11 ( .D(pgm_inhi_bias), .B(vddp_), .G(vdd_tieh), .S(net0259));
pch_25  M14_1_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M14_0_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M5 ( .D(net0164), .B(vddp_), .G(dec_bias_p), .S(net0241));
pch_25  M7_1_ ( .D(net0241), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M7_0_ ( .D(net0241), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M4 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p), .S(net0241));
nor2_hvt I121 ( .A(net086), .B(fsm_pgmien_b_buf), .Y(pgm_trim0_en));
nor2_hvt I114 ( .B(tm_dma), .Y(net0116), .A(tm_dma));
nor4_hvt I105 ( .D(fsm_trim_ipp[0]), .B(fsm_trim_ipp[2]), .Y(net086),
     .A(fsm_trim_ipp[3]), .C(fsm_trim_ipp[1]));
nand2_hvt I71 ( .B(fsm_din), .A(fsm_pgmien), .Y(fsm_pgmien_b_buf));
inv_hvt I115 ( .A(net0116), .Y(net0187));
inv_hvt I58 ( .A(pgmen_b), .Y(pgmen));
inv_hvt I131 ( .A(fsm_pgm), .Y(pgmen_b));
inv_hvt I72 ( .A(fsm_pgmien_b_buf), .Y(fsm_pgmien_buf));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_ls_vdd2vdd25 I56 ( .in(pgmen), .sup(vddp_),
     .out_vddio_b(pgmen_b_25), .out_vddio(pgmen_25), .in_b(pgmen_b));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_wr_sup, View - schematic
// LAST TIME SAVED: Aug 10 11:01:54 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_wr_sup ( wr_sup_25, wrsup_2vdd, wrsup_2vdd_25 );
inout  wr_sup_25;

input  wrsup_2vdd, wrsup_2vdd_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M5 ( .D(net17), .B(vddp_), .G(wrsup_2vdd_25), .S(vddp_));
pch_25  M0 ( .D(net17), .B(wr_sup_25), .G(wrsup_2vdd), .S(wr_sup_25));
nch_na25  M13 ( .D(vdd_), .B(GND_), .G(wrsup_2vdd_25), .S(wr_sup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_ls25_1b, View - schematic
// LAST TIME SAVED: Oct  1 12:09:28 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25_1b ( out_25, in );
output  out_25;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I145 ( .A(in), .Y(net45));
inv_25 I153 ( .IN(out_b_25), .OUT(out_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I112 ( .in(in), .sup(vddp_), .out_vddio_b(out_b_25),
     .out_vddio(net025), .in_b(net45));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_ls25, View - schematic
// LAST TIME SAVED: Sep  7 15:15:51 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25 ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25,
     gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25, s_25,
     testdec_even_b_25, testdec_odd_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, wrsup_2vdd_25, fsm_gwlbdis, gnv, gred,
     gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en, gwlbsup_vddp,
     gwlbsup_vpxa, gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, s,
     testdec_even_b, testdec_odd_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25,
     testdec_even_b_25, testdec_odd_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, wrsup_2vdd_25;

input  fsm_gwlbdis, gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, testdec_even_b, testdec_odd_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

output [5:0]  gnv_b_25;
output [3:0]  s_25;
output [5:0]  gnv_25;
output [1:0]  gred_25;
output [1:0]  gred_b_25;

input [5:0]  gnv;
input [3:0]  s;
input [1:0]  gred;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I_1_ ( .IN(gred_25[1]), .OUT(gred_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I_0_ ( .IN(gred_25[0]), .OUT(gred_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_5_ ( .IN(gnv_25[5]), .OUT(gnv_b_25[5]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_4_ ( .IN(gnv_25[4]), .OUT(gnv_b_25[4]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_3_ ( .IN(gnv_25[3]), .OUT(gnv_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_2_ ( .IN(gnv_25[2]), .OUT(gnv_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_1_ ( .IN(gnv_25[1]), .OUT(gnv_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_0_ ( .IN(gnv_25[0]), .OUT(gnv_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I143 ( .IN(net101), .OUT(fsm_gwlbdis_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_gwlwr_ctrl_ls25_1b I139 ( .in(gwlb_dis), .out_25(gwlb_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_frcen ( .in(wr_frcen),
     .out_25(wr_frcen_25));
ml_gwlwr_ctrl_ls25_1b I144 ( .in(gwlb_en), .out_25(gwlb_en_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vpp ( .in(gwphv_vppint),
     .out_25(gwphv_vppint_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwlb_vddp ( .in(gwlbsup_vddp),
     .out_25(gwlbsup_vddp_25));
ml_gwlwr_ctrl_ls25_1b ls25_gwlb_vpp ( .in(gwlbsup_vpxa),
     .out_25(gwlbsup_vpxa_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_vdd ( .in(wrsup_2vdd),
     .out_25(wrsup_2vdd_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_dis ( .in(wr_dis), .out_25(wr_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vddp ( .in(gwphv_vddp),
     .out_25(gwphv_vddp_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_frcen ( .in(wp_frcen),
     .out_25(wp_frcen_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_dis ( .in(wp_dis), .out_25(wp_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwl_red ( .in(gwl_red),
     .out_25(gwl_red_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_nvcm ( .in(gwl_nvcm),
     .out_25(gwl_nvcm_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_misc ( .in(gwl_misc),
     .out_25(gwl_misc_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_1_ ( .in(gred[1]),
     .out_25(gred_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_0_ ( .in(gred[0]),
     .out_25(gred_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_5_ ( .in(gnv[5]), .out_25(gnv_25[5]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_4_ ( .in(gnv[4]), .out_25(gnv_25[4]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_3_ ( .in(gnv[3]), .out_25(gnv_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_2_ ( .in(gnv[2]), .out_25(gnv_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_1_ ( .in(gnv[1]), .out_25(gnv_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_0_ ( .in(gnv[0]), .out_25(gnv_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_3_ ( .in(s[3]), .out_25(s_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_2_ ( .in(s[2]), .out_25(s_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_1_ ( .in(s[1]), .out_25(s_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_0_ ( .in(s[0]), .out_25(s_25[0]));
ml_gwlwr_ctrl_ls25_1b I136 ( .in(pgminhi_dmmy_b),
     .out_25(pgminhi_dmmy_b_25));
ml_gwlwr_ctrl_ls25_1b I140 ( .in(fsm_gwlbdis), .out_25(net101));
ml_gwlwr_ctrl_ls25_1b I137 ( .in(testdec_even_b),
     .out_25(testdec_even_b_25));
ml_gwlwr_ctrl_ls25_1b I138 ( .in(testdec_odd_b),
     .out_25(testdec_odd_b_25));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_npgate_gen, View - schematic
// LAST TIME SAVED: Sep  2 17:11:20 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_core_sa_npgate_gen ( sa_ngate, saen_25, saen_b_vpxa,
     saprd_b_vpxa, sdiode_en_vpxa, vpxa, fsm_tm_rprd, fsm_tm_sdiode,
     fsm_tm_testdec, saen, satrim, vddp_tieh );
output  saen_25, saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa;

inout  vpxa;

input  fsm_tm_rprd, fsm_tm_sdiode, fsm_tm_testdec, saen, vddp_tieh;

output [4:1]  sa_ngate;

input [2:0]  satrim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  ydec_b;

wire  [2:0]  ydec;

wire  [4:1]  trim;

wire  [7:0]  dec_trim;

wire  [7:0]  dec_trim_b;

wire  [0:3]  net48;



nand2_hvt I183 ( .Y(net037), .B(fsm_tm_rprd), .A(net078));
inv_25 I149 ( .IN(net052), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nor4_hvt I102 ( .D(fsm_tm_testdec), .C(dec_trim[7]), .A(dec_trim[5]),
     .B(dec_trim[6]), .Y(net47));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_4_ ( .Y(dec_trim_b[4]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_3_ ( .Y(dec_trim_b[3]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_2_ ( .Y(dec_trim_b[2]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nand3_hvt I37_1_ ( .Y(dec_trim_b[1]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_0_ ( .Y(dec_trim_b[0]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nor2_hvt I75_4_ ( .Y(net48[0]), .B(dec_trim[4]), .A(sa_high_res));
nor2_hvt I75_3_ ( .Y(net48[1]), .B(dec_trim[3]), .A(trim[4]));
nor2_hvt I75_2_ ( .Y(net48[2]), .B(dec_trim[2]), .A(trim[3]));
nor2_hvt I75_1_ ( .Y(net48[3]), .B(dec_trim[1]), .A(trim[2]));
inv_hvt I158_2_ ( .A(satrim[2]), .Y(ydec_b[2]));
inv_hvt I158_1_ ( .A(satrim[1]), .Y(ydec_b[1]));
inv_hvt I158_0_ ( .A(satrim[0]), .Y(ydec_b[0]));
inv_hvt I160_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I160_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I160_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I160_4_ ( .A(dec_trim_b[4]), .Y(dec_trim[4]));
inv_hvt I160_3_ ( .A(dec_trim_b[3]), .Y(dec_trim[3]));
inv_hvt I160_2_ ( .A(dec_trim_b[2]), .Y(dec_trim[2]));
inv_hvt I160_1_ ( .A(dec_trim_b[1]), .Y(dec_trim[1]));
inv_hvt I160_0_ ( .A(dec_trim_b[0]), .Y(dec_trim[0]));
inv_hvt I163 ( .A(net078), .Y(net080));
inv_hvt I162 ( .A(net076), .Y(net078));
inv_hvt I165 ( .A(net073), .Y(net071));
inv_hvt I166 ( .A(net075), .Y(net073));
inv_hvt I167 ( .A(fsm_tm_sdiode), .Y(net075));
inv_hvt I175 ( .A(net059), .Y(net061));
inv_hvt I176 ( .A(net037), .Y(net059));
inv_hvt I114 ( .A(net47), .Y(sa_high_res));
inv_hvt I161 ( .A(saen), .Y(net076));
inv_hvt I159_2_ ( .A(ydec_b[2]), .Y(ydec[2]));
inv_hvt I159_1_ ( .A(ydec_b[1]), .Y(ydec[1]));
inv_hvt I159_0_ ( .A(ydec_b[0]), .Y(ydec[0]));
inv_hvt I76_4_ ( .A(net48[0]), .Y(trim[4]));
inv_hvt I76_3_ ( .A(net48[1]), .Y(trim[3]));
inv_hvt I76_2_ ( .A(net48[2]), .Y(trim[2]));
inv_hvt I76_1_ ( .A(net48[3]), .Y(trim[1]));
inv_hvt I78_4_ ( .A(trim[4]), .Y(sa_ngate[4]));
inv_hvt I78_3_ ( .A(trim[3]), .Y(sa_ngate[3]));
inv_hvt I78_2_ ( .A(trim[2]), .Y(sa_ngate[2]));
inv_hvt I78_1_ ( .A(trim[1]), .Y(sa_ngate[1]));
ml_hv_invx3 I135 ( .sel_hv(net048), .sel_25(net048),
     .vddp_tieh(vddp_tieh), .out_b_hv(saen_b_vpxa), .in_hv(vpxa));
ml_hv_invx3 I168 ( .sel_hv(net0123), .sel_25(net0123),
     .vddp_tieh(vddp_tieh), .out_b_hv(sdiode_en_vpxa), .in_hv(vpxa));
ml_hv_invx3 I178 ( .sel_hv(net0109), .sel_25(net0109),
     .vddp_tieh(vddp_tieh), .out_b_hv(saprd_b_vpxa), .in_hv(vpxa));
ml_ls_vdd2vdd25 I136 ( .in(net053), .sup(vpxa), .out_vddio_b(net047),
     .out_vddio(net048), .in_b(net052));
ml_ls_vdd2vdd25 I137 ( .in(net078), .sup(vddp_), .out_vddio_b(net052),
     .out_vddio(net053), .in_b(net080));
ml_ls_vdd2vdd25 I172 ( .in(net0129), .sup(vpxa), .out_vddio_b(net0123),
     .out_vddio(net0124), .in_b(net0128));
ml_ls_vdd2vdd25 I173 ( .in(net073), .sup(vddp_), .out_vddio_b(net0128),
     .out_vddio(net0129), .in_b(net071));
ml_ls_vdd2vdd25 I180 ( .in(net0104), .sup(vpxa), .out_vddio_b(net0108),
     .out_vddio(net0109), .in_b(net0103));
ml_ls_vdd2vdd25 I181 ( .in(net059), .sup(vddp_), .out_vddio_b(net0103),
     .out_vddio(net0104), .in_b(net061));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl, View - schematic
// LAST TIME SAVED: Nov 22 16:36:48 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25, gred_25,
     gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25,
     gwlb_en_25, pgminhi_dmmy_b_25, s_25, s_rd_b_hv, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, bgr, bl_pgm_glb,
     gwl_b_sup_25, gwp_sup_hv, srdsup_hv, vddp_tieh, vpp_int, vpxa,
     wr_sup_25, fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rprd, fsm_tm_trow,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, s_rdin_hv, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25;

inout  bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv, srdsup_hv, vddp_tieh,
     vpp_int, vpxa, wr_sup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [3:0]  s_rd_b_hv;
output [3:0]  s_25;
output [1:0]  gred_b_25;
output [1:0]  gred_25;
output [5:0]  gnv_b_25;
output [4:1]  sa_ngate;
output [5:0]  gnv_25;

input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_trim_rrefpgm;
input [7:0]  fsm_rowadd;
input [0:0]  fsm_coladd;
input [3:0]  s_rdin_hv;
input [2:0]  fsm_trim_rrefrd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  gred;

wire  [2:0]  sa_trim;

wire  [5:0]  gnv;

wire  [3:0]  s;



vdd_tielow I204 ( .gnd_tiel(net0165));
nch_hvt  M2 ( .D(net0159), .B(GND_), .G(net0159), .S(gnd_));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net0159), .S(vddp_));
ml_rdhv_inv Iml_rdhv_inv_3_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[3]), .s_rd_b_hv(s_rd_b_hv[3]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_2_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[2]), .s_rd_b_hv(s_rd_b_hv[2]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_1_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[1]), .s_rd_b_hv(s_rd_b_hv[1]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_0_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[0]), .s_rd_b_hv(s_rd_b_hv[0]),
     .vddp_tieh(vddp_tieh));
ml_hvmux_hotswitch_enhance Ihvmux_gwpsup_hv ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwphv_vppint_25), .sel_hv_a_25(gwphv_vddp_25),
     .out_hv(gwp_sup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_gwlwr_ctrl_logic Igwlwr_ctrl_logic ( .fsm_tm_rprd(fsm_tm_rprd),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_pgmdisc(fsm_pgmdisc), .gwlb_en(gwlb_en),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_rd(fsm_rd), .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[0]), .wrsup_2vdd(wrsup_2vdd),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .testdec_prec_b(testdec_prec_b),
     .testdec_odd_b(testdec_odd_b), .testdec_even_b(testdec_even_b),
     .testdec_en_b(testdec_en_b), .saen(saen), .sa_trim(sa_trim[2:0]),
     .s(s[3:0]), .pgminhi_dmmy_b(net179), .gwphv_vppint(gwphv_vppint),
     .gwphv_vddp(gwphv_vddp), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vddp(gwlbsup_vddp), .gwlb_dis(gwlb_dis),
     .gwl_misc(gwl_misc), .gred(gred[1:0]), .gnv(gnv[5:0]));
ml_hvmux_hotswitch Ihvmux_gwlbsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwlbsup_vpxa_25), .sel_hv_a_25(gwlbsup_vddp_25),
     .out_hv(gwl_b_sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_gwlwr_bldrv Igwlwr_bldrv ( .fsm_din(fsm_din), .tm_dma(tm_dma),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .bl_frc_gnd(gnd_), .bgr(bgr),
     .bl_pgm_glb(bl_pgm_glb));
ml_gwlwr_ctrl_wr_sup Igwlwr_ctrl_wr_sup ( .wrsup_2vdd(wrsup_2vdd),
     .wrsup_2vdd_25(wrsup_2vdd_25), .wr_sup_25(wr_sup_25));
ml_gwlwr_ctrl_ls25 Igwlwr_ctrl_ls25 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_en(gwlb_en), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwlb_dis(gwlb_dis), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vpxa_25(gwlbsup_vpxa_25), .wrsup_2vdd_25(wrsup_2vdd_25),
     .wrsup_2vdd(wrsup_2vdd), .testdec_odd_b(testdec_odd_b),
     .testdec_even_b(testdec_even_b),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .pgminhi_dmmy_b(net179),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwphv_vddp(gwphv_vddp),
     .gwlbsup_vddp(gwlbsup_vddp), .gwphv_vppint(gwphv_vppint),
     .gwlbsup_vddp_25(gwlbsup_vddp_25),
     .gwphv_vppint_25(gwphv_vppint_25), .gwphv_vddp_25(gwphv_vddp_25),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .s(s[3:0]), .gwl_red(fsm_nv_rrow),
     .gwl_nvcm(fsm_nv_bstream), .gwl_misc(gwl_misc), .gred(gred[1:0]),
     .gnv(gnv[5:0]), .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]));
ml_core_sa_npgate_gen Icore_sa_npgate_gen ( .fsm_tm_sdiode(net0165),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .sdiode_en_vpxa(sdiode_en_vpxa), .sa_ngate(sa_ngate[4:1]),
     .fsm_tm_testdec(tm_testdec), .satrim(sa_trim[2:0]),
     .vddp_tieh(vddp_tieh), .saen(saen), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .vpxa(vpxa));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_top_1f, View - schematic
// LAST TIME SAVED: Mar  7 17:51:21 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_gwlwr_top_1f ( fsm_gwlbdis_b_25, gwl_b_25, gwl_b_sup_25,
     gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b, wr, bgr,
     bl_pgm_glb, srdsup_hv, vpp_int, vpxa, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     s_rdin_hv, tm_dma, tm_testdec, tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_b_sup_25, pgminhi_dmmy_b_25, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b;

inout  bgr, bl_pgm_glb, srdsup_hv, vpp_int, vpxa;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [107:0]  wr;
output [26:0]  gwl_b_25;
output [3:0]  s_rd_b_hv;
output [26:0]  gwp_hv;
output [4:1]  sa_ngate;

input [7:0]  fsm_rowadd;
input [3:0]  s_rdin_hv;
input [2:0]  fsm_trim_rrefpgm;
input [0:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_trim_ipp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_25;

wire  [1:0]  gred_b_25;

wire  [1:0]  gred_25;

wire  [5:0]  gnv_b_25;

wire  [5:0]  gnv_25;



ml_gwlwr_1f Igwlwr ( .gwp_hv(gwp_hv[26:0]), .gwl_b_25(gwl_b_25[26:0]),
     .wr(wr[107:0]), .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .wr_sup_25(wr_sup_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));
ml_gwlwr_ctrl Igwlwr_ctrl ( .saprd_b_vpxa(saprd_b_vpxa),
     .sdiode_en_vpxa(sdiode_en_vpxa), .srdsup_hv(srdsup_hv),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rdin_hv(s_rdin_hv[3:0]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_en_b(testdec_en_b), .testdec_prec_b(testdec_prec_b),
     .fsm_pgmdisc(fsm_pgmdisc), .gwlb_en_25(gwlb_en_25),
     .fsm_din(fsm_din), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_allwl_l(fsm_tm_allwl_l), .fsm_tm_allwl_h(fsm_tm_allwl_h),
     .fsm_tm_allbl_l(fsm_tm_allbl_l), .fsm_tm_allbl_h(fsm_tm_allbl_h),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .s_25(s_25[3:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_red_25(gwl_red_25), .gwl_nvcm_25(gwl_nvcm_25),
     .gwl_misc_25(gwl_misc_25), .gred_b_25(gred_b_25[1:0]),
     .gred_25(gred_25[1:0]), .gnv_b_25(gnv_b_25[5:0]),
     .gnv_25(gnv_25[5:0]), .wr_sup_25(wr_sup_25), .vpxa(vpxa),
     .vpp_int(vpp_int), .vddp_tieh(vddp_tieh), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr));

endmodule
// Library - xpmem, Cell - cram2x2, View - schematic
// LAST TIME SAVED: Jun 24 18:02:08 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module cram2x2 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [3:0]  q_b;
output [3:0]  q;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  r_vdd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



eh_cram_cell_4 I_1_10 ( .q_b(q_b[1]), .q(q[1]), .wl(wl[0]), .bl(bl[1]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I_2_01 ( .q_b(q_b[2]), .q(q[2]), .wl(wl[1]), .bl(bl[0]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));
eh_cram_cell_4 I_0_00 ( .q_b(q_b[0]), .q(q[0]), .wl(wl[0]), .bl(bl[0]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I_3_11 ( .q_b(q_b[3]), .q(q[3]), .wl(wl[1]), .bl(bl[1]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_core_1f, View - schematic
// LAST TIME SAVED: Dec 31 15:08:48 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_chip_nvcm_core_1f ( nv_dataout, s_rd, bgr, ngate_25,
     sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi, vpp_int, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_multibl_read, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_ref,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_trim_ipp,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, s_rdin_hv, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi,
     vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [8:0]  nv_dataout;
output [3:0]  s_rd;

input [2:0]  fsm_trim_rrefpgm;
input [1:0]  fsm_tm_ref;
input [3:0]  fsm_trim_ipp;
input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_blkadd;
input [9:0]  fsm_coladd;
input [3:0]  s_rdin_hv;
input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [26:0]  gwl_b_25;

wire  [107:0]  wr;

wire  [3:0]  s_rd_b_hv;

wire  [26:0]  gwp_hv;

wire  [4:1]  sa_ngate;



ml_core_bank_1_1f Ibank_1 ( .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .gwl_b_25(gwl_b_25[26:0]), .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .tm_allbank_sel(tm_allbank_sel),
     .saprd_b_vpxa(saprd_b_vxpa), .gwl_b_sup_25(gwl_b_sup_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .ngate_25(ngate_25),
     .s_rd(s_rd[3:0]), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .bl_pgm_glb(bl_pgm_glb),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd(fsm_blkadd[3:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_rprd(fsm_tm_rprd), .nv_dataout(nv_dataout[8:4]));
ml_core_bank_0_1f Ibank_0 ( .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .gwl_b_25(gwl_b_25[26:0]), .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .saen_25(saen_25), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .saen_b_vpxa(saen_b_vpxa),
     .saprd_b_vpxa(saprd_b_vxpa), .gwl_b_sup_25(gwl_b_sup_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .fsm_nvcmen(fsm_nvcmen), .fsm_pgm(fsm_pgm),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd(fsm_blkadd[3:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_tm_trow(fsm_tm_trow), .ngate_25(ngate_25),
     .nv_dataout(nv_dataout[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .tm_allbank_sel(tm_allbank_sel));
ml_gwlwr_top_1f Igwlwr_top_1f ( .gwl_b_25(gwl_b_25[26:0]),
     .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wgnden(fsm_wgnden), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_tm_allbl_h(tm_allbl_h),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .saprd_b_vpxa(saprd_b_vxpa),
     .fsm_lshven(fsm_lshven), .fsm_wren(fsm_wren),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .testdec_en_b(testdec_en_b), .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .sdiode_en_vpxa(net335), .srdsup_hv(srdsup_hv), .vpxa(vpxa),
     .vpp_int(vpp_int), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr),
     .gwl_b_sup_25(gwl_b_sup_25), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rdin_hv(s_rdin_hv[3:0]), .tm_testdec(fsm_tm_testdec),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .sa_ngate(sa_ngate[4:1]), .testdec_prec_b(testdec_prec_b),
     .fsm_wpen(fsm_wpen), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_tm_allwl_l(tm_allwl_l), .fsm_tm_allbl_l(tm_allbl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .fsm_din(fsm_din), .tm_dma(tm_dma));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_buf, View - schematic
// LAST TIME SAVED: Sep 30 11:47:35 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_chip_buf ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(in), .Y(net120));
inv_hvt I45 ( .A(net120), .Y(out));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_buf_hvsw_8f, View - schematic
// LAST TIME SAVED: Sep 10 14:09:50 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_chip_buf_hvsw_8f ( fsm_bgr_dis_buf, fsm_nvcmen_buf,
     fsm_pumpen_buf, fsm_tm_xforce_buf, fsm_tm_xvpxaint_buf,
     fsm_trim_vbg_buf, fsm_vrdwl_buf, fsm_bgr_dis, fsm_nvcmen,
     fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint, fsm_trim_vbg,
     fsm_vrdwl );
output  fsm_bgr_dis_buf, fsm_nvcmen_buf, fsm_pumpen_buf,
     fsm_tm_xforce_buf, fsm_tm_xvpxaint_buf;

input  fsm_bgr_dis, fsm_nvcmen, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint;

output [2:0]  fsm_vrdwl_buf;
output [3:0]  fsm_trim_vbg_buf;

input [2:0]  fsm_vrdwl;
input [3:0]  fsm_trim_vbg;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net256;



mux2_hvt I158 ( .in1(net153), .in0(net153), .out(net263),
     .sel(gnd_in));
mux2_hvt I206 ( .in1(gnd_in), .in0(gnd_in), .out(net161),
     .sel(gnd_in));
mux2_hvt I156 ( .in1(net161), .in0(net161), .out(net157),
     .sel(gnd_in));
mux2_hvt I157 ( .in1(net157), .in0(net157), .out(net153),
     .sel(gnd_in));
nor3_hvt I137 ( .B(net203), .Y(net199), .A(net203), .C(net203));
nor3_hvt I138 ( .B(net199), .Y(net195), .A(net199), .C(net199));
nor3_hvt I141 ( .B(net195), .Y(net191), .A(net195), .C(net195));
nor3_hvt I142 ( .B(net191), .Y(net187), .A(net191), .C(net191));
nor3_hvt I152 ( .B(net175), .Y(net171), .A(net175), .C(net175));
nor3_hvt I151 ( .B(net179), .Y(net175), .A(net179), .C(net179));
nor3_hvt I148 ( .B(net183), .Y(net179), .A(net183), .C(net183));
nor3_hvt I147 ( .B(net187), .Y(net183), .A(net187), .C(net187));
nor3_hvt I129 ( .B(net207), .Y(net203), .A(net207), .C(net207));
nor3_hvt I155 ( .B(net171), .Y(net262), .A(net171), .C(net171));
nand3_hvt I154 ( .Y(net261), .B(net212), .C(net212), .A(net212));
nand3_hvt I246 ( .Y(net244), .B(net248), .C(net248), .A(net248));
nand3_hvt I143 ( .Y(net228), .B(net232), .C(net232), .A(net232));
nand3_hvt I140 ( .Y(net232), .B(net236), .C(net236), .A(net236));
nand3_hvt I139 ( .Y(net236), .B(net240), .C(net240), .A(net240));
nand3_hvt I136 ( .Y(net240), .B(net244), .C(net244), .A(net244));
nand3_hvt I146 ( .Y(net224), .B(net228), .C(net228), .A(net228));
nand3_hvt I149 ( .Y(net220), .B(net224), .C(net224), .A(net224));
nand3_hvt I150 ( .Y(net216), .B(net220), .C(net220), .A(net220));
nand3_hvt I153 ( .Y(net212), .B(net216), .C(net216), .A(net216));
ml_chip_buf I120_3_ ( .in(vdd_spare), .out(net256[0]));
ml_chip_buf I120_2_ ( .in(vdd_spare), .out(net256[1]));
ml_chip_buf I120_1_ ( .in(vdd_spare), .out(net256[2]));
ml_chip_buf I120_0_ ( .in(vdd_spare), .out(net256[3]));
ml_chip_buf I159 ( .in(fsm_pumpen), .out(fsm_pumpen_buf));
ml_chip_buf I50_3_ ( .in(fsm_trim_vbg[3]), .out(fsm_trim_vbg_buf[3]));
ml_chip_buf I50_2_ ( .in(fsm_trim_vbg[2]), .out(fsm_trim_vbg_buf[2]));
ml_chip_buf I50_1_ ( .in(fsm_trim_vbg[1]), .out(fsm_trim_vbg_buf[1]));
ml_chip_buf I50_0_ ( .in(fsm_trim_vbg[0]), .out(fsm_trim_vbg_buf[0]));
ml_chip_buf I163 ( .in(fsm_bgr_dis), .out(fsm_bgr_dis_buf));
ml_chip_buf I49_2_ ( .in(fsm_vrdwl[2]), .out(fsm_vrdwl_buf[2]));
ml_chip_buf I49_1_ ( .in(fsm_vrdwl[1]), .out(fsm_vrdwl_buf[1]));
ml_chip_buf I49_0_ ( .in(fsm_vrdwl[0]), .out(fsm_vrdwl_buf[0]));
ml_chip_buf I53 ( .in(fsm_nvcmen), .out(fsm_nvcmen_buf));
ml_chip_buf I161 ( .in(fsm_tm_xvpxaint), .out(fsm_tm_xvpxaint_buf));
ml_chip_buf I160 ( .in(fsm_tm_xforce), .out(fsm_tm_xforce_buf));
vdd_tielow I135 ( .gnd_tiel(gnd_in));
vdd_tielow I145 ( .gnd_tiel(net248));
vdd_tielow I144 ( .gnd_tiel(net207));
vdd_tiehigh I117 ( .vdd_tieh(vdd_spare));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_buf, View - schematic
// LAST TIME SAVED: Oct  6 16:26:13 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_bgr_buf ( sa_out, en_25, inn, inp, sa_bias_25 );
inout  sa_out;

input  en_25, inn, inp, sa_bias_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M0 ( .D(sa_mirr_25), .B(GND_), .G(inp), .S(net436));
nch_na25  M1 ( .D(sa_out), .B(GND_), .G(inn), .S(net436));
nch_na25  M2 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_na25  M4 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_na25  M8 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_na25  M7 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M46 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M92 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M97 ( .D(tie_low), .B(GND_), .G(net0239), .S(GND_));
nch_25  M3 ( .D(net436), .B(GND_), .G(sa_bias_25), .S(GND_));
pch_25  M93 ( .D(net0123), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M95 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M94 ( .D(net0119), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M96 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M71 ( .D(sa_mirr_25), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M101 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M102 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M98 ( .D(net0239), .B(vddp_), .G(net0239), .S(vddp_));
pch_25  M10 ( .D(sa_mirr_25), .B(vddp_), .G(en_25), .S(vddp_));
pch_25  M91 ( .D(sa_out), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M25 ( .D(sa_out), .B(vddp_), .G(en_25), .S(vddp_));

endmodule
// Library - tsmcN40, Cell - nand4_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:24 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module nand4_25 ( Y, A, B, C, D, G, Gb, P, Pb );
output  Y;

input  A, B, C, D, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M6 ( .D(net14), .B(Gb), .G(C), .S(net10));
nch_25  M7 ( .D(net10), .B(Gb), .G(D), .S(G));
nch_25  M4 ( .D(Y), .B(Gb), .G(A), .S(net18));
nch_25  M5 ( .D(net18), .B(Gb), .G(B), .S(net14));
pch_25  M2 ( .D(Y), .B(Pb), .G(C), .S(P));
pch_25  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(P));
pch_25  M3 ( .D(Y), .B(Pb), .G(D), .S(P));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ref_sw, View - schematic
// LAST TIME SAVED: Jul  9 15:54:44 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpp_ref_sw ( in, out, sel_b_25 );
inout  in, out;

input  sel_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I281 ( .IN(sel_b_25), .OUT(net122), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M12 ( .D(out), .B(GND_), .G(net122), .S(in));
pch_25  M14 ( .D(in), .B(vddp_), .G(sel_b_25), .S(out));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_res_100_ohm, View - schematic
// LAST TIME SAVED: May 28 16:29:33 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_bgr_res_100_ohm ( b, t );
inout  b, t;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo  R9 ( .MINUS(net7), .PLUS(net7));
rppolywo  R3 ( .MINUS(b), .PLUS(t));
rppolywo  R2 ( .MINUS(b), .PLUS(t));
rppolywo  R4 ( .MINUS(b), .PLUS(t));
rppolywo  R5 ( .MINUS(b), .PLUS(t));
rppolywo  R6 ( .MINUS(b), .PLUS(t));
rppolywo  R8 ( .MINUS(b), .PLUS(t));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr, View - schematic
// LAST TIME SAVED: Jan  3 16:50:37 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_bgr ( bgr, bgr_bias, sa_bias_25, en_25 );
inout  bgr, bgr_bias, sa_bias_25;

input  en_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M75 ( .D(sa_mirr_25), .B(GND_), .G(in_pnpx8), .S(net436));
nch_na25  M60 ( .D(bgr_bias), .B(GND_), .G(in_pnpx1), .S(net436));
inv_25 I186 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nch_na25_macx  M76 ( .D(GND_), .G(tie_low), .S(GND_));
nch_na25_macx  M79 ( .D(GND_), .G(tie_low), .S(GND_));
nch_na25_macx  M78 ( .D(GND_), .G(tie_low), .S(GND_));
nch_na25_macx  M77 ( .D(GND_), .G(tie_low), .S(GND_));
pnp  QQ8 ( .C(GND_), .B(GND_), .E(net423));
pnp  QQ1 ( .C(GND_), .B(GND_), .E(in_pnpx1));
rppolywo  R4 ( .MINUS(sa_bias_25), .PLUS(net0209));
rppolywo  R0 ( .MINUS(net0209), .PLUS(net0303));
rppolywo  R3 ( .MINUS(in_pnpx1), .PLUS(bgr));
rppolywo  R1 ( .MINUS(in_pnpx8), .PLUS(bgr));
rppolywo  R2 ( .MINUS(net423), .PLUS(in_pnpx8));
rppolywo  R5 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R6 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R7 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R8 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R10 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R11 ( .MINUS(GND_), .PLUS(GND_));
nch_25  M97 ( .D(tie_low), .B(GND_), .G(net0309), .S(GND_));
nch_25  M82 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M58 ( .D(net0224), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M59 ( .D(net0224), .B(GND_), .G(en_b_25), .S(GND_));
nch_25  M85 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M100 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M96 ( .D(net0224), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M86 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M91 ( .D(GND_), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M94 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M23 ( .D(bgr), .B(GND_), .G(en_b_25), .S(GND_));
nch_25  M46 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M27 ( .D(sa_bias_25), .B(GND_), .G(en_b_25), .S(GND_));
nch_25  M92 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M81 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M95 ( .D(net0224), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M93 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M3 ( .D(net436), .B(GND_), .G(sa_bias_25), .S(GND_));
pch_25  M88 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M22 ( .D(vddp_), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M62 ( .D(in_pnpx1), .B(vddp_), .G(net0224), .S(net0303));
pch_25  M83 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M98 ( .D(net0309), .B(vddp_), .G(net0309), .S(vddp_));
pch_25  M71 ( .D(sa_mirr_25), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M89 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M99 ( .D(net0323), .B(vddp_), .G(en_b_25), .S(vddp_));
pch_25  M74 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M40 ( .D(net0303), .B(vddp_), .G(en_b_25), .S(vddp_));
pch_25  M90 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M10 ( .D(sa_mirr_25), .B(vddp_), .G(en_25), .S(vddp_));
pch_25  M72 ( .D(net0224), .B(vddp_), .G(bgr_bias), .S(net0303));
pch_25  M80 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M73 ( .D(bgr), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M84 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M64 ( .D(bgr_bias), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M87 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M25 ( .D(bgr_bias), .B(vddp_), .G(en_25), .S(vddp_));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_top, View - schematic
// LAST TIME SAVED: Sep 10 14:19:39 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_bgr_top ( bgr_int, fsm_bgr_dis_buf, fsm_nvcmen_buf,
     fsm_trim_vbg_buf );
inout  bgr_int;

input  fsm_bgr_dis_buf, fsm_nvcmen_buf;

input [3:0]  fsm_trim_vbg_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net0169;

wire  [0:3]  net190;

wire  [0:3]  net192;

wire  [0:1]  net0170;

wire  [0:3]  net200;

wire  [0:3]  net201;

wire  [3:0]  bgrtrim_25;

wire  [15:0]  bgr_dec_b_25;

wire  [0:15]  vref;

wire  [3:0]  bgrtrim_b_25;



vdd_tiehigh I205 ( .vdd_tieh(net0167));
nand2_hvt I323 ( .B(fsm_nvcmen_buf), .A(net0281), .Y(net188));
ml_bgr_buf Iml_bgr_buf ( .sa_bias_25(sa_bias_25), .inp(bgr),
     .inn(vref[8]), .en_25(bgr_en_25), .sa_out(vref_reg));
nand4_25 I135_7_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[7]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_6_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[6]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_5_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[5]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_4_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[4]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_3_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[3]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_2_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[2]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_1_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[1]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_0_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[0]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_15_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[15]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_14_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[14]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_13_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[13]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_12_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[12]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_11_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[11]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_10_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[10]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_9_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[9]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_8_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[8]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
pch_25  M6_1_ ( .D(net0169[0]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M6_0_ ( .D(net0169[1]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M7_1_ ( .D(net0170[0]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M7_0_ ( .D(net0170[1]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M3 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M73 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M4 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M2 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M5 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M25 ( .D(net113), .B(vddp_), .G(bgr_en_b), .S(vddp_));
nch_na25_macx  M10 ( .D(gnd_), .G(vref_reg), .S(gnd_));
nch_na25_macx  M8 ( .D(gnd_), .G(vref_reg), .S(gnd_));
nch_na25_macx  M11 ( .D(gnd_), .G(bgr_int), .S(gnd_));
nch_na25_macx  M60 ( .D(net124), .G(vref_reg), .S(net0155));
nch_na25_macx  M0 ( .D(gnd_), .G(vref_reg), .S(gnd_));
ml_vpp_ref_sw I169 ( .in(bgr_int), .out(net0238), .sel_b_25(bgr_en_b));
ml_vpp_ref_sw I170 ( .in(bgr_int), .out(vref_vdd),
     .sel_b_25(bgr_en_25));
ml_vpp_ref_sw ref_sw_7_ ( .in(net0238), .out(vref[7]),
     .sel_b_25(bgr_dec_b_25[7]));
ml_vpp_ref_sw ref_sw_6_ ( .in(net0238), .out(vref[6]),
     .sel_b_25(bgr_dec_b_25[6]));
ml_vpp_ref_sw ref_sw_5_ ( .in(net0238), .out(vref[5]),
     .sel_b_25(bgr_dec_b_25[5]));
ml_vpp_ref_sw ref_sw_4_ ( .in(net0238), .out(vref[4]),
     .sel_b_25(bgr_dec_b_25[4]));
ml_vpp_ref_sw ref_sw_3_ ( .in(net0238), .out(vref[3]),
     .sel_b_25(bgr_dec_b_25[3]));
ml_vpp_ref_sw ref_sw_2_ ( .in(net0238), .out(vref[2]),
     .sel_b_25(bgr_dec_b_25[2]));
ml_vpp_ref_sw ref_sw_1_ ( .in(net0238), .out(vref[1]),
     .sel_b_25(bgr_dec_b_25[1]));
ml_vpp_ref_sw ref_sw_0_ ( .in(net0238), .out(vref[0]),
     .sel_b_25(bgr_dec_b_25[0]));
ml_vpp_ref_sw ref_sw_15_ ( .in(net0238), .out(vref[15]),
     .sel_b_25(bgr_dec_b_25[15]));
ml_vpp_ref_sw ref_sw_14_ ( .in(net0238), .out(vref[14]),
     .sel_b_25(bgr_dec_b_25[14]));
ml_vpp_ref_sw ref_sw_13_ ( .in(net0238), .out(vref[13]),
     .sel_b_25(bgr_dec_b_25[13]));
ml_vpp_ref_sw ref_sw_12_ ( .in(net0238), .out(vref[12]),
     .sel_b_25(bgr_dec_b_25[12]));
ml_vpp_ref_sw ref_sw_11_ ( .in(net0238), .out(vref[11]),
     .sel_b_25(bgr_dec_b_25[11]));
ml_vpp_ref_sw ref_sw_10_ ( .in(net0238), .out(vref[10]),
     .sel_b_25(bgr_dec_b_25[10]));
ml_vpp_ref_sw ref_sw_9_ ( .in(net0238), .out(vref[9]),
     .sel_b_25(bgr_dec_b_25[9]));
ml_vpp_ref_sw ref_sw_8_ ( .in(net0238), .out(vref[8]),
     .sel_b_25(bgr_dec_b_25[8]));
rppolywo  R0 ( .MINUS(vref[15]), .PLUS(net0147));
rppolywo  R8 ( .MINUS(gnd_), .PLUS(vref[0]));
rppolywo  R2 ( .MINUS(net0147), .PLUS(net124));
ml_bgr_res_100_ohm I90 ( .t(vref[8]), .b(vref[7]));
ml_bgr_res_100_ohm I91 ( .t(vref[7]), .b(vref[6]));
ml_bgr_res_100_ohm I92 ( .t(vref[6]), .b(vref[5]));
ml_bgr_res_100_ohm I93 ( .t(vref[4]), .b(vref[3]));
ml_bgr_res_100_ohm I94 ( .t(vref[5]), .b(vref[4]));
ml_bgr_res_100_ohm I95 ( .t(vref[1]), .b(vref[0]));
ml_bgr_res_100_ohm I97 ( .t(vref[2]), .b(vref[1]));
ml_bgr_res_100_ohm I100 ( .t(vref[3]), .b(vref[2]));
ml_bgr_res_100_ohm I101 ( .t(vref[13]), .b(vref[14]));
ml_bgr_res_100_ohm I102 ( .t(vref[14]), .b(vref[15]));
ml_bgr_res_100_ohm I104 ( .t(vref[11]), .b(vref[12]));
ml_bgr_res_100_ohm I105 ( .t(vref[12]), .b(vref[13]));
ml_bgr_res_100_ohm I106 ( .t(vref[10]), .b(vref[11]));
ml_bgr_res_100_ohm I107 ( .t(vref[9]), .b(vref[10]));
ml_bgr_res_100_ohm I108 ( .t(vref[8]), .b(vref[9]));
ml_bgr Iml_bgr ( .bgr_bias(bgr_bias), .sa_bias_25(sa_bias_25),
     .en_25(bgr_en_25), .bgr(bgr));
inv_25 I186 ( .IN(net195), .OUT(bgr_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I139 ( .IN(net196), .OUT(bgr_en_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I198_3_ ( .IN(net201[0]), .OUT(bgrtrim_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_2_ ( .IN(net201[1]), .OUT(bgrtrim_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_1_ ( .IN(net201[2]), .OUT(bgrtrim_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_0_ ( .IN(net201[3]), .OUT(bgrtrim_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_3_ ( .IN(net200[0]), .OUT(bgrtrim_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_2_ ( .IN(net200[1]), .OUT(bgrtrim_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_1_ ( .IN(net200[2]), .OUT(bgrtrim_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_0_ ( .IN(net200[3]), .OUT(bgrtrim_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I192 ( .IN(net0313), .OUT(bgr2vdd_25_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I189 ( .IN(net0312), .OUT(bgr2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I88_3_ ( .A(fsm_trim_vbg_buf[3]), .Y(net190[0]));
inv_hvt I88_2_ ( .A(fsm_trim_vbg_buf[2]), .Y(net190[1]));
inv_hvt I88_1_ ( .A(fsm_trim_vbg_buf[1]), .Y(net190[2]));
inv_hvt I88_0_ ( .A(fsm_trim_vbg_buf[0]), .Y(net190[3]));
inv_hvt I167 ( .A(net188), .Y(net186));
inv_hvt I183 ( .A(net0167), .Y(net0326));
inv_hvt I168 ( .A(fsm_bgr_dis_buf), .Y(net0281));
inv_hvt I174 ( .A(net0326), .Y(vref_vdd));
inv_hvt I87_3_ ( .A(net190[0]), .Y(net192[0]));
inv_hvt I87_2_ ( .A(net190[1]), .Y(net192[1]));
inv_hvt I87_1_ ( .A(net190[2]), .Y(net192[2]));
inv_hvt I87_0_ ( .A(net190[3]), .Y(net192[3]));
ml_ls_vdd2vdd25 I80_3_ ( .in(net192[0]), .sup(vddp_),
     .out_vddio_b(net200[0]), .out_vddio(net201[0]), .in_b(net190[0]));
ml_ls_vdd2vdd25 I80_2_ ( .in(net192[1]), .sup(vddp_),
     .out_vddio_b(net200[1]), .out_vddio(net201[1]), .in_b(net190[1]));
ml_ls_vdd2vdd25 I80_1_ ( .in(net192[2]), .sup(vddp_),
     .out_vddio_b(net200[2]), .out_vddio(net201[2]), .in_b(net190[2]));
ml_ls_vdd2vdd25 I80_0_ ( .in(net192[3]), .sup(vddp_),
     .out_vddio_b(net200[3]), .out_vddio(net201[3]), .in_b(net190[3]));
ml_ls_vdd2vdd25 I177 ( .in(vref_vdd), .sup(vddp_),
     .out_vddio_b(net0312), .out_vddio(net0313), .in_b(net0326));
ml_ls_vdd2vdd25 I335 ( .in(net186), .sup(vddp_), .out_vddio_b(net195),
     .out_vddio(net196), .in_b(net188));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_buf, View - schematic
// LAST TIME SAVED: Sep  3 15:27:07 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_pump_vpxa_buf ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I38 ( .IN(in), .OUT(net15), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
inv_25 I195 ( .IN(net15), .OUT(out), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - ice8chip, Cell - cram_2x2x2_ice8p, View - schematic
// LAST TIME SAVED: Jun 24 17:55:16 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module cram_2x2x2_ice8p ( q, q_b, bl, pgate_l, pgate_r, r_gnd_l,
     r_gnd_r, reset_l, reset_r, wl_l, wl_r );



output [7:0]  q_b;
output [7:0]  q;

inout [3:0]  bl;

input [1:0]  r_gnd_r;
input [1:0]  pgate_l;
input [1:0]  reset_r;
input [1:0]  wl_r;
input [1:0]  reset_l;
input [1:0]  pgate_r;
input [1:0]  r_gnd_l;
input [1:0]  wl_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 I_mem_r ( .bl(bl[3:2]), .q_b(q_b[7:4]), .reset(reset_r[1:0]),
     .q(q[7:4]), .wl(wl_r[1:0]), .r_vdd(r_gnd_r[1:0]),
     .pgate(pgate_r[1:0]));
cram2x2 I_mem_l ( .bl(bl[1:0]), .q_b(q_b[3:0]), .reset(reset_l[1:0]),
     .q(q[3:0]), .wl(wl_l[1:0]), .r_vdd(r_gnd_l[1:0]),
     .pgate(pgate_l[1:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_pump, View - schematic
// LAST TIME SAVED: Aug 30 18:07:52 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpp_pump ( pump_in, clkin_25, en_25 );
inout  pump_in;

input  clkin_25, en_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));
nmoscap_25  C1 ( .MINUS(clk_b_25), .PLUS(s_3));
nch_na25  M1 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
nch_na25  M2 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
nch_na25  M3 ( .D(s_2), .B(GND_), .G(s_2), .S(s_3));
nch_na25  M22 ( .D(net23), .B(GND_), .G(net23), .S(s_0));
nch_na25  M4 ( .D(s_3), .B(GND_), .G(s_3), .S(pump_in));
pch_25  M0 ( .D(net23), .B(vddp_), .G(net64), .S(vddp_));
inv_25 I230 ( .IN(clkin_25), .OUT(net0124), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I232 ( .IN(net088), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I233 ( .IN(net0100), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I234 ( .IN(net094), .OUT(net0106), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I235 ( .IN(net0106), .OUT(net0100), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I236 ( .IN(clkin_25), .OUT(net094), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I237 ( .IN(net0124), .OUT(net088), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I231 ( .IN(en_25), .OUT(net64), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd2vdd25_vpxa, View - schematic
// LAST TIME SAVED: Nov  6 18:00:25 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25_vpxa ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
nch_25  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));
pch_25  M0 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
pch_25  M1 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
pch_25  M2 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
pch_25  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));

endmodule
// Library - NVCM_40nm, Cell - ml_hv2vddp_sw, View - schematic
// LAST TIME SAVED: Nov 30 14:58:28 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hv2vddp_sw ( out_hv, hv2vddp, vddp_tieh, vpxa );
inout  out_hv;

input  hv2vddp, vddp_tieh, vpxa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ls_vdd2vdd25_vpxa I64 ( .in(net44), .sup(vddp_),
     .out_vddio_b(net060), .out_vddio(net37), .in_b(net46));
pch_25  M1 ( .D(net27), .B(out_hv), .G(sw_vpp_b), .S(out_hv));
pch_25  M0 ( .D(net27), .B(vddp_), .G(sw_vddp_b), .S(vddp_));
inv_25 I62 ( .IN(net37), .OUT(sw_vddp_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I71 ( .IN(net060), .OUT(net035), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I65 ( .A(hv2vddp), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(sw_vddp_b),
     .sel_25(net035), .out_b_hv(sw_vpp_b), .in_hv(out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ref, View - schematic
// LAST TIME SAVED: Oct  8 16:18:32 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpp_ref ( vref_25, bgr, pumpen_25, vppwl_25 );
inout  vref_25;

input  bgr, pumpen_25;

input [2:0]  vppwl_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_b_25;

wire  [7:0]  red_dec_25;



nand3_25 I44_7_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[7]),
     .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_6_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[6]),
     .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_5_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[5]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_4_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[4]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_3_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[3]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_2_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[2]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_1_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[1]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_0_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[0]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nch_25  M10 ( .D(net163), .B(GND_), .G(bgr), .S(gnd_));
nch_25  M14 ( .D(net0113), .B(GND_), .G(vppref_en_b_25), .S(gnd_));
nch_25  M15 ( .D(ctrl_gate_25), .B(GND_), .G(vppref_en_b_25),
     .S(gnd_));
nch_25  M8 ( .D(ctrl_gate_25), .B(GND_), .G(bgr_mirror_25),
     .S(net163));
nch_25  M13 ( .D(net0113), .B(GND_), .G(bgr), .S(net163));
nch_na25  M0 ( .D(net179), .B(GND_), .G(ctrl_gate_25),
     .S(bgr_mirror_25));
nmoscap_25  C3 ( .MINUS(net0129), .PLUS(net0113));
nmoscap_25  C2 ( .MINUS(gnd_), .PLUS(ctrl_gate_25));
rppolywo_m  R14 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R15 ( .MINUS(net104), .PLUS(net0216), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net0216), .PLUS(net139), .BULK(GND_));
rppolywo_m  R19 ( .MINUS(net139), .PLUS(net0213), .BULK(GND_));
rppolywo_m  R22 ( .MINUS(net0213), .PLUS(net98), .BULK(GND_));
rppolywo_m  R25 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R24 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(net0100), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(net0100), .PLUS(net0100), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(net0100), .PLUS(net0193), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net0193), .PLUS(net110), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(bgr_mirror_25), .PLUS(net0129), .BULK(GND_));
pch_25  M1 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(net175));
pch_25  M18 ( .D(net179), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
pch_25  M5 ( .D(ctrl_gate_25), .B(vddp_), .G(net0113), .S(net175));
pch_25  M6 ( .D(net0113), .B(vddp_), .G(net0113), .S(net175));
pch_25  M7 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
inv_25 I38 ( .IN(pumpen_25), .OUT(vppref_en_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_2_ ( .IN(vppwl_25[2]), .OUT(vppwl_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_1_ ( .IN(vppwl_25[1]), .OUT(vppwl_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_0_ ( .IN(vppwl_25[0]), .OUT(vppwl_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_vpp_ref_sw I281 ( .in(net0213), .out(vref_25),
     .sel_b_25(red_dec_25[6]));
ml_vpp_ref_sw I287 ( .in(net0216), .out(vref_25),
     .sel_b_25(red_dec_25[4]));
ml_vpp_ref_sw I283 ( .in(net98), .out(vref_25),
     .sel_b_25(red_dec_25[7]));
ml_vpp_ref_sw I290 ( .in(net0193), .out(vref_25),
     .sel_b_25(red_dec_25[0]));
ml_vpp_ref_sw I288 ( .in(net104), .out(vref_25),
     .sel_b_25(red_dec_25[3]));
ml_vpp_ref_sw I284 ( .in(net139), .out(vref_25),
     .sel_b_25(red_dec_25[5]));
ml_vpp_ref_sw I291 ( .in(net110), .out(vref_25),
     .sel_b_25(red_dec_25[1]));
ml_vpp_ref_sw I292 ( .in(net113), .out(vref_25),
     .sel_b_25(red_dec_25[2]));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ctrl, View - schematic
// LAST TIME SAVED: Nov  6 18:30:47 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpp_ctrl ( pumpen_25, vpint_en, vpp_2_vdd, vppdisc_vpxa,
     vppwl_25, vpxa, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_vpgmwl_buf, fsm_wgnden );
output  pumpen_25, vpint_en, vpp_2_vdd, vppdisc_vpxa;

inout  vpxa;

input  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint, fsm_wgnden;

output [2:0]  vppwl_25;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  net082;

wire  [0:2]  net092;

wire  [0:2]  net038;

wire  [0:2]  net068;



ml_ls_vdd2vdd25_vpxa I173 ( .in(fsm_pgmdisc_buf), .sup(vpxa),
     .out_vddio_b(net088), .out_vddio(net048), .in_b(net0106));
ml_dff_nvcm I77 ( .CLK(net084), .QN(vpp_pumpen_b), .R(pgm_dis),
     .D(vdd_tieh), .Q(vpp_pumpen));
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(net0122));
inv_25 I95_2_ ( .IN(net068[0]), .OUT(vppwl_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_1_ ( .IN(net068[1]), .OUT(vppwl_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_0_ ( .IN(net068[2]), .OUT(vppwl_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I81 ( .IN(net073), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(net088), .OUT(vppdisc_vpxa), .P(vpxa), .Pb(vpxa),
     .G(gnd_), .Gb(gnd_));
nand3_hvt I79 ( .C(net086), .A(fsm_pgm_buf), .Y(pgm_dis),
     .B(fsm_nvcmen_buf));
nor2_hvt I111 ( .A(vpp_pumpen_b), .B(net080), .Y(net0133));
nor2_hvt I87 ( .A(vpp_pumpen), .Y(net036), .B(fsm_pgmdisc_buf));
nand4_hvt I75 ( .D(fsm_pgm_buf), .C(fsm_lshven_buf), .A(net0127),
     .Y(net046), .B(net0127));
inv_hvt I107 ( .A(net0122), .Y(net0124));
inv_hvt I109 ( .A(fsm_pgmvfy_buf), .Y(net0127));
inv_hvt I131 ( .A(net049), .Y(net080));
inv_hvt I110_2_ ( .A(net092[0]), .Y(net082[0]));
inv_hvt I110_1_ ( .A(net092[1]), .Y(net082[1]));
inv_hvt I110_0_ ( .A(net092[2]), .Y(net082[2]));
inv_hvt I76 ( .A(net046), .Y(net084));
inv_hvt I108 ( .A(fsm_pgmdisc_buf), .Y(net0122));
inv_hvt I78 ( .A(net0124), .Y(net086));
inv_hvt I113 ( .A(vpp_pumpen_b), .Y(vpint_en));
inv_hvt I91 ( .A(net036), .Y(net089));
inv_hvt I90 ( .A(net089), .Y(vpp_2_vdd));
inv_hvt I98_2_ ( .A(fsm_vpgmwl_buf[2]), .Y(net092[0]));
inv_hvt I98_1_ ( .A(fsm_vpgmwl_buf[1]), .Y(net092[1]));
inv_hvt I98_0_ ( .A(fsm_vpgmwl_buf[0]), .Y(net092[2]));
inv_hvt I112 ( .A(net0133), .Y(net0134));
inv_hvt I101 ( .A(fsm_pgmdisc_buf), .Y(net0106));
nand2_hvt I104 ( .A(fsm_tm_xforce), .Y(net049), .B(fsm_tm_xvppint));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_ls_vdd2vdd25 I96_2_ ( .in(net082[0]), .sup(vddp_),
     .out_vddio_b(net068[0]), .out_vddio(net038[0]), .in_b(net092[0]));
ml_ls_vdd2vdd25 I96_1_ ( .in(net082[1]), .sup(vddp_),
     .out_vddio_b(net068[1]), .out_vddio(net038[1]), .in_b(net092[1]));
ml_ls_vdd2vdd25 I96_0_ ( .in(net082[2]), .sup(vddp_),
     .out_vddio_b(net068[2]), .out_vddio(net038[2]), .in_b(net092[2]));
ml_ls_vdd2vdd25 I84 ( .in(net0133), .sup(vddp_), .out_vddio_b(net073),
     .out_vddio(net074), .in_b(net0134));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_reg, View - schematic
// LAST TIME SAVED: Nov  8 10:29:35 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpp_reg ( slow_25, bgr, pbias_25, pump_in, vpp_int, vpxa,
     pumpen_25, vppdisc_vpxa, vref_25 );
output  slow_25;

inout  bgr, pbias_25, pump_in, vpp_int, vpxa;

input  pumpen_25, vppdisc_vpxa, vref_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I211 ( .IN(en_buf_b_25), .OUT(en_buf_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I212 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R5 ( .MINUS(net0165), .PLUS(vpp_int), .BULK(GND_));
rppolywo_m  R6 ( .MINUS(gnd_), .PLUS(net0178), .BULK(GND_));
rppolywo_m  R14 ( .MINUS(net0271), .PLUS(vdd_), .BULK(GND_));
rppolywo_m  R15 ( .MINUS(net0271), .PLUS(vdd_), .BULK(GND_));
rppolywo_m  R16 ( .MINUS(net0271), .PLUS(vdd_), .BULK(GND_));
rppolywo_m  R11 ( .MINUS(vdd_), .PLUS(net0271), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(vdd_), .PLUS(net0271), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(pump_gate), .PLUS(pump_in), .BULK(GND_));
rppolywo_m  R7 ( .MINUS(net0178), .PLUS(net0175), .BULK(GND_));
rppolywo_m  R13 ( .MINUS(vdd_), .PLUS(net0271), .BULK(GND_));
pch_25  M31 ( .D(net0203), .B(net0165), .G(dis_pgate_25), .S(net0165));
pch_25  M2 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
pch_25  M9 ( .D(net0200), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
pch_25  M8_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
pch_25  M8_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
pch_25  M14 ( .D(pump_opamp_out), .B(net125), .G(vref_25), .S(net125));
pch_25  M18 ( .D(net122), .B(vpp_int), .G(net122), .S(vpp_int));
pch_25  M13 ( .D(net124), .B(net125), .G(vdiv), .S(net125));
pch_25  M32 ( .D(dis_pgate_25), .B(vpxa), .G(dis_pgate_25), .S(vpxa));
pch_25  M33 ( .D(dis_pgate_25), .B(vpxa), .G(vppdisc_vpxa), .S(vpxa));
pch_25  M12 ( .D(net125), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M19 ( .D(net134), .B(net122), .G(net134), .S(net122));
pch_25  M21 ( .D(net138), .B(net134), .G(net138), .S(net134));
pch_25  M23 ( .D(net142), .B(net138), .G(net142), .S(net138));
pch_25  M24 ( .D(vdiv), .B(net142), .G(vdiv), .S(net142));
pch_25  M25 ( .D(net0224), .B(vdiv), .G(net0224), .S(vdiv));
nch_25  M40 ( .D(net0264), .B(GND_), .G(vppdisc_vpxa), .S(gnd_));
nch_25  M16 ( .D(net124), .B(GND_), .G(net124), .S(net155));
nch_25  M17 ( .D(net155), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M6 ( .D(vpp_int), .B(GND_), .G(en_buf_25), .S(net168));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
nch_25  M20 ( .D(slow_25), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M7 ( .D(net168), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M4 ( .D(dis_pgate_25), .B(GND_), .G(net0208), .S(net0264));
nch_25  M41 ( .D(net0224), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M15 ( .D(pump_opamp_out), .B(GND_), .G(net124), .S(net155));
nch_25  M0 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net0175));
nch_na25  M11 ( .D(net0199), .B(GND_), .G(vppdisc_vpxa), .S(net0271));
nch_na25  M22 ( .D(vpp_int), .B(GND_), .G(pump_gate), .S(pump_in));
nch_na25  M1 ( .D(GND_), .B(GND_), .G(pump_gate), .S(GND_));
nch_na25  M10 ( .D(net0203), .B(GND_), .G(net0208), .S(net0199));
nch_na25  M5 ( .D(pump_opamp_out), .B(GND_), .G(vpp_int),
     .S(pump_opamp_out));
vddp_tiehigh I261 ( .vddp_tieh(net0208));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_vco, View - schematic
// LAST TIME SAVED: Aug 25 11:10:03 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpp_vco ( clk_25_0, clk_25_1, pbias_25, slow_25, en_25,
     freq_25 );
output  clk_25_0, clk_25_1;

inout  pbias_25, slow_25;

input  en_25;

input [1:0]  freq_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:1]  freq_b_25;



nch_na25  M4 ( .D(GND_), .B(GND_), .G(net173), .S(GND_));
nch_na25  M15 ( .D(GND_), .B(GND_), .G(net185), .S(GND_));
nch_na25  M16 ( .D(GND_), .B(GND_), .G(net193), .S(GND_));
nch_na25  M2 ( .D(GND_), .B(GND_), .G(net189), .S(GND_));
nch_25  M5 ( .D(net173), .B(GND_), .G(net185), .S(net177));
nch_25  M6 ( .D(net177), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M13 ( .D(net181), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M14 ( .D(net185), .B(GND_), .G(net193), .S(net181));
nch_25  M8 ( .D(net189), .B(GND_), .G(net173), .S(net201));
nch_25  M17 ( .D(net193), .B(GND_), .G(net195), .S(net197));
nch_25  M18 ( .D(net197), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M1 ( .D(net201), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M23 ( .D(pbias_osc_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M24 ( .D(slow_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M25 ( .D(nbias_osc_25), .B(GND_), .G(en_25), .S(slow_25));
nand2_25 I96 ( .G(GND_), .Pb(vddp_), .A(net189), .Y(net195), .P(vddp_),
     .B(en_25), .Gb(GND_));
nand2_25 I205 ( .G(GND_), .Pb(vddp_), .A(net185), .Y(net0205),
     .P(vddp_), .B(en_25), .Gb(GND_));
pch_25  M7 ( .D(net173), .B(vddp_), .G(net185), .S(net236));
pch_25  M10 ( .D(net236), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M9 ( .D(net248), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M3 ( .D(net189), .B(vddp_), .G(net173), .S(net248));
pch_25  M11 ( .D(net256), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M12 ( .D(net185), .B(vddp_), .G(net193), .S(net256));
pch_25  M19 ( .D(net193), .B(vddp_), .G(net195), .S(net260));
pch_25  M20 ( .D(net260), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M22 ( .D(pbias_osc_25), .B(vddp_), .G(en_b_25), .S(net228));
pch_25  M26_1_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M26_0_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_1_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_0_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M28 ( .D(net212), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M29 ( .D(nbias_osc_25), .B(vddp_), .G(freq_25[0]), .S(net212));
pch_25  M30 ( .D(nbias_osc_25), .B(vddp_), .G(freq_b_25[1]),
     .S(net208));
pch_25  M21 ( .D(net228), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
inv_25 I201 ( .IN(net195), .OUT(clk_25_0), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(net0205), .OUT(clk_25_1), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I188 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I199 ( .IN(freq_25[1]), .OUT(freq_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));

endmodule
// Library - NVCM_40nm, Cell - ml_vppint_top, View - schematic
// LAST TIME SAVED: Nov  6 18:24:09 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vppint_top ( vpint_en, vpp_int, vpxa, bgr, fsm_lshven_buf,
     fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf, fsm_pgmvfy_buf,
     fsm_tm_xforce, fsm_tm_xvppint, fsm_vpgmwl_buf, fsm_wgnden_buf );
output  vpint_en;

inout  vpp_int, vpxa;

input  bgr, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_wgnden_buf;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_25;

wire  [1:0]  freq_25;



ml_pump_vpxa_buf I95 ( .in(clkin_0_25), .out(net52));
ml_pump_vpxa_buf I81 ( .in(clkin_1_25), .out(net061));
ml_vpp_pump Ivpp_pump_0 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(clkin_1_25));
ml_vpp_pump Ivpp_pump_1 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net061));
ml_vpp_pump Ivpp_pump_2 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net52));
inv_25 I38 ( .IN(vddp_tieh), .OUT(freq_25[1]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I91 ( .IN(vddp_tieh), .OUT(freq_25[0]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpp_int));
ml_hv2vddp_sw Ivpxa_2vddp_sw ( .vpxa(vpxa), .hv2vddp(vpp_2_vdd),
     .vddp_tieh(vddp_tieh), .out_hv(vpp_int));
ml_vpp_ref Ivpp_ref ( .vref_25(vref_25), .vppwl_25(vppwl_25[2:0]),
     .pumpen_25(pumpen_25), .bgr(bgr));
ml_vpp_ctrl Ivpp_ctrl ( .vppdisc_vpxa(vppdisc_vpxa), .vpxa(vpxa),
     .vpint_en(vpint_en), .fsm_pgmvfy_buf(fsm_pgmvfy_buf),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .fsm_wgnden(fsm_wgnden_buf),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf), .vppwl_25(vppwl_25[2:0]),
     .vpp_2_vdd(vpp_2_vdd), .pumpen_25(pumpen_25));
ml_vpp_reg Ivpp_reg ( .vpxa(vpxa), .vppdisc_vpxa(vppdisc_vpxa),
     .bgr(bgr), .slow_25(slow_25), .pbias_25(pbias_25),
     .vref_25(vref_25), .pumpen_25(pumpen_25), .pump_in(pump_in),
     .vpp_int(vpp_int));
ml_vpp_vco Ivpp_vco ( .clk_25_1(clkin_1_25), .pbias_25(pbias_25),
     .slow_25(slow_25), .freq_25(freq_25[1:0]), .en_25(pumpen_25),
     .clk_25_0(clkin_0_25));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_3.3v, View - schematic
// LAST TIME SAVED: Aug 30 18:07:58 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_pump_vpxa_3_3v ( out, clkin_25, en_25 );
inout  out;

input  clkin_25, en_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C1 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C2 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C3 ( .MINUS(clk_25), .PLUS(s_2));
nch_na25  M1 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
nch_na25  M2 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
nch_na25  M3 ( .D(s_2), .B(GND_), .G(s_2), .S(out));
nch_na25  M4 ( .D(net73), .B(GND_), .G(net73), .S(s_0));
pch_25  M6 ( .D(net73), .B(vddp_), .G(net114), .S(vddp_));
inv_25 I230 ( .IN(clkin_25), .OUT(net120), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I231 ( .IN(en_25), .OUT(net114), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I232 ( .IN(net78), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I233 ( .IN(net90), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I234 ( .IN(net84), .OUT(net96), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I235 ( .IN(net96), .OUT(net90), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I236 ( .IN(clkin_25), .OUT(net84), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I237 ( .IN(net120), .OUT(net78), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));

endmodule
// Library - sbtlibn65lp, Cell - ml_dlatch_25, View - schematic
// LAST TIME SAVED: Aug 30 17:06:09 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_dlatch_25 ( Q_25, D_25, EN_25, R_25 );
output  Q_25;

input  D_25, EN_25, R_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_25 I161 ( .A(net52), .Y(Q_25), .Gb(GND_), .G(GND_), .Pb(vddp_),
     .P(vddp_), .B(R_25));
inv_25 I156 ( .IN(EN_25), .OUT(EN_B_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nch_25  M0 ( .D(net52), .B(GND_), .G(D_25), .S(net48));
nch_25  M1 ( .D(net48), .B(GND_), .G(EN_25), .S(GND_));
nch_25  M5 ( .D(net40), .B(GND_), .G(EN_B_25), .S(GND_));
nch_25  M6 ( .D(net52), .B(GND_), .G(Q_25), .S(net40));
pch_25  M2 ( .D(net52), .B(vddp_), .G(Q_25), .S(net31));
pch_25  M8 ( .D(net31), .B(vddp_), .G(EN_25), .S(vddp_));
pch_25  M7 ( .D(net39), .B(vddp_), .G(EN_B_25), .S(vddp_));
pch_25  M3 ( .D(net52), .B(vddp_), .G(D_25), .S(net39));

endmodule
// Library - ice1chip, Cell - ice1f_cram_row142col4, View - schematic
// LAST TIME SAVED: Mar 10 12:33:59 2011
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module ice1f_cram_row142col4 ( bl, pgate_l, pgate_r, reset_l, reset_r,
     vdd_cntl_l, vdd_cntl_r, wl_l, wl_r );


inout [3:0]  bl;

input [141:0]  wl_r;
input [141:0]  pgate_l;
input [141:0]  wl_l;
input [141:0]  reset_r;
input [141:0]  vdd_cntl_r;
input [141:0]  pgate_r;
input [141:0]  reset_l;
input [141:0]  vdd_cntl_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:567]  net35;

wire  [0:567]  net36;

wire  [141:0]  r_gnd_r;

wire  [141:0]  r_gnd_l;



pch_hvt  M0_141_ ( .D(r_gnd_r[141]), .B(vdd_), .G(vdd_cntl_r[141]),
     .S(vdd_));
pch_hvt  M0_140_ ( .D(r_gnd_r[140]), .B(vdd_), .G(vdd_cntl_r[140]),
     .S(vdd_));
pch_hvt  M0_139_ ( .D(r_gnd_r[139]), .B(vdd_), .G(vdd_cntl_r[139]),
     .S(vdd_));
pch_hvt  M0_138_ ( .D(r_gnd_r[138]), .B(vdd_), .G(vdd_cntl_r[138]),
     .S(vdd_));
pch_hvt  M0_137_ ( .D(r_gnd_r[137]), .B(vdd_), .G(vdd_cntl_r[137]),
     .S(vdd_));
pch_hvt  M0_136_ ( .D(r_gnd_r[136]), .B(vdd_), .G(vdd_cntl_r[136]),
     .S(vdd_));
pch_hvt  M0_135_ ( .D(r_gnd_r[135]), .B(vdd_), .G(vdd_cntl_r[135]),
     .S(vdd_));
pch_hvt  M0_134_ ( .D(r_gnd_r[134]), .B(vdd_), .G(vdd_cntl_r[134]),
     .S(vdd_));
pch_hvt  M0_133_ ( .D(r_gnd_r[133]), .B(vdd_), .G(vdd_cntl_r[133]),
     .S(vdd_));
pch_hvt  M0_132_ ( .D(r_gnd_r[132]), .B(vdd_), .G(vdd_cntl_r[132]),
     .S(vdd_));
pch_hvt  M0_131_ ( .D(r_gnd_r[131]), .B(vdd_), .G(vdd_cntl_r[131]),
     .S(vdd_));
pch_hvt  M0_130_ ( .D(r_gnd_r[130]), .B(vdd_), .G(vdd_cntl_r[130]),
     .S(vdd_));
pch_hvt  M0_129_ ( .D(r_gnd_r[129]), .B(vdd_), .G(vdd_cntl_r[129]),
     .S(vdd_));
pch_hvt  M0_128_ ( .D(r_gnd_r[128]), .B(vdd_), .G(vdd_cntl_r[128]),
     .S(vdd_));
pch_hvt  M0_127_ ( .D(r_gnd_r[127]), .B(vdd_), .G(vdd_cntl_r[127]),
     .S(vdd_));
pch_hvt  M0_126_ ( .D(r_gnd_r[126]), .B(vdd_), .G(vdd_cntl_r[126]),
     .S(vdd_));
pch_hvt  M0_125_ ( .D(r_gnd_r[125]), .B(vdd_), .G(vdd_cntl_r[125]),
     .S(vdd_));
pch_hvt  M0_124_ ( .D(r_gnd_r[124]), .B(vdd_), .G(vdd_cntl_r[124]),
     .S(vdd_));
pch_hvt  M0_123_ ( .D(r_gnd_r[123]), .B(vdd_), .G(vdd_cntl_r[123]),
     .S(vdd_));
pch_hvt  M0_122_ ( .D(r_gnd_r[122]), .B(vdd_), .G(vdd_cntl_r[122]),
     .S(vdd_));
pch_hvt  M0_121_ ( .D(r_gnd_r[121]), .B(vdd_), .G(vdd_cntl_r[121]),
     .S(vdd_));
pch_hvt  M0_120_ ( .D(r_gnd_r[120]), .B(vdd_), .G(vdd_cntl_r[120]),
     .S(vdd_));
pch_hvt  M0_119_ ( .D(r_gnd_r[119]), .B(vdd_), .G(vdd_cntl_r[119]),
     .S(vdd_));
pch_hvt  M0_118_ ( .D(r_gnd_r[118]), .B(vdd_), .G(vdd_cntl_r[118]),
     .S(vdd_));
pch_hvt  M0_117_ ( .D(r_gnd_r[117]), .B(vdd_), .G(vdd_cntl_r[117]),
     .S(vdd_));
pch_hvt  M0_116_ ( .D(r_gnd_r[116]), .B(vdd_), .G(vdd_cntl_r[116]),
     .S(vdd_));
pch_hvt  M0_115_ ( .D(r_gnd_r[115]), .B(vdd_), .G(vdd_cntl_r[115]),
     .S(vdd_));
pch_hvt  M0_114_ ( .D(r_gnd_r[114]), .B(vdd_), .G(vdd_cntl_r[114]),
     .S(vdd_));
pch_hvt  M0_113_ ( .D(r_gnd_r[113]), .B(vdd_), .G(vdd_cntl_r[113]),
     .S(vdd_));
pch_hvt  M0_112_ ( .D(r_gnd_r[112]), .B(vdd_), .G(vdd_cntl_r[112]),
     .S(vdd_));
pch_hvt  M0_111_ ( .D(r_gnd_r[111]), .B(vdd_), .G(vdd_cntl_r[111]),
     .S(vdd_));
pch_hvt  M0_110_ ( .D(r_gnd_r[110]), .B(vdd_), .G(vdd_cntl_r[110]),
     .S(vdd_));
pch_hvt  M0_109_ ( .D(r_gnd_r[109]), .B(vdd_), .G(vdd_cntl_r[109]),
     .S(vdd_));
pch_hvt  M0_108_ ( .D(r_gnd_r[108]), .B(vdd_), .G(vdd_cntl_r[108]),
     .S(vdd_));
pch_hvt  M0_107_ ( .D(r_gnd_r[107]), .B(vdd_), .G(vdd_cntl_r[107]),
     .S(vdd_));
pch_hvt  M0_106_ ( .D(r_gnd_r[106]), .B(vdd_), .G(vdd_cntl_r[106]),
     .S(vdd_));
pch_hvt  M0_105_ ( .D(r_gnd_r[105]), .B(vdd_), .G(vdd_cntl_r[105]),
     .S(vdd_));
pch_hvt  M0_104_ ( .D(r_gnd_r[104]), .B(vdd_), .G(vdd_cntl_r[104]),
     .S(vdd_));
pch_hvt  M0_103_ ( .D(r_gnd_r[103]), .B(vdd_), .G(vdd_cntl_r[103]),
     .S(vdd_));
pch_hvt  M0_102_ ( .D(r_gnd_r[102]), .B(vdd_), .G(vdd_cntl_r[102]),
     .S(vdd_));
pch_hvt  M0_101_ ( .D(r_gnd_r[101]), .B(vdd_), .G(vdd_cntl_r[101]),
     .S(vdd_));
pch_hvt  M0_100_ ( .D(r_gnd_r[100]), .B(vdd_), .G(vdd_cntl_r[100]),
     .S(vdd_));
pch_hvt  M0_99_ ( .D(r_gnd_r[99]), .B(vdd_), .G(vdd_cntl_r[99]),
     .S(vdd_));
pch_hvt  M0_98_ ( .D(r_gnd_r[98]), .B(vdd_), .G(vdd_cntl_r[98]),
     .S(vdd_));
pch_hvt  M0_97_ ( .D(r_gnd_r[97]), .B(vdd_), .G(vdd_cntl_r[97]),
     .S(vdd_));
pch_hvt  M0_96_ ( .D(r_gnd_r[96]), .B(vdd_), .G(vdd_cntl_r[96]),
     .S(vdd_));
pch_hvt  M0_95_ ( .D(r_gnd_r[95]), .B(vdd_), .G(vdd_cntl_r[95]),
     .S(vdd_));
pch_hvt  M0_94_ ( .D(r_gnd_r[94]), .B(vdd_), .G(vdd_cntl_r[94]),
     .S(vdd_));
pch_hvt  M0_93_ ( .D(r_gnd_r[93]), .B(vdd_), .G(vdd_cntl_r[93]),
     .S(vdd_));
pch_hvt  M0_92_ ( .D(r_gnd_r[92]), .B(vdd_), .G(vdd_cntl_r[92]),
     .S(vdd_));
pch_hvt  M0_91_ ( .D(r_gnd_r[91]), .B(vdd_), .G(vdd_cntl_r[91]),
     .S(vdd_));
pch_hvt  M0_90_ ( .D(r_gnd_r[90]), .B(vdd_), .G(vdd_cntl_r[90]),
     .S(vdd_));
pch_hvt  M0_89_ ( .D(r_gnd_r[89]), .B(vdd_), .G(vdd_cntl_r[89]),
     .S(vdd_));
pch_hvt  M0_88_ ( .D(r_gnd_r[88]), .B(vdd_), .G(vdd_cntl_r[88]),
     .S(vdd_));
pch_hvt  M0_87_ ( .D(r_gnd_r[87]), .B(vdd_), .G(vdd_cntl_r[87]),
     .S(vdd_));
pch_hvt  M0_86_ ( .D(r_gnd_r[86]), .B(vdd_), .G(vdd_cntl_r[86]),
     .S(vdd_));
pch_hvt  M0_85_ ( .D(r_gnd_r[85]), .B(vdd_), .G(vdd_cntl_r[85]),
     .S(vdd_));
pch_hvt  M0_84_ ( .D(r_gnd_r[84]), .B(vdd_), .G(vdd_cntl_r[84]),
     .S(vdd_));
pch_hvt  M0_83_ ( .D(r_gnd_r[83]), .B(vdd_), .G(vdd_cntl_r[83]),
     .S(vdd_));
pch_hvt  M0_82_ ( .D(r_gnd_r[82]), .B(vdd_), .G(vdd_cntl_r[82]),
     .S(vdd_));
pch_hvt  M0_81_ ( .D(r_gnd_r[81]), .B(vdd_), .G(vdd_cntl_r[81]),
     .S(vdd_));
pch_hvt  M0_80_ ( .D(r_gnd_r[80]), .B(vdd_), .G(vdd_cntl_r[80]),
     .S(vdd_));
pch_hvt  M0_79_ ( .D(r_gnd_r[79]), .B(vdd_), .G(vdd_cntl_r[79]),
     .S(vdd_));
pch_hvt  M0_78_ ( .D(r_gnd_r[78]), .B(vdd_), .G(vdd_cntl_r[78]),
     .S(vdd_));
pch_hvt  M0_77_ ( .D(r_gnd_r[77]), .B(vdd_), .G(vdd_cntl_r[77]),
     .S(vdd_));
pch_hvt  M0_76_ ( .D(r_gnd_r[76]), .B(vdd_), .G(vdd_cntl_r[76]),
     .S(vdd_));
pch_hvt  M0_75_ ( .D(r_gnd_r[75]), .B(vdd_), .G(vdd_cntl_r[75]),
     .S(vdd_));
pch_hvt  M0_74_ ( .D(r_gnd_r[74]), .B(vdd_), .G(vdd_cntl_r[74]),
     .S(vdd_));
pch_hvt  M0_73_ ( .D(r_gnd_r[73]), .B(vdd_), .G(vdd_cntl_r[73]),
     .S(vdd_));
pch_hvt  M0_72_ ( .D(r_gnd_r[72]), .B(vdd_), .G(vdd_cntl_r[72]),
     .S(vdd_));
pch_hvt  M0_71_ ( .D(r_gnd_r[71]), .B(vdd_), .G(vdd_cntl_r[71]),
     .S(vdd_));
pch_hvt  M0_70_ ( .D(r_gnd_r[70]), .B(vdd_), .G(vdd_cntl_r[70]),
     .S(vdd_));
pch_hvt  M0_69_ ( .D(r_gnd_r[69]), .B(vdd_), .G(vdd_cntl_r[69]),
     .S(vdd_));
pch_hvt  M0_68_ ( .D(r_gnd_r[68]), .B(vdd_), .G(vdd_cntl_r[68]),
     .S(vdd_));
pch_hvt  M0_67_ ( .D(r_gnd_r[67]), .B(vdd_), .G(vdd_cntl_r[67]),
     .S(vdd_));
pch_hvt  M0_66_ ( .D(r_gnd_r[66]), .B(vdd_), .G(vdd_cntl_r[66]),
     .S(vdd_));
pch_hvt  M0_65_ ( .D(r_gnd_r[65]), .B(vdd_), .G(vdd_cntl_r[65]),
     .S(vdd_));
pch_hvt  M0_64_ ( .D(r_gnd_r[64]), .B(vdd_), .G(vdd_cntl_r[64]),
     .S(vdd_));
pch_hvt  M0_63_ ( .D(r_gnd_r[63]), .B(vdd_), .G(vdd_cntl_r[63]),
     .S(vdd_));
pch_hvt  M0_62_ ( .D(r_gnd_r[62]), .B(vdd_), .G(vdd_cntl_r[62]),
     .S(vdd_));
pch_hvt  M0_61_ ( .D(r_gnd_r[61]), .B(vdd_), .G(vdd_cntl_r[61]),
     .S(vdd_));
pch_hvt  M0_60_ ( .D(r_gnd_r[60]), .B(vdd_), .G(vdd_cntl_r[60]),
     .S(vdd_));
pch_hvt  M0_59_ ( .D(r_gnd_r[59]), .B(vdd_), .G(vdd_cntl_r[59]),
     .S(vdd_));
pch_hvt  M0_58_ ( .D(r_gnd_r[58]), .B(vdd_), .G(vdd_cntl_r[58]),
     .S(vdd_));
pch_hvt  M0_57_ ( .D(r_gnd_r[57]), .B(vdd_), .G(vdd_cntl_r[57]),
     .S(vdd_));
pch_hvt  M0_56_ ( .D(r_gnd_r[56]), .B(vdd_), .G(vdd_cntl_r[56]),
     .S(vdd_));
pch_hvt  M0_55_ ( .D(r_gnd_r[55]), .B(vdd_), .G(vdd_cntl_r[55]),
     .S(vdd_));
pch_hvt  M0_54_ ( .D(r_gnd_r[54]), .B(vdd_), .G(vdd_cntl_r[54]),
     .S(vdd_));
pch_hvt  M0_53_ ( .D(r_gnd_r[53]), .B(vdd_), .G(vdd_cntl_r[53]),
     .S(vdd_));
pch_hvt  M0_52_ ( .D(r_gnd_r[52]), .B(vdd_), .G(vdd_cntl_r[52]),
     .S(vdd_));
pch_hvt  M0_51_ ( .D(r_gnd_r[51]), .B(vdd_), .G(vdd_cntl_r[51]),
     .S(vdd_));
pch_hvt  M0_50_ ( .D(r_gnd_r[50]), .B(vdd_), .G(vdd_cntl_r[50]),
     .S(vdd_));
pch_hvt  M0_49_ ( .D(r_gnd_r[49]), .B(vdd_), .G(vdd_cntl_r[49]),
     .S(vdd_));
pch_hvt  M0_48_ ( .D(r_gnd_r[48]), .B(vdd_), .G(vdd_cntl_r[48]),
     .S(vdd_));
pch_hvt  M0_47_ ( .D(r_gnd_r[47]), .B(vdd_), .G(vdd_cntl_r[47]),
     .S(vdd_));
pch_hvt  M0_46_ ( .D(r_gnd_r[46]), .B(vdd_), .G(vdd_cntl_r[46]),
     .S(vdd_));
pch_hvt  M0_45_ ( .D(r_gnd_r[45]), .B(vdd_), .G(vdd_cntl_r[45]),
     .S(vdd_));
pch_hvt  M0_44_ ( .D(r_gnd_r[44]), .B(vdd_), .G(vdd_cntl_r[44]),
     .S(vdd_));
pch_hvt  M0_43_ ( .D(r_gnd_r[43]), .B(vdd_), .G(vdd_cntl_r[43]),
     .S(vdd_));
pch_hvt  M0_42_ ( .D(r_gnd_r[42]), .B(vdd_), .G(vdd_cntl_r[42]),
     .S(vdd_));
pch_hvt  M0_41_ ( .D(r_gnd_r[41]), .B(vdd_), .G(vdd_cntl_r[41]),
     .S(vdd_));
pch_hvt  M0_40_ ( .D(r_gnd_r[40]), .B(vdd_), .G(vdd_cntl_r[40]),
     .S(vdd_));
pch_hvt  M0_39_ ( .D(r_gnd_r[39]), .B(vdd_), .G(vdd_cntl_r[39]),
     .S(vdd_));
pch_hvt  M0_38_ ( .D(r_gnd_r[38]), .B(vdd_), .G(vdd_cntl_r[38]),
     .S(vdd_));
pch_hvt  M0_37_ ( .D(r_gnd_r[37]), .B(vdd_), .G(vdd_cntl_r[37]),
     .S(vdd_));
pch_hvt  M0_36_ ( .D(r_gnd_r[36]), .B(vdd_), .G(vdd_cntl_r[36]),
     .S(vdd_));
pch_hvt  M0_35_ ( .D(r_gnd_r[35]), .B(vdd_), .G(vdd_cntl_r[35]),
     .S(vdd_));
pch_hvt  M0_34_ ( .D(r_gnd_r[34]), .B(vdd_), .G(vdd_cntl_r[34]),
     .S(vdd_));
pch_hvt  M0_33_ ( .D(r_gnd_r[33]), .B(vdd_), .G(vdd_cntl_r[33]),
     .S(vdd_));
pch_hvt  M0_32_ ( .D(r_gnd_r[32]), .B(vdd_), .G(vdd_cntl_r[32]),
     .S(vdd_));
pch_hvt  M0_31_ ( .D(r_gnd_r[31]), .B(vdd_), .G(vdd_cntl_r[31]),
     .S(vdd_));
pch_hvt  M0_30_ ( .D(r_gnd_r[30]), .B(vdd_), .G(vdd_cntl_r[30]),
     .S(vdd_));
pch_hvt  M0_29_ ( .D(r_gnd_r[29]), .B(vdd_), .G(vdd_cntl_r[29]),
     .S(vdd_));
pch_hvt  M0_28_ ( .D(r_gnd_r[28]), .B(vdd_), .G(vdd_cntl_r[28]),
     .S(vdd_));
pch_hvt  M0_27_ ( .D(r_gnd_r[27]), .B(vdd_), .G(vdd_cntl_r[27]),
     .S(vdd_));
pch_hvt  M0_26_ ( .D(r_gnd_r[26]), .B(vdd_), .G(vdd_cntl_r[26]),
     .S(vdd_));
pch_hvt  M0_25_ ( .D(r_gnd_r[25]), .B(vdd_), .G(vdd_cntl_r[25]),
     .S(vdd_));
pch_hvt  M0_24_ ( .D(r_gnd_r[24]), .B(vdd_), .G(vdd_cntl_r[24]),
     .S(vdd_));
pch_hvt  M0_23_ ( .D(r_gnd_r[23]), .B(vdd_), .G(vdd_cntl_r[23]),
     .S(vdd_));
pch_hvt  M0_22_ ( .D(r_gnd_r[22]), .B(vdd_), .G(vdd_cntl_r[22]),
     .S(vdd_));
pch_hvt  M0_21_ ( .D(r_gnd_r[21]), .B(vdd_), .G(vdd_cntl_r[21]),
     .S(vdd_));
pch_hvt  M0_20_ ( .D(r_gnd_r[20]), .B(vdd_), .G(vdd_cntl_r[20]),
     .S(vdd_));
pch_hvt  M0_19_ ( .D(r_gnd_r[19]), .B(vdd_), .G(vdd_cntl_r[19]),
     .S(vdd_));
pch_hvt  M0_18_ ( .D(r_gnd_r[18]), .B(vdd_), .G(vdd_cntl_r[18]),
     .S(vdd_));
pch_hvt  M0_17_ ( .D(r_gnd_r[17]), .B(vdd_), .G(vdd_cntl_r[17]),
     .S(vdd_));
pch_hvt  M0_16_ ( .D(r_gnd_r[16]), .B(vdd_), .G(vdd_cntl_r[16]),
     .S(vdd_));
pch_hvt  M0_15_ ( .D(r_gnd_r[15]), .B(vdd_), .G(vdd_cntl_r[15]),
     .S(vdd_));
pch_hvt  M0_14_ ( .D(r_gnd_r[14]), .B(vdd_), .G(vdd_cntl_r[14]),
     .S(vdd_));
pch_hvt  M0_13_ ( .D(r_gnd_r[13]), .B(vdd_), .G(vdd_cntl_r[13]),
     .S(vdd_));
pch_hvt  M0_12_ ( .D(r_gnd_r[12]), .B(vdd_), .G(vdd_cntl_r[12]),
     .S(vdd_));
pch_hvt  M0_11_ ( .D(r_gnd_r[11]), .B(vdd_), .G(vdd_cntl_r[11]),
     .S(vdd_));
pch_hvt  M0_10_ ( .D(r_gnd_r[10]), .B(vdd_), .G(vdd_cntl_r[10]),
     .S(vdd_));
pch_hvt  M0_9_ ( .D(r_gnd_r[9]), .B(vdd_), .G(vdd_cntl_r[9]),
     .S(vdd_));
pch_hvt  M0_8_ ( .D(r_gnd_r[8]), .B(vdd_), .G(vdd_cntl_r[8]),
     .S(vdd_));
pch_hvt  M0_7_ ( .D(r_gnd_r[7]), .B(vdd_), .G(vdd_cntl_r[7]),
     .S(vdd_));
pch_hvt  M0_6_ ( .D(r_gnd_r[6]), .B(vdd_), .G(vdd_cntl_r[6]),
     .S(vdd_));
pch_hvt  M0_5_ ( .D(r_gnd_r[5]), .B(vdd_), .G(vdd_cntl_r[5]),
     .S(vdd_));
pch_hvt  M0_4_ ( .D(r_gnd_r[4]), .B(vdd_), .G(vdd_cntl_r[4]),
     .S(vdd_));
pch_hvt  M0_3_ ( .D(r_gnd_r[3]), .B(vdd_), .G(vdd_cntl_r[3]),
     .S(vdd_));
pch_hvt  M0_2_ ( .D(r_gnd_r[2]), .B(vdd_), .G(vdd_cntl_r[2]),
     .S(vdd_));
pch_hvt  M0_1_ ( .D(r_gnd_r[1]), .B(vdd_), .G(vdd_cntl_r[1]),
     .S(vdd_));
pch_hvt  M0_0_ ( .D(r_gnd_r[0]), .B(vdd_), .G(vdd_cntl_r[0]),
     .S(vdd_));
pch_hvt  M3_141_ ( .D(r_gnd_l[141]), .B(vdd_), .G(vdd_cntl_l[141]),
     .S(vdd_));
pch_hvt  M3_140_ ( .D(r_gnd_l[140]), .B(vdd_), .G(vdd_cntl_l[140]),
     .S(vdd_));
pch_hvt  M3_139_ ( .D(r_gnd_l[139]), .B(vdd_), .G(vdd_cntl_l[139]),
     .S(vdd_));
pch_hvt  M3_138_ ( .D(r_gnd_l[138]), .B(vdd_), .G(vdd_cntl_l[138]),
     .S(vdd_));
pch_hvt  M3_137_ ( .D(r_gnd_l[137]), .B(vdd_), .G(vdd_cntl_l[137]),
     .S(vdd_));
pch_hvt  M3_136_ ( .D(r_gnd_l[136]), .B(vdd_), .G(vdd_cntl_l[136]),
     .S(vdd_));
pch_hvt  M3_135_ ( .D(r_gnd_l[135]), .B(vdd_), .G(vdd_cntl_l[135]),
     .S(vdd_));
pch_hvt  M3_134_ ( .D(r_gnd_l[134]), .B(vdd_), .G(vdd_cntl_l[134]),
     .S(vdd_));
pch_hvt  M3_133_ ( .D(r_gnd_l[133]), .B(vdd_), .G(vdd_cntl_l[133]),
     .S(vdd_));
pch_hvt  M3_132_ ( .D(r_gnd_l[132]), .B(vdd_), .G(vdd_cntl_l[132]),
     .S(vdd_));
pch_hvt  M3_131_ ( .D(r_gnd_l[131]), .B(vdd_), .G(vdd_cntl_l[131]),
     .S(vdd_));
pch_hvt  M3_130_ ( .D(r_gnd_l[130]), .B(vdd_), .G(vdd_cntl_l[130]),
     .S(vdd_));
pch_hvt  M3_129_ ( .D(r_gnd_l[129]), .B(vdd_), .G(vdd_cntl_l[129]),
     .S(vdd_));
pch_hvt  M3_128_ ( .D(r_gnd_l[128]), .B(vdd_), .G(vdd_cntl_l[128]),
     .S(vdd_));
pch_hvt  M3_127_ ( .D(r_gnd_l[127]), .B(vdd_), .G(vdd_cntl_l[127]),
     .S(vdd_));
pch_hvt  M3_126_ ( .D(r_gnd_l[126]), .B(vdd_), .G(vdd_cntl_l[126]),
     .S(vdd_));
pch_hvt  M3_125_ ( .D(r_gnd_l[125]), .B(vdd_), .G(vdd_cntl_l[125]),
     .S(vdd_));
pch_hvt  M3_124_ ( .D(r_gnd_l[124]), .B(vdd_), .G(vdd_cntl_l[124]),
     .S(vdd_));
pch_hvt  M3_123_ ( .D(r_gnd_l[123]), .B(vdd_), .G(vdd_cntl_l[123]),
     .S(vdd_));
pch_hvt  M3_122_ ( .D(r_gnd_l[122]), .B(vdd_), .G(vdd_cntl_l[122]),
     .S(vdd_));
pch_hvt  M3_121_ ( .D(r_gnd_l[121]), .B(vdd_), .G(vdd_cntl_l[121]),
     .S(vdd_));
pch_hvt  M3_120_ ( .D(r_gnd_l[120]), .B(vdd_), .G(vdd_cntl_l[120]),
     .S(vdd_));
pch_hvt  M3_119_ ( .D(r_gnd_l[119]), .B(vdd_), .G(vdd_cntl_l[119]),
     .S(vdd_));
pch_hvt  M3_118_ ( .D(r_gnd_l[118]), .B(vdd_), .G(vdd_cntl_l[118]),
     .S(vdd_));
pch_hvt  M3_117_ ( .D(r_gnd_l[117]), .B(vdd_), .G(vdd_cntl_l[117]),
     .S(vdd_));
pch_hvt  M3_116_ ( .D(r_gnd_l[116]), .B(vdd_), .G(vdd_cntl_l[116]),
     .S(vdd_));
pch_hvt  M3_115_ ( .D(r_gnd_l[115]), .B(vdd_), .G(vdd_cntl_l[115]),
     .S(vdd_));
pch_hvt  M3_114_ ( .D(r_gnd_l[114]), .B(vdd_), .G(vdd_cntl_l[114]),
     .S(vdd_));
pch_hvt  M3_113_ ( .D(r_gnd_l[113]), .B(vdd_), .G(vdd_cntl_l[113]),
     .S(vdd_));
pch_hvt  M3_112_ ( .D(r_gnd_l[112]), .B(vdd_), .G(vdd_cntl_l[112]),
     .S(vdd_));
pch_hvt  M3_111_ ( .D(r_gnd_l[111]), .B(vdd_), .G(vdd_cntl_l[111]),
     .S(vdd_));
pch_hvt  M3_110_ ( .D(r_gnd_l[110]), .B(vdd_), .G(vdd_cntl_l[110]),
     .S(vdd_));
pch_hvt  M3_109_ ( .D(r_gnd_l[109]), .B(vdd_), .G(vdd_cntl_l[109]),
     .S(vdd_));
pch_hvt  M3_108_ ( .D(r_gnd_l[108]), .B(vdd_), .G(vdd_cntl_l[108]),
     .S(vdd_));
pch_hvt  M3_107_ ( .D(r_gnd_l[107]), .B(vdd_), .G(vdd_cntl_l[107]),
     .S(vdd_));
pch_hvt  M3_106_ ( .D(r_gnd_l[106]), .B(vdd_), .G(vdd_cntl_l[106]),
     .S(vdd_));
pch_hvt  M3_105_ ( .D(r_gnd_l[105]), .B(vdd_), .G(vdd_cntl_l[105]),
     .S(vdd_));
pch_hvt  M3_104_ ( .D(r_gnd_l[104]), .B(vdd_), .G(vdd_cntl_l[104]),
     .S(vdd_));
pch_hvt  M3_103_ ( .D(r_gnd_l[103]), .B(vdd_), .G(vdd_cntl_l[103]),
     .S(vdd_));
pch_hvt  M3_102_ ( .D(r_gnd_l[102]), .B(vdd_), .G(vdd_cntl_l[102]),
     .S(vdd_));
pch_hvt  M3_101_ ( .D(r_gnd_l[101]), .B(vdd_), .G(vdd_cntl_l[101]),
     .S(vdd_));
pch_hvt  M3_100_ ( .D(r_gnd_l[100]), .B(vdd_), .G(vdd_cntl_l[100]),
     .S(vdd_));
pch_hvt  M3_99_ ( .D(r_gnd_l[99]), .B(vdd_), .G(vdd_cntl_l[99]),
     .S(vdd_));
pch_hvt  M3_98_ ( .D(r_gnd_l[98]), .B(vdd_), .G(vdd_cntl_l[98]),
     .S(vdd_));
pch_hvt  M3_97_ ( .D(r_gnd_l[97]), .B(vdd_), .G(vdd_cntl_l[97]),
     .S(vdd_));
pch_hvt  M3_96_ ( .D(r_gnd_l[96]), .B(vdd_), .G(vdd_cntl_l[96]),
     .S(vdd_));
pch_hvt  M3_95_ ( .D(r_gnd_l[95]), .B(vdd_), .G(vdd_cntl_l[95]),
     .S(vdd_));
pch_hvt  M3_94_ ( .D(r_gnd_l[94]), .B(vdd_), .G(vdd_cntl_l[94]),
     .S(vdd_));
pch_hvt  M3_93_ ( .D(r_gnd_l[93]), .B(vdd_), .G(vdd_cntl_l[93]),
     .S(vdd_));
pch_hvt  M3_92_ ( .D(r_gnd_l[92]), .B(vdd_), .G(vdd_cntl_l[92]),
     .S(vdd_));
pch_hvt  M3_91_ ( .D(r_gnd_l[91]), .B(vdd_), .G(vdd_cntl_l[91]),
     .S(vdd_));
pch_hvt  M3_90_ ( .D(r_gnd_l[90]), .B(vdd_), .G(vdd_cntl_l[90]),
     .S(vdd_));
pch_hvt  M3_89_ ( .D(r_gnd_l[89]), .B(vdd_), .G(vdd_cntl_l[89]),
     .S(vdd_));
pch_hvt  M3_88_ ( .D(r_gnd_l[88]), .B(vdd_), .G(vdd_cntl_l[88]),
     .S(vdd_));
pch_hvt  M3_87_ ( .D(r_gnd_l[87]), .B(vdd_), .G(vdd_cntl_l[87]),
     .S(vdd_));
pch_hvt  M3_86_ ( .D(r_gnd_l[86]), .B(vdd_), .G(vdd_cntl_l[86]),
     .S(vdd_));
pch_hvt  M3_85_ ( .D(r_gnd_l[85]), .B(vdd_), .G(vdd_cntl_l[85]),
     .S(vdd_));
pch_hvt  M3_84_ ( .D(r_gnd_l[84]), .B(vdd_), .G(vdd_cntl_l[84]),
     .S(vdd_));
pch_hvt  M3_83_ ( .D(r_gnd_l[83]), .B(vdd_), .G(vdd_cntl_l[83]),
     .S(vdd_));
pch_hvt  M3_82_ ( .D(r_gnd_l[82]), .B(vdd_), .G(vdd_cntl_l[82]),
     .S(vdd_));
pch_hvt  M3_81_ ( .D(r_gnd_l[81]), .B(vdd_), .G(vdd_cntl_l[81]),
     .S(vdd_));
pch_hvt  M3_80_ ( .D(r_gnd_l[80]), .B(vdd_), .G(vdd_cntl_l[80]),
     .S(vdd_));
pch_hvt  M3_79_ ( .D(r_gnd_l[79]), .B(vdd_), .G(vdd_cntl_l[79]),
     .S(vdd_));
pch_hvt  M3_78_ ( .D(r_gnd_l[78]), .B(vdd_), .G(vdd_cntl_l[78]),
     .S(vdd_));
pch_hvt  M3_77_ ( .D(r_gnd_l[77]), .B(vdd_), .G(vdd_cntl_l[77]),
     .S(vdd_));
pch_hvt  M3_76_ ( .D(r_gnd_l[76]), .B(vdd_), .G(vdd_cntl_l[76]),
     .S(vdd_));
pch_hvt  M3_75_ ( .D(r_gnd_l[75]), .B(vdd_), .G(vdd_cntl_l[75]),
     .S(vdd_));
pch_hvt  M3_74_ ( .D(r_gnd_l[74]), .B(vdd_), .G(vdd_cntl_l[74]),
     .S(vdd_));
pch_hvt  M3_73_ ( .D(r_gnd_l[73]), .B(vdd_), .G(vdd_cntl_l[73]),
     .S(vdd_));
pch_hvt  M3_72_ ( .D(r_gnd_l[72]), .B(vdd_), .G(vdd_cntl_l[72]),
     .S(vdd_));
pch_hvt  M3_71_ ( .D(r_gnd_l[71]), .B(vdd_), .G(vdd_cntl_l[71]),
     .S(vdd_));
pch_hvt  M3_70_ ( .D(r_gnd_l[70]), .B(vdd_), .G(vdd_cntl_l[70]),
     .S(vdd_));
pch_hvt  M3_69_ ( .D(r_gnd_l[69]), .B(vdd_), .G(vdd_cntl_l[69]),
     .S(vdd_));
pch_hvt  M3_68_ ( .D(r_gnd_l[68]), .B(vdd_), .G(vdd_cntl_l[68]),
     .S(vdd_));
pch_hvt  M3_67_ ( .D(r_gnd_l[67]), .B(vdd_), .G(vdd_cntl_l[67]),
     .S(vdd_));
pch_hvt  M3_66_ ( .D(r_gnd_l[66]), .B(vdd_), .G(vdd_cntl_l[66]),
     .S(vdd_));
pch_hvt  M3_65_ ( .D(r_gnd_l[65]), .B(vdd_), .G(vdd_cntl_l[65]),
     .S(vdd_));
pch_hvt  M3_64_ ( .D(r_gnd_l[64]), .B(vdd_), .G(vdd_cntl_l[64]),
     .S(vdd_));
pch_hvt  M3_63_ ( .D(r_gnd_l[63]), .B(vdd_), .G(vdd_cntl_l[63]),
     .S(vdd_));
pch_hvt  M3_62_ ( .D(r_gnd_l[62]), .B(vdd_), .G(vdd_cntl_l[62]),
     .S(vdd_));
pch_hvt  M3_61_ ( .D(r_gnd_l[61]), .B(vdd_), .G(vdd_cntl_l[61]),
     .S(vdd_));
pch_hvt  M3_60_ ( .D(r_gnd_l[60]), .B(vdd_), .G(vdd_cntl_l[60]),
     .S(vdd_));
pch_hvt  M3_59_ ( .D(r_gnd_l[59]), .B(vdd_), .G(vdd_cntl_l[59]),
     .S(vdd_));
pch_hvt  M3_58_ ( .D(r_gnd_l[58]), .B(vdd_), .G(vdd_cntl_l[58]),
     .S(vdd_));
pch_hvt  M3_57_ ( .D(r_gnd_l[57]), .B(vdd_), .G(vdd_cntl_l[57]),
     .S(vdd_));
pch_hvt  M3_56_ ( .D(r_gnd_l[56]), .B(vdd_), .G(vdd_cntl_l[56]),
     .S(vdd_));
pch_hvt  M3_55_ ( .D(r_gnd_l[55]), .B(vdd_), .G(vdd_cntl_l[55]),
     .S(vdd_));
pch_hvt  M3_54_ ( .D(r_gnd_l[54]), .B(vdd_), .G(vdd_cntl_l[54]),
     .S(vdd_));
pch_hvt  M3_53_ ( .D(r_gnd_l[53]), .B(vdd_), .G(vdd_cntl_l[53]),
     .S(vdd_));
pch_hvt  M3_52_ ( .D(r_gnd_l[52]), .B(vdd_), .G(vdd_cntl_l[52]),
     .S(vdd_));
pch_hvt  M3_51_ ( .D(r_gnd_l[51]), .B(vdd_), .G(vdd_cntl_l[51]),
     .S(vdd_));
pch_hvt  M3_50_ ( .D(r_gnd_l[50]), .B(vdd_), .G(vdd_cntl_l[50]),
     .S(vdd_));
pch_hvt  M3_49_ ( .D(r_gnd_l[49]), .B(vdd_), .G(vdd_cntl_l[49]),
     .S(vdd_));
pch_hvt  M3_48_ ( .D(r_gnd_l[48]), .B(vdd_), .G(vdd_cntl_l[48]),
     .S(vdd_));
pch_hvt  M3_47_ ( .D(r_gnd_l[47]), .B(vdd_), .G(vdd_cntl_l[47]),
     .S(vdd_));
pch_hvt  M3_46_ ( .D(r_gnd_l[46]), .B(vdd_), .G(vdd_cntl_l[46]),
     .S(vdd_));
pch_hvt  M3_45_ ( .D(r_gnd_l[45]), .B(vdd_), .G(vdd_cntl_l[45]),
     .S(vdd_));
pch_hvt  M3_44_ ( .D(r_gnd_l[44]), .B(vdd_), .G(vdd_cntl_l[44]),
     .S(vdd_));
pch_hvt  M3_43_ ( .D(r_gnd_l[43]), .B(vdd_), .G(vdd_cntl_l[43]),
     .S(vdd_));
pch_hvt  M3_42_ ( .D(r_gnd_l[42]), .B(vdd_), .G(vdd_cntl_l[42]),
     .S(vdd_));
pch_hvt  M3_41_ ( .D(r_gnd_l[41]), .B(vdd_), .G(vdd_cntl_l[41]),
     .S(vdd_));
pch_hvt  M3_40_ ( .D(r_gnd_l[40]), .B(vdd_), .G(vdd_cntl_l[40]),
     .S(vdd_));
pch_hvt  M3_39_ ( .D(r_gnd_l[39]), .B(vdd_), .G(vdd_cntl_l[39]),
     .S(vdd_));
pch_hvt  M3_38_ ( .D(r_gnd_l[38]), .B(vdd_), .G(vdd_cntl_l[38]),
     .S(vdd_));
pch_hvt  M3_37_ ( .D(r_gnd_l[37]), .B(vdd_), .G(vdd_cntl_l[37]),
     .S(vdd_));
pch_hvt  M3_36_ ( .D(r_gnd_l[36]), .B(vdd_), .G(vdd_cntl_l[36]),
     .S(vdd_));
pch_hvt  M3_35_ ( .D(r_gnd_l[35]), .B(vdd_), .G(vdd_cntl_l[35]),
     .S(vdd_));
pch_hvt  M3_34_ ( .D(r_gnd_l[34]), .B(vdd_), .G(vdd_cntl_l[34]),
     .S(vdd_));
pch_hvt  M3_33_ ( .D(r_gnd_l[33]), .B(vdd_), .G(vdd_cntl_l[33]),
     .S(vdd_));
pch_hvt  M3_32_ ( .D(r_gnd_l[32]), .B(vdd_), .G(vdd_cntl_l[32]),
     .S(vdd_));
pch_hvt  M3_31_ ( .D(r_gnd_l[31]), .B(vdd_), .G(vdd_cntl_l[31]),
     .S(vdd_));
pch_hvt  M3_30_ ( .D(r_gnd_l[30]), .B(vdd_), .G(vdd_cntl_l[30]),
     .S(vdd_));
pch_hvt  M3_29_ ( .D(r_gnd_l[29]), .B(vdd_), .G(vdd_cntl_l[29]),
     .S(vdd_));
pch_hvt  M3_28_ ( .D(r_gnd_l[28]), .B(vdd_), .G(vdd_cntl_l[28]),
     .S(vdd_));
pch_hvt  M3_27_ ( .D(r_gnd_l[27]), .B(vdd_), .G(vdd_cntl_l[27]),
     .S(vdd_));
pch_hvt  M3_26_ ( .D(r_gnd_l[26]), .B(vdd_), .G(vdd_cntl_l[26]),
     .S(vdd_));
pch_hvt  M3_25_ ( .D(r_gnd_l[25]), .B(vdd_), .G(vdd_cntl_l[25]),
     .S(vdd_));
pch_hvt  M3_24_ ( .D(r_gnd_l[24]), .B(vdd_), .G(vdd_cntl_l[24]),
     .S(vdd_));
pch_hvt  M3_23_ ( .D(r_gnd_l[23]), .B(vdd_), .G(vdd_cntl_l[23]),
     .S(vdd_));
pch_hvt  M3_22_ ( .D(r_gnd_l[22]), .B(vdd_), .G(vdd_cntl_l[22]),
     .S(vdd_));
pch_hvt  M3_21_ ( .D(r_gnd_l[21]), .B(vdd_), .G(vdd_cntl_l[21]),
     .S(vdd_));
pch_hvt  M3_20_ ( .D(r_gnd_l[20]), .B(vdd_), .G(vdd_cntl_l[20]),
     .S(vdd_));
pch_hvt  M3_19_ ( .D(r_gnd_l[19]), .B(vdd_), .G(vdd_cntl_l[19]),
     .S(vdd_));
pch_hvt  M3_18_ ( .D(r_gnd_l[18]), .B(vdd_), .G(vdd_cntl_l[18]),
     .S(vdd_));
pch_hvt  M3_17_ ( .D(r_gnd_l[17]), .B(vdd_), .G(vdd_cntl_l[17]),
     .S(vdd_));
pch_hvt  M3_16_ ( .D(r_gnd_l[16]), .B(vdd_), .G(vdd_cntl_l[16]),
     .S(vdd_));
pch_hvt  M3_15_ ( .D(r_gnd_l[15]), .B(vdd_), .G(vdd_cntl_l[15]),
     .S(vdd_));
pch_hvt  M3_14_ ( .D(r_gnd_l[14]), .B(vdd_), .G(vdd_cntl_l[14]),
     .S(vdd_));
pch_hvt  M3_13_ ( .D(r_gnd_l[13]), .B(vdd_), .G(vdd_cntl_l[13]),
     .S(vdd_));
pch_hvt  M3_12_ ( .D(r_gnd_l[12]), .B(vdd_), .G(vdd_cntl_l[12]),
     .S(vdd_));
pch_hvt  M3_11_ ( .D(r_gnd_l[11]), .B(vdd_), .G(vdd_cntl_l[11]),
     .S(vdd_));
pch_hvt  M3_10_ ( .D(r_gnd_l[10]), .B(vdd_), .G(vdd_cntl_l[10]),
     .S(vdd_));
pch_hvt  M3_9_ ( .D(r_gnd_l[9]), .B(vdd_), .G(vdd_cntl_l[9]),
     .S(vdd_));
pch_hvt  M3_8_ ( .D(r_gnd_l[8]), .B(vdd_), .G(vdd_cntl_l[8]),
     .S(vdd_));
pch_hvt  M3_7_ ( .D(r_gnd_l[7]), .B(vdd_), .G(vdd_cntl_l[7]),
     .S(vdd_));
pch_hvt  M3_6_ ( .D(r_gnd_l[6]), .B(vdd_), .G(vdd_cntl_l[6]),
     .S(vdd_));
pch_hvt  M3_5_ ( .D(r_gnd_l[5]), .B(vdd_), .G(vdd_cntl_l[5]),
     .S(vdd_));
pch_hvt  M3_4_ ( .D(r_gnd_l[4]), .B(vdd_), .G(vdd_cntl_l[4]),
     .S(vdd_));
pch_hvt  M3_3_ ( .D(r_gnd_l[3]), .B(vdd_), .G(vdd_cntl_l[3]),
     .S(vdd_));
pch_hvt  M3_2_ ( .D(r_gnd_l[2]), .B(vdd_), .G(vdd_cntl_l[2]),
     .S(vdd_));
pch_hvt  M3_1_ ( .D(r_gnd_l[1]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  M3_0_ ( .D(r_gnd_l[0]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));
cram_2x2x2_ice8p I_mem2x2x2t_70_ ( .wl_r(wl_r[141:140]),
     .wl_l(wl_l[141:140]), .reset_r(reset_r[141:140]),
     .reset_l(reset_l[141:140]), .pgate_r(pgate_r[141:140]),
     .pgate_l(pgate_l[141:140]), .q_b(net35[0:7]), .q(net36[0:7]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[141:140]),
     .r_gnd_r(r_gnd_r[141:140]));
cram_2x2x2_ice8p I_mem2x2x2t_69_ ( .wl_r(wl_r[139:138]),
     .wl_l(wl_l[139:138]), .reset_r(reset_r[139:138]),
     .reset_l(reset_l[139:138]), .pgate_r(pgate_r[139:138]),
     .pgate_l(pgate_l[139:138]), .q_b(net35[8:15]), .q(net36[8:15]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[139:138]),
     .r_gnd_r(r_gnd_r[139:138]));
cram_2x2x2_ice8p I_mem2x2x2t_68_ ( .wl_r(wl_r[137:136]),
     .wl_l(wl_l[137:136]), .reset_r(reset_r[137:136]),
     .reset_l(reset_l[137:136]), .pgate_r(pgate_r[137:136]),
     .pgate_l(pgate_l[137:136]), .q_b(net35[16:23]), .q(net36[16:23]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[137:136]),
     .r_gnd_r(r_gnd_r[137:136]));
cram_2x2x2_ice8p I_mem2x2x2t_67_ ( .wl_r(wl_r[135:134]),
     .wl_l(wl_l[135:134]), .reset_r(reset_r[135:134]),
     .reset_l(reset_l[135:134]), .pgate_r(pgate_r[135:134]),
     .pgate_l(pgate_l[135:134]), .q_b(net35[24:31]), .q(net36[24:31]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[135:134]),
     .r_gnd_r(r_gnd_r[135:134]));
cram_2x2x2_ice8p I_mem2x2x2t_66_ ( .wl_r(wl_r[133:132]),
     .wl_l(wl_l[133:132]), .reset_r(reset_r[133:132]),
     .reset_l(reset_l[133:132]), .pgate_r(pgate_r[133:132]),
     .pgate_l(pgate_l[133:132]), .q_b(net35[32:39]), .q(net36[32:39]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[133:132]),
     .r_gnd_r(r_gnd_r[133:132]));
cram_2x2x2_ice8p I_mem2x2x2t_65_ ( .wl_r(wl_r[131:130]),
     .wl_l(wl_l[131:130]), .reset_r(reset_r[131:130]),
     .reset_l(reset_l[131:130]), .pgate_r(pgate_r[131:130]),
     .pgate_l(pgate_l[131:130]), .q_b(net35[40:47]), .q(net36[40:47]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[131:130]),
     .r_gnd_r(r_gnd_r[131:130]));
cram_2x2x2_ice8p I_mem2x2x2t_64_ ( .wl_r(wl_r[129:128]),
     .wl_l(wl_l[129:128]), .reset_r(reset_r[129:128]),
     .reset_l(reset_l[129:128]), .pgate_r(pgate_r[129:128]),
     .pgate_l(pgate_l[129:128]), .q_b(net35[48:55]), .q(net36[48:55]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[129:128]),
     .r_gnd_r(r_gnd_r[129:128]));
cram_2x2x2_ice8p I_mem2x2x2t_63_ ( .wl_r(wl_r[127:126]),
     .wl_l(wl_l[127:126]), .reset_r(reset_r[127:126]),
     .reset_l(reset_l[127:126]), .pgate_r(pgate_r[127:126]),
     .pgate_l(pgate_l[127:126]), .q_b(net35[56:63]), .q(net36[56:63]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[127:126]),
     .r_gnd_r(r_gnd_r[127:126]));
cram_2x2x2_ice8p I_mem2x2x2t_62_ ( .wl_r(wl_r[125:124]),
     .wl_l(wl_l[125:124]), .reset_r(reset_r[125:124]),
     .reset_l(reset_l[125:124]), .pgate_r(pgate_r[125:124]),
     .pgate_l(pgate_l[125:124]), .q_b(net35[64:71]), .q(net36[64:71]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[125:124]),
     .r_gnd_r(r_gnd_r[125:124]));
cram_2x2x2_ice8p I_mem2x2x2t_61_ ( .wl_r(wl_r[123:122]),
     .wl_l(wl_l[123:122]), .reset_r(reset_r[123:122]),
     .reset_l(reset_l[123:122]), .pgate_r(pgate_r[123:122]),
     .pgate_l(pgate_l[123:122]), .q_b(net35[72:79]), .q(net36[72:79]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[123:122]),
     .r_gnd_r(r_gnd_r[123:122]));
cram_2x2x2_ice8p I_mem2x2x2t_60_ ( .wl_r(wl_r[121:120]),
     .wl_l(wl_l[121:120]), .reset_r(reset_r[121:120]),
     .reset_l(reset_l[121:120]), .pgate_r(pgate_r[121:120]),
     .pgate_l(pgate_l[121:120]), .q_b(net35[80:87]), .q(net36[80:87]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[121:120]),
     .r_gnd_r(r_gnd_r[121:120]));
cram_2x2x2_ice8p I_mem2x2x2t_59_ ( .wl_r(wl_r[119:118]),
     .wl_l(wl_l[119:118]), .reset_r(reset_r[119:118]),
     .reset_l(reset_l[119:118]), .pgate_r(pgate_r[119:118]),
     .pgate_l(pgate_l[119:118]), .q_b(net35[88:95]), .q(net36[88:95]),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[119:118]),
     .r_gnd_r(r_gnd_r[119:118]));
cram_2x2x2_ice8p I_mem2x2x2t_58_ ( .wl_r(wl_r[117:116]),
     .wl_l(wl_l[117:116]), .reset_r(reset_r[117:116]),
     .reset_l(reset_l[117:116]), .pgate_r(pgate_r[117:116]),
     .pgate_l(pgate_l[117:116]), .q_b(net35[96:103]),
     .q(net36[96:103]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[117:116]),
     .r_gnd_r(r_gnd_r[117:116]));
cram_2x2x2_ice8p I_mem2x2x2t_57_ ( .wl_r(wl_r[115:114]),
     .wl_l(wl_l[115:114]), .reset_r(reset_r[115:114]),
     .reset_l(reset_l[115:114]), .pgate_r(pgate_r[115:114]),
     .pgate_l(pgate_l[115:114]), .q_b(net35[104:111]),
     .q(net36[104:111]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[115:114]),
     .r_gnd_r(r_gnd_r[115:114]));
cram_2x2x2_ice8p I_mem2x2x2t_56_ ( .wl_r(wl_r[113:112]),
     .wl_l(wl_l[113:112]), .reset_r(reset_r[113:112]),
     .reset_l(reset_l[113:112]), .pgate_r(pgate_r[113:112]),
     .pgate_l(pgate_l[113:112]), .q_b(net35[112:119]),
     .q(net36[112:119]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[113:112]),
     .r_gnd_r(r_gnd_r[113:112]));
cram_2x2x2_ice8p I_mem2x2x2t_55_ ( .wl_r(wl_r[111:110]),
     .wl_l(wl_l[111:110]), .reset_r(reset_r[111:110]),
     .reset_l(reset_l[111:110]), .pgate_r(pgate_r[111:110]),
     .pgate_l(pgate_l[111:110]), .q_b(net35[120:127]),
     .q(net36[120:127]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[111:110]),
     .r_gnd_r(r_gnd_r[111:110]));
cram_2x2x2_ice8p I_mem2x2x2t_54_ ( .wl_r(wl_r[109:108]),
     .wl_l(wl_l[109:108]), .reset_r(reset_r[109:108]),
     .reset_l(reset_l[109:108]), .pgate_r(pgate_r[109:108]),
     .pgate_l(pgate_l[109:108]), .q_b(net35[128:135]),
     .q(net36[128:135]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[109:108]),
     .r_gnd_r(r_gnd_r[109:108]));
cram_2x2x2_ice8p I_mem2x2x2t_53_ ( .wl_r(wl_r[107:106]),
     .wl_l(wl_l[107:106]), .reset_r(reset_r[107:106]),
     .reset_l(reset_l[107:106]), .pgate_r(pgate_r[107:106]),
     .pgate_l(pgate_l[107:106]), .q_b(net35[136:143]),
     .q(net36[136:143]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[107:106]),
     .r_gnd_r(r_gnd_r[107:106]));
cram_2x2x2_ice8p I_mem2x2x2t_52_ ( .wl_r(wl_r[105:104]),
     .wl_l(wl_l[105:104]), .reset_r(reset_r[105:104]),
     .reset_l(reset_l[105:104]), .pgate_r(pgate_r[105:104]),
     .pgate_l(pgate_l[105:104]), .q_b(net35[144:151]),
     .q(net36[144:151]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[105:104]),
     .r_gnd_r(r_gnd_r[105:104]));
cram_2x2x2_ice8p I_mem2x2x2t_51_ ( .wl_r(wl_r[103:102]),
     .wl_l(wl_l[103:102]), .reset_r(reset_r[103:102]),
     .reset_l(reset_l[103:102]), .pgate_r(pgate_r[103:102]),
     .pgate_l(pgate_l[103:102]), .q_b(net35[152:159]),
     .q(net36[152:159]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[103:102]),
     .r_gnd_r(r_gnd_r[103:102]));
cram_2x2x2_ice8p I_mem2x2x2t_50_ ( .wl_r(wl_r[101:100]),
     .wl_l(wl_l[101:100]), .reset_r(reset_r[101:100]),
     .reset_l(reset_l[101:100]), .pgate_r(pgate_r[101:100]),
     .pgate_l(pgate_l[101:100]), .q_b(net35[160:167]),
     .q(net36[160:167]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[101:100]),
     .r_gnd_r(r_gnd_r[101:100]));
cram_2x2x2_ice8p I_mem2x2x2t_49_ ( .wl_r(wl_r[99:98]),
     .wl_l(wl_l[99:98]), .reset_r(reset_r[99:98]),
     .reset_l(reset_l[99:98]), .pgate_r(pgate_r[99:98]),
     .pgate_l(pgate_l[99:98]), .q_b(net35[168:175]),
     .q(net36[168:175]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[99:98]),
     .r_gnd_r(r_gnd_r[99:98]));
cram_2x2x2_ice8p I_mem2x2x2t_48_ ( .wl_r(wl_r[97:96]),
     .wl_l(wl_l[97:96]), .reset_r(reset_r[97:96]),
     .reset_l(reset_l[97:96]), .pgate_r(pgate_r[97:96]),
     .pgate_l(pgate_l[97:96]), .q_b(net35[176:183]),
     .q(net36[176:183]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[97:96]),
     .r_gnd_r(r_gnd_r[97:96]));
cram_2x2x2_ice8p I_mem2x2x2t_47_ ( .wl_r(wl_r[95:94]),
     .wl_l(wl_l[95:94]), .reset_r(reset_r[95:94]),
     .reset_l(reset_l[95:94]), .pgate_r(pgate_r[95:94]),
     .pgate_l(pgate_l[95:94]), .q_b(net35[184:191]),
     .q(net36[184:191]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[95:94]),
     .r_gnd_r(r_gnd_r[95:94]));
cram_2x2x2_ice8p I_mem2x2x2t_46_ ( .wl_r(wl_r[93:92]),
     .wl_l(wl_l[93:92]), .reset_r(reset_r[93:92]),
     .reset_l(reset_l[93:92]), .pgate_r(pgate_r[93:92]),
     .pgate_l(pgate_l[93:92]), .q_b(net35[192:199]),
     .q(net36[192:199]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[93:92]),
     .r_gnd_r(r_gnd_r[93:92]));
cram_2x2x2_ice8p I_mem2x2x2t_45_ ( .wl_r(wl_r[91:90]),
     .wl_l(wl_l[91:90]), .reset_r(reset_r[91:90]),
     .reset_l(reset_l[91:90]), .pgate_r(pgate_r[91:90]),
     .pgate_l(pgate_l[91:90]), .q_b(net35[200:207]),
     .q(net36[200:207]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[91:90]),
     .r_gnd_r(r_gnd_r[91:90]));
cram_2x2x2_ice8p I_mem2x2x2t_44_ ( .wl_r(wl_r[89:88]),
     .wl_l(wl_l[89:88]), .reset_r(reset_r[89:88]),
     .reset_l(reset_l[89:88]), .pgate_r(pgate_r[89:88]),
     .pgate_l(pgate_l[89:88]), .q_b(net35[208:215]),
     .q(net36[208:215]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[89:88]),
     .r_gnd_r(r_gnd_r[89:88]));
cram_2x2x2_ice8p I_mem2x2x2t_43_ ( .wl_r(wl_r[87:86]),
     .wl_l(wl_l[87:86]), .reset_r(reset_r[87:86]),
     .reset_l(reset_l[87:86]), .pgate_r(pgate_r[87:86]),
     .pgate_l(pgate_l[87:86]), .q_b(net35[216:223]),
     .q(net36[216:223]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[87:86]),
     .r_gnd_r(r_gnd_r[87:86]));
cram_2x2x2_ice8p I_mem2x2x2t_42_ ( .wl_r(wl_r[85:84]),
     .wl_l(wl_l[85:84]), .reset_r(reset_r[85:84]),
     .reset_l(reset_l[85:84]), .pgate_r(pgate_r[85:84]),
     .pgate_l(pgate_l[85:84]), .q_b(net35[224:231]),
     .q(net36[224:231]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[85:84]),
     .r_gnd_r(r_gnd_r[85:84]));
cram_2x2x2_ice8p I_mem2x2x2t_41_ ( .wl_r(wl_r[83:82]),
     .wl_l(wl_l[83:82]), .reset_r(reset_r[83:82]),
     .reset_l(reset_l[83:82]), .pgate_r(pgate_r[83:82]),
     .pgate_l(pgate_l[83:82]), .q_b(net35[232:239]),
     .q(net36[232:239]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[83:82]),
     .r_gnd_r(r_gnd_r[83:82]));
cram_2x2x2_ice8p I_mem2x2x2t_40_ ( .wl_r(wl_r[81:80]),
     .wl_l(wl_l[81:80]), .reset_r(reset_r[81:80]),
     .reset_l(reset_l[81:80]), .pgate_r(pgate_r[81:80]),
     .pgate_l(pgate_l[81:80]), .q_b(net35[240:247]),
     .q(net36[240:247]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[81:80]),
     .r_gnd_r(r_gnd_r[81:80]));
cram_2x2x2_ice8p I_mem2x2x2t_39_ ( .wl_r(wl_r[79:78]),
     .wl_l(wl_l[79:78]), .reset_r(reset_r[79:78]),
     .reset_l(reset_l[79:78]), .pgate_r(pgate_r[79:78]),
     .pgate_l(pgate_l[79:78]), .q_b(net35[248:255]),
     .q(net36[248:255]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[79:78]),
     .r_gnd_r(r_gnd_r[79:78]));
cram_2x2x2_ice8p I_mem2x2x2t_38_ ( .wl_r(wl_r[77:76]),
     .wl_l(wl_l[77:76]), .reset_r(reset_r[77:76]),
     .reset_l(reset_l[77:76]), .pgate_r(pgate_r[77:76]),
     .pgate_l(pgate_l[77:76]), .q_b(net35[256:263]),
     .q(net36[256:263]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[77:76]),
     .r_gnd_r(r_gnd_r[77:76]));
cram_2x2x2_ice8p I_mem2x2x2t_37_ ( .wl_r(wl_r[75:74]),
     .wl_l(wl_l[75:74]), .reset_r(reset_r[75:74]),
     .reset_l(reset_l[75:74]), .pgate_r(pgate_r[75:74]),
     .pgate_l(pgate_l[75:74]), .q_b(net35[264:271]),
     .q(net36[264:271]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[75:74]),
     .r_gnd_r(r_gnd_r[75:74]));
cram_2x2x2_ice8p I_mem2x2x2t_36_ ( .wl_r(wl_r[73:72]),
     .wl_l(wl_l[73:72]), .reset_r(reset_r[73:72]),
     .reset_l(reset_l[73:72]), .pgate_r(pgate_r[73:72]),
     .pgate_l(pgate_l[73:72]), .q_b(net35[272:279]),
     .q(net36[272:279]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[73:72]),
     .r_gnd_r(r_gnd_r[73:72]));
cram_2x2x2_ice8p I_mem2x2x2t_35_ ( .wl_r(wl_r[71:70]),
     .wl_l(wl_l[71:70]), .reset_r(reset_r[71:70]),
     .reset_l(reset_l[71:70]), .pgate_r(pgate_r[71:70]),
     .pgate_l(pgate_l[71:70]), .q_b(net35[280:287]),
     .q(net36[280:287]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[71:70]),
     .r_gnd_r(r_gnd_r[71:70]));
cram_2x2x2_ice8p I_mem2x2x2t_34_ ( .wl_r(wl_r[69:68]),
     .wl_l(wl_l[69:68]), .reset_r(reset_r[69:68]),
     .reset_l(reset_l[69:68]), .pgate_r(pgate_r[69:68]),
     .pgate_l(pgate_l[69:68]), .q_b(net35[288:295]),
     .q(net36[288:295]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[69:68]),
     .r_gnd_r(r_gnd_r[69:68]));
cram_2x2x2_ice8p I_mem2x2x2t_33_ ( .wl_r(wl_r[67:66]),
     .wl_l(wl_l[67:66]), .reset_r(reset_r[67:66]),
     .reset_l(reset_l[67:66]), .pgate_r(pgate_r[67:66]),
     .pgate_l(pgate_l[67:66]), .q_b(net35[296:303]),
     .q(net36[296:303]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[67:66]),
     .r_gnd_r(r_gnd_r[67:66]));
cram_2x2x2_ice8p I_mem2x2x2t_32_ ( .wl_r(wl_r[65:64]),
     .wl_l(wl_l[65:64]), .reset_r(reset_r[65:64]),
     .reset_l(reset_l[65:64]), .pgate_r(pgate_r[65:64]),
     .pgate_l(pgate_l[65:64]), .q_b(net35[304:311]),
     .q(net36[304:311]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[65:64]),
     .r_gnd_r(r_gnd_r[65:64]));
cram_2x2x2_ice8p I_mem2x2x2t_31_ ( .wl_r(wl_r[63:62]),
     .wl_l(wl_l[63:62]), .reset_r(reset_r[63:62]),
     .reset_l(reset_l[63:62]), .pgate_r(pgate_r[63:62]),
     .pgate_l(pgate_l[63:62]), .q_b(net35[312:319]),
     .q(net36[312:319]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[63:62]),
     .r_gnd_r(r_gnd_r[63:62]));
cram_2x2x2_ice8p I_mem2x2x2t_30_ ( .wl_r(wl_r[61:60]),
     .wl_l(wl_l[61:60]), .reset_r(reset_r[61:60]),
     .reset_l(reset_l[61:60]), .pgate_r(pgate_r[61:60]),
     .pgate_l(pgate_l[61:60]), .q_b(net35[320:327]),
     .q(net36[320:327]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[61:60]),
     .r_gnd_r(r_gnd_r[61:60]));
cram_2x2x2_ice8p I_mem2x2x2t_29_ ( .wl_r(wl_r[59:58]),
     .wl_l(wl_l[59:58]), .reset_r(reset_r[59:58]),
     .reset_l(reset_l[59:58]), .pgate_r(pgate_r[59:58]),
     .pgate_l(pgate_l[59:58]), .q_b(net35[328:335]),
     .q(net36[328:335]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[59:58]),
     .r_gnd_r(r_gnd_r[59:58]));
cram_2x2x2_ice8p I_mem2x2x2t_28_ ( .wl_r(wl_r[57:56]),
     .wl_l(wl_l[57:56]), .reset_r(reset_r[57:56]),
     .reset_l(reset_l[57:56]), .pgate_r(pgate_r[57:56]),
     .pgate_l(pgate_l[57:56]), .q_b(net35[336:343]),
     .q(net36[336:343]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[57:56]),
     .r_gnd_r(r_gnd_r[57:56]));
cram_2x2x2_ice8p I_mem2x2x2t_27_ ( .wl_r(wl_r[55:54]),
     .wl_l(wl_l[55:54]), .reset_r(reset_r[55:54]),
     .reset_l(reset_l[55:54]), .pgate_r(pgate_r[55:54]),
     .pgate_l(pgate_l[55:54]), .q_b(net35[344:351]),
     .q(net36[344:351]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[55:54]),
     .r_gnd_r(r_gnd_r[55:54]));
cram_2x2x2_ice8p I_mem2x2x2t_26_ ( .wl_r(wl_r[53:52]),
     .wl_l(wl_l[53:52]), .reset_r(reset_r[53:52]),
     .reset_l(reset_l[53:52]), .pgate_r(pgate_r[53:52]),
     .pgate_l(pgate_l[53:52]), .q_b(net35[352:359]),
     .q(net36[352:359]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[53:52]),
     .r_gnd_r(r_gnd_r[53:52]));
cram_2x2x2_ice8p I_mem2x2x2t_25_ ( .wl_r(wl_r[51:50]),
     .wl_l(wl_l[51:50]), .reset_r(reset_r[51:50]),
     .reset_l(reset_l[51:50]), .pgate_r(pgate_r[51:50]),
     .pgate_l(pgate_l[51:50]), .q_b(net35[360:367]),
     .q(net36[360:367]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[51:50]),
     .r_gnd_r(r_gnd_r[51:50]));
cram_2x2x2_ice8p I_mem2x2x2t_24_ ( .wl_r(wl_r[49:48]),
     .wl_l(wl_l[49:48]), .reset_r(reset_r[49:48]),
     .reset_l(reset_l[49:48]), .pgate_r(pgate_r[49:48]),
     .pgate_l(pgate_l[49:48]), .q_b(net35[368:375]),
     .q(net36[368:375]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[49:48]),
     .r_gnd_r(r_gnd_r[49:48]));
cram_2x2x2_ice8p I_mem2x2x2t_23_ ( .wl_r(wl_r[47:46]),
     .wl_l(wl_l[47:46]), .reset_r(reset_r[47:46]),
     .reset_l(reset_l[47:46]), .pgate_r(pgate_r[47:46]),
     .pgate_l(pgate_l[47:46]), .q_b(net35[376:383]),
     .q(net36[376:383]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[47:46]),
     .r_gnd_r(r_gnd_r[47:46]));
cram_2x2x2_ice8p I_mem2x2x2t_22_ ( .wl_r(wl_r[45:44]),
     .wl_l(wl_l[45:44]), .reset_r(reset_r[45:44]),
     .reset_l(reset_l[45:44]), .pgate_r(pgate_r[45:44]),
     .pgate_l(pgate_l[45:44]), .q_b(net35[384:391]),
     .q(net36[384:391]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[45:44]),
     .r_gnd_r(r_gnd_r[45:44]));
cram_2x2x2_ice8p I_mem2x2x2t_21_ ( .wl_r(wl_r[43:42]),
     .wl_l(wl_l[43:42]), .reset_r(reset_r[43:42]),
     .reset_l(reset_l[43:42]), .pgate_r(pgate_r[43:42]),
     .pgate_l(pgate_l[43:42]), .q_b(net35[392:399]),
     .q(net36[392:399]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[43:42]),
     .r_gnd_r(r_gnd_r[43:42]));
cram_2x2x2_ice8p I_mem2x2x2t_20_ ( .wl_r(wl_r[41:40]),
     .wl_l(wl_l[41:40]), .reset_r(reset_r[41:40]),
     .reset_l(reset_l[41:40]), .pgate_r(pgate_r[41:40]),
     .pgate_l(pgate_l[41:40]), .q_b(net35[400:407]),
     .q(net36[400:407]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[41:40]),
     .r_gnd_r(r_gnd_r[41:40]));
cram_2x2x2_ice8p I_mem2x2x2t_19_ ( .wl_r(wl_r[39:38]),
     .wl_l(wl_l[39:38]), .reset_r(reset_r[39:38]),
     .reset_l(reset_l[39:38]), .pgate_r(pgate_r[39:38]),
     .pgate_l(pgate_l[39:38]), .q_b(net35[408:415]),
     .q(net36[408:415]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[39:38]),
     .r_gnd_r(r_gnd_r[39:38]));
cram_2x2x2_ice8p I_mem2x2x2t_18_ ( .wl_r(wl_r[37:36]),
     .wl_l(wl_l[37:36]), .reset_r(reset_r[37:36]),
     .reset_l(reset_l[37:36]), .pgate_r(pgate_r[37:36]),
     .pgate_l(pgate_l[37:36]), .q_b(net35[416:423]),
     .q(net36[416:423]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[37:36]),
     .r_gnd_r(r_gnd_r[37:36]));
cram_2x2x2_ice8p I_mem2x2x2t_17_ ( .wl_r(wl_r[35:34]),
     .wl_l(wl_l[35:34]), .reset_r(reset_r[35:34]),
     .reset_l(reset_l[35:34]), .pgate_r(pgate_r[35:34]),
     .pgate_l(pgate_l[35:34]), .q_b(net35[424:431]),
     .q(net36[424:431]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[35:34]),
     .r_gnd_r(r_gnd_r[35:34]));
cram_2x2x2_ice8p I_mem2x2x2t_16_ ( .wl_r(wl_r[33:32]),
     .wl_l(wl_l[33:32]), .reset_r(reset_r[33:32]),
     .reset_l(reset_l[33:32]), .pgate_r(pgate_r[33:32]),
     .pgate_l(pgate_l[33:32]), .q_b(net35[432:439]),
     .q(net36[432:439]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[33:32]),
     .r_gnd_r(r_gnd_r[33:32]));
cram_2x2x2_ice8p I_mem2x2x2t_15_ ( .wl_r(wl_r[31:30]),
     .wl_l(wl_l[31:30]), .reset_r(reset_r[31:30]),
     .reset_l(reset_l[31:30]), .pgate_r(pgate_r[31:30]),
     .pgate_l(pgate_l[31:30]), .q_b(net35[440:447]),
     .q(net36[440:447]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[31:30]),
     .r_gnd_r(r_gnd_r[31:30]));
cram_2x2x2_ice8p I_mem2x2x2t_14_ ( .wl_r(wl_r[29:28]),
     .wl_l(wl_l[29:28]), .reset_r(reset_r[29:28]),
     .reset_l(reset_l[29:28]), .pgate_r(pgate_r[29:28]),
     .pgate_l(pgate_l[29:28]), .q_b(net35[448:455]),
     .q(net36[448:455]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[29:28]),
     .r_gnd_r(r_gnd_r[29:28]));
cram_2x2x2_ice8p I_mem2x2x2t_13_ ( .wl_r(wl_r[27:26]),
     .wl_l(wl_l[27:26]), .reset_r(reset_r[27:26]),
     .reset_l(reset_l[27:26]), .pgate_r(pgate_r[27:26]),
     .pgate_l(pgate_l[27:26]), .q_b(net35[456:463]),
     .q(net36[456:463]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[27:26]),
     .r_gnd_r(r_gnd_r[27:26]));
cram_2x2x2_ice8p I_mem2x2x2t_12_ ( .wl_r(wl_r[25:24]),
     .wl_l(wl_l[25:24]), .reset_r(reset_r[25:24]),
     .reset_l(reset_l[25:24]), .pgate_r(pgate_r[25:24]),
     .pgate_l(pgate_l[25:24]), .q_b(net35[464:471]),
     .q(net36[464:471]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[25:24]),
     .r_gnd_r(r_gnd_r[25:24]));
cram_2x2x2_ice8p I_mem2x2x2t_11_ ( .wl_r(wl_r[23:22]),
     .wl_l(wl_l[23:22]), .reset_r(reset_r[23:22]),
     .reset_l(reset_l[23:22]), .pgate_r(pgate_r[23:22]),
     .pgate_l(pgate_l[23:22]), .q_b(net35[472:479]),
     .q(net36[472:479]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[23:22]),
     .r_gnd_r(r_gnd_r[23:22]));
cram_2x2x2_ice8p I_mem2x2x2t_10_ ( .wl_r(wl_r[21:20]),
     .wl_l(wl_l[21:20]), .reset_r(reset_r[21:20]),
     .reset_l(reset_l[21:20]), .pgate_r(pgate_r[21:20]),
     .pgate_l(pgate_l[21:20]), .q_b(net35[480:487]),
     .q(net36[480:487]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[21:20]),
     .r_gnd_r(r_gnd_r[21:20]));
cram_2x2x2_ice8p I_mem2x2x2t_9_ ( .wl_r(wl_r[19:18]),
     .wl_l(wl_l[19:18]), .reset_r(reset_r[19:18]),
     .reset_l(reset_l[19:18]), .pgate_r(pgate_r[19:18]),
     .pgate_l(pgate_l[19:18]), .q_b(net35[488:495]),
     .q(net36[488:495]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[19:18]),
     .r_gnd_r(r_gnd_r[19:18]));
cram_2x2x2_ice8p I_mem2x2x2t_8_ ( .wl_r(wl_r[17:16]),
     .wl_l(wl_l[17:16]), .reset_r(reset_r[17:16]),
     .reset_l(reset_l[17:16]), .pgate_r(pgate_r[17:16]),
     .pgate_l(pgate_l[17:16]), .q_b(net35[496:503]),
     .q(net36[496:503]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[17:16]),
     .r_gnd_r(r_gnd_r[17:16]));
cram_2x2x2_ice8p I_mem2x2x2t_7_ ( .wl_r(wl_r[15:14]),
     .wl_l(wl_l[15:14]), .reset_r(reset_r[15:14]),
     .reset_l(reset_l[15:14]), .pgate_r(pgate_r[15:14]),
     .pgate_l(pgate_l[15:14]), .q_b(net35[504:511]),
     .q(net36[504:511]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[15:14]),
     .r_gnd_r(r_gnd_r[15:14]));
cram_2x2x2_ice8p I_mem2x2x2t_6_ ( .wl_r(wl_r[13:12]),
     .wl_l(wl_l[13:12]), .reset_r(reset_r[13:12]),
     .reset_l(reset_l[13:12]), .pgate_r(pgate_r[13:12]),
     .pgate_l(pgate_l[13:12]), .q_b(net35[512:519]),
     .q(net36[512:519]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[13:12]),
     .r_gnd_r(r_gnd_r[13:12]));
cram_2x2x2_ice8p I_mem2x2x2t_5_ ( .wl_r(wl_r[11:10]),
     .wl_l(wl_l[11:10]), .reset_r(reset_r[11:10]),
     .reset_l(reset_l[11:10]), .pgate_r(pgate_r[11:10]),
     .pgate_l(pgate_l[11:10]), .q_b(net35[520:527]),
     .q(net36[520:527]), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[11:10]),
     .r_gnd_r(r_gnd_r[11:10]));
cram_2x2x2_ice8p I_mem2x2x2t_4_ ( .wl_r(wl_r[9:8]), .wl_l(wl_l[9:8]),
     .reset_r(reset_r[9:8]), .reset_l(reset_l[9:8]),
     .pgate_r(pgate_r[9:8]), .pgate_l(pgate_l[9:8]),
     .q_b(net35[528:535]), .q(net36[528:535]), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[9:8]), .r_gnd_r(r_gnd_r[9:8]));
cram_2x2x2_ice8p I_mem2x2x2t_3_ ( .wl_r(wl_r[7:6]), .wl_l(wl_l[7:6]),
     .reset_r(reset_r[7:6]), .reset_l(reset_l[7:6]),
     .pgate_r(pgate_r[7:6]), .pgate_l(pgate_l[7:6]),
     .q_b(net35[536:543]), .q(net36[536:543]), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[7:6]), .r_gnd_r(r_gnd_r[7:6]));
cram_2x2x2_ice8p I_mem2x2x2t_2_ ( .wl_r(wl_r[5:4]), .wl_l(wl_l[5:4]),
     .reset_r(reset_r[5:4]), .reset_l(reset_l[5:4]),
     .pgate_r(pgate_r[5:4]), .pgate_l(pgate_l[5:4]),
     .q_b(net35[544:551]), .q(net36[544:551]), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[5:4]), .r_gnd_r(r_gnd_r[5:4]));
cram_2x2x2_ice8p I_mem2x2x2t_1_ ( .wl_r(wl_r[3:2]), .wl_l(wl_l[3:2]),
     .reset_r(reset_r[3:2]), .reset_l(reset_l[3:2]),
     .pgate_r(pgate_r[3:2]), .pgate_l(pgate_l[3:2]),
     .q_b(net35[552:559]), .q(net36[552:559]), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[3:2]), .r_gnd_r(r_gnd_r[3:2]));
cram_2x2x2_ice8p I_mem2x2x2t_0_ ( .wl_r(wl_r[1:0]), .wl_l(wl_l[1:0]),
     .reset_r(reset_r[1:0]), .reset_l(reset_l[1:0]),
     .pgate_r(pgate_r[1:0]), .pgate_l(pgate_l[1:0]),
     .q_b(net35[560:567]), .q(net36[560:567]), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[1:0]), .r_gnd_r(r_gnd_r[1:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_clk_reg, View - schematic
// LAST TIME SAVED: Aug 30 17:59:46 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_pump_clk_reg ( clk_out_25, clk_in_25, pump_chrg_25,
     pump_on_25 );
output  clk_out_25;

input  clk_in_25, pump_chrg_25, pump_on_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I78 ( .G(GND_), .Pb(vddp_), .A(pump_chrg_25), .Y(clk_freeze),
     .P(vddp_), .B(pump_on_25), .Gb(GND_));
inv_25 I72 ( .IN(net020), .OUT(clk_equal), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(vddp_tieh), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
exor2_25 I85 ( .A(clk_in_25), .Y(net020), .B(clk_out_25));
vddp_tiehigh I117 ( .vddp_tieh(vddp_tieh));
ml_dlatch_25 I63 ( .D_25(clk_in_25), .EN_25(clk_go), .R_25(net34),
     .Q_25(clk_out_25));
ml_dlatch_25 I64 ( .D_25(vddp_tieh), .EN_25(clk_equal),
     .R_25(clk_freeze), .Q_25(clk_go));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_x2, View - schematic
// LAST TIME SAVED: Sep  1 14:53:51 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_pump_vpxa_x2 ( vpxa_int, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, pumpen_25, vpxa_clk_25, vpxa_clk_b_25 );
inout  vpxa_int;

input  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25, pumpen_25,
     vpxa_clk_25, vpxa_clk_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_pump_vpxa_buf I80 ( .in(net43), .out(clkin_2_25));
ml_pump_vpxa_buf I79 ( .in(net47), .out(net22));
ml_pump_vpxa_buf I78 ( .in(net39), .out(clkin_0_25));
ml_pump_vpxa_buf I81 ( .in(net22), .out(clkin_1_25));
ml_pump_vpxa_3_3v Ivpxa_pump_0 ( .en_25(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_0_25));
ml_pump_vpxa_3_3v Ivpxa_pump_2 ( .en_25(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_2_25));
ml_pump_vpxa_3_3v Ivpxa_pump_1 ( .en_25(pumpen_25),
     .clkin_25(clkin_1_25), .out(vpxa_int));
ml_pump_clk_reg Iclk_reg_0 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_0_25), .pump_on_25(pumpen_25),
     .clk_out_25(net39));
ml_pump_clk_reg Iclk_reg_2 ( .clk_in_25(vpxa_clk_b_25),
     .pump_chrg_25(pump_chrg_2_25), .pump_on_25(pumpen_25),
     .clk_out_25(net43));
ml_pump_clk_reg Iclk_reg_1 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_1_25), .pump_on_25(pumpen_25),
     .clk_out_25(net47));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_osc, View - schematic
// LAST TIME SAVED: Sep  2 15:47:56 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpxa_osc ( vpxa_clk_25, bgr, freq_25, pumpen_25 );
output  vpxa_clk_25;

inout  bgr;

input  pumpen_25;

input [1:0]  freq_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  freq_buf_b_25;



rppolywo_m  R6 ( .MINUS(gnd_), .PLUS(net043), .BULK(GND_));
rppolywo_m  R7 ( .MINUS(net043), .PLUS(net044), .BULK(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
pch_25  M9 ( .D(net061), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
pch_25  M10 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
pch_25  M8_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
pch_25  M8_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
nch_25  M12 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
nch_25  M11 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net044));
inv_25 I227 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I226 ( .IN(freq_25[0]), .OUT(freq_buf_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_vpp_vco Ivpx_vpp_vco ( .clk_25_1(net040), .pbias_25(pbias_25),
     .slow_25(net86), .freq_25({freq_25[1], freq_buf_b_25[0]}),
     .en_25(pumpen_25), .clk_25_0(vpxa_clk_25));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_ctrl, View - schematic
// LAST TIME SAVED: Sep  1 14:08:10 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpxa_ctrl ( pumpen, pumpen_25, vpxa_2_vdd, fsm_pumpen,
     fsm_tm_xforce, fsm_tm_xvpxaint );
output  pumpen, pumpen_25, vpxa_2_vdd;

input  fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I103 ( .A(vpxa_2_vdd), .B(net065), .Y(pumpen));
nand2_hvt I73 ( .A(fsm_tm_xvpxaint), .B(fsm_tm_xforce), .Y(net042));
inv_hvt I78 ( .A(pumpen), .Y(net075));
inv_hvt I77 ( .A(net042), .Y(net065));
inv_hvt I131 ( .A(fsm_pumpen), .Y(vpxa_2_vdd));
inv_25 I38 ( .IN(net045), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I173 ( .in(pumpen), .sup(vddp_), .out_vddio_b(net045),
     .out_vddio(net046), .in_b(net075));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff_25, View - schematic
// LAST TIME SAVED: Aug 30 17:06:17 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_dff_25 ( Q_25, Q_B_25, CLK_25, D_25, R_25 );
output  Q_25, Q_B_25;

input  CLK_25, D_25, R_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I96 ( .IN(Q_25), .OUT(Q_B_25), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I72 ( .IN(CLK_25), .OUT(net044), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I95 ( .IN(net044), .OUT(net038), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
ml_dlatch_25 Ilatch2 ( .D_25(net053), .EN_25(net038), .R_25(R_25),
     .Q_25(Q_25));
ml_dlatch_25 Ilatch1 ( .Q_25(net053), .EN_25(net044), .D_25(D_25),
     .R_25(R_25));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_n, View - schematic
// LAST TIME SAVED: Aug 30 15:13:05 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp_n ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M8 ( .D(out_ref), .B(GND_), .G(in_ref), .S(net049));
nch_25  M3 ( .D(out_div), .B(GND_), .G(in_div), .S(net049));
nch_25  M6_1_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
pch_25  M1 ( .D(out_ref), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M0 ( .D(out_div), .B(vddp_), .G(out_ref), .S(vddp_));
pch_25  M5 ( .D(out_div), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M7 ( .D(out_ref), .B(vddp_), .G(out_ref), .S(vddp_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_top_n, View - schematic
// LAST TIME SAVED: Aug 30 15:12:30 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp_top_n ( pump_chrg_25, in_div, in_ref, sa_bias,
     saen_25 );
output  pump_chrg_25;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I103 ( .G(gnd_), .Pb(vddp_), .A(saen_25), .Y(chrg_b_25),
     .P(vddp_), .B(net27), .Gb(gnd_));
nch_25  M6_1_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
inv_25 I102 ( .IN(chrg_b_25), .OUT(pump_chrg_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I104 ( .IN(out_div2), .OUT(net27), .P(vddp_), .Pb(vddp_),
     .G(net087), .Gb(gnd_));
ml_core_sa_comp_n Icore_sa_comp_n0 ( .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp_n Iml_core_sa_comp_n1 ( .out_div(out_div2),
     .out_ref(out_ref2), .in_div(in_div2), .in_ref(in_ref2),
     .sa_bias(sa_bias), .saen_25(saen_25));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_reg, View - schematic
// LAST TIME SAVED: Nov  6 18:01:31 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpxa_reg ( freq_25, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, vpxa_int, bgr, fsm_vrdwl, pumpen, vpxa_clk_25 );
output  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25;

inout  vpxa_int;

input  bgr, pumpen, vpxa_clk_25;

output [1:0]  freq_25;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  vrdwl_b_vpxa;

wire  [0:2]  vrdwl_vpxa;

wire  [0:1]  freq_in_25;



ml_ls_vdd2vdd25_vpxa I191 ( .in(saen_25), .sup(vpxa_int),
     .out_vddio_b(saen_b_vpxa), .out_vddio(net0210), .in_b(saen_b_25));
ml_ls_vdd2vdd25_vpxa I87 ( .in(net171), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[2]), .out_vddio(vrdwl_b_vpxa[2]),
     .in_b(net175));
ml_ls_vdd2vdd25_vpxa I98 ( .in(net176), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[1]), .out_vddio(vrdwl_b_vpxa[1]),
     .in_b(net180));
ml_ls_vdd2vdd25_vpxa I99 ( .in(net181), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[0]), .out_vddio(vrdwl_b_vpxa[0]),
     .in_b(net185));
rppolywo_m  R29 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R28 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R27 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(in_div_0), .PLUS(net202), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net232), .PLUS(net223), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(net270), .PLUS(net226), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net226), .PLUS(net229), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(sa_bias), .PLUS(net232), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net202), .PLUS(net237), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(net237), .PLUS(net270), .BULK(GND_));
rppolywo_m  R30 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(gnd_), .PLUS(in_div_2), .BULK(GND_));
rppolywo_m  R31 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
nch_25  M2 ( .D(sa_bias), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M32 ( .D(net229), .B(GND_), .G(vrdwl_b_vpxa[2]), .S(net226));
nch_25  M0_3_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_2_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_1_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_0_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M7 ( .D(net270), .B(GND_), .G(vrdwl_b_vpxa[0]), .S(net237));
nch_25  M4 ( .D(net226), .B(GND_), .G(vrdwl_b_vpxa[1]), .S(net270));
nand2_25 I194 ( .G(GND_), .Pb(vddp_), .A(net0179), .Y(freq_in_25[1]),
     .P(vddp_), .B(net0234), .Gb(GND_));
nand2_25 I145 ( .G(GND_), .Pb(vddp_), .A(net0171), .Y(freq_in_25[0]),
     .P(vddp_), .B(net0179), .Gb(GND_));
nand3_25 I193 ( .B(pump_chrg_1_b_25), .A(pump_chrg_2_25), .Y(net0171),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I192 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0179),
     .C(pump_chrg_0_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I159 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0234),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
pch_25  M3 ( .D(net229), .B(vpxa_int), .G(saen_b_vpxa), .S(vpxa_int));
pch_25  M11_1_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M11_0_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M37 ( .D(net226), .B(vpxa_int), .G(vrdwl_vpxa[2]), .S(net229));
pch_25  M1 ( .D(net223), .B(vddp_), .G(saen_b_25), .S(vddp_));
pch_25  M5 ( .D(net270), .B(vpxa_int), .G(vrdwl_vpxa[1]), .S(net226));
pch_25  M6 ( .D(net237), .B(vpxa_int), .G(vrdwl_vpxa[0]), .S(net270));
pch_25  M8_1_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
pch_25  M8_0_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
inv_25 I196 ( .IN(net169), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I197 ( .IN(net168), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I195 ( .IN(pump_chrg_0_25), .OUT(pump_chrg_0_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
inv_25 I154 ( .IN(pump_chrg_1_25), .OUT(pump_chrg_1_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_dff_25 I125 ( .Q_B_25(net0187), .R_25(saen_b_25),
     .D_25(freq_in_25[1]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[1]));
ml_dff_25 I126 ( .Q_B_25(net0192), .R_25(saen_b_25),
     .D_25(freq_in_25[0]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[0]));
inv_hvt I85 ( .A(net171), .Y(net175));
inv_hvt I183 ( .A(fsm_vrdwl[2]), .Y(net171));
inv_hvt I83 ( .A(pumpen), .Y(net143));
inv_hvt I82 ( .A(net143), .Y(net145));
inv_hvt I184 ( .A(fsm_vrdwl[1]), .Y(net176));
inv_hvt I187 ( .A(fsm_vrdwl[0]), .Y(net181));
inv_hvt I186 ( .A(net181), .Y(net185));
inv_hvt I185 ( .A(net176), .Y(net180));
ml_ls_vdd2vdd25 I335 ( .in(net145), .sup(vddp_), .out_vddio_b(net168),
     .out_vddio(net169), .in_b(net143));
ml_core_sa_comp_top_n Icore_sa_comp_top_n2 (
     .pump_chrg_25(pump_chrg_2_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_2));
ml_core_sa_comp_top_n core_sa_comp_top_n0 (
     .pump_chrg_25(pump_chrg_0_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_0));
ml_core_sa_comp_top_n Icore_sa_comp_top_n1 (
     .pump_chrg_25(pump_chrg_1_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_1));

endmodule
// Library - NVCM_40nm, Cell - ml_hv2vdd_sw, View - schematic
// LAST TIME SAVED: Aug 30 15:14:40 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hv2vdd_sw ( out_hv, hv2vdd, vddp_tieh );
inout  out_hv;

input  hv2vdd, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M2 ( .D(vdd_), .B(GND_), .G(hv2vdd_25), .S(net27));
nch_na25  M0 ( .D(net27), .B(GND_), .G(vddp_tieh), .S(out_hv));
inv_25 I62 ( .IN(net40), .OUT(hv2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I71 ( .A(net46), .Y(net44));
inv_hvt I72 ( .A(hv2vdd), .Y(net46));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net40),
     .out_vddio(net37), .in_b(net46));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_top, View - schematic
// LAST TIME SAVED: Nov  8 10:18:53 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_vpxa_top ( vpxa_int, bgr, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint, fsm_vrdwl );
inout  vpxa_int;

input  bgr, fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  freq_25;



nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpxa_int));
inv_25 I73 ( .IN(vpxa_clk_25), .OUT(vpxa_clk_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_pump_vpxa_x2 Ipump_vpxa_x3 ( .vpxa_clk_b_25(vpxa_clk_b_25),
     .vpxa_clk_25(vpxa_clk_25), .pumpen_25(pumpen_25),
     .pump_chrg_2_25(pump_chrg_2_25), .pump_chrg_1_25(pump_chrg_1_25),
     .pump_chrg_0_25(pump_chrg_0_25), .vpxa_int(vpxa_int));
ml_vpxa_osc Ivpxa_osc ( .freq_25(freq_25[1:0]), .bgr(bgr),
     .pumpen_25(pumpen_25), .vpxa_clk_25(vpxa_clk_25));
ml_vpxa_ctrl Ivpxa_ctrl ( .fsm_pumpen(fsm_pumpen), .pumpen(pumpen),
     .pumpen_25(pumpen_25), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .vpxa_2_vdd(vpxa_2_vdd));
vddp_tiehigh I118 ( .vddp_tieh(vddp_tieh));
ml_vpxa_reg Ivpxa_reg ( .pump_chrg_0_25(pump_chrg_0_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_2_25(pump_chrg_2_25),
     .freq_25(freq_25[1:0]), .vpxa_clk_25(vpxa_clk_25),
     .pumpen(pumpen), .fsm_vrdwl(fsm_vrdwl[2:0]), .bgr(bgr),
     .vpxa_int(vpxa_int));
ml_hv2vdd_sw Ivpxa_2vdd_sw ( .vddp_tieh(vddp_tieh),
     .hv2vdd(vpxa_2_vdd), .out_hv(vpxa_int));

endmodule
// Library - xpmem, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Aug 20 09:48:05 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - NVCM_40nm, Cell - ml_rdhv_gen, View - schematic
// LAST TIME SAVED: Jul 27 12:15:43 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_rdhv_gen ( s_rdin_hv, srdsup_hv, s_rdin, vddp_tieh );
output  s_rdin_hv;

inout  srdsup_hv;

input  s_rdin, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_s_b_hv_sw Iml_s_b_25_sw ( .sbout_high_25(s_rdin_high_25),
     .sbout_gnd_25(net31), .sbout_hv(s_rdin_hv), .ssup_hv(srdsup_hv),
     .vddp_tieh(vddp_tieh));
ml_ls_vdd2vdd25 Iml_ls_vdd2vdd25 ( .in(s_rdin), .sup(vddp_),
     .out_vddio_b(net31), .out_vddio(s_rdin_high_25), .in_b(net35));
inv_hvt I439 ( .A(s_rdin), .Y(net35));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_top_ctrl, View - schematic
// LAST TIME SAVED: Nov  5 16:32:34 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hvmux_top_ctrl ( bgrext_en, bgrint_en, en_vblinhi,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp, fsm_lshven,
     fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en );
output  bgrext_en, bgrint_en, en_vblinhi, ngate_vddp, ngate_vpxa,
     sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint,
     vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint, vpxaint_ext,
     vtmode, ysup25_2vdd, ysup25_2vddp;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor4_hvt I186 ( .D(fsm_tm_rprd), .C(fsm_rd), .A(fsm_tm_rd_mode),
     .B(fsm_pgmvfy), .Y(net0349));
nand4_hvt I322 ( .D(fsm_lshven), .A(fsm_pgm), .C(fsm_lshven),
     .Y(pgmpulse_b), .B(net0236));
nand4_hvt I35 ( .D(fsm_lshven), .C(net0318), .A(fsm_pgm), .Y(net0196),
     .B(net0327));
anor21_hvt I245 ( .A(net0189), .B(net0193), .Y(vppint_ext),
     .C(net0190));
anor21_hvt I109 ( .A(net0201), .B(net0199), .Y(vpxa_ext), .C(net0190));
nand3_hvt I288 ( .Y(net0193), .B(pmprd), .C(pmprd),
     .A(fsm_tm_xvppint));
nand3_hvt I291 ( .Y(net0201), .B(vddp_rd_b), .C(gnd_tiel),
     .A(fsm_tm_xforce));
nand3_hvt I292 ( .Y(net0213), .B(net0321), .C(net0196), .A(net0321));
nand3_hvt I290 ( .Y(net0199), .B(pmprd), .C(pmprd), .A(gnd_tiel));
nand3_hvt I289 ( .Y(net0189), .B(vpint_en), .C(fsm_tm_xvppint),
     .A(fsm_tm_xforce));
nor3_hvt I286 ( .B(net0240), .Y(rd_vddp), .A(net0240),
     .C(fsm_nvcmen_b));
nor3_hvt I285 ( .B(tm_testdec), .Y(en_vblinhi), .A(fsm_nvcmen_b),
     .C(tm_allbl_l));
mux2_hvt I260 ( .in1(fsm_wgnden), .in0(fsm_wpen), .out(net0217),
     .sel(pgmpulse_b));
nor2_hvt I272 ( .A(net75), .B(net93), .Y(ysup25_2vdd));
nor2_hvt I279 ( .A(net0251), .B(net0266), .Y(sbhvsup_vppint));
nor2_hvt I283 ( .A(vddp_rd_b), .B(net0258), .Y(vpxa_vppd));
nor2_hvt I271 ( .A(net87), .B(net73), .Y(ysup25_2vddp));
nor2_hvt I273 ( .A(net0349), .B(net0240), .Y(vddp_rd));
nor2_hvt I281 ( .A(net0324), .B(fsm_nvcmen_b), .Y(net0251));
nor2_hvt I276 ( .A(net0272), .B(rd_vddp), .Y(ngate_vpxa));
nor2_hvt I280 ( .A(net0268), .B(net0213), .Y(sb25sup_vpxa));
nor2_hvt I275 ( .A(net0331), .B(net0270), .Y(ngate_vddp));
nor2_hvt I274 ( .A(fsm_tm_rprd), .B(gnd_tiel), .Y(net0240));
nor2_hvt I278 ( .A(net0264), .B(net0311), .Y(sbhvsup_vddp));
nor2_hvt I282 ( .A(net0256), .B(vddp_rd), .Y(vpxa_vpxaint));
nor2_hvt I277 ( .A(net0325), .B(net0260), .Y(sb25sup_vddp));
inv_hvt I294 ( .A(net77), .Y(vtmode));
inv_hvt I323 ( .A(fsm_pgmvfy), .Y(net0236));
inv_hvt I319 ( .A(ngate_vpxa), .Y(net0339));
inv_hvt I304 ( .A(net0251), .Y(net0311));
inv_hvt I315 ( .A(vddp_rd), .Y(vddp_rd_b));
inv_hvt I318 ( .A(ysup25_2vdd), .Y(ysup25_2vdd_b));
inv_hvt I314 ( .A(vpxa_vppd), .Y(net0297));
inv_hvt I309 ( .A(net0277), .Y(bgrext_en));
inv_hvt I317 ( .A(fsm_pgmvfy), .Y(net0327));
inv_hvt I316 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I297 ( .A(ysup25_2vddp), .Y(ysup25_2vddp_b));
inv_hvt I298 ( .A(rd_vddp), .Y(net0331));
inv_hvt I310 ( .A(fsm_pumpen), .Y(net0190));
inv_hvt I307 ( .A(sbhvsup_vddp), .Y(net0309));
inv_hvt I305 ( .A(sb25sup_vpxa), .Y(net0323));
inv_hvt I308 ( .A(sbhvsup_vppint), .Y(net0313));
inv_hvt I296 ( .A(net93), .Y(net87));
inv_hvt I295 ( .A(net80), .Y(net93));
inv_hvt I321 ( .A(fsm_tm_rprd), .Y(net0318));
inv_hvt I303 ( .A(pgmpulse_b), .Y(net0324));
inv_hvt I306 ( .A(pgmpulse_b), .Y(pgmpulse));
inv_hvt I300 ( .A(sb25sup_vddp), .Y(net0329));
inv_hvt I302 ( .A(rd_vddp), .Y(net0321));
inv_hvt I301 ( .A(net0213), .Y(net0325));
inv_hvt I311 ( .A(net0286), .Y(vpxaint_ext));
inv_hvt I312 ( .A(fsm_tm_xforce), .Y(pmprd));
inv_hvt I299 ( .A(ngate_vddp), .Y(net0335));
inv_hvt I313 ( .A(vpxa_vpxaint), .Y(net0319));
inv_hvt I233 ( .A(fsm_nvcmen_b), .Y(fsm_nvcmen_buf));
nand2_hvt I268 ( .A(fsm_nvcmen_buf), .Y(net0277), .B(fsm_tm_xvbg));
nand2_hvt I266 ( .A(fsm_nvcmen), .Y(net80), .B(net0217));
nand2_hvt I269 ( .A(bgrext_en), .Y(bgrint_en), .B(fsm_tm_xforce));
nand2_hvt I267 ( .A(fsm_pumpen), .Y(net0286), .B(fsm_tm_xvpxaint));
nand2_hvt I104 ( .A(fsm_nvcmen), .Y(net77), .B(tm_wleqbl));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
ml_pump_a_clkdly I219 ( .in(ysup25_2vddp_b), .out(net75));
ml_pump_a_clkdly I227 ( .in(net0297), .out(net0256));
ml_pump_a_clkdly I226 ( .in(net0319), .out(net0258));
ml_pump_a_clkdly I209 ( .in(net0323), .out(net0260));
ml_pump_a_clkdly I184 ( .in(ysup25_2vdd_b), .out(net73));
ml_pump_a_clkdly I217 ( .in(net0313), .out(net0264));
ml_pump_a_clkdly I216 ( .in(net0309), .out(net0266));
ml_pump_a_clkdly I208 ( .in(net0329), .out(net0268));
ml_pump_a_clkdly I198 ( .in(net0339), .out(net0270));
ml_pump_a_clkdly I197 ( .in(net0335), .out(net0272));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_ls25, View - schematic
// LAST TIME SAVED: Sep  7 10:34:50 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hvmux_ls25 ( bgrext_en_25, bgrint_en_25, ngate_vddp_25,
     ngate_vpxa_25, sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25, bgrext_en, bgrint_en,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp );
output  bgrext_en_25, bgrint_en_25, ngate_vddp_25, ngate_vpxa_25,
     sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25;

input  bgrext_en, bgrint_en, ngate_vddp, ngate_vpxa, sb25sup_vddp,
     sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint, vppint_ext, vpxa_ext,
     vpxa_vppd, vpxa_vpxaint, vpxaint_ext, vtmode, ysup25_2vdd,
     ysup25_2vddp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I471 ( .IN(net0138), .OUT(bgrint_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I472 ( .IN(net0148), .OUT(bgrext_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I473 ( .IN(net0128), .OUT(vppint_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I474 ( .IN(net0123), .OUT(vpxa_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I475 ( .IN(net0158), .OUT(vpxaint_ext_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I476 ( .IN(net0133), .OUT(vpxa_vppd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I477 ( .IN(net0163), .OUT(vpxa_vpxaint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I406 ( .IN(net077), .OUT(ysup25_2vddp_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I463 ( .IN(net0168), .OUT(ysup25_2vdd_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I464 ( .IN(net0193), .OUT(vtmode_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I465 ( .IN(net0173), .OUT(ngate_vddp_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I466 ( .IN(net0183), .OUT(ngate_vpxa_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I467 ( .IN(net0188), .OUT(sb25sup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I468 ( .IN(net0153), .OUT(sb25sup_vpxa_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I469 ( .IN(net0203), .OUT(sbhvsup_vppint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I470 ( .IN(net0198), .OUT(sbhvsup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_hvt I457 ( .A(vpxa_vppd), .Y(net054));
inv_hvt I435 ( .A(vpxa_vpxaint), .Y(net0112));
inv_hvt I462 ( .A(bgrint_en), .Y(net058));
inv_hvt I461 ( .A(bgrext_en), .Y(net068));
inv_hvt I460 ( .A(vppint_ext), .Y(net066));
inv_hvt I455 ( .A(ysup25_2vddp), .Y(net0328));
inv_hvt I454 ( .A(ysup25_2vdd), .Y(net0312));
inv_hvt I447 ( .A(ngate_vpxa), .Y(net0318));
inv_hvt I439 ( .A(sbhvsup_vppint), .Y(net0326));
inv_hvt I446 ( .A(sb25sup_vddp), .Y(net0320));
inv_hvt I216 ( .A(ysup25_2vdd), .Y(net092));
inv_hvt I458 ( .A(vpxaint_ext), .Y(net060));
inv_hvt I442 ( .A(sbhvsup_vddp), .Y(net0324));
inv_hvt I443 ( .A(sb25sup_vpxa), .Y(net0322));
inv_hvt I450 ( .A(ngate_vddp), .Y(net0316));
inv_hvt I217 ( .A(net092), .Y(ysup25_2vdd_buf));
inv_hvt I451 ( .A(vtmode), .Y(net0314));
inv_hvt I459 ( .A(vpxa_ext), .Y(net082));
ml_ls_vdd2vdd25 I336 ( .in(vpxa_ext), .sup(vddp_),
     .out_vddio_b(net0123), .out_vddio(net0207), .in_b(net082));
ml_ls_vdd2vdd25 I337 ( .in(vppint_ext), .sup(vddp_),
     .out_vddio_b(net0128), .out_vddio(net0208), .in_b(net066));
ml_ls_vdd2vdd25 I338 ( .in(vpxa_vppd), .sup(vddp_),
     .out_vddio_b(net0133), .out_vddio(net0211), .in_b(net054));
ml_ls_vdd2vdd25 I339 ( .in(bgrint_en), .sup(vddp_),
     .out_vddio_b(net0138), .out_vddio(net0209), .in_b(net058));
ml_ls_vdd2vdd25 I332 ( .in(bgrext_en), .sup(vddp_),
     .out_vddio_b(net0148), .out_vddio(net0149), .in_b(net068));
ml_ls_vdd2vdd25 I238 ( .in(sb25sup_vpxa), .sup(vddp_),
     .out_vddio_b(net0153), .out_vddio(net0154), .in_b(net0322));
ml_ls_vdd2vdd25 I334 ( .in(vpxaint_ext), .sup(vddp_),
     .out_vddio_b(net0158), .out_vddio(net0214), .in_b(net060));
ml_ls_vdd2vdd25 I335 ( .in(vpxa_vpxaint), .sup(vddp_),
     .out_vddio_b(net0163), .out_vddio(net0206), .in_b(net0112));
ml_ls_vdd2vdd25 I212 ( .in(ysup25_2vdd), .sup(vddp_),
     .out_vddio_b(net0168), .out_vddio(net0169), .in_b(net0312));
ml_ls_vdd2vdd25 I226 ( .in(ngate_vddp), .sup(vddp_),
     .out_vddio_b(net0173), .out_vddio(net0174), .in_b(net0316));
ml_ls_vdd2vdd25 I203 ( .in(net0328), .sup(vddp_), .out_vddio_b(net077),
     .out_vddio(net078), .in_b(ysup25_2vddp));
ml_ls_vdd2vdd25 I221 ( .in(ngate_vpxa), .sup(vddp_),
     .out_vddio_b(net0183), .out_vddio(net0184), .in_b(net0318));
ml_ls_vdd2vdd25 I233 ( .in(sb25sup_vddp), .sup(vddp_),
     .out_vddio_b(net0188), .out_vddio(net0219), .in_b(net0320));
ml_ls_vdd2vdd25 I207 ( .in(vtmode), .sup(vddp_), .out_vddio_b(net0193),
     .out_vddio(net0194), .in_b(net0314));
ml_ls_vdd2vdd25 I260 ( .in(sbhvsup_vddp), .sup(vddp_),
     .out_vddio_b(net0198), .out_vddio(net0220), .in_b(net0324));
ml_ls_vdd2vdd25 I261 ( .in(sbhvsup_vppint), .sup(vddp_),
     .out_vddio_b(net0203), .out_vddio(net0204), .in_b(net0326));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_bgrxcvr, View - schematic
// LAST TIME SAVED: Sep  3 09:50:30 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hvmux_bgrxcvr ( bgr, bgr_int, bgrint_en_25, vpp,
     bgrext_en_25, vddp_tieh );
inout  bgr, bgr_int, bgrint_en_25, vpp;

input  bgrext_en_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M2 ( .D(vpp), .B(GND_), .G(vddp_tieh), .S(net53));
nch_25  M1 ( .D(net53), .B(GND_), .G(bgrext_en_25), .S(bgr));
nch_na25  M0 ( .D(bgr), .B(GND_), .G(bgrint_en_25), .S(bgr_int));

endmodule
// Library - NVCM_40nm, Cell - ml_ysup_25_switch, View - schematic
// LAST TIME SAVED: Sep  3 09:40:13 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_ysup_25_switch ( vdd, vddp, ysup_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25 );
inout  vdd, vddp, ysup_25;

input  ysup25_2vdd_25, ysup25_2vdd_buf, ysup25_2vddp_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd), .B(GND_), .G(ysup25_2vdd_25), .S(ysup_25));
pch_25  M5 ( .D(net73), .B(vddp), .G(ysup25_2vddp_b_25), .S(vddp));
pch_25  M0 ( .D(ysup_25), .B(ysup_25), .G(ysup25_2vdd_buf), .S(net73));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_vblinhi, View - schematic
// LAST TIME SAVED: Nov  8 18:40:26 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_vblinhi ( vblinhi, vpxa, en_vblinhi, vtmode,
     vtmode_25 );
inout  vblinhi, vpxa;

input  en_vblinhi, vtmode, vtmode_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M0_9_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_8_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_7_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_6_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_5_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_4_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_3_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_2_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_1_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_0_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
pch_hvt  M7_9_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_8_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_7_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_6_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_5_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_4_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_3_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_2_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_1_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_0_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
nch_25  M9 ( .D(net035), .B(GND_), .G(net035), .S(vblinhi));
nch_25  M8 ( .D(vpxa), .B(GND_), .G(vtmode_25), .S(net035));
nor2_hvt I191 ( .A(en_vblinhi), .B(vtmode_buf), .Y(ngate_inhi_lv));
inv_hvt I192 ( .A(net063), .Y(vtmode_buf));
inv_hvt I190 ( .A(vtmode), .Y(net063));
nand2_hvt I104 ( .A(net063), .Y(pgate_inhi_lv), .B(en_vblinhi));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_top, View - schematic
// LAST TIME SAVED: Nov 24 19:40:38 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_hvmux_top ( s_rdin_hv, bgr, bgr_int, ngate_25, sb25sup_25,
     sbhvsup_hv, srdsup_hv, vblinhi, vpp, vpp_int, vpxa, vpxa_int,
     ysup_25, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen,
     fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, s_rd,
     tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );

inout  bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv,
     vblinhi, vpp, vpp_int, vpxa, vpxa_int, ysup_25;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en;

output [3:0]  s_rdin_hv;

input [3:0]  s_rd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_rdin;

wire  [0:3]  net294;



nch_hvt  M1 ( .D(net299), .B(GND_), .G(net299), .S(gnd_));
inv_hvt I210_3_ ( .A(s_rd[3]), .Y(net294[0]));
inv_hvt I210_2_ ( .A(s_rd[2]), .Y(net294[1]));
inv_hvt I210_1_ ( .A(s_rd[1]), .Y(net294[2]));
inv_hvt I210_0_ ( .A(s_rd[0]), .Y(net294[3]));
inv_hvt I211_3_ ( .A(net294[0]), .Y(s_rdin[3]));
inv_hvt I211_2_ ( .A(net294[1]), .Y(s_rdin[2]));
inv_hvt I211_1_ ( .A(net294[2]), .Y(s_rdin[1]));
inv_hvt I211_0_ ( .A(net294[3]), .Y(s_rdin[0]));
ml_rdhv_gen Iml_rdhv_inv_3_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[3]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[3]));
ml_rdhv_gen Iml_rdhv_inv_2_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[2]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[2]));
ml_rdhv_gen Iml_rdhv_inv_1_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[1]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[1]));
ml_rdhv_gen Iml_rdhv_inv_0_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[0]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[0]));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net299), .S(vddp_));
ml_hv_hotswitch_enhance Ixcvr_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(vppint_ext_25), .hv_in_hv(vpp_int), .hv_out_hv(vpp));
ml_hvmux_top_ctrl Ihvmux_top_ctrl ( .fsm_tm_rprd(fsm_tm_rprd),
     .vpint_en(vpint_en), .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl),
     .tm_testdec(tm_testdec), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_lshven(fsm_lshven), .ysup25_2vddp(ysup25_2vddp),
     .ysup25_2vdd(ysup25_2vdd), .vtmode(vtmode),
     .vpxaint_ext(vpxaint_ext), .vpxa_vpxaint(vpxa_vpxaint),
     .vpxa_vppd(vpxa_vppd), .vpxa_ext(vpxa_ext),
     .vppint_ext(vppint_ext), .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .en_vblinhi(en_vblinhi),
     .bgrint_en(bgrint_en), .bgrext_en(bgrext_en));
ml_hvmux_ls25 Ihvmux_ls25 ( .ysup25_2vddp(ysup25_2vddp),
     .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vppint_25(sbhvsup_vppint_25), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en), .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vtmode_25(vtmode_25),
     .vpxaint_ext_25(vpxaint_ext_25),
     .vpxa_vpxaint_25(vpxa_vpxaint_25), .vpxa_vppd_25(vpxa_vppd_25),
     .vpxa_ext_25(net309), .vppint_ext_25(vppint_ext_25),
     .sbhvsup_vddp_25(sbhvsup_vddp_25),
     .sb25sup_vpxa_25(sb25sup_vpxa_25),
     .sb25sup_vddp_25(sb25sup_vddp_25), .ngate_vpxa_25(ngate_vpxa_25),
     .ngate_vddp_25(ngate_vddp_25), .bgrint_en_25(bgrint_en_25),
     .bgrext_en_25(bgrext_en_25));
ml_hvmux_bgrxcvr Ixcvr_bgr ( .vddp_tieh(vddp_tieh),
     .bgrext_en_25(bgrext_en_25), .vpp(vpp),
     .bgrint_en_25(bgrint_en_25), .bgr_int(bgr_int), .bgr(bgr));
ml_hv_hotswitch Ixcvr_vpxa_int ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa_int), .hv_out_hv(vpp));
ml_hvmux_hotswitch I212 ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(srdsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sbhvsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(sbhvsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sb25sup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sb25sup_vpxa_25), .sel_hv_a_25(sb25sup_vddp_25),
     .out_hv(sb25sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_ngate ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(ngate_vpxa_25), .sel_hv_a_25(ngate_vddp_25),
     .out_hv(ngate_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_1_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vddp_), .hvin_a_hv(vpxa_int));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_0_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vddp_), .hvin_a_hv(vpxa_int));
ml_ysup_25_switch Isw_ysup25_1_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ysup_25_switch Isw_ysup25_0_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_1_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_0_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_hvsw_8f, View - schematic
// LAST TIME SAVED: Nov  6 17:49:25 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_chip_nvcm_hvsw_8f ( s_rdin_hv, bgr, ngate_25, sb25sup_25,
     sbhvsup_hv, srdsup_hv, vblinhi, vpp, vpp_int, vpxa, ysup_25,
     fsm_bgr_dis, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint,
     fsm_tm_xvpxaint, fsm_trim_vbg, fsm_vpgmwl, fsm_vrdwl, fsm_wgnden,
     fsm_wpen, s_rd, tm_allbl_l, tm_wleqbl );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi, vpp,
     vpp_int, vpxa, ysup_25;

input  fsm_bgr_dis, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_wleqbl;

output [3:0]  s_rdin_hv;

input [2:0]  fsm_vrdwl;
input [3:0]  fsm_trim_vbg;
input [3:0]  s_rd;
input [2:0]  fsm_vpgmwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  fsm_vrdw_buf;

wire  [3:0]  fsm_trim_vbg_buf;



ml_chip_buf_hvsw_8f Ichip_buf_top ( .fsm_bgr_dis(fsm_bgr_dis),
     .fsm_pumpen_buf(fsm_pumpen_buf),
     .fsm_vrdwl_buf(fsm_vrdw_buf[2:0]), .fsm_vrdwl(fsm_vrdwl[2:0]),
     .fsm_tm_xvpxaint_buf(net193),
     .fsm_tm_xforce_buf(fsm_tm_xforce_buf),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_bgr_dis_buf(fsm_bgr_dis_buf), .fsm_pumpen(fsm_pumpen),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]), .fsm_nvcmen(fsm_nvcmen),
     .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen_buf));
ml_bgr_top Ibgr_top ( .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .fsm_bgr_dis_buf(fsm_bgr_dis_buf), .bgr_int(bgr_int));
ml_vppint_top Ivppint_top ( .vpxa(vpxa),
     .fsm_vpgmwl_buf(fsm_vpgmwl[2:0]), .fsm_pgmdisc_buf(fsm_pgmdisc),
     .fsm_pgm_buf(fsm_pgm), .fsm_lshven_buf(fsm_lshven),
     .vpint_en(vpint_en), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmvfy_buf(fsm_pgmvfy), .fsm_wgnden_buf(fsm_wgnden),
     .fsm_nvcmen_buf(fsm_nvcmen), .bgr(bgr), .vpp_int(vpp_int),
     .fsm_tm_xvppint(fsm_tm_xvppint));
ml_vpxa_top Ivpxa_top ( .fsm_vrdwl(fsm_vrdw_buf[2:0]),
     .fsm_tm_xvpxaint(net193), .fsm_tm_xforce(fsm_tm_xforce_buf),
     .bgr(bgr), .vpxa_int(vpxa_int), .fsm_pumpen(fsm_pumpen_buf));
ml_hvmux_top Ihvmux_top ( .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_lshven(fsm_lshven), .bgr(bgr), .bgr_int(bgr_int),
     .ngate_25(ngate_25), .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .vpp(vpp), .vpp_int(vpp_int),
     .vpxa(vpxa), .ysup_25(ysup_25), .vblinhi(vblinhi),
     .tm_testdec(fsm_tm_testdec), .srdsup_hv(srdsup_hv),
     .s_rd(s_rd[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rdin_hv(s_rdin_hv[3:0]), .vpint_en(vpint_en),
     .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl), .vpxa_int(vpxa_int));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_1f, View - schematic
// LAST TIME SAVED: May 26 11:17:02 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_chip_nvcm_1f ( nv_dataout, vpp, fsm_bgr_dis, fsm_blkadd,
     fsm_blkadd_b, fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven,
     fsm_multibl_read, fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rowadd, fsm_rst_b,
     fsm_sample, fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_trim_ipp, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_trim_vbg, fsm_vpgmwl, fsm_vpxaset, fsm_vrdwl,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr, tm_wleqbl );

inout  vpp;

input  fsm_bgr_dis, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxaint,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl;

output [8:0]  nv_dataout;

input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_trim_vbg;
input [2:0]  fsm_vpgmwl;
input [2:0]  fsm_vrdwl;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_trim_ipp;
input [9:0]  fsm_coladd;
input [1:0]  fsm_tm_ref;
input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_rdin_hv;

wire  [3:0]  s_rd;



ml_chip_nvcm_core_1f Iml_chip_nvcm_core_1f (
     .fsm_tm_ref(fsm_tm_ref[1:0]), .fsm_wren(fsm_wren),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rdin_hv(s_rdin_hv[3:0]),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[8:0]),
     .fsm_pgmhv(fsm_pgmhv), .fsm_gwlbdis(fsm_gwlbdis),
     .vpp_int(vpp_int), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_pgm(fsm_pgm),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_din(fsm_din), .fsm_rd(fsm_rd), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_pgmdisc(fsm_pgmdisc),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ngate_25(ngate_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol), .bgr(bgr),
     .fsm_blkadd(fsm_blkadd[3:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi(vblinhi), .s_rd(s_rd[3:0]), .srdsup_hv(srdsup_hv),
     .ysup_25(ysup_25), .vpxa(vpxa));
ml_chip_nvcm_hvsw_8f Ihvsw ( .bgr(bgr),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .vpp_int(vpp_int), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd), .fsm_wpen(fsm_wpen),
     .s_rdin_hv(s_rdin_hv[3:0]), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .srdsup_hv(srdsup_hv), .s_rd(s_rd[3:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .tm_allbl_l(tm_allbl_l),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_pumpen(fsm_pumpen), .sb25sup_25(sb25sup_25),
     .fsm_lshven(fsm_lshven), .sbhvsup_hv(sbhvsup_hv), .vpxa(vpxa),
     .ysup_25(ysup_25), .ngate_25(ngate_25), .fsm_wgnden(fsm_wgnden),
     .vblinhi(vblinhi), .tm_wleqbl(tm_wleqbl), .vpp(vpp),
     .fsm_vrdwl(fsm_vrdwl[2:0]), .fsm_bgr_dis(fsm_bgr_dis),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_vpgmwl(fsm_vpgmwl[2:0]), .fsm_tm_testdec(fsm_tm_testdec));
nmoscap_25  C0 ( .MINUS(GND_), .PLUS(vddp_));
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(vddp_));

endmodule
// Library - ice8chip, Cell - sg_bufx10_ice8p, View - schematic
// LAST TIME SAVED: Sep  1 14:14:18 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module sg_bufx10_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - bram_bufferx16_2inv, View - schematic
// LAST TIME SAVED: May 13 10:13:11 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_bufferx16_2inv ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I4 ( .A(net6), .Y(out));
inv I3 ( .A(in), .Y(net6));

endmodule
// Library - ice1chip, Cell - nvcm_ml_block_ice1f_june, View -
//schematic
// LAST TIME SAVED: Jun 29 10:02:26 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module nvcm_ml_block_ice1f_june ( bp0, fsm_recall, fsm_tm_margin0_read,
     nvcm_boot, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b,
     tgnd_fsm, tvdd_fsm, vpp, clk, nvcm_ce_b, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b, tgnd_fsm, tvdd_fsm;

inout  vpp;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [8:0]  nv_dataout;

wire  [3:0]  fsm_blkadd;

wire  [2:0]  fsm_trim_vrdwl;

wire  [2:0]  fsm_trim_vpgmwl;

wire  [3:0]  fsm_trim_vbg;

wire  [2:0]  fsm_trim_rrefrd;

wire  [2:0]  fsm_trim_rrefpgm;

wire  [3:0]  fsm_trim_ipp;

wire  [3:0]  fsm_blkadd_b;

wire  [1:0]  fsm_tm_ref_buf;

wire  [11:0]  fsm_coladd;

wire  [8:0]  fsm_rowadd;


/*
nvcm_top_ice8p I_nvcm_top_ice8p ( .fsm_tm_bgr_dis(fsm_bgr_dis),
     .fsm_tm_allbank_sel(fsm_tm_allbank_sel),
     .fsm_coladd(fsm_coladd[11:0]), .nvcm_max_coladd({tgnd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tgnd_fsm, tvdd_fsm, tgnd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm, tvdd_fsm}),
     .nvcm_max_rowadd({tgnd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm, tvdd_fsm}),
     .status_wip(net249), .fsm_tm_ref(fsm_tm_ref_buf[1:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .nvcm_boot(nvcm_boot),
     .spi_ss_b(spi_ss_b), .spi_sdi(spi_sdi),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_ce_b(nvcm_ce_b), .nv_dataout(nv_dataout[8:0]), .clk(clk),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .nvcm_relextspi(nvcm_relextspi), .nvcm_rdy(nvcm_rdy),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_trim_vrdwl(fsm_trim_vrdwl[2:0]),
     .fsm_trim_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_multibl_read(fsm_trim_multibl_read),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxa_int(fsm_tm_xvpxa_int), .fsm_tm_xvpp(fsm_tm_xvpp),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_vwleqbl(fsm_tm_vwleqbl),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_testdec_wr(fsm_tm_testdec_wr),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_tcol(fsm_tm_tcol),
     .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_margin0_read(fsm_tm_margin0_read),
     .fsm_tm_dma(fsm_tm_dma), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_sample(fsm_sample),
     .fsm_rowadd(fsm_rowadd[8:0]), .fsm_recall(fsm_recall),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_redrow(fsm_nv_redrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .bp0(bp0));
ml_chip_nvcm_1f I_ml_chip_nvcm ( .fsm_tm_ref(fsm_tm_ref_buf[1:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .fsm_bgr_dis(fsm_bgr_dis),
     .tm_allbank_sel(fsm_tm_allbank_sel), .fsm_coladd(fsm_coladd[9:0]),
     .tm_wleqbl(fsm_tm_vwleqbl), .tm_testdec_wr(fsm_tm_testdec_wr),
     .tm_tcol(fsm_tm_tcol), .tm_dma(fsm_tm_dma),
     .tm_allwl_l(fsm_tm_allwl_l), .tm_allwl_h(fsm_tm_allwl_h),
     .tm_allbl_l(fsm_tm_allbl_l), .tm_allbl_h(fsm_tm_allbl_h),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vrdwl(fsm_trim_vrdwl[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxaint(fsm_tm_xvpxa_int), .fsm_tm_xvppint(fsm_tm_xvpp),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(rst_bd), .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rrow(fsm_nv_redrow), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_multibl_read(fsm_trim_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .nv_dataout(nv_dataout[8:0]), .vpp(vpp));
tiehi I442 ( .tiehi(tvdd_fsm));
tielo I369 ( .tielo(tgnd_fsm));
sg_bufx10_ice8p I541 ( .in(rst_b), .out(rst_bd));
*/
endmodule
// Library - ice8chip, Cell - smc_and_jtag_ice8p, View - schematic
// LAST TIME SAVED: Sep 30 15:13:23 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module smc_and_jtag_ice8p ( bm_bank_sdi, bm_banksel, bm_clk, bm_init,
     bm_rcapmux_en, bm_sa, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_banksel, cm_clk, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2, cm_sdi_u3, data_muxsel, data_muxsel1,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0, j_hiz_b,
     j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck, j_tdi,
     j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, psdo, rst_b,
     smc_load_nvcm_bstream, smc_osc_fsel, smc_oscoff_b, smc_podt_off,
     smc_podt_rst, smc_read, smc_row_inc, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rsr_rst, smc_rwl_en, smc_seq_rst,
     smc_wcram_rst, smc_wdis_dclk, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, tdo_oe_pad, tdo_pad,
     bm_bank_sdo, boot, bp0, bschain_sdo, cdone_in, cm_last_rsr,
     cm_monitor_cell, cm_sdo_u0, cm_sdo_u1, cm_sdo_u2, cm_sdo_u3,
     cnt_podt_out, coldboot_sel, creset_b, idcode_msb20bits, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     osc_clk, por_b, psdi, spi_clk_in, spi_sdi, spi_ss_in_b, tck_pad,
     tdi_pad, tms_pad, trst_pad, warmboot_sel );
output  bm_clk, bm_init, bm_rcapmux_en, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_clk, data_muxsel,
     data_muxsel1, en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0,
     j_hiz_b, j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck,
     j_tdi, j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, rst_b,
     smc_load_nvcm_bstream, smc_oscoff_b, smc_podt_off, smc_podt_rst,
     smc_read, smc_row_inc, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rsr_rst, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_wdis_dclk, smc_write, smc_wset_prec, smc_wset_precgnd,
     smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_oe_pad, tdo_pad;

input  boot, bp0, bschain_sdo, cdone_in, cm_last_rsr, cnt_podt_out,
     creset_b, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, osc_clk, por_b, spi_clk_in, spi_sdi,
     spi_ss_in_b, tck_pad, tdi_pad, tms_pad, trst_pad;

output [10:0]  bm_sa;
output [1:0]  cm_sdi_u2;
output [1:0]  smc_osc_fsel;
output [3:0]  bm_banksel;
output [3:0]  cm_banksel;
output [7:1]  psdo;
output [1:0]  cm_sdi_u3;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_sdi_u0;
output [3:0]  bm_bank_sdi;

input [3:0]  cm_monitor_cell;
input [1:0]  cm_sdo_u0;
input [7:1]  psdi;
input [1:0]  coldboot_sel;
input [1:0]  warmboot_sel;
input [19:0]  idcode_msb20bits;
input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdo_u2;
input [3:0]  bm_bank_sdo;
input [1:0]  cm_sdo_u3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - xpmem, Cell - ml_buf_ice5_2, View - schematic
// LAST TIME SAVED: Jun 14 11:22:45 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_buf_ice5_2 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_rowdrv2_last, View - schematic
// LAST TIME SAVED: Aug 18 15:57:39 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_rowdrv2_last ( pgate, reset, smc_rsr_out, vddctrl, wl,
     wl_rd_sup, wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write
     );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
ml_dff I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));

endmodule
// Library - xpmem, Cell - ml_rowdrvsup2, View - schematic
// LAST TIME SAVED: Jul 23 17:04:42 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_rowdrvsup2 ( wl_rd_sup, wl_rden_b );
inout  wl_rd_sup, wl_rden_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R2 ( .MINUS(net089), .PLUS(net095), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net0104), .PLUS(net0110), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net095), .PLUS(net0158), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(wl_rd_sup), .PLUS(net0104), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(net080), .PLUS(net092), .BULK(gnd_));
rppolywo_m  R3 ( .MINUS(net092), .PLUS(net089), .BULK(gnd_));
rppolywo_m  R9 ( .MINUS(net083), .PLUS(net086), .BULK(gnd_));
rppolywo_m  R8 ( .MINUS(net086), .PLUS(net080), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(net077), .PLUS(net083), .BULK(gnd_));
rppolywo_m  R13 ( .MINUS(net0108), .PLUS(net0107), .BULK(gnd_));
rppolywo_m  R11 ( .MINUS(net071), .PLUS(net077), .BULK(gnd_));
rppolywo_m  R12 ( .MINUS(net0108), .PLUS(net071), .BULK(gnd_));
rppolywo_m  R15 ( .MINUS(net0113), .PLUS(wl_rd_sup), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net0110), .PLUS(net045), .BULK(gnd_));
rppolywo_m  R14 ( .MINUS(net0107), .PLUS(net0113), .BULK(gnd_));
nch_hvt  MN16 ( .D(wl_rd_sup), .B(gnd_), .G(act_rd_b), .S(gnd_));
nch_hvt  MN14 ( .D(net0158), .B(gnd_), .G(act_rd), .S(gnd_));
pch_hvt  MP13 ( .D(wl_rden_b), .B(vdd_), .G(net059), .S(vdd_));
pch_hvt  MP15 ( .D(net045), .B(vdd_), .G(act_rd_b), .S(vdd_));
inv_hvt I217 ( .A(wl_rden_b), .Y(net0142));
inv_hvt I220 ( .A(net0142), .Y(act_rd_b));
inv_hvt I180 ( .A(act_rd_b), .Y(act_rd));
tielo I223 ( .tielo(net059));

endmodule
// Library - xpmem, Cell - ml_rowdrv2, View - schematic
// LAST TIME SAVED: Jul 14 10:46:41 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_rowdrv2 ( pgate, reset, smc_rsr_out, vddctrl, wl, wl_rd_sup,
     wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
ml_dff I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile_last, View - schematic
// LAST TIME SAVED: Jan 24 11:25:01 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_rowdrv_tile_last ( pgate, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  reset;
output [15:0]  wl;
output [15:0]  vddctrl;
output [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  smc_rsr_out;



nor2_hvt I211 ( .A(smc_rsr_out[15]), .Y(net049), .B(smc_rsr_inc_out));
inv_hvt I215 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I216 ( .A(net041), .Y(por_rst_buf));
inv_hvt I217 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I391 ( .A(net049), .Y(smc_rsr_inc_last));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I213 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net079));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I214 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I212 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I190 ( .A(net079), .Y(smc_rsr_1st_out));
ml_rowdrv2_last Iml_rowdrv2_last ( .smc_rsr_inc(smc_rsr_inc_last),
     .smc_rsr_in(smc_rsr_out[14]), .rsr_rst(rsr_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_rst(cram_rst_buf),
     .smc_rsr_out(smc_rsr_out[15]), .reset(reset[15]), .wl(wl[15]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile, View - schematic
// LAST TIME SAVED: Jul 23 16:59:38 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_rowdrv_tile ( pgate, por_rst_out, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  por_rst_out, smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  vddctrl;
output [15:0]  pgate;
output [15:0]  wl;
output [15:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



inv_hvt I223 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I216 ( .A(cram_rst), .Y(net057));
inv_hvt I218 ( .A(net069), .Y(smc_write_buf));
inv_hvt I215 ( .A(cram_vddoff), .Y(net061));
inv_hvt I219 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I220 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I214 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I213 ( .A(smc_write), .Y(net069));
inv_hvt I221 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I212 ( .A(cram_wl_en), .Y(net055));
inv_hvt I217 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I190 ( .A(net037), .Y(smc_rsr_1st_out));
inv_hvt I211 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net037));
inv_hvt I210 ( .A(rsr_rst), .Y(net047));
inv_hvt I192 ( .A(por_rst), .Y(net041));
inv_hvt I222 ( .A(net041), .Y(por_rst_out));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I224 ( .A(net055), .Y(cram_wl_en_buf));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_15_ ( .reset(reset[15]), .wl(wl[15]),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[14]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[15]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_bank_ice1f, View - schematic
// LAST TIME SAVED: Mar  8 10:01:50 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_rowdrv_bank_ice1f ( jtag_rowtest_mode_b, last_rsr, pgate,
     reset, vddctrl, wl, banksel, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst,
     smc_rsr_inc, smc_write, trst_b );
output  jtag_rowtest_mode_b, last_rsr;

input  banksel, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst, smc_rsr_inc,
     smc_write, trst_b;

output [143:0]  reset;
output [143:0]  vddctrl;
output [143:0]  wl;
output [143:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  smc_rsr_1st_out_buf;

wire  [8:0]  smc_rsr_out;

wire  [7:0]  por_rst_out;

wire  [7:0]  smc_rsr_inc_out;

wire  [0:8]  smc_rsr_1st_out;



tielo I252 ( .tielo(net0130));
nand3_hvt I231 ( .Y(net186), .B(net190), .C(net190), .A(net190));
nand3_hvt I230 ( .Y(net190), .B(net195), .C(net195), .A(net195));
nand3_hvt I224 ( .B(net131), .Y(net195), .A(net131), .C(net131));
nand2_hvt I233 ( .A(smc_rsr_inc), .B(banksel), .Y(net181));
mux2_hvt I161 ( .in1(jtag_clk), .in0(net263), .out(net184),
     .sel(net256));
nor3_hvt I238 ( .B(por_rst), .Y(net248), .A(net208), .C(trst));
nor3_hvt I232 ( .C(rsr_rst), .A(jtag_rowtest_rst), .B(net0130),
     .Y(net213));
nor3_hvt I218 ( .B(net225), .Y(net215), .A(net225), .C(net225));
nor3_hvt I220 ( .B(net215), .Y(net219), .A(net215), .C(net215));
nor3_hvt I217 ( .C(net131), .A(net131), .B(net131), .Y(net225));
nor3_hvt I244 ( .B(por_rst), .Y(net227), .A(net276),
     .C(smc_rsr_1st_out_buf[0]));
nor2_hvt I239 ( .A(jtag_rowtest_rst), .B(net248), .Y(net208));
nor2_hvt I193 ( .A(por_rst), .B(rsr_set_1st), .Y(net252));
nor2_hvt I245 ( .A(rsr_set_1st), .B(net227), .Y(net276));
inv_hvt I247 ( .A(net256), .Y(jtag_rowtest_mode_b));
inv_hvt I241 ( .A(net208), .Y(net256));
inv_hvt I192 ( .A(net213), .Y(rsr_set_1st));
inv_hvt I234 ( .A(net181), .Y(net263));
inv_hvt I35 ( .A(net264), .Y(smc_rsr_1st_out_buf[0]));
inv_hvt I240 ( .A(trst_b), .Y(trst));
inv_hvt I210 ( .A(net268), .Y(last_rsr));
inv_hvt I391 ( .A(net252), .Y(rst_row_reg));
inv_hvt I36 ( .A(smc_rsr_1st_out[0]), .Y(net264));
inv_hvt I209 ( .A(smc_rsr_out[8]), .Y(net268));
inv_hvt I205 ( .A(net276), .Y(smc_rsr_in_1st));
tiehi I269 ( .tiehi(net162));
tiehi I249 ( .tiehi(net131));
tiehi I250 ( .tiehi(net132));
ml_buf_ice5_2 I227 ( .in(net131), .o(net134), .sel(net131));
ml_buf_ice5_2 I216 ( .in(net131), .o(net137), .sel(net131));
ml_buf_ice5_2 I198 ( .sel(banksel), .in(cram_wl_en),
     .o(cram_wl_en_buf));
ml_buf_ice5_2 I196 ( .sel(banksel), .in(cram_rst), .o(cram_rst_buf));
ml_buf_ice5_2 I199 ( .sel(net132), .in(por_rst), .o(por_rst_buf));
ml_buf_ice5_2 I197 ( .sel(banksel), .in(cram_vddoff),
     .o(cram_vddoff_buf));
ml_buf_ice5_2 I195 ( .sel(banksel), .in(cram_pgateoff),
     .o(cram_pgateoff_buf));
ml_buf_ice5_2 I201 ( .sel(banksel), .in(smc_write), .o(smc_write_buf));
ml_buf_ice5_2 I203 ( .sel(net184), .in(net184), .o(smc_rsr_inc_buf));
ml_buf_ice5_2 I213 ( .in(net162), .o(net161), .sel(net162));
ml_rowdrv_tile_last I_ml_rowdrv_tile_last (
     .smc_rsr_inc_out(smc_rsr_inc_out_last), .pgate(pgate[143:128]),
     .wl(wl[143:128]), .vddctrl(vddctrl[143:128]),
     .reset(reset[143:128]), .smc_rsr_1st_out(smc_rsr_1st_out[8]),
     .smcc_rsr_out(smc_rsr_out[8]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_buf), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[7]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf));
ml_rowdrv_tile I_ml_rowdrv_tile_7_ ( .por_rst_out(por_rst_out[7]),
     .smc_rsr_inc_out(smc_rsr_inc_out[7]),
     .smcc_rsr_out(smc_rsr_out[7]),
     .smc_rsr_1st_out(smc_rsr_1st_out[7]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out_last), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[6]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[127:112]), .vddctrl(vddctrl[127:112]),
     .reset(reset[127:112]), .pgate(pgate[127:112]));
ml_rowdrv_tile I_ml_rowdrv_tile_6_ ( .por_rst_out(por_rst_out[6]),
     .smc_rsr_inc_out(smc_rsr_inc_out[6]),
     .smcc_rsr_out(smc_rsr_out[6]),
     .smc_rsr_1st_out(smc_rsr_1st_out[6]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[7]), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[5]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[111:96]), .vddctrl(vddctrl[111:96]), .reset(reset[111:96]),
     .pgate(pgate[111:96]));
ml_rowdrv_tile I_ml_rowdrv_tile_5_ ( .por_rst_out(por_rst_out[5]),
     .smc_rsr_inc_out(smc_rsr_inc_out[5]),
     .smcc_rsr_out(smc_rsr_out[5]),
     .smc_rsr_1st_out(smc_rsr_1st_out[5]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[6]), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[4]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[95:80]), .vddctrl(vddctrl[95:80]), .reset(reset[95:80]),
     .pgate(pgate[95:80]));
ml_rowdrv_tile I_ml_rowdrv_tile_4_ ( .por_rst_out(por_rst_out[4]),
     .smc_rsr_inc_out(smc_rsr_inc_out[4]),
     .smcc_rsr_out(smc_rsr_out[4]),
     .smc_rsr_1st_out(smc_rsr_1st_out[4]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[5]), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[3]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[79:64]), .vddctrl(vddctrl[79:64]), .reset(reset[79:64]),
     .pgate(pgate[79:64]));
ml_rowdrv_tile I_ml_rowdrv_tile_3_ ( .por_rst_out(por_rst_out[3]),
     .smc_rsr_inc_out(smc_rsr_inc_out[3]),
     .smcc_rsr_out(smc_rsr_out[3]),
     .smc_rsr_1st_out(smc_rsr_1st_out[3]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[4]), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[2]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[63:48]), .vddctrl(vddctrl[63:48]), .reset(reset[63:48]),
     .pgate(pgate[63:48]));
ml_rowdrv_tile I_ml_rowdrv_tile_2_ ( .por_rst_out(por_rst_out[2]),
     .smc_rsr_inc_out(smc_rsr_inc_out[2]),
     .smcc_rsr_out(smc_rsr_out[2]),
     .smc_rsr_1st_out(smc_rsr_1st_out[2]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[3]), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[1]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[47:32]), .vddctrl(vddctrl[47:32]), .reset(reset[47:32]),
     .pgate(pgate[47:32]));
ml_rowdrv_tile I_ml_rowdrv_tile_1_ ( .por_rst_out(por_rst_out[1]),
     .smc_rsr_inc_out(smc_rsr_inc_out[1]),
     .smcc_rsr_out(smc_rsr_out[1]),
     .smc_rsr_1st_out(smc_rsr_1st_out[1]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[2]), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[0]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[31:16]), .vddctrl(vddctrl[31:16]), .reset(reset[31:16]),
     .pgate(pgate[31:16]));
ml_rowdrv_tile I_ml_rowdrv_tile_0_ ( .por_rst_out(por_rst_out[0]),
     .smc_rsr_inc_out(smc_rsr_inc_out[0]),
     .smcc_rsr_out(smc_rsr_out[0]),
     .smc_rsr_1st_out(smc_rsr_1st_out[0]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[1]), .smc_rsr_in(smc_rsr_in_1st),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[15:0]), .vddctrl(vddctrl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]));

endmodule
// Library - ice8chip, Cell - sg_dffbuf_modified, View - schematic
// LAST TIME SAVED: Aug 19 09:09:59 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module sg_dffbuf_modified ( dffout, clk, d, r );
output  dffout;

input  clk, d, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff I0 ( .R(r), .D(d), .CLK(clk), .QN(net9), .Q(net10));
sg_bufx10_ice8p I5 ( .in(net10), .out(dffout));

endmodule
// Library - leafcell, Cell - bram_sdo_reg, View - schematic
// LAST TIME SAVED: Jul  8 11:50:49 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_sdo_reg ( do, tielo, clk, di );
output  do, tielo;

input  clk, di;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff I_bm_sdo_dff ( .R(tielo), .D(di), .CLK(clk), .QN(net11),
     .Q(net018));
bram_bufferx16_2inv I51 ( .in(net018), .out(do));
tielo I_tielo ( .tielo(tielo));

endmodule
// Library - leafcell, Cell - bram_bufferx4, View - schematic
// LAST TIME SAVED: Aug 12 09:08:27 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module bram_bufferx4 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - ice1chip, Cell - CHIP_route_lft_ice1f, View - schematic
// LAST TIME SAVED: Apr 22 10:30:29 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module CHIP_route_lft_ice1f ( cm_banksel_bltld3_1_, cm_clk_bltld3,
     cm_sdi_u1d3, cm_sdo_u1d1, core_por_b_rowu1, cram_prec_bltld3,
     cram_pullup_bltld3, cram_write_bltld3, data_muxsel1_bltld3,
     data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     last_rsr, pgate_l, reset_l, smc_wdis_dclk_bltld3,
     smc_write_bltld3, vdd_cntl_l, wl_l, cm_banksel_blbld1,
     cm_banksel_blbld, cm_clk_blbld, cm_sdi_u1d, cm_sdo_u1,
     core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0 );
output  cm_banksel_bltld3_1_, cm_clk_bltld3, core_por_b_rowu1,
     cram_prec_bltld3, cram_pullup_bltld3, cram_write_bltld3,
     data_muxsel1_bltld3, data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     smc_wdis_dclk_bltld3, smc_write_bltld3;

input  cm_clk_blbld, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;

output [1:0]  cm_sdo_u1d1;
output [287:0]  reset_l;
output [287:0]  wl_l;
output [1:0]  cm_sdi_u1d3;
output [287:0]  vdd_cntl_l;
output [1:0]  last_rsr;
output [287:0]  pgate_l;

input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdi_u1d;
input [1:1]  cm_banksel_blbld;
input [0:0]  cm_banksel_blbld1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdi_u1d0;

wire  [0:1]  net299;

wire  [1:1]  cm_banksel_bltld;

wire  [1:0]  cm_sdo_u1d0;

wire  [1:0]  dff_out;



ml_rowdrv_bank_ice1f I_ml_rowdrv_bank1f_bot ( .wl(wl_l[143:0]),
     .pgate(pgate_l[143:0]), .reset(reset_l[143:0]),
     .vddctrl(vdd_cntl_l[143:0]), .trst_b(j_rst_bl0),
     .smc_write(smc_writel0),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu0_b),
     .last_rsr(last_rsr[0]), .banksel(cm_banksel_blbld1[0]),
     .cram_pgateoff(cram_pgateoffl0), .cram_rst(cram_rstl0),
     .cram_vddoff(cram_vddoffl0), .cram_wl_en(cram_wl_enl0),
     .jtag_clk(tck_padl0), .jtag_rowtest_rst(row_testl1),
     .por_rst(core_por_bbl0), .rsr_rst(smc_rsr_rstl0),
     .smc_rsr_inc(smc_row_incl0));
ml_rowdrv_bank_ice1f I_ml_rowdrv_bank1f_top ( .wl({wl_l[144],
     wl_l[145], wl_l[146], wl_l[147], wl_l[148], wl_l[149], wl_l[150],
     wl_l[151], wl_l[152], wl_l[153], wl_l[154], wl_l[155], wl_l[156],
     wl_l[157], wl_l[158], wl_l[159], wl_l[160], wl_l[161], wl_l[162],
     wl_l[163], wl_l[164], wl_l[165], wl_l[166], wl_l[167], wl_l[168],
     wl_l[169], wl_l[170], wl_l[171], wl_l[172], wl_l[173], wl_l[174],
     wl_l[175], wl_l[176], wl_l[177], wl_l[178], wl_l[179], wl_l[180],
     wl_l[181], wl_l[182], wl_l[183], wl_l[184], wl_l[185], wl_l[186],
     wl_l[187], wl_l[188], wl_l[189], wl_l[190], wl_l[191], wl_l[192],
     wl_l[193], wl_l[194], wl_l[195], wl_l[196], wl_l[197], wl_l[198],
     wl_l[199], wl_l[200], wl_l[201], wl_l[202], wl_l[203], wl_l[204],
     wl_l[205], wl_l[206], wl_l[207], wl_l[208], wl_l[209], wl_l[210],
     wl_l[211], wl_l[212], wl_l[213], wl_l[214], wl_l[215], wl_l[216],
     wl_l[217], wl_l[218], wl_l[219], wl_l[220], wl_l[221], wl_l[222],
     wl_l[223], wl_l[224], wl_l[225], wl_l[226], wl_l[227], wl_l[228],
     wl_l[229], wl_l[230], wl_l[231], wl_l[232], wl_l[233], wl_l[234],
     wl_l[235], wl_l[236], wl_l[237], wl_l[238], wl_l[239], wl_l[240],
     wl_l[241], wl_l[242], wl_l[243], wl_l[244], wl_l[245], wl_l[246],
     wl_l[247], wl_l[248], wl_l[249], wl_l[250], wl_l[251], wl_l[252],
     wl_l[253], wl_l[254], wl_l[255], wl_l[256], wl_l[257], wl_l[258],
     wl_l[259], wl_l[260], wl_l[261], wl_l[262], wl_l[263], wl_l[264],
     wl_l[265], wl_l[266], wl_l[267], wl_l[268], wl_l[269], wl_l[270],
     wl_l[271], wl_l[272], wl_l[273], wl_l[274], wl_l[275], wl_l[276],
     wl_l[277], wl_l[278], wl_l[279], wl_l[280], wl_l[281], wl_l[282],
     wl_l[283], wl_l[284], wl_l[285], wl_l[286], wl_l[287]}),
     .pgate({pgate_l[144], pgate_l[145], pgate_l[146], pgate_l[147],
     pgate_l[148], pgate_l[149], pgate_l[150], pgate_l[151],
     pgate_l[152], pgate_l[153], pgate_l[154], pgate_l[155],
     pgate_l[156], pgate_l[157], pgate_l[158], pgate_l[159],
     pgate_l[160], pgate_l[161], pgate_l[162], pgate_l[163],
     pgate_l[164], pgate_l[165], pgate_l[166], pgate_l[167],
     pgate_l[168], pgate_l[169], pgate_l[170], pgate_l[171],
     pgate_l[172], pgate_l[173], pgate_l[174], pgate_l[175],
     pgate_l[176], pgate_l[177], pgate_l[178], pgate_l[179],
     pgate_l[180], pgate_l[181], pgate_l[182], pgate_l[183],
     pgate_l[184], pgate_l[185], pgate_l[186], pgate_l[187],
     pgate_l[188], pgate_l[189], pgate_l[190], pgate_l[191],
     pgate_l[192], pgate_l[193], pgate_l[194], pgate_l[195],
     pgate_l[196], pgate_l[197], pgate_l[198], pgate_l[199],
     pgate_l[200], pgate_l[201], pgate_l[202], pgate_l[203],
     pgate_l[204], pgate_l[205], pgate_l[206], pgate_l[207],
     pgate_l[208], pgate_l[209], pgate_l[210], pgate_l[211],
     pgate_l[212], pgate_l[213], pgate_l[214], pgate_l[215],
     pgate_l[216], pgate_l[217], pgate_l[218], pgate_l[219],
     pgate_l[220], pgate_l[221], pgate_l[222], pgate_l[223],
     pgate_l[224], pgate_l[225], pgate_l[226], pgate_l[227],
     pgate_l[228], pgate_l[229], pgate_l[230], pgate_l[231],
     pgate_l[232], pgate_l[233], pgate_l[234], pgate_l[235],
     pgate_l[236], pgate_l[237], pgate_l[238], pgate_l[239],
     pgate_l[240], pgate_l[241], pgate_l[242], pgate_l[243],
     pgate_l[244], pgate_l[245], pgate_l[246], pgate_l[247],
     pgate_l[248], pgate_l[249], pgate_l[250], pgate_l[251],
     pgate_l[252], pgate_l[253], pgate_l[254], pgate_l[255],
     pgate_l[256], pgate_l[257], pgate_l[258], pgate_l[259],
     pgate_l[260], pgate_l[261], pgate_l[262], pgate_l[263],
     pgate_l[264], pgate_l[265], pgate_l[266], pgate_l[267],
     pgate_l[268], pgate_l[269], pgate_l[270], pgate_l[271],
     pgate_l[272], pgate_l[273], pgate_l[274], pgate_l[275],
     pgate_l[276], pgate_l[277], pgate_l[278], pgate_l[279],
     pgate_l[280], pgate_l[281], pgate_l[282], pgate_l[283],
     pgate_l[284], pgate_l[285], pgate_l[286], pgate_l[287]}),
     .reset({reset_l[144], reset_l[145], reset_l[146], reset_l[147],
     reset_l[148], reset_l[149], reset_l[150], reset_l[151],
     reset_l[152], reset_l[153], reset_l[154], reset_l[155],
     reset_l[156], reset_l[157], reset_l[158], reset_l[159],
     reset_l[160], reset_l[161], reset_l[162], reset_l[163],
     reset_l[164], reset_l[165], reset_l[166], reset_l[167],
     reset_l[168], reset_l[169], reset_l[170], reset_l[171],
     reset_l[172], reset_l[173], reset_l[174], reset_l[175],
     reset_l[176], reset_l[177], reset_l[178], reset_l[179],
     reset_l[180], reset_l[181], reset_l[182], reset_l[183],
     reset_l[184], reset_l[185], reset_l[186], reset_l[187],
     reset_l[188], reset_l[189], reset_l[190], reset_l[191],
     reset_l[192], reset_l[193], reset_l[194], reset_l[195],
     reset_l[196], reset_l[197], reset_l[198], reset_l[199],
     reset_l[200], reset_l[201], reset_l[202], reset_l[203],
     reset_l[204], reset_l[205], reset_l[206], reset_l[207],
     reset_l[208], reset_l[209], reset_l[210], reset_l[211],
     reset_l[212], reset_l[213], reset_l[214], reset_l[215],
     reset_l[216], reset_l[217], reset_l[218], reset_l[219],
     reset_l[220], reset_l[221], reset_l[222], reset_l[223],
     reset_l[224], reset_l[225], reset_l[226], reset_l[227],
     reset_l[228], reset_l[229], reset_l[230], reset_l[231],
     reset_l[232], reset_l[233], reset_l[234], reset_l[235],
     reset_l[236], reset_l[237], reset_l[238], reset_l[239],
     reset_l[240], reset_l[241], reset_l[242], reset_l[243],
     reset_l[244], reset_l[245], reset_l[246], reset_l[247],
     reset_l[248], reset_l[249], reset_l[250], reset_l[251],
     reset_l[252], reset_l[253], reset_l[254], reset_l[255],
     reset_l[256], reset_l[257], reset_l[258], reset_l[259],
     reset_l[260], reset_l[261], reset_l[262], reset_l[263],
     reset_l[264], reset_l[265], reset_l[266], reset_l[267],
     reset_l[268], reset_l[269], reset_l[270], reset_l[271],
     reset_l[272], reset_l[273], reset_l[274], reset_l[275],
     reset_l[276], reset_l[277], reset_l[278], reset_l[279],
     reset_l[280], reset_l[281], reset_l[282], reset_l[283],
     reset_l[284], reset_l[285], reset_l[286], reset_l[287]}),
     .vddctrl({vdd_cntl_l[144], vdd_cntl_l[145], vdd_cntl_l[146],
     vdd_cntl_l[147], vdd_cntl_l[148], vdd_cntl_l[149],
     vdd_cntl_l[150], vdd_cntl_l[151], vdd_cntl_l[152],
     vdd_cntl_l[153], vdd_cntl_l[154], vdd_cntl_l[155],
     vdd_cntl_l[156], vdd_cntl_l[157], vdd_cntl_l[158],
     vdd_cntl_l[159], vdd_cntl_l[160], vdd_cntl_l[161],
     vdd_cntl_l[162], vdd_cntl_l[163], vdd_cntl_l[164],
     vdd_cntl_l[165], vdd_cntl_l[166], vdd_cntl_l[167],
     vdd_cntl_l[168], vdd_cntl_l[169], vdd_cntl_l[170],
     vdd_cntl_l[171], vdd_cntl_l[172], vdd_cntl_l[173],
     vdd_cntl_l[174], vdd_cntl_l[175], vdd_cntl_l[176],
     vdd_cntl_l[177], vdd_cntl_l[178], vdd_cntl_l[179],
     vdd_cntl_l[180], vdd_cntl_l[181], vdd_cntl_l[182],
     vdd_cntl_l[183], vdd_cntl_l[184], vdd_cntl_l[185],
     vdd_cntl_l[186], vdd_cntl_l[187], vdd_cntl_l[188],
     vdd_cntl_l[189], vdd_cntl_l[190], vdd_cntl_l[191],
     vdd_cntl_l[192], vdd_cntl_l[193], vdd_cntl_l[194],
     vdd_cntl_l[195], vdd_cntl_l[196], vdd_cntl_l[197],
     vdd_cntl_l[198], vdd_cntl_l[199], vdd_cntl_l[200],
     vdd_cntl_l[201], vdd_cntl_l[202], vdd_cntl_l[203],
     vdd_cntl_l[204], vdd_cntl_l[205], vdd_cntl_l[206],
     vdd_cntl_l[207], vdd_cntl_l[208], vdd_cntl_l[209],
     vdd_cntl_l[210], vdd_cntl_l[211], vdd_cntl_l[212],
     vdd_cntl_l[213], vdd_cntl_l[214], vdd_cntl_l[215],
     vdd_cntl_l[216], vdd_cntl_l[217], vdd_cntl_l[218],
     vdd_cntl_l[219], vdd_cntl_l[220], vdd_cntl_l[221],
     vdd_cntl_l[222], vdd_cntl_l[223], vdd_cntl_l[224],
     vdd_cntl_l[225], vdd_cntl_l[226], vdd_cntl_l[227],
     vdd_cntl_l[228], vdd_cntl_l[229], vdd_cntl_l[230],
     vdd_cntl_l[231], vdd_cntl_l[232], vdd_cntl_l[233],
     vdd_cntl_l[234], vdd_cntl_l[235], vdd_cntl_l[236],
     vdd_cntl_l[237], vdd_cntl_l[238], vdd_cntl_l[239],
     vdd_cntl_l[240], vdd_cntl_l[241], vdd_cntl_l[242],
     vdd_cntl_l[243], vdd_cntl_l[244], vdd_cntl_l[245],
     vdd_cntl_l[246], vdd_cntl_l[247], vdd_cntl_l[248],
     vdd_cntl_l[249], vdd_cntl_l[250], vdd_cntl_l[251],
     vdd_cntl_l[252], vdd_cntl_l[253], vdd_cntl_l[254],
     vdd_cntl_l[255], vdd_cntl_l[256], vdd_cntl_l[257],
     vdd_cntl_l[258], vdd_cntl_l[259], vdd_cntl_l[260],
     vdd_cntl_l[261], vdd_cntl_l[262], vdd_cntl_l[263],
     vdd_cntl_l[264], vdd_cntl_l[265], vdd_cntl_l[266],
     vdd_cntl_l[267], vdd_cntl_l[268], vdd_cntl_l[269],
     vdd_cntl_l[270], vdd_cntl_l[271], vdd_cntl_l[272],
     vdd_cntl_l[273], vdd_cntl_l[274], vdd_cntl_l[275],
     vdd_cntl_l[276], vdd_cntl_l[277], vdd_cntl_l[278],
     vdd_cntl_l[279], vdd_cntl_l[280], vdd_cntl_l[281],
     vdd_cntl_l[282], vdd_cntl_l[283], vdd_cntl_l[284],
     vdd_cntl_l[285], vdd_cntl_l[286], vdd_cntl_l[287]}),
     .smc_write(smc_write_bltld3), .smc_rsr_inc(net303),
     .rsr_rst(net289), .por_rst(core_por_b_rowu1),
     .jtag_rowtest_rst(net345), .jtag_clk(net305), .cram_wl_en(net273),
     .cram_vddoff(net335), .cram_rst(net319), .cram_pgateoff(net295),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu1_b),
     .last_rsr(last_rsr[1]), .banksel(net231), .trst_b(net311));
tielo I74 ( .tielo(net219));
sg_bufx10_ice8p I28 ( .in(smc_writel0), .out(net221));
sg_bufx10_ice8p I35 ( .in(net291), .out(net223));
sg_bufx10_ice8p I45 ( .in(row_testl1), .out(net225));
sg_bufx10_ice8p I44 ( .in(net225), .out(net227));
sg_bufx10_ice8p I2 ( .in(cram_write_bltld), .out(net229));
sg_bufx10_ice8p I67 ( .in(cm_banksel_bltld[1]), .out(net231));
sg_bufx10_ice8p I39 ( .in(net237), .out(net233));
sg_bufx10_ice8p I4 ( .in(data_muxsel1_blbld),
     .out(data_muxsel1_bltld));
sg_bufx10_ice8p I40 ( .in(cram_wl_enl0), .out(net237));
sg_bufx10_ice8p I37 ( .in(cram_vddoffl0), .out(net239));
sg_bufx10_ice8p I22 ( .in(core_por_bbl0), .out(net241));
sg_bufx10_ice8p I5 ( .in(data_muxsel1_bltld), .out(net243));
sg_bufx10_ice8p I527 ( .in(net327), .out(en_8bconfig_b_bltld3));
sg_bufx10_ice8p I523 ( .in(net283), .out(data_muxsel_bltld3));
sg_bufx10_ice8p I524 ( .in(net243), .out(data_muxsel1_bltld3));
sg_bufx10_ice8p I526 ( .in(net343), .out(cram_prec_bltld3));
sg_bufx10_ice8p I33 ( .in(cram_rstl0), .out(net253));
sg_bufx10_ice8p I70_1_ ( .in(cm_sdo_u1[1]), .out(cm_sdo_u1d0[1]));
sg_bufx10_ice8p I70_0_ ( .in(cm_sdo_u1[0]), .out(cm_sdo_u1d0[0]));
sg_bufx10_ice8p I528 ( .in(net337), .out(smc_wdis_dclk_bltld3));
sg_bufx10_ice8p I18 ( .in(smc_rsr_rstl0), .out(net259));
sg_bufx10_ice8p I529 ( .in(net293), .out(cram_pullup_bltld3));
sg_bufx10_ice8p I3 ( .in(cram_write_blbld), .out(cram_write_bltld));
sg_bufx10_ice8p I532 ( .in(net363), .out(cm_clk_bltld3));
sg_bufx10_ice8p I79 ( .in(cm_clk_blbld), .out(cm_clk_bltld));
sg_bufx10_ice8p I8 ( .in(cram_pullup_blbld), .out(cram_pullup_bltld));
sg_bufx10_ice8p I7 ( .in(data_muxsel_blbld), .out(data_muxsel_bltld));
sg_bufx10_ice8p I554 ( .in(net233), .out(net273));
sg_bufx10_ice8p I27 ( .in(net221), .out(net275));
sg_bufx10_ice8p I25 ( .in(smc_row_incl0), .out(net277));
sg_bufx10_ice8p I47 ( .in(net357), .out(net279));
sg_bufx10_ice8p I68_1_ ( .in(cm_sdi_u1d[1]), .out(cm_sdi_u1d0[1]));
sg_bufx10_ice8p I68_0_ ( .in(cm_sdi_u1d[0]), .out(cm_sdi_u1d0[0]));
sg_bufx10_ice8p I6 ( .in(data_muxsel_bltld), .out(net283));
sg_bufx10_ice8p I38 ( .in(net239), .out(net285));
sg_bufx10_ice8p I19 ( .in(net259), .out(net287));
sg_bufx10_ice8p I546 ( .in(net287), .out(net289));
sg_bufx10_ice8p I36 ( .in(cram_pgateoffl0), .out(net291));
sg_bufx10_ice8p I9 ( .in(cram_pullup_bltld), .out(net293));
sg_bufx10_ice8p I547 ( .in(net223), .out(net295));
sg_bufx10_ice8p I552 ( .in(net275), .out(smc_write_bltld3));
sg_bufx10_ice8p I69_1_ ( .in(cm_sdi_u1d0[1]), .out(net299[0]));
sg_bufx10_ice8p I69_0_ ( .in(cm_sdi_u1d0[0]), .out(net299[1]));
sg_bufx10_ice8p I549 ( .in(net349), .out(net303));
sg_bufx10_ice8p I544 ( .in(net279), .out(net305));
sg_bufx10_ice8p I530_1_ ( .in(net299[0]), .out(cm_sdi_u1d3[1]));
sg_bufx10_ice8p I530_0_ ( .in(net299[1]), .out(cm_sdi_u1d3[0]));
sg_bufx10_ice8p I545 ( .in(net353), .out(net311));
sg_bufx10_ice8p I531 ( .in(net231), .out(cm_banksel_bltld3_1_));
sg_bufx10_ice8p I551 ( .in(net331), .out(net319));
sg_bufx10_ice8p I553 ( .in(net355), .out(core_por_b_rowu1));
sg_bufx10_ice8p I81 ( .in(cm_clk_bltld), .out(net363));
sg_bufx10_ice8p I15 ( .in(en_8bconfig_b_blbld),
     .out(en_8bconfig_b_bltld));
sg_bufx10_ice8p I14 ( .in(en_8bconfig_b_bltld), .out(net327));
sg_bufx10_ice8p I0 ( .in(cram_prec_blbld), .out(cram_prec_bltld));
sg_bufx10_ice8p I34 ( .in(net253), .out(net331));
sg_bufx10_ice8p I49 ( .in(j_rst_bl0), .out(net333));
sg_bufx10_ice8p I550 ( .in(net285), .out(net335));
sg_bufx10_ice8p I13 ( .in(smc_wdis_dclk_bltld), .out(net337));
sg_bufx10_ice8p I66 ( .in(cm_banksel_blbld[1]),
     .out(cm_banksel_bltld[1]));
sg_bufx10_ice8p I80_1_ ( .in(dff_out[1]), .out(cm_sdo_u1d1[1]));
sg_bufx10_ice8p I80_0_ ( .in(dff_out[0]), .out(cm_sdo_u1d1[0]));
sg_bufx10_ice8p I1 ( .in(cram_prec_bltld), .out(net343));
sg_bufx10_ice8p I548 ( .in(net227), .out(net345));
sg_bufx10_ice8p I525 ( .in(net229), .out(cram_write_bltld3));
sg_bufx10_ice8p I26 ( .in(net277), .out(net349));
sg_bufx10_ice8p I12 ( .in(smc_wdis_dclk_blbld),
     .out(smc_wdis_dclk_bltld));
sg_bufx10_ice8p I48 ( .in(net333), .out(net353));
sg_bufx10_ice8p I21 ( .in(net241), .out(net355));
sg_bufx10_ice8p I46 ( .in(tck_padl0), .out(net357));
sg_dffbuf_modified I73_1_ ( .d(cm_sdo_u1d0[1]), .clk(net363),
     .dffout(dff_out[1]), .r(net219));
sg_dffbuf_modified I73_0_ ( .d(cm_sdo_u1d0[0]), .clk(net363),
     .dffout(dff_out[0]), .r(net219));
sg_dffbuf_modified I77 ( .d(last_rsr[0]), .clk(net363),
     .dffout(last_rsr0), .r(net219));

endmodule
// Library - leafcell, Cell - creset_filter, View - schematic
// LAST TIME SAVED: Sep 30 15:04:05 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module creset_filter ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I11 ( .in(net042), .out(out));
nch_hvt  M0 ( .D(net13), .B(gnd_), .G(in), .S(gnd_));
nch_hvt  MN31 ( .D(net17), .B(gnd_), .G(net9), .S(gnd_));
rppolywo_m  R0 ( .MINUS(net17), .PLUS(pbias), .BULK(gnd_));
pch_hvt  M3 ( .D(net13), .B(vdd_), .G(net042), .S(vdd_));
pch_hvt  M2 ( .D(net13), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  M1 ( .D(vdd_), .B(vdd_), .G(net13), .S(vdd_));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(net9), .S(vdd_));
inv_hvt I6 ( .A(net13), .Y(net042));
inv_hvt I4 ( .A(in), .Y(net9));

endmodule
// Library - ice8chip, Cell - bram_bufferx16_ice8p, View - schematic
// LAST TIME SAVED: Aug  6 14:53:07 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module bram_bufferx16_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I5 ( .A(net07), .Y(net09));
inv_hvt I2 ( .A(in), .Y(net07));
inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(net09), .Y(net6));

endmodule
// Library - ice8chip, Cell - eh_io_pup_2_new_ice8p, View - schematic
// LAST TIME SAVED: Aug 25 11:50:10 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module eh_io_pup_2_new_ice8p ( por_b, core_por_b, vdd_io );
output  por_b;

input  core_por_b, vdd_io;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M8 ( .D(net104), .B(gnd_), .G(v_in), .S(net104));
nch_lvt  M23 ( .D(net104), .B(gnd_), .G(v_in), .S(net0196));
sg_bufx10_ice8p I_clkbuf ( .in(net84), .out(por_b));
nch_na25  M27 ( .D(net0224), .B(gnd_), .G(net0224), .S(net0132));
nch_na25  M24 ( .D(net0132), .B(gnd_), .G(net0132), .S(net0220));
nch_na25  M25 ( .D(net0220), .B(gnd_), .G(net0220), .S(net0216));
nch_na25  M9 ( .D(net158), .B(gnd_), .G(net158), .S(net154));
nch_na25  M13 ( .D(net150), .B(gnd_), .G(net150), .S(net162));
nch_na25  M16 ( .D(v_in), .B(gnd_), .G(net147), .S(net0195));
nch_na25  M20 ( .D(net162), .B(gnd_), .G(net162), .S(net0112));
nch_na25  M12 ( .D(net154), .B(gnd_), .G(net154), .S(net150));
nch_na25  M26 ( .D(net0216), .B(gnd_), .G(net0216), .S(gnd_));
nch_na25  M21 ( .D(net0112), .B(gnd_), .G(net0112), .S(gnd_));
rppolywo_m  R66 ( .MINUS(gnd_), .PLUS(net145), .BULK(gnd_));
nch_25  MN6 ( .D(net0195), .B(gnd_), .G(net145), .S(gnd_));
nch_25  M10 ( .D(net0195), .B(gnd_), .G(net147), .S(net158));
nch_25  M14 ( .D(v_in), .B(gnd_), .G(net147), .S(net0224));
nch_hvt  M22 ( .D(net104), .B(gnd_), .G(v_in), .S(net104));
nch_hvt  MN1 ( .D(net0196), .B(gnd_), .G(core_por_b), .S(gnd_));
nch_hvt  M2 ( .D(net84), .B(gnd_), .G(net104), .S(gnd_));
pch_hvt  M17 ( .D(net104), .B(vdd_), .G(v_in), .S(vdd_));
pch_hvt  MP8 ( .D(net104), .B(vdd_), .G(core_por_b), .S(vdd_));
pch_hvt  M0 ( .D(net84), .B(vdd_), .G(net104), .S(vdd_));
pch_25  M1 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
pch_25  M5 ( .D(net0195), .B(vdd_io), .G(net0195), .S(vdd_io));
pch_25  M3 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
pch_25  M7 ( .D(net0195), .B(vdd_io), .G(net145), .S(net0195));
pch_25  M6 ( .D(net0195), .B(vdd_io), .G(net0195), .S(vdd_io));
pch_25  M4 ( .D(net0195), .B(vdd_io), .G(net0195), .S(vdd_io));
vdd_tiehigh I96 ( .vdd_tieh(net147));

endmodule
// Library - ice8chip, Cell - eh_core_pup_2, View - schematic
// LAST TIME SAVED: Sep  7 10:17:18 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module eh_core_pup_2 ( por_b );
output  por_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I7 ( .A(out_1), .Y(out_2));
inv_hvt I9 ( .A(out_2), .Y(out_3));
inv_hvt I11 ( .A(out_3), .Y(por_b));
nch_hvt  M3 ( .D(gnd_), .B(gnd_), .G(out_2), .S(gnd_));
nch_hvt  M4 ( .D(gnd_), .B(gnd_), .G(net148), .S(gnd_));
nch_hvt  M0 ( .D(out_1), .B(gnd_), .G(net148), .S(gnd_));
nch_hvt  M5 ( .D(gnd_), .B(gnd_), .G(net148), .S(gnd_));
nch_hvt  M1 ( .D(out_1), .B(gnd_), .G(out_2), .S(gnd_));
rppolywo  R10 ( .MINUS(net130), .PLUS(net109));
rppolywo  R12 ( .MINUS(net154), .PLUS(net157));
rppolywo  R6 ( .MINUS(out_1), .PLUS(net124));
rppolywo  R9 ( .MINUS(net118), .PLUS(net130));
rppolywo  R15 ( .MINUS(net166), .PLUS(div_1));
rppolywo  R13 ( .MINUS(net157), .PLUS(net145));
rppolywo  R1 ( .MINUS(net068), .PLUS(net048));
rppolywo  R2 ( .MINUS(net067), .PLUS(net068));
rppolywo  R4 ( .MINUS(net142), .PLUS(net148));
rppolywo  R5 ( .MINUS(div_1), .PLUS(net142));
rppolywo  R41 ( .MINUS(net039), .PLUS(net042));
rppolywo  R40 ( .MINUS(net042), .PLUS(vdd_));
rppolywo  R11 ( .MINUS(net109), .PLUS(net154));
rppolywo  R0 ( .MINUS(net048), .PLUS(net039));
rppolywo  R8 ( .MINUS(net127), .PLUS(net118));
rppolywo  R14 ( .MINUS(net145), .PLUS(net166));
rppolywo  R3 ( .MINUS(net148), .PLUS(net067));
rppolywo  R7 ( .MINUS(net124), .PLUS(net127));

endmodule
// Library - ice8chip, Cell - SMC_CORE_POR_right_ice8p, View -
//schematic
// LAST TIME SAVED: Sep 29 09:25:02 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module SMC_CORE_POR_right_ice8p ( core_por_b0, core_por_bb, smc_por_b,
     creset_b, smc_core_por_bottom1, smc_core_por_bottom2,
     vddio_rightbank );
output  core_por_b0, core_por_bb, smc_por_b;

input  creset_b, smc_core_por_bottom1, smc_core_por_bottom2,
     vddio_rightbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



sg_bufx10_ice8p I500 ( .in(net032), .out(core_por_bb));
eh_io_pup_2_new_ice8p Ieh_io_pup_2_new_ice8p ( .core_por_b(net026),
     .vdd_io(vddio_rightbank), .por_b(net3));
eh_core_pup_2 Ieh_core_pup_2 ( .por_b(net026));
nand2_hvt I6 ( .A(net026), .Y(net021), .B(creset_b));
inv_hvt I11 ( .A(net04), .Y(smc_por_b));
inv_hvt I701 ( .A(core_por_b0), .Y(net032));
inv_hvt I7 ( .A(net021), .Y(core_por_b0));
nand4_hvt I2 ( .D(core_por_b0), .C(smc_core_por_bottom2), .A(net3),
     .Y(net04), .B(smc_core_por_bottom1));

endmodule
// Library - ice8chip, Cell - ml_cram_logic_ice8p, View - schematic
// LAST TIME SAVED: Oct 22 15:51:24 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_cram_logic_ice8p ( cram_pgateoff, cram_prec, cram_pullup_b,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, smc_clk_out, por,
     smc_clk, smc_read, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rwl_en, smc_seq_rst, smc_wcram_rst, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en );
output  cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, smc_clk_out;

input  por, smc_clk, smc_read, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_write, smc_wset_prec, smc_wset_precgnd, smc_wwlwrt_dis,
     smc_wwlwrt_en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C2 ( .MINUS(GND_), .PLUS(net326));
nmoscap_25  C1 ( .MINUS(GND_), .PLUS(net306));
nmoscap_25  C0 ( .MINUS(GND_), .PLUS(net314));
tielo I480 ( .tielo(net235));
sg_bufx10_ice8p I461 ( .in(net321), .out(cram_pullup_b));
sg_bufx10_ice8p I446 ( .in(net245), .out(cram_prec));
sg_bufx10_ice8p I457 ( .in(net234), .out(cram_wl_en));
sg_bufx10_ice8p I467 ( .in(net226), .out(cram_pgateoff));
sg_bufx10_ice8p I447 ( .in(cram_write_int), .out(cram_write));
sg_bufx10_ice8p I526 ( .in(net295), .out(cram_vddoff));
nand2_hvt I213 ( .A(net285), .Y(net222), .B(net311));
mux2_hvt I430 ( .in1(net407), .in0(net254), .out(net226),
     .sel(net235));
mux2_hvt I428 ( .in1(cram_write_int), .in0(net319), .out(net230),
     .sel(net285));
mux2_hvt I429 ( .in1(net254), .in0(net230), .out(net234),
     .sel(net235));
mux2_hvt I295 ( .in1(net255), .in0(net293), .out(net238),
     .sel(net285));
nor2_hvt I402 ( .A(net240), .B(smc_wset_precgnd), .Y(net242));
nor2_hvt I329 ( .A(net287), .B(smc_seq_rst), .Y(net245));
nor2_hvt I398 ( .A(smc_rpull_b), .B(net247), .Y(net248));
nor2_hvt I393 ( .A(set_wl_write), .B(reset_logic), .Y(net251));
nor2_hvt I364 ( .A(net426), .B(smc_seq_rst), .Y(net254));
nor2_hvt I400 ( .A(net255), .B(smc_wset_prec), .Y(net257));
nor2_hvt I366 ( .A(reset_logic), .B(net417), .Y(net260));
nor2_hvt I223 ( .A(net359), .B(por), .Y(net263));
nor2_hvt I390 ( .A(smc_write), .B(smc_seq_rst), .Y(net266));
nor2_hvt I392 ( .A(net240), .B(cram_rst), .Y(net269));
nor2_hvt I389 ( .A(net442), .B(reset_logic), .Y(net272));
nor2_hvt I385 ( .A(smc_rprec), .B(net274), .Y(net368));
nor2_hvt I414 ( .A(net276), .B(smc_wwlwrt_en), .Y(net278));
nor2_hvt I391 ( .A(cram_rst), .B(reset_logic), .Y(net281));
inv_hvt I458 ( .A(net272), .Y(rst_rpull_rwl));
inv_hvt I452 ( .A(net266), .Y(net285));
inv_hvt I451 ( .A(net238), .Y(net287));
inv_hvt I459 ( .A(smc_rwl_en), .Y(net289));
inv_hvt I373 ( .A(set_wl_write), .Y(net314));
inv_hvt I346 ( .A(net368), .Y(net293));
inv_hvt I464 ( .A(net222), .Y(net295));
inv_hvt I468 ( .A(net456), .Y(net297));
inv_hvt I454 ( .A(net260), .Y(dis_pgatewrt));
inv_hvt I403 ( .A(net242), .Y(net444));
inv_hvt I450 ( .A(net257), .Y(net303));
inv_hvt I448 ( .A(net281), .Y(net443));
inv_hvt I442 ( .A(net306), .Y(net307));
inv_hvt I444 ( .A(net315), .Y(net306));
inv_hvt I453 ( .A(net269), .Y(net311));
inv_hvt I445 ( .A(net307), .Y(net326));
inv_hvt I435 ( .A(net314), .Y(net315));
inv_hvt I4 ( .A(sm_clk_b), .Y(smc_clk_out));
inv_hvt I421 ( .A(net421), .Y(net319));
inv_hvt I462 ( .A(net247), .Y(net321));
inv_hvt I3 ( .A(smc_clk), .Y(sm_clk_b));
inv_hvt I449 ( .A(net251), .Y(net325));
inv_hvt I443 ( .A(net326), .Y(cram_write_int));
inv_hvt I465 ( .A(cram_rst_int_b), .Y(cram_rst));
inv_hvt I456 ( .A(net263), .Y(reset_logic));
inv_hvt I463 ( .A(net451), .Y(net247));
inv_hvt I460 ( .A(net248), .Y(net335));
inv_hvt I466 ( .A(net297), .Y(cram_rst_int_b));
inv_hvt I256 ( .A(net436), .Y(set_wl_write));
inv_hvt I455 ( .A(net278), .Y(net341));
nor3_hvt I472 ( .B(net347), .Y(net343), .A(net347), .C(net347));
nor3_hvt I471 ( .B(net351), .Y(net347), .A(net351), .C(net351));
nor3_hvt I470 ( .B(net363), .Y(net351), .A(net363), .C(net363));
nor3_hvt I217 ( .B(vdd_tieh), .Y(net355), .A(vdd_tieh), .C(vdd_tieh));
nor3_hvt I386 ( .B(smc_seq_rst), .Y(net359), .A(smc_write),
     .C(smc_read));
nor3_hvt I469 ( .B(net355), .Y(net363), .A(net355), .C(net355));
nor3_hvt I387 ( .B(smc_rwl_en), .Y(net274), .A(net368),
     .C(reset_logic));
nand3_hvt I476 ( .Y(net370), .B(net386), .C(net386), .A(net386));
nand3_hvt I477 ( .Y(net374), .B(net370), .C(net370), .A(net370));
nand3_hvt I478 ( .Y(net378), .B(net374), .C(net374), .A(net374));
nand3_hvt I479 ( .Y(net382), .B(net378), .C(net378), .A(net378));
nand3_hvt I426 ( .Y(net386), .B(vdd_tieh), .C(vdd_tieh), .A(vdd_tieh));
ml_dff I432 ( .R(dis_pgatewrt), .D(net412), .CLK(smc_clk_out),
     .QN(net406), .Q(net407));
ml_dff I431 ( .R(dis_pgatewrt), .D(net254), .CLK(sm_clk_b),
     .QN(net411), .Q(net412));
ml_dff I411 ( .R(reset_logic), .D(smc_wwlwrt_dis), .CLK(smc_clk),
     .QN(net416), .Q(net417));
ml_dff I408 ( .R(rst_rpull_rwl), .D(vdd_tieh), .CLK(net289),
     .QN(net421), .Q(net400));
ml_dff I405 ( .R(dis_pgatewrt), .D(vdd_tieh), .CLK(set_wl_write),
     .QN(net426), .Q(net399));
ml_dff I412 ( .R(net325), .D(net303), .CLK(smc_clk_out), .QN(net394),
     .Q(net255));
ml_dff I410 ( .R(dis_pgatewrt), .D(net341), .CLK(smc_clk_out),
     .QN(net436), .Q(net276));
ml_dff I108 ( .R(reset_logic), .D(smc_rrst_pullwlen),
     .CLK(smc_clk_out), .QN(net402), .Q(net442));
ml_dff I413 ( .R(net443), .D(net444), .CLK(smc_clk_out), .QN(net446),
     .Q(net240));
ml_dff I407 ( .R(rst_rpull_rwl), .D(net335), .CLK(smc_clk_out),
     .QN(net451), .Q(net397));
ml_dff I406 ( .R(reset_logic), .D(smc_wcram_rst), .CLK(smc_clk_out),
     .QN(net456), .Q(net457));
tiehi I427 ( .tiehi(vdd_tieh));

endmodule
// Library - xpmem, Cell - ml_dff_osc, View - schematic
// LAST TIME SAVED: Oct  7 11:47:56 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_dff_osc ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - misc, Cell - ml_mux3_hvt, View - schematic
// LAST TIME SAVED: May 13 15:14:37 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_mux3_hvt ( out, in0, in1, in2, sel );
output  out;

input  in0, in1, in2;

input [3:0]  sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I21 ( .A(sel[0]), .Y(net30));
inv_hvt I24 ( .A(sel[1]), .Y(net28));
inv_hvt I25 ( .A(sel[2]), .Y(net26));
txgate_hvt I23 ( .in(in1), .out(out), .pp(net28), .nn(sel[1]));
txgate_hvt I20 ( .in(in0), .out(out), .pp(net30), .nn(sel[0]));
txgate_hvt I26 ( .in(in2), .out(out), .pp(net26), .nn(sel[2]));
nch_hvt  MN19 ( .D(out), .B(gnd_), .G(sel[3]), .S(gnd_));

endmodule
// Library - misc, Cell - ml_osc_stage, View - schematic
// LAST TIME SAVED: Sep 30 16:59:25 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_osc_stage ( out, clkin, oscen_b, pbias, sel_trim );
output  out;

input  clkin, oscen_b, pbias;

input [3:0]  sel_trim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C5 ( .MINUS(gnd_), .PLUS(loadbot_0));
nmoscap_25  C6 ( .MINUS(gnd_), .PLUS(loadbot_1));
nmoscap_25  C4 ( .MINUS(gnd_), .PLUS(loadbot_2));
nch_hvt  MN41 ( .D(loadbot_0), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN39 ( .D(loadbot_2), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN29 ( .D(out), .B(gnd_), .G(in_bot), .S(gnd_));
nch_hvt  MN42 ( .D(loadbot_1), .B(gnd_), .G(net419), .S(gnd_));
pch_hvt  M3 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net456));
pch_hvt  M2 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net452));
pch_hvt  MP30 ( .D(net452), .B(vdd_), .G(oscen_b), .S(vdd_));
pch_hvt  MP72 ( .D(net456), .B(vdd_), .G(sel_trim[2]), .S(net452));
pch_hvt  MP33 ( .D(out), .B(vdd_), .G(in_bot), .S(vdd_));
inv_hvt I229 ( .A(net403), .Y(net419));
nor2_hvt I228 ( .A(clkin), .B(oscen_b), .Y(net403));
ml_mux3_hvt Iml_mux3_hvt_bot ( .in1(loadbot_1), .in0(loadbot_0),
     .out(in_bot), .sel(sel_trim[3:0]), .in2(loadbot_2));

endmodule
// Library - ice8chip, Cell - clk_mux_2to1_ice8p, View - schematic
// LAST TIME SAVED: Nov  5 16:41:18 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module clk_mux_2to1_ice8p ( clk, cbit, cbitb, min, prog );
output  clk;

input  cbit, cbitb, prog;

input [1:0]  min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I_inv0 ( .A(prog), .Y(net030));
nand2_lvt I_nand2_1 ( .A(st2), .Y(clkb), .B(net030));
inv_lvt I_inv2 ( .A(clkb), .Y(clk));
txgate_lvt I_txgate_hvt0 ( .in(min[0]), .out(st2), .pp(cbit),
     .nn(cbitb));
txgate_lvt I_txgate_hvt1 ( .in(min[1]), .out(st2), .pp(cbitb),
     .nn(cbit));

endmodule
// Library - misc, Cell - ml_osc_logic, View - schematic
// LAST TIME SAVED: Oct  7 11:48:52 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_osc_logic ( sel_trim, clkin, smc_osc_fsel, smc_oscen );

input  clkin, smc_oscen;

output [3:0]  sel_trim;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:2]  in_sel;



ml_dff_osc I174 ( .R(reset_ff), .D(net050), .CLK(clkin_buf_b),
     .QN(net150), .Q(net172));
ml_dff_osc I238 ( .R(reset_ff), .D(net050), .CLK(clkin_buf),
     .QN(net154), .Q(net177));
ml_dff_osc I244 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf),
     .QN(net155), .Q(net182));
ml_dff_osc I245 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf_b),
     .QN(net153), .Q(net187));
ml_dff_osc I242 ( .R(reset_ff), .D(net048), .CLK(clkin_buf_b),
     .QN(net191), .Q(net192));
ml_dff_osc I243 ( .R(reset_ff), .D(net048), .CLK(clkin_buf),
     .QN(net152), .Q(net197));
nor2_hvt I256 ( .A(smc_osc_fsel[1]), .B(smc_osc_fsel[0]),
     .Y(in_sel[2]));
inv_hvt I293 ( .A(net197), .Y(net052));
inv_hvt I263 ( .A(clkin_buf), .Y(net065));
inv_hvt I283 ( .A(clkin_buf_b), .Y(clkin_buf));
inv_hvt I284 ( .A(smc_oscen), .Y(reset_ff));
inv_hvt I282 ( .A(clkin), .Y(clkin_buf_b));
inv_hvt I255 ( .A(smc_osc_fsel[1]), .Y(in_sel[1]));
inv_hvt I294 ( .A(net192), .Y(net054));
inv_hvt I295 ( .A(net177), .Y(net057));
inv_hvt I296 ( .A(net172), .Y(net061));
inv_hvt I261 ( .A(in_sel[2]), .Y(net050));
inv_hvt I262 ( .A(in_sel[1]), .Y(net048));
inv_hvt I299 ( .A(net059), .Y(net0143));
inv_hvt I297 ( .A(net065), .Y(net063));
inv_hvt I302 ( .A(net094), .Y(net096));
inv_hvt I298 ( .A(net063), .Y(net059));
inv_hvt I304 ( .A(net0143), .Y(net092));
inv_hvt I303 ( .A(net092), .Y(net094));
inv_hvt I301 ( .A(net096), .Y(clkin_buf_delay));
inv_hvt I285 ( .A(net058), .Y(sel_trim[3]));
tiehis I281 ( .tiehi(net058));
ml_mux2_hvt I279 ( .in1(net182), .in0(net187), .out(sel_trim[0]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I277 ( .in1(net057), .in0(net061), .out(sel_trim[2]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I278 ( .in1(net052), .in0(net054), .out(sel_trim[1]),
     .sel(clkin_buf_delay));

endmodule
// Library - misc, Cell - ml_osc, View - schematic
// LAST TIME SAVED: Oct  7 11:48:19 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_osc ( clk_out, smc_osc_fsel, smc_oscen );
output  clk_out;

input  smc_oscen;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sel_trim;



ml_dff_osc I174 ( .R(oscen_b), .D(clkby2_b), .CLK(clk_dffin),
     .QN(clkby2_b), .Q(clkby2));
ml_dff_osc I279 ( .R(oscen_b), .D(net063), .CLK(net0115), .QN(net063),
     .Q(net066));
rppolywo_m  R18 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net437), .PLUS(net383), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R3 ( .MINUS(net366), .PLUS(net076), .BULK(gnd_));
rppolywo_m  R2 ( .MINUS(net383), .PLUS(net366), .BULK(gnd_));
rppolywo_m  R5 ( .MINUS(net070), .PLUS(pbias), .BULK(gnd_));
rppolywo_m  R4 ( .MINUS(net076), .PLUS(net070), .BULK(gnd_));
nch_hvt  MN31 ( .D(net437), .B(gnd_), .G(smc_oscen), .S(gnd_));
pch_hvt  M0 ( .D(net0101), .B(vdd_), .G(oscen_b), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(net0101));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(smc_oscen), .S(vdd_));
nand2_hvt I175 ( .A(out_bot), .Y(clk_dffin), .B(out_top));
inv_hvt I280 ( .A(clkby2), .Y(net0115));
inv_hvt I222 ( .A(clkby2), .Y(clkby2_b_buf));
inv_hvt I220 ( .A(clkby2_b), .Y(clkby2_buf));
inv_hvt I176 ( .A(net063), .Y(clk_out));
inv_hvt I198 ( .A(smc_oscen), .Y(oscen_b));
ml_osc_stage Istage_bot ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_b_buf), .out(out_bot), .sel_trim(sel_trim[3:0]));
ml_osc_stage Istage_top ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_buf), .out(out_top), .sel_trim(sel_trim[3:0]));
ml_osc_logic Iosc_logic ( .sel_trim(sel_trim[3:0]),
     .smc_oscen(smc_oscen), .smc_osc_fsel(smc_osc_fsel[1:0]),
     .clkin(clk_out));

endmodule
// Library - misc, Cell - ml_osc_top, View - schematic
// LAST TIME SAVED: Oct 13 10:43:19 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_osc_top ( cnt_podt_out, smc_clk, crst_b, por_b, smc_osc_fsel,
     smc_oscoff_b, smc_podt_off, smc_podt_rst );
output  cnt_podt_out, smc_clk;

input  crst_b, por_b, smc_oscoff_b, smc_podt_off, smc_podt_rst;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  q_b;

wire  [10:0]  q;



ml_dff_osc I230 ( .R(cnt_rst), .D(net076), .CLK(q_b[10]), .QN(net067),
     .Q(net063));
ml_dff_osc I243 ( .R(rst_off_latch), .D(net0174), .CLK(clk_out_b),
     .QN(smc_off_b), .Q(net0152));
ml_dff_osc I228_10_ ( .R(cnt_rst), .D(q_b[10]), .CLK(q[9]),
     .QN(q_b[10]), .Q(q[10]));
ml_dff_osc I228_9_ ( .R(cnt_rst), .D(q_b[9]), .CLK(q[8]), .QN(q_b[9]),
     .Q(q[9]));
ml_dff_osc I228_8_ ( .R(cnt_rst), .D(q_b[8]), .CLK(q[7]), .QN(q_b[8]),
     .Q(q[8]));
ml_dff_osc I228_7_ ( .R(cnt_rst), .D(q_b[7]), .CLK(q[6]), .QN(q_b[7]),
     .Q(q[7]));
ml_dff_osc I228_6_ ( .R(cnt_rst), .D(q_b[6]), .CLK(q[5]), .QN(q_b[6]),
     .Q(q[6]));
ml_dff_osc I228_5_ ( .R(cnt_rst), .D(q_b[5]), .CLK(q[4]), .QN(q_b[5]),
     .Q(q[5]));
ml_dff_osc I228_4_ ( .R(cnt_rst), .D(q_b[4]), .CLK(q[3]), .QN(q_b[4]),
     .Q(q[4]));
ml_dff_osc I228_3_ ( .R(cnt_rst), .D(q_b[3]), .CLK(q[2]), .QN(q_b[3]),
     .Q(q[3]));
ml_dff_osc I228_2_ ( .R(cnt_rst), .D(q_b[2]), .CLK(q[1]), .QN(q_b[2]),
     .Q(q[2]));
ml_dff_osc I228_1_ ( .R(cnt_rst), .D(q_b[1]), .CLK(q[0]), .QN(q_b[1]),
     .Q(q[1]));
ml_dff_osc I228_0_ ( .R(cnt_rst), .D(q_b[0]), .CLK(clk_in),
     .QN(q_b[0]), .Q(q[0]));
nand2_hvt I227 ( .A(smc_off_b), .B(rst_osc_b), .Y(disable_osc));
nand2_hvt I270 ( .A(crst_b), .Y(net064), .B(por_b));
inv_hvt I233 ( .A(clk_out), .Y(clk_out_b));
inv_hvt I271 ( .A(net064), .Y(rst_osc_b));
inv_hvt I267 ( .A(net078), .Y(clk_in));
inv_hvt I262 ( .A(net067), .Y(cnt_podt_out));
inv_hvt I275 ( .A(smc_oscoff_b), .Y(net0174));
inv_hvt I277 ( .A(net054), .Y(cnt_rst));
inv_hvt I229 ( .A(rst_osc_b), .Y(net090));
inv_hvt I253 ( .A(net0124), .Y(rst_off_latch));
inv_hvt I232 ( .A(clk_out_b), .Y(smc_clk));
nor2_hvt I272 ( .A(net066), .B(disable_osc), .Y(smc_oscen));
nor2_hvt I266 ( .A(clk_out), .B(smc_podt_off), .Y(net078));
nor2_hvt I273 ( .A(smc_oscoff_b), .B(rst_osc_b), .Y(net066));
nor2_hvt I276 ( .A(net090), .B(smc_podt_rst), .Y(net054));
nor2_hvt I274 ( .A(smc_oscoff_b), .B(cnt_rst), .Y(net0124));
tiehis I179 ( .tiehi(net076));
ml_osc Iml_osc ( .smc_osc_fsel(smc_osc_fsel[1:0]), .clk_out(clk_out),
     .smc_oscen(smc_oscen));

endmodule
// Library - ice1chip, Cell - CHIP_route_lft2rgt_ice1f_june, View -
//schematic
// LAST TIME SAVED: Jun 29 09:58:31 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module CHIP_route_lft2rgt_ice1f_june ( bm_banksel_i[3:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa[7:0], bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i[3:0], bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0,
     cdone_out, ceb0, cm_banksel_blbrd_2_, cm_banksel_bldld[1:0],
     cm_banksel_bltrd1_3_, cm_clk_blbrd, cm_clk_bltrd1, cm_sdi_u0[1:0],
     cm_sdi_u1[1:0], cm_sdi_u2d[1:0], cm_sdi_u3d2[1:0], core_por_b0,
     core_por_b1, core_por_b_rowu3, core_por_bb, cram_pgateoff,
     cram_prec, cram_prec_bltrd1, cram_pullup_b, cram_pullup_b_bltrd1,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, cram_write_bltrd1,
     data_muxsel1_blbrd, data_muxsel1_bltrd1, data_muxsel_blbrd,
     data_muxsel_bltrd1, en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1,
     end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     last_rsr[1:0], md_spi_b, mode0, mux_jtag_sel, nvcm_spi_sdi,
     nvcm_spi_ss_b, pgate_r[287:0], reset_b_r[287:0], row_test0, rst_b,
     sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1,
     smc_write0, smc_write_bltl1d1, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, update0, vdd_cntl_r[287:0], wl_r[287:0],
     bm_sdo_o[3:0], bp0, cdone_in, cm_sdo_u0d1[1:0], cm_sdo_u1d3[1:0],
     cm_sdo_u2d1[1:0], cm_sdo_u3[1:0], creset_b_int, fabric_out_12_00,
     fabric_out_13_01, fabric_out_13_02, fromsdo,
     idcode_msb20bits[19:0], last_rsr3, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, spi_ss_in_bbank[4:0],
     tck_pad, tdi_pad, tms_pad, trstb_pad, vddio_rightbank );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bltrd1_3_, cm_clk_blbrd,
     cm_clk_bltrd1, core_por_b0, core_por_b1, core_por_b_rowu3,
     core_por_bb, cram_pgateoff, cram_prec, cram_prec_bltrd1,
     cram_pullup_b, cram_pullup_b_bltrd1, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, cram_write_bltrd1, data_muxsel1_blbrd,
     data_muxsel1_bltrd1, data_muxsel_blbrd, data_muxsel_bltrd1,
     en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1, end_of_startup,
     gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, mux_jtag_sel, nvcm_spi_sdi, nvcm_spi_ss_b, row_test0,
     rst_b, sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1,
     smc_write0, smc_write_bltl1d1, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, update0;

input  bp0, cdone_in, creset_b_int, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fromsdo, last_rsr3, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, tck_pad, tdi_pad,
     tms_pad, trstb_pad, vddio_rightbank;

output [287:0]  vdd_cntl_r;
output [1:0]  cm_banksel_bldld;
output [287:0]  reset_b_r;
output [3:0]  bm_sdi_i;
output [287:0]  pgate_r;
output [1:0]  cm_sdi_u2d;
output [1:0]  last_rsr;
output [10:0]  bm_sa;
output [1:0]  cm_sdi_u0;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_sdi_u3d2;
output [287:0]  wl_r;
output [3:0]  bm_banksel_i;

input [1:0]  cm_sdo_u3;
input [1:0]  cm_sdo_u1d3;
input [1:0]  cm_sdo_u2d1;
input [19:0]  idcode_msb20bits;
input [1:0]  cm_sdo_u0d1;
input [3:0]  bm_sdo_o;
input [4:0]  spi_ss_in_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net350;

wire  [1:0]  cdsbus0;

wire  [1:0]  smc_osco_fsel;

wire  [3:0]  cm_banksel;

wire  [1:0]  dff_out_top;

wire  [0:1]  net332;

wire  [0:6]  net0409;

wire  [0:1]  net336;

wire  [0:1]  net447;

wire  [0:1]  net448;

wire  [0:1]  net354;

wire  [0:1]  net334;

wire  [0:1]  net446;

wire  [0:1]  net346;



smc_and_jtag_ice8p I_smc_and_jtag_ice8p ( .bm_sa(bm_sa[10:0]),
     .warmboot_sel({fabric_out_13_02, fabric_out_13_01}),
     .trst_pad(trstb_pad), .tms_pad(tms_pad), .tdi_pad(tdi_pad),
     .tck_pad(tck_pad), .spi_ss_in_b(spi_ss_in_bbank[4]),
     .cdone_in(cdone_in), .spi_sdi(spi_ss_in_bbank[2]),
     .spi_clk_in(spi_ss_in_bbank[3]), .psdi({net497, net497, net497,
     net497, net497, net497, net497}), .por_b(smc_por_b0),
     .osc_clk(osc_clk), .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .idcode_msb20bits(idcode_msb20bits[19:0]),
     .creset_b(crst_filterout), .coldboot_sel(spi_ss_in_bbank[1:0]),
     .cnt_podt_out(cnt_podt_out), .cm_sdo_u3(dff_out_top[1:0]),
     .cm_sdo_u2(cm_sdo_u2d1[1:0]), .cm_sdo_u1(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0(cm_sdo_u0d1[1:0]), .cm_monitor_cell({net497, net497,
     net497, net497}), .cm_last_rsr(last_rsr3), .bschain_sdo(fromsdo),
     .bp0(bp0), .boot(fabric_out_12_00), .bm_bank_sdo(bm_sdo_o[3:0]),
     .tdo_pad(totdopad), .tdo_oe_pad(sdo_enable),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out),
     .smc_wwlwrt_en(smc_wwlwrt_en), .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wdis_dclk(smc_wdis_dclk_blbrd),
     .smc_wcram_rst(smc_wcram_rst), .smc_seq_rst(smc_seq_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rsr_rst(smc_rsr_rst),
     .smc_rrst_pullwlen(smc_rrst_pullwlen), .smc_rpull_b(smc_rpull_b),
     .smc_rprec(smc_rprec), .smc_row_inc(smc_row_inc),
     .smc_read(smc_read), .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .psdo(net0409[0:6]), .nvcm_spi_ss_b(nvcm_spi_ss_b),
     .nvcm_spi_sdi(nvcm_spi_sdi), .md_spi_b(md_spi_b),
     .j_upd_dr(update0), .j_tdi(j_tdi), .j_tck(j_tck),
     .j_shift0(shift0), .j_sft_dr(shiftromsmc), .j_rst_b(j_rst_b),
     .j_row_test(row_test0), .j_mode(mode0), .j_hiz_b(hiz_b0),
     .j_ceb0(ceb0), .gsr(net439), .gint_hz(net440),
     .end_of_startup(net441), .en_8bconfig_b(en_8bconfig_b_blbrd),
     .data_muxsel1(data_muxsel1_blbrd),
     .data_muxsel(data_muxsel_blbrd), .cm_sdi_u3(cdsbus0[1:0]),
     .cm_sdi_u2(net446[0:1]), .cm_sdi_u1(net447[0:1]),
     .cm_sdi_u0(net448[0:1]), .cm_clk(cm_clk),
     .cm_banksel(cm_banksel[3:0]), .cdone_out(cdone_out),
     .bs_en(bs_en0), .bm_wdummymux_en(bm_wdummymux_en_i),
     .bm_sweb(bm_sweb_i), .bm_sreb(bm_sreb_i), .bm_sclkrw(bm_sclkrw_i),
     .bm_rcapmux_en(bm_rcapmux_en_i), .bm_init(bm_init_i),
     .bm_clk(bm_sclk_i), .bm_banksel(bm_banksel_i[3:0]),
     .bm_bank_sdi(bm_sdi_i[3:0]));
CHIP_route_lft_ice1f I_chip_route_lft2rgt_ice1f (
     .pgate_l(pgate_r[287:0]), .reset_l(reset_b_r[287:0]),
     .vdd_cntl_l(vdd_cntl_r[287:0]), .wl_l(wl_r[287:0]),
     .tck_padl0(j_tck), .smc_writel0(smc_write0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbrd),
     .smc_rsr_rstl0(smc_rsr_rst), .smc_row_incl0(smc_row_inc),
     .row_testl1(row_test0), .j_rst_bl0(j_rst_b),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbrd),
     .data_muxsel_blbld(data_muxsel_blbrd),
     .data_muxsel1_blbld(data_muxsel1_blbrd),
     .cram_write_blbld(cram_write), .cram_wl_enl0(cram_wl_en),
     .cram_vddoffl0(cram_vddoff), .cram_rstl0(cram_rst),
     .cram_pullup_blbld(cram_pullup_b), .cram_prec_blbld(cram_prec),
     .cram_pgateoffl0(cram_pgateoff), .core_por_bbl0(core_por_bb),
     .cm_sdo_u1(cm_sdo_u3[1:0]), .cm_sdi_u1d(cdsbus0[1:0]),
     .cm_clk_blbld(cm_clk_blbrd), .cm_banksel_blbld(cm_banksel[3]),
     .cm_banksel_blbld1(cm_banksel_blbrd_2_),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltrd1),
     .last_rsr(last_rsr[1:0]), .last_rsr0(net485),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu2_b),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltrd1),
     .data_muxsel1_bltld3(data_muxsel1_bltrd1),
     .cram_write_bltld3(cram_write_bltrd1),
     .cram_pullup_bltld3(cram_pullup_b_bltrd1),
     .cram_prec_bltld3(cram_prec_bltrd1),
     .core_por_b_rowu1(core_por_b_rowu3),
     .smc_write_bltld3(smc_write_bltl1d1),
     .cm_sdo_u1d1(dff_out_top[1:0]), .cm_sdi_u1d3(cm_sdi_u3d2[1:0]),
     .cm_clk_bltld3(cm_clk_bltrd1),
     .cm_banksel_bltld3_1_(cm_banksel_bltrd1_3_));
creset_filter I561 ( .in(creset_b_int), .out(crst_filterout));
bram_bufferx16_ice8p I702 ( .in(core_por_b0), .out(core_por_b1));
sg_bufx10_ice8p I558 ( .in(net441), .out(end_of_startup));
sg_bufx10_ice8p I559 ( .in(net439), .out(gsr));
sg_bufx10_ice8p I560 ( .in(net440), .out(gint_hz));
sg_bufx10_ice8p I550_1_ ( .in(net346[0]), .out(net332[0]));
sg_bufx10_ice8p I550_0_ ( .in(net346[1]), .out(net332[1]));
sg_bufx10_ice8p I476_1_ ( .in(net350[0]), .out(net334[0]));
sg_bufx10_ice8p I476_0_ ( .in(net350[1]), .out(net334[1]));
sg_bufx10_ice8p I478_1_ ( .in(net354[0]), .out(net336[0]));
sg_bufx10_ice8p I478_0_ ( .in(net354[1]), .out(net336[1]));
sg_bufx10_ice8p I479_1_ ( .in(net334[0]), .out(cm_sdi_u0[1]));
sg_bufx10_ice8p I479_0_ ( .in(net334[1]), .out(cm_sdi_u0[0]));
sg_bufx10_ice8p I480_1_ ( .in(net336[0]), .out(cm_sdi_u2d[1]));
sg_bufx10_ice8p I480_0_ ( .in(net336[1]), .out(cm_sdi_u2d[0]));
sg_bufx10_ice8p I481_1_ ( .in(net332[0]), .out(cm_sdi_u1[1]));
sg_bufx10_ice8p I481_0_ ( .in(net332[1]), .out(cm_sdi_u1[0]));
sg_bufx10_ice8p I551 ( .in(en_8bconfig_b_blbrd), .out(net0327));
sg_bufx10_ice8p I722_1_ ( .in(net447[0]), .out(net346[0]));
sg_bufx10_ice8p I722_0_ ( .in(net447[1]), .out(net346[1]));
sg_bufx10_ice8p I683_1_ ( .in(cm_banksel[1]),
     .out(cm_banksel_bldld[1]));
sg_bufx10_ice8p I683_0_ ( .in(cm_banksel[0]),
     .out(cm_banksel_bldld[0]));
sg_bufx10_ice8p I664_1_ ( .in(net448[0]), .out(net350[0]));
sg_bufx10_ice8p I664_0_ ( .in(net448[1]), .out(net350[1]));
sg_bufx10_ice8p I681 ( .in(cm_banksel[2]), .out(cm_banksel_blbrd_2_));
sg_bufx10_ice8p I723_1_ ( .in(net446[0]), .out(net354[0]));
sg_bufx10_ice8p I723_0_ ( .in(net446[1]), .out(net354[1]));
SMC_CORE_POR_right_ice8p I_SMC_CORE_POR_right (
     .core_por_b0(core_por_b0), .core_por_bb(core_por_bb),
     .vddio_rightbank(vddio_rightbank), .smc_por_b(smc_por_b0),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .creset_b(crst_filterout));
ml_cram_logic_ice8p ml_cram_logic_ice8p_1f (
     .smc_wwlwrt_en(smc_wwlwrt_en), .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wcram_rst(smc_wcram_rst), .smc_seq_rst(smc_seq_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rrst_pullwlen(smc_rrst_pullwlen),
     .smc_rpull_b(smc_rpull_b), .smc_rprec(smc_rprec),
     .smc_read(smc_read), .smc_clk(cm_clk), .por(core_por_bb),
     .smc_clk_out(cm_clk_blbrd), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff));
inv_hvt Imux4jtag_sel ( .A(trstb_pad), .Y(mux_jtag_sel));
ml_osc_top I_ml_osc_top ( .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]), .por_b(core_por_b0),
     .crst_b(crst_filterout), .smc_clk(osc_clk),
     .cnt_podt_out(cnt_podt_out));
tielo I553 ( .tielo(net497));

endmodule
// Library - xpmem, Cell - ml_dff_bl, View - schematic
// LAST TIME SAVED: May 11 18:38:30 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_dff_bl ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_clk_buf, View - schematic
// LAST TIME SAVED: Aug  9 18:57:25 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blsa_clk_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_powersurg_buf, View - schematic
// LAST TIME SAVED: Jun 18 17:30:09 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_powersurg_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I404 ( .A(net016), .Y(net012));
inv_hvt I405 ( .A(net012), .Y(o));
inv_hvt I391 ( .A(net77), .Y(net016));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_sch, View - schematic
// LAST TIME SAVED: Nov  8 11:11:57 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blsa_sch ( dataout, bl, prec_sup, cram_prec, cram_pullup_b,
     cram_write, data_muxsel, datain, latch_clock, latch_reset,
     prec_hold_b, smc_wdic_clk );
output  dataout;

inout  bl, prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, datain,
     latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff Idff ( .R(latch_reset), .D(dff_in), .CLK(latch_clock),
     .QN(write_data_b), .Q(dff_data));
pch_hvt  MP8 ( .D(net0148), .B(vdd_), .G(dataout), .S(vdd_));
pch_hvt  MP9 ( .D(bl), .B(vdd_), .G(net084), .S(net0148));
pch_hvt  M0 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  M3 ( .D(net0110), .B(vdd_), .G(cram_write), .S(prec_sup));
pch_hvt  MP12 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  M2 ( .D(bl), .B(vdd_), .G(prec_hold_b), .S(net0110));
pch_hvt  MP4 ( .D(net0143), .B(vdd_), .G(cram_pullup_b), .S(vdd_));
pch_hvt  MP5 ( .D(sa_out), .B(vdd_), .G(bl), .S(net0143));
nch_hvt  MN12 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN8 ( .D(sa_out), .B(gnd_), .G(cram_pullup_b), .S(gnd_));
nch_hvt  M1 ( .D(net0166), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN3 ( .D(sa_out), .B(gnd_), .G(bl), .S(gnd_));
nch_hvt  MN6 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
nor2_hvt I223 ( .A(net084), .B(write_data_b), .Y(n_gate));
inv_hvt I163 ( .A(write_data_b), .Y(dataout));
inv_hvt I159 ( .A(cram_prec), .Y(net0161));
inv_hvt I160 ( .A(cram_write), .Y(net084));
mux2_hvt I161 ( .in1(sa_out), .in0(datain), .out(latch_in),
     .sel(data_muxsel));
mux2_hvt I164 ( .in1(dff_data), .in0(latch_in), .out(dff_in),
     .sel(smc_wdic_clk));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_bram10k, View - schematic
// LAST TIME SAVED: Aug  4 18:43:48 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blsa_tile_bram10k ( cram_prec_out, cram_write_out, data_out,
     para_out, bl, prec_sup, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, datain, latch_clock, latch_reset,
     para_en, para_in, prec_hold_b, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out, para_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, para_en, para_in, prec_hold_b,
     smc_wdic_clk;

inout [41:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:5]  data_in;

wire  [1:4]  data_dummy_in;

wire  [0:14]  ck;

wire  [0:41]  dataout;



mux2_hvt I216 ( .in1(net119), .in0(dataout[6]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I208 ( .in1(data_dummy_in[2]), .in0(dataout[3]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I209 ( .in1(data_dummy_in[3]), .in0(dataout[4]),
     .out(data_in[3]), .sel(data_muxsel1));
mux2_hvt I196 ( .in1(data_dummy_in[1]), .in0(dataout[2]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I210 ( .in1(data_dummy_in[4]), .in0(dataout[5]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I217 ( .in1(para_in), .in0(dataout[1]), .out(data_out_mux),
     .sel(para_en));
inv_hvt I262 ( .A(data_out_mux), .Y(net151));
inv_hvt I261 ( .A(net151), .Y(data_in[0]));
inv_hvt I175 ( .A(dataout[1]), .Y(net154));
inv_hvt I176 ( .A(net154), .Y(para_out));
inv_hvt I172 ( .A(net160), .Y(data_out));
inv_hvt I171 ( .A(dataout[41]), .Y(net160));
inv_hvt I201 ( .A(latch_clock), .Y(net0133));
inv_hvt I207 ( .A(net0105), .Y(ck[14]));
inv_hvt I206 ( .A(net0107), .Y(net0105));
inv_hvt I205 ( .A(net0133), .Y(net0107));
ml_dff_bl I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net97), .Q(net119));
ml_dff_bl I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net92), .Q(data_dummy_in[4]));
ml_dff_bl I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net87), .Q(data_dummy_in[2]));
ml_dff_bl I179 ( .R(latch_reset), .D(data_in[0]), .CLK(ck[14]),
     .QN(net82), .Q(data_dummy_in[1]));
ml_dff_bl I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net77), .Q(data_dummy_in[3]));
ml_blsa_clk_buf I192_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I192_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I192_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I192_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I192_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I192_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I192_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I192_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I192_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I192_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I192_0_ ( .in(latch_clock), .o(ck[0]));
ml_powersurg_buf I165 ( .in(cram_prec), .o(net162));
ml_powersurg_buf I163 ( .in(net162), .o(net164));
ml_powersurg_buf I162 ( .in(net170), .o(net166));
ml_powersurg_buf I169 ( .in(net166), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(cram_write), .o(net170));
ml_powersurg_buf I168 ( .in(net164), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[14]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[15]),
     .dataout(dataout[15]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[13]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[14]),
     .dataout(dataout[14]), .cram_prec(net164));

endmodule
// Library - xpmem, Cell - ml_blsa_tile, View - schematic
// LAST TIME SAVED: Jan  7 13:26:29 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blsa_tile ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [53:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [53:0]  dataout;

wire  [13:0]  ck;



inv_hvt I172 ( .A(net48), .Y(data_out));
inv_hvt I171 ( .A(dataout[53]), .Y(net48));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_powersurg_buf I161 ( .in(cram_write), .o(net53));
ml_powersurg_buf I165 ( .in(net57), .o(net55));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net57));
ml_powersurg_buf I163 ( .in(net55), .o(net59));
ml_powersurg_buf I162 ( .in(net65), .o(net61));
ml_powersurg_buf I169 ( .in(net61), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net53), .o(net65));
ml_powersurg_buf I168 ( .in(net59), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_47_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[47]),
     .dataout(dataout[47]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_46_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[46]),
     .dataout(dataout[46]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_45_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[45]),
     .dataout(dataout[45]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_44_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[44]),
     .dataout(dataout[44]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_43_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[43]),
     .dataout(dataout[43]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_42_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[42]),
     .dataout(dataout[42]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net55));
ml_blsa_sch I170_53_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[53]), .dataout(dataout[53]),
     .cram_prec(net57));
ml_blsa_sch I170_52_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[52]), .dataout(dataout[52]),
     .cram_prec(net57));
ml_blsa_sch I170_51_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[51]), .dataout(dataout[51]),
     .cram_prec(net57));
ml_blsa_sch I170_50_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[50]), .dataout(dataout[50]),
     .cram_prec(net57));
ml_blsa_sch I170_49_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[49]), .dataout(dataout[49]),
     .cram_prec(net57));
ml_blsa_sch I170_48_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[48]), .dataout(dataout[48]),
     .cram_prec(net57));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net59));

endmodule
// Library - ice8chip, Cell - clk_mux2to1_ice8p, View - schematic
// LAST TIME SAVED: Nov  9 10:58:23 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module clk_mux2to1_ice8p ( gnet, bl, min0, min1, min2, min3, pgate_l,
     pgate_r, prog, reset_l, reset_r, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r );


input  prog;

output [3:0]  gnet;

inout [3:0]  bl;

input [1:0]  min2;
input [1:0]  pgate_l;
input [1:0]  reset_l;
input [1:0]  min0;
input [1:0]  reset_r;
input [1:0]  min1;
input [1:0]  min3;
input [1:0]  vdd_cntl_r;
input [1:0]  wl_l;
input [1:0]  vdd_cntl_l;
input [1:0]  pgate_r;
input [1:0]  wl_r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [7:0]  cbitb;

wire  [7:0]  cbit;

wire  [0:1]  l_vdd;



clk_mux_2to1_ice8p I_clkmux3 ( .prog(prog), .cbit(cbit[3]),
     .cbitb(cbitb[3]), .min(min3[1:0]), .clk(gnet[3]));
clk_mux_2to1_ice8p I_clkmux1 ( .prog(prog), .cbit(cbit[1]),
     .cbitb(cbitb[1]), .min(min1[1:0]), .clk(gnet[1]));
clk_mux_2to1_ice8p I_clkmux2 ( .prog(prog), .cbit(cbit[2]),
     .cbitb(cbitb[2]), .min(min2[1:0]), .clk(gnet[2]));
clk_mux_2to1_ice8p I_clkmux0 ( .prog(prog), .cbit(cbit[0]),
     .cbitb(cbitb[0]), .min(min0[1:0]), .clk(gnet[0]));
pch_hvt  I_pch_hvt_l_1_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(l_vdd[0]));
pch_hvt  I_pch_hvt_l_0_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(l_vdd[1]));
pch_hvt  M0_1_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_r[1]), .S(r_vdd[1]));
pch_hvt  M0_0_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_r[0]), .S(r_vdd[0]));
cram2x2 I_cram2x2_lft ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset_l[1:0]), .q(cbit[3:0]), .wl(wl_l[1:0]),
     .r_vdd(l_vdd[0:1]), .pgate(pgate_l[1:0]));
cram2x2 I_cram2x2_rgt ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset_r[1:0]), .q(cbit[7:4]), .wl(wl_r[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate_r[1:0]));

endmodule
// Library - xpmem, Cell - ml_blprecwrt_en, View - schematic
// LAST TIME SAVED: Aug  5 16:47:07 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blprecwrt_en ( data_out, action, clkin, data_in, rst );
output  data_out;

input  action, clkin, data_in, rst;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor3_hvt I105 ( .B(net86), .Y(net94), .A(net98), .C(rst));
nor2_hvt I103 ( .A(net88), .B(net94), .Y(net98));
inv_hvt I66 ( .A(net89), .Y(net88));
inv_hvt I168 ( .A(action), .Y(net86));
inv_hvt I165 ( .A(net98), .Y(data_out));
nand3_hvt I160 ( .Y(net89), .B(data_in), .C(action), .A(clkin));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_bram10k, View - schematic
// LAST TIME SAVED: Oct 20 17:35:57 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex2_bram10k ( data_out, latch_clock_out, para_out,
     prec_out, wrt_out, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, datain, latch_clock_in, latch_reset,
     para_en, para_in, prec_in, smc_clk_dpr, smc_wdic_clk, smc_write,
     wrt_in );
output  data_out, latch_clock_out, para_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, para_en, para_in, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in;

inout [95:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



tiehi I284 ( .tiehi(prec_hold_b));
pch_hvt  M3 ( .D(prec_sup), .B(vdd_), .G(net095), .S(vdd_));
nor2_hvt I385 ( .A(latch_reset), .B(net092), .Y(net067));
inv_hvt I198 ( .A(prec_hold_b), .Y(net095));
inv_hvt I189 ( .A(net100), .Y(latch_clock_out));
inv_hvt I191 ( .A(latch_clock_in), .Y(net100));
inv_hvt I193 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I196 ( .A(net067), .Y(net068));
inv_hvt I197 ( .A(net0130), .Y(net0105));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));
inv_hvt I187 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I188 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I192 ( .A(latch_reset), .Y(net94));
inv_hvt I194 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I190 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I195 ( .A(smc_wdic_clk), .Y(net088));
ml_blsa_tile_bram10k tile0 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .para_en(para_en), .para_in(para_in),
     .para_out(para_out), .bl(bl[41:0]),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_out),
     .cram_prec_out(prec_en_last));
ml_blsa_tile tile1 ( .prec_sup(prec_sup), .prec_hold_b(prec_hold_b),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[95:42]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net092));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net068), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net0130));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));

endmodule
// Library - xpmem, Cell - ml_buf_ice5, View - schematic
// LAST TIME SAVED: Aug  4 15:14:20 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_buf_ice5 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_last, View - schematic
// LAST TIME SAVED: Aug  4 18:09:54 2010
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blsa_tile_last ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [17:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:0]  ck;

wire  [17:0]  dataout;



ml_dff Idff ( .R(latch_reset), .D(dataout[16]), .CLK(ck[0]),
     .QN(net50), .Q(net45));
ml_dff I179 ( .R(latch_reset), .D(net58), .CLK(ck[0]), .QN(net49),
     .Q(net61));
mux2_hvt I174 ( .in1(net45), .in0(dataout[17]), .out(net58),
     .sel(data_muxsel));
tiehis I185 ( .tiehi(net040));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_buf_ice5 I205 ( .in(net61), .o(data_out), .sel(net040));
ml_powersurg_buf I169 ( .in(cram_write), .o(cram_write_out));
ml_powersurg_buf I168 ( .in(cram_prec), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[16]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[17]), .dataout(dataout[17]));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[15]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[16]), .dataout(dataout[16]));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex1_last_ice1f, View - schematic
// LAST TIME SAVED: Jan 20 18:04:52 2011
// NETLIST TIME: Jun 29 10:32:27 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex1_last_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [71:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I385 ( .A(net0111), .B(latch_reset), .Y(net0121));
ml_blsa_tile_last Iml_blsa_tile_last ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .bl(bl[71:54]),
     .latch_reset(latch_reset_buf), .datain(datain_io),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_1st), .cram_prec_out(prec_en_1st),
     .latch_clock(latch_clock_out), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blsa_tile Iml_blsa_tile_0 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_dic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_1st), .cram_prec(prec_en_1st),
     .data_out(datain_io), .cram_write_out(wrt_out),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
tiehi I284 ( .tiehi(prec_hold_b));
pch_hvt  M0 ( .D(prec_sup), .B(vdd_), .G(vdd_), .S(vdd_));
inv_hvt I197 ( .A(prec_hold_b), .Y(vdd_));
inv_hvt I194 ( .A(smc_wdic_clk), .Y(net0125));
inv_hvt I196 ( .A(net0124), .Y(net066));
inv_hvt I187 ( .A(net0121), .Y(net068));
inv_hvt I193 ( .A(latch_reset), .Y(net0127));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net0133));
inv_hvt I204 ( .A(net0137), .Y(latch_clock_out));
inv_hvt I208 ( .A(net0125), .Y(smc_dic_clk_buf));
inv_hvt I192 ( .A(latch_clock_in), .Y(net0137));
inv_hvt I190 ( .A(net0139), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net0139));
inv_hvt I203 ( .A(net0133), .Y(cram_pullup_b_buf));
inv_hvt I207 ( .A(net0127), .Y(latch_reset_buf));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net068), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net0124));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net0111));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex1_ice1f, View - schematic
// LAST TIME SAVED: Jan 20 17:58:11 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex1_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [53:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_0 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_out), .cram_prec_out(prec_en_last),
     .bl(bl[53:0]));
tiehi I284 ( .tiehi(prec_hold_b));
pch_hvt  M3 ( .D(prec_sup), .B(vdd_), .G(net075), .S(vdd_));
nor2_hvt I385 ( .A(latch_reset), .B(net049), .Y(net051));
inv_hvt I186 ( .A(data_muxsel), .Y(net084));
inv_hvt I190 ( .A(net084), .Y(data_muxsel_buf));
inv_hvt I199 ( .A(latch_clock_in), .Y(net0100));
inv_hvt I200 ( .A(prec_hold_b), .Y(net075));
inv_hvt I221 ( .A(net096), .Y(net054));
inv_hvt I201 ( .A(net051), .Y(net052));
inv_hvt I198 ( .A(net0100), .Y(latch_clock_out));
inv_hvt I197 ( .A(net090), .Y(cram_pullup_b_buf));
inv_hvt I205 ( .A(smc_wdic_clk), .Y(net094));
inv_hvt I204 ( .A(net094), .Y(smc_wdic_clk_buf));
inv_hvt I196 ( .A(cram_pullup_b), .Y(net090));
inv_hvt I203 ( .A(net086), .Y(latch_reset_buf));
inv_hvt I202 ( .A(latch_reset), .Y(net086));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net052), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net096));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net049));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_1st, View - schematic
// LAST TIME SAVED: Aug  4 18:53:38 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ml_blsa_tile_1st ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [55:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:4]  data_dummy_in;

wire  [0:55]  dataout;

wire  [1:5]  data_in;

wire  [0:14]  ck;



ml_dff I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net132), .Q(net154));
ml_dff I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net137), .Q(data_dummy_in[4]));
ml_dff I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net142), .Q(data_dummy_in[2]));
ml_dff I179 ( .R(latch_reset), .D(datain), .CLK(ck[14]), .QN(net147),
     .Q(data_dummy_in[1]));
ml_dff I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net152), .Q(data_dummy_in[3]));
inv_hvt I171 ( .A(dataout[55]), .Y(net121));
inv_hvt I172 ( .A(net121), .Y(data_out));
inv_hvt I224 ( .A(net0130), .Y(ck[14]));
inv_hvt I225 ( .A(net0129), .Y(net0130));
inv_hvt I226 ( .A(net0126), .Y(net0129));
inv_hvt I229 ( .A(latch_clock), .Y(net0122));
inv_hvt I227 ( .A(net0124), .Y(net0126));
inv_hvt I228 ( .A(net0122), .Y(net0124));
mux2_hvt I197 ( .in1(net154), .in0(dataout[4]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I232 ( .in1(data_dummy_in[2]), .in0(dataout[1]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I230 ( .in1(data_dummy_in[4]), .in0(dataout[3]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I233 ( .in1(data_dummy_in[1]), .in0(dataout[0]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I231 ( .in1(data_dummy_in[3]), .in0(dataout[2]),
     .out(data_in[3]), .sel(data_muxsel1));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[14]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[13]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[12]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[11]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[10]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[9]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[8]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[7]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[6]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[4]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[3]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[2]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[1]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(datain), .cram_prec(cram_prec_out),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_47_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[47]),
     .dataout(dataout[47]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_46_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[46]),
     .dataout(dataout[46]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_45_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[45]),
     .dataout(dataout[45]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_44_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[44]),
     .dataout(dataout[44]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_43_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[43]),
     .dataout(dataout[43]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_42_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[42]),
     .dataout(dataout[42]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[41]),
     .dataout(dataout[41]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[40]),
     .dataout(dataout[40]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[39]),
     .dataout(dataout[39]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[38]),
     .dataout(dataout[38]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[37]),
     .dataout(dataout[37]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[36]),
     .dataout(dataout[36]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[35]),
     .dataout(dataout[35]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[34]),
     .dataout(dataout[34]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[33]),
     .dataout(dataout[33]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[32]),
     .dataout(dataout[32]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_55_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[54]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[55]),
     .dataout(dataout[55]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_54_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[53]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[54]),
     .dataout(dataout[54]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_53_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[53]),
     .dataout(dataout[53]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_52_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[52]),
     .dataout(dataout[52]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_51_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[51]),
     .dataout(dataout[51]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_50_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[50]),
     .dataout(dataout[50]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_49_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[49]),
     .dataout(dataout[49]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_48_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[48]),
     .dataout(dataout[48]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[31]),
     .dataout(dataout[31]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[30]),
     .dataout(dataout[30]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[29]),
     .dataout(dataout[29]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[28]),
     .dataout(dataout[28]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[27]),
     .dataout(dataout[27]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[26]),
     .dataout(dataout[26]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[25]),
     .dataout(dataout[25]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[24]),
     .dataout(dataout[24]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[23]),
     .dataout(dataout[23]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[22]),
     .dataout(dataout[22]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[21]),
     .dataout(dataout[21]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[20]),
     .dataout(dataout[20]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[19]),
     .dataout(dataout[19]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[18]),
     .dataout(dataout[18]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[17]),
     .dataout(dataout[17]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[16]),
     .dataout(dataout[16]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_powersurg_buf I161 ( .in(cram_write), .o(net104));
ml_powersurg_buf I165 ( .in(net108), .o(net106));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net108));
ml_powersurg_buf I163 ( .in(net106), .o(net110));
ml_powersurg_buf I162 ( .in(net116), .o(net112));
ml_powersurg_buf I169 ( .in(net112), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net104), .o(net116));
ml_powersurg_buf I168 ( .in(net110), .o(cram_prec_out));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_1st_ice1f, View - schematic
// LAST TIME SAVED: Jan 20 17:52:04 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex2_1st_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [109:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_1 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_wdic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[109:56]));
ml_blsa_tile_1st Iml_blsa_tile_1st_0 ( .prec_sup(prec_sup),
     .prec_hold_b(prec_hold_b), .bl(bl[55:0]),
     .cram_pullup_b(cram_pullup_buf), .latch_clock(latch_clock_out),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .datain(datain), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_mid),
     .cram_prec(prec_en_mid), .data_out(data_tile),
     .cram_write_out(wrt_out), .cram_prec_out(prec_en_last));
nor2_hvt I385 ( .A(latch_reset), .B(net86), .Y(net117));
pch_hvt  M3 ( .D(prec_sup), .B(vdd_), .G(net106), .S(vdd_));
tiehi I284 ( .tiehi(prec_hold_b));
inv_hvt I190 ( .A(net095), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net095));
inv_hvt I202 ( .A(latch_reset), .Y(net0113));
inv_hvt I203 ( .A(net0113), .Y(latch_reset_buf));
inv_hvt I196 ( .A(cram_pullup_b), .Y(net0109));
inv_hvt I204 ( .A(net0105), .Y(smc_wdic_clk_buf));
inv_hvt I200 ( .A(prec_hold_b), .Y(net106));
inv_hvt I205 ( .A(smc_wdic_clk), .Y(net0105));
inv_hvt I221 ( .A(net138), .Y(net110));
inv_hvt I197 ( .A(net0109), .Y(cram_pullup_buf));
inv_hvt I198 ( .A(net099), .Y(latch_clock_out));
inv_hvt I199 ( .A(latch_clock_in), .Y(net099));
inv_hvt I201 ( .A(net117), .Y(net118));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net118), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net138));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net86));

endmodule
// Library - xpmem, Cell - ml_buf_ice1f, View - schematic
// LAST TIME SAVED: Jan  7 14:21:36 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ml_buf_ice1f ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_bank_ice1f, View - schematic
// LAST TIME SAVED: Mar  8 09:38:22 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ml_blsa_bank_ice1f ( cm_sdo_u, bl, banksel, cm_sdi_u,
     cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk,
     smc_write );


input  banksel, cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk,
     smc_write;

output [1:0]  cm_sdo_u;

inout [331:0]  bl;

input [1:0]  cm_sdi_u;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tilex2_bram10k I_lt_34 ( .smc_write(smc_write_buf),
     .para_en(cor_en_8bpcfg_buf), .para_in(sdi1_buf),
     .para_out(para_out), .bl(bl[259:164]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net0137),
     .latch_clock_out(net0171), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret), .wrt_in(wrt_out_5),
     .prec_in(prec_out_5), .latch_reset(latch_reset_buf),
     .datain(data_out_2), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_34),
     .prec_out(prec_out_34), .data_out(data_out_34));
ml_blsa_tilex1_last_ice1f I_lt_5 ( .smc_write(smc_write_buf),
     .bl(bl[331:260]), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(smc_clk), .latch_clock_out(net0137),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf),
     .wrt_in(cram_write_buf), .prec_in(net377),
     .latch_reset(latch_reset_buf), .datain(data_out_34),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_5), .prec_out(prec_out_5),
     .data_out(cm_sdo_u[1]));
ml_blsa_tilex1_ice1f I_lt_2 ( .smc_write(smc_write_buf),
     .bl(bl[163:110]), .cram_pullup_b(net0161),
     .latch_clock_in(net0171), .latch_clock_out(net393),
     .smc_wdic_clk(net0158), .smc_clk_dpr(net0165),
     .wrt_in(wrt_out_34), .prec_in(prec_out_34),
     .latch_reset(latch_reset_buf), .datain(data_out_01),
     .data_muxsel1(net0152), .data_muxsel(net0149),
     .cram_write(net0146), .cram_prec(net0155), .wrt_out(wrt_out_2),
     .prec_out(prec_out_2), .data_out(data_out_2));
ml_blsa_tilex2_1st_ice1f I_lt_01 ( .smc_write(smc_write_buf),
     .wrt_in(wrt_out_2), .prec_in(prec_out_2),
     .latch_reset(latch_reset_buf), .datain(net0140),
     .data_muxsel1(net0152), .data_muxsel(net0149),
     .cram_write(net0146), .bl(bl[109:0]), .cram_prec(net0155),
     .wrt_out(wrt_out_01), .prec_out(prec_out_01),
     .data_out(data_out_01), .latch_clock_in(net393),
     .cram_pullup_b(net0161), .latch_clock_out(net440),
     .smc_wdic_clk(net0158), .smc_clk_dpr(net0354));
ml_buf_ice1f I291 ( .in(net0160), .o(net0165),
     .sel(smc_clk_buf_b_ret));
ml_buf_ice1f I292 ( .in(net0160), .o(net0354), .sel(smc_clk_buf));
ml_buf_ice1f I284 ( .in(net0160), .o(net0140), .sel(sdi0_buf));
ml_buf_ice1f I247 ( .in(cm_sdi_u[1]), .o(sdi1_buf), .sel(net527));
ml_buf_ice1f I249 ( .in(net519), .o(cor_en_8bpcfg_buf), .sel(net527));
ml_buf_ice1f I285 ( .in(net0160), .o(net0146), .sel(cram_write_buf));
ml_buf_ice1f I265 ( .in(net527), .o(cm_sdo_u[0]), .sel(net451));
ml_buf_ice1f I257 ( .in(smc_wdic_clk), .o(smc_wdic_clk_buf),
     .sel(banksel));
ml_buf_ice1f I203 ( .in(data_muxsel1), .o(data_muxsel1_buf),
     .sel(banksel));
ml_buf_ice1f I205 ( .in(latch_reset), .o(latch_reset_buf),
     .sel(net529));
ml_buf_ice1f I207 ( .in(cram_write), .o(cram_write_buf),
     .sel(banksel));
ml_buf_ice1f I208 ( .in(cram_pullup_logic_b), .o(cram_pullup_b_buf),
     .sel(cram_pullup_logic_b));
ml_buf_ice1f I288 ( .in(net0160), .o(net0149), .sel(data_muxsel_buf));
ml_buf_ice1f I201 ( .in(cram_prec), .o(cram_prec_buf), .sel(banksel));
ml_buf_ice1f I289 ( .in(net0160), .o(net0152), .sel(data_muxsel1_buf));
ml_buf_ice1f I294b ( .in(banksel), .o(smc_write_buf), .sel(smc_write));
ml_buf_ice1f I216 ( .in(net528), .o(net474), .sel(net528));
ml_buf_ice1f I286 ( .in(net0160), .o(net0155), .sel(cram_prec_buf));
ml_buf_ice1f I8 ( .in(net0160), .o(net0158), .sel(smc_wdic_clk_buf));
ml_buf_ice1f I290 ( .in(net0160), .o(net0161),
     .sel(cram_pullup_b_buf));
ml_buf_ice1f I245 ( .in(cm_sdi_u[0]), .o(sdi0_buf), .sel(net527));
ml_buf_ice1f I187 ( .in(smc_clk), .o(smc_clk_buf), .sel(smc_clk));
ml_buf_ice1f I188 ( .in(net525), .o(smc_clk_buf_b_ret), .sel(net525));
ml_buf_ice1f I204 ( .in(data_muxsel), .o(data_muxsel_buf),
     .sel(banksel));
ml_buf_ice1f I227 ( .in(net532), .o(net489), .sel(net532));
nor3_hvt I217 ( .B(net531), .Y(net492), .A(net531), .C(net531));
nor3_hvt I220 ( .B(net500), .Y(net496), .A(net500), .C(net500));
nor3_hvt I218 ( .B(net492), .Y(net500), .A(net492), .C(net492));
nand3_hvt I231 ( .Y(net503), .B(net507), .C(net507), .A(net507));
nand3_hvt I230 ( .Y(net507), .B(net511), .C(net511), .A(net511));
nand3_hvt I224 ( .Y(net511), .B(net526), .C(net526), .A(net526));
nor2_hvt I254 ( .B(net515), .Y(net522), .A(cram_pullup_b));
inv_hvt I253 ( .A(cor_en_8bpcfg_b), .Y(net519));
inv_hvt I256 ( .A(banksel), .Y(net515));
inv_hvt I255 ( .A(net522), .Y(cram_pullup_logic_b));
inv_hvt I189 ( .A(smc_clk), .Y(net525));
tiehi I268 ( .tiehi(net526));
tiehi I272 ( .tiehi(net527));
tiehi I287 ( .tiehi(net0160));
tiehi I271 ( .tiehi(net528));
tiehi I273 ( .tiehi(net529));
tiehi I267 ( .tiehi(net377));
tiehi I270 ( .tiehi(net531));
tiehi I269 ( .tiehi(net532));
ml_dff_bl I_ml_dff_bl ( .R(latch_reset_buf), .D(para_out),
     .CLK(smc_clk), .QN(net536), .Q(net451));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev0, View - schematic
// LAST TIME SAVED: Jun 23 08:48:28 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module clkmandcmuxrev0 ( clk, clkb, glb2local, s_r, cbit, cbitb,
     glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, min0, min1,
     min2, min3, prog );
output  clk, clkb, s_r;

input  prog;

output [3:0]  glb2local;

input [7:0]  min2;
input [7:0]  min0;
input [7:0]  min3;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g0;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g3;
input [7:0]  min1;
input [31:0]  cbit;
input [31:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_mux12to1_icc I_clkmux12to1 ( .prog(prog), .min({lc_trk_g3[1],
     lc_trk_g2[0], lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}),
     .clk(clk), .clkb(clkb), .cbitb({cbitb[31], cbitb[4], cbitb[3],
     cbitb[2], cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3],
     cbit[2], cbit[1], cbit[0]}), .cenb(ceb));
clk_mux8to1 I_clkmux8to1_0 ( .prog(prog), .inmuxo(glb2local[0]),
     .min(min3[7:0]), .cbit(cbit[16:13]), .cbitb(cbitb[16:13]));
clk_mux8to1 I_clkmux8to1_1 ( .prog(prog), .inmuxo(glb2local[1]),
     .min(min2[7:0]), .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I_clkmux8to1_3 ( .prog(prog), .inmuxo(glb2local[3]),
     .min(min0[7:0]), .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));
clk_mux8to1 I_clkmux8to1_2 ( .prog(prog), .inmuxo(glb2local[2]),
     .min(min1[7:0]), .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
ce_clkm8to1 I_cemux8to1 ( .cbitb(cbitb[8:5]), .min({lc_trk_g3[3],
     lc_trk_g2[2], lc_trk_g1[3], lc_trk_g0[2], glb_netwk[7],
     glb_netwk[5], glb_netwk[3], glb_netwk[1]}), .cbit(cbit[8:5]),
     .moutb(ceb), .prog(prog));
sr_clkm8to1 I_srmux8to1 ( .cbitb(cbitb[12:9]), .min({lc_trk_g3[5],
     lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4], glb_netwk[6],
     glb_netwk[4], glb_netwk[2], glb_netwk[0]}), .cbit(cbit[12:9]),
     .mout(s_r), .prog(prog));

endmodule
// Library - ice1chip, Cell - CHIP_route_top_ice1f, View - schematic
// LAST TIME SAVED: Mar  7 16:46:33 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module CHIP_route_top_ice1f ( cm_sdo_u1, cm_sdo_u3, bl_top,
     cm_banksel_bltld3, cm_banksel_bltrd1, cm_clk_bltld3,
     cm_clk_bltrd1, cm_prec_bltld3, cm_sdi_u1d3, cm_sdi_u3d2,
     core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1r,
     smc_write_bltl1d1, smc_write_bltld3 );


input  cm_clk_bltld3, cm_clk_bltrd1, cm_prec_bltld3, core_por_b_rowu1,
     core_por_b_rowu3, cram_prec_bltrd1, cram_pullup_b_bltrd1,
     cram_pullup_bltld3, cram_write_bltld3, cram_write_bltrd1,
     data_muxsel1_bltld3, data_muxsel1_bltrd1, data_muxsel_bltld3,
     data_muxsel_bltrd1, en_8bconfig_b_bltld3, en_8bconfig_b_bltrd1,
     smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1r, smc_write_bltl1d1,
     smc_write_bltld3;

output [1:0]  cm_sdo_u1;
output [1:0]  cm_sdo_u3;

inout [663:0]  bl_top;

input [3:3]  cm_banksel_bltrd1;
input [1:0]  cm_sdi_u1d3;
input [1:0]  cm_sdi_u3d2;
input [1:1]  cm_banksel_bltld3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_bank_ice1f I_bltr ( .smc_write(smc_write_bltl1d1),
     .bl(bl_top[663:332]), .smc_wdic_clk(smc_wdis_dclk_bltrd1r),
     .smc_clk(cm_clk_bltrd1), .cm_sdi_u(cm_sdi_u3d2[1:0]),
     .latch_reset(core_por_b_rowu3), .cm_sdo_u(cm_sdo_u3[1:0]),
     .data_muxsel1(data_muxsel1_bltrd1),
     .data_muxsel(data_muxsel_bltrd1), .cram_write(cram_write_bltrd1),
     .cram_prec(cram_prec_bltrd1),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltrd1),
     .cram_pullup_b(cram_pullup_b_bltrd1),
     .banksel(cm_banksel_bltrd1[3]));
ml_blsa_bank_ice1f I_bltlu1 ( .smc_write(smc_write_bltld3),
     .bl({bl_top[0], bl_top[1], bl_top[2], bl_top[3], bl_top[4],
     bl_top[5], bl_top[6], bl_top[7], bl_top[8], bl_top[9], bl_top[10],
     bl_top[11], bl_top[12], bl_top[13], bl_top[14], bl_top[15],
     bl_top[16], bl_top[17], bl_top[18], bl_top[19], bl_top[20],
     bl_top[21], bl_top[22], bl_top[23], bl_top[24], bl_top[25],
     bl_top[26], bl_top[27], bl_top[28], bl_top[29], bl_top[30],
     bl_top[31], bl_top[32], bl_top[33], bl_top[34], bl_top[35],
     bl_top[36], bl_top[37], bl_top[38], bl_top[39], bl_top[40],
     bl_top[41], bl_top[42], bl_top[43], bl_top[44], bl_top[45],
     bl_top[46], bl_top[47], bl_top[48], bl_top[49], bl_top[50],
     bl_top[51], bl_top[52], bl_top[53], bl_top[54], bl_top[55],
     bl_top[56], bl_top[57], bl_top[58], bl_top[59], bl_top[60],
     bl_top[61], bl_top[62], bl_top[63], bl_top[64], bl_top[65],
     bl_top[66], bl_top[67], bl_top[68], bl_top[69], bl_top[70],
     bl_top[71], bl_top[72], bl_top[73], bl_top[74], bl_top[75],
     bl_top[76], bl_top[77], bl_top[78], bl_top[79], bl_top[80],
     bl_top[81], bl_top[82], bl_top[83], bl_top[84], bl_top[85],
     bl_top[86], bl_top[87], bl_top[88], bl_top[89], bl_top[90],
     bl_top[91], bl_top[92], bl_top[93], bl_top[94], bl_top[95],
     bl_top[96], bl_top[97], bl_top[98], bl_top[99], bl_top[100],
     bl_top[101], bl_top[102], bl_top[103], bl_top[104], bl_top[105],
     bl_top[106], bl_top[107], bl_top[108], bl_top[109], bl_top[110],
     bl_top[111], bl_top[112], bl_top[113], bl_top[114], bl_top[115],
     bl_top[116], bl_top[117], bl_top[118], bl_top[119], bl_top[120],
     bl_top[121], bl_top[122], bl_top[123], bl_top[124], bl_top[125],
     bl_top[126], bl_top[127], bl_top[128], bl_top[129], bl_top[130],
     bl_top[131], bl_top[132], bl_top[133], bl_top[134], bl_top[135],
     bl_top[136], bl_top[137], bl_top[138], bl_top[139], bl_top[140],
     bl_top[141], bl_top[142], bl_top[143], bl_top[144], bl_top[145],
     bl_top[146], bl_top[147], bl_top[148], bl_top[149], bl_top[150],
     bl_top[151], bl_top[152], bl_top[153], bl_top[154], bl_top[155],
     bl_top[156], bl_top[157], bl_top[158], bl_top[159], bl_top[160],
     bl_top[161], bl_top[162], bl_top[163], bl_top[164], bl_top[165],
     bl_top[166], bl_top[167], bl_top[168], bl_top[169], bl_top[170],
     bl_top[171], bl_top[172], bl_top[173], bl_top[174], bl_top[175],
     bl_top[176], bl_top[177], bl_top[178], bl_top[179], bl_top[180],
     bl_top[181], bl_top[182], bl_top[183], bl_top[184], bl_top[185],
     bl_top[186], bl_top[187], bl_top[188], bl_top[189], bl_top[190],
     bl_top[191], bl_top[192], bl_top[193], bl_top[194], bl_top[195],
     bl_top[196], bl_top[197], bl_top[198], bl_top[199], bl_top[200],
     bl_top[201], bl_top[202], bl_top[203], bl_top[204], bl_top[205],
     bl_top[206], bl_top[207], bl_top[208], bl_top[209], bl_top[210],
     bl_top[211], bl_top[212], bl_top[213], bl_top[214], bl_top[215],
     bl_top[216], bl_top[217], bl_top[218], bl_top[219], bl_top[220],
     bl_top[221], bl_top[222], bl_top[223], bl_top[224], bl_top[225],
     bl_top[226], bl_top[227], bl_top[228], bl_top[229], bl_top[230],
     bl_top[231], bl_top[232], bl_top[233], bl_top[234], bl_top[235],
     bl_top[236], bl_top[237], bl_top[238], bl_top[239], bl_top[240],
     bl_top[241], bl_top[242], bl_top[243], bl_top[244], bl_top[245],
     bl_top[246], bl_top[247], bl_top[248], bl_top[249], bl_top[250],
     bl_top[251], bl_top[252], bl_top[253], bl_top[254], bl_top[255],
     bl_top[256], bl_top[257], bl_top[258], bl_top[259], bl_top[260],
     bl_top[261], bl_top[262], bl_top[263], bl_top[264], bl_top[265],
     bl_top[266], bl_top[267], bl_top[268], bl_top[269], bl_top[270],
     bl_top[271], bl_top[272], bl_top[273], bl_top[274], bl_top[275],
     bl_top[276], bl_top[277], bl_top[278], bl_top[279], bl_top[280],
     bl_top[281], bl_top[282], bl_top[283], bl_top[284], bl_top[285],
     bl_top[286], bl_top[287], bl_top[288], bl_top[289], bl_top[290],
     bl_top[291], bl_top[292], bl_top[293], bl_top[294], bl_top[295],
     bl_top[296], bl_top[297], bl_top[298], bl_top[299], bl_top[300],
     bl_top[301], bl_top[302], bl_top[303], bl_top[304], bl_top[305],
     bl_top[306], bl_top[307], bl_top[308], bl_top[309], bl_top[310],
     bl_top[311], bl_top[312], bl_top[313], bl_top[314], bl_top[315],
     bl_top[316], bl_top[317], bl_top[318], bl_top[319], bl_top[320],
     bl_top[321], bl_top[322], bl_top[323], bl_top[324], bl_top[325],
     bl_top[326], bl_top[327], bl_top[328], bl_top[329], bl_top[330],
     bl_top[331]}), .smc_wdic_clk(smc_wdis_dclk_bltld3),
     .smc_clk(cm_clk_bltld3), .cm_sdi_u(cm_sdi_u1d3[1:0]),
     .latch_reset(core_por_b_rowu1), .cm_sdo_u(cm_sdo_u1[1:0]),
     .data_muxsel1(data_muxsel1_bltld3),
     .data_muxsel(data_muxsel_bltld3), .cram_write(cram_write_bltld3),
     .cram_prec(cm_prec_bltld3),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltld3),
     .cram_pullup_b(cram_pullup_bltld3),
     .banksel(cm_banksel_bltld3[1]));

endmodule
// Library - ice1chip, Cell - CHIP_route_bot_ice1f_blbank, View -
//schematic
// LAST TIME SAVED: Mar  8 09:53:19 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module CHIP_route_bot_ice1f_blbank ( cm_sdo_u0, cm_sdo_u2, bl_bot,
     cm_banksel_blbld1_0_, cm_banksel_blbrd_2_, cm_clk_blbld,
     cm_clk_blbrd, cm_sdi_u0d1, cm_sdi_u2d, core_por_bb, core_por_bbl0,
     cram_prec, cram_prec_blbld, cram_pullup_b, cram_pullup_blbld,
     cram_write, cram_write_blbld, data_muxsel1_blbld,
     data_muxsel1_blbrd, data_muxsel_blbld, data_muxsel_blbrd,
     en_8bconfig_b_blbld, en_8bconfig_b_blbrd, smc_wdis_dclk_blbld,
     smc_wdis_dclk_blbrd, smc_write, smc_writel0 );


input  cm_banksel_blbld1_0_, cm_banksel_blbrd_2_, cm_clk_blbld,
     cm_clk_blbrd, core_por_bb, core_por_bbl0, cram_prec,
     cram_prec_blbld, cram_pullup_b, cram_pullup_blbld, cram_write,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel1_blbrd,
     data_muxsel_blbld, data_muxsel_blbrd, en_8bconfig_b_blbld,
     en_8bconfig_b_blbrd, smc_wdis_dclk_blbld, smc_wdis_dclk_blbrd,
     smc_write, smc_writel0;

output [1:0]  cm_sdo_u2;
output [1:0]  cm_sdo_u0;

inout [663:0]  bl_bot;

input [1:0]  cm_sdi_u2d;
input [1:0]  cm_sdi_u0d1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



CHIP_route_top_ice1f I_CHIP_route_top_ice1f ( .bl_top(bl_bot[663:0]),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_blbld),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_blbrd),
     .en_8bconfig_b_bltld3(en_8bconfig_b_blbld),
     .data_muxsel_bltrd1(data_muxsel_blbrd),
     .data_muxsel_bltld3(data_muxsel_blbld),
     .data_muxsel1_bltrd1(data_muxsel1_blbrd),
     .data_muxsel1_bltld3(data_muxsel1_blbld),
     .cram_write_bltrd1(cram_write),
     .cram_write_bltld3(cram_write_blbld),
     .cram_pullup_bltld3(cram_pullup_blbld),
     .cram_pullup_b_bltrd1(cram_pullup_b),
     .cram_prec_bltrd1(cram_prec), .core_por_b_rowu3(core_por_bb),
     .core_por_b_rowu1(core_por_bbl0), .cm_sdi_u3d2(cm_sdi_u2d[1:0]),
     .cm_sdi_u1d3(cm_sdi_u0d1[1:0]), .cm_prec_bltld3(cram_prec_blbld),
     .cm_clk_bltrd1(cm_clk_blbrd), .cm_clk_bltld3(cm_clk_blbld),
     .cm_banksel_bltrd1(cm_banksel_blbrd_2_),
     .cm_banksel_bltld3(cm_banksel_blbld1_0_),
     .cm_sdo_u3(cm_sdo_u2[1:0]), .cm_sdo_u1(cm_sdo_u0[1:0]),
     .smc_write_bltld3(smc_writel0), .smc_write_bltl1d1(smc_write));

endmodule
// Library - ice1chip, Cell - CHIP_route_bot_ice1f, View - schematic
// LAST TIME SAVED: Apr 22 10:25:51 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module CHIP_route_bot_ice1f ( cm_banksel_blbld1_0_,
     cm_banksel_blbld_1_, cm_clk_blbld, cm_sdi_u1d, cm_sdo_u0d1,
     cm_sdo_u1d3, cm_sdo_u2d1, core_por_b2, core_por_bbl0,
     cram_pgateoffl0, cram_prec_blbld, cram_pullup_blbld, cram_rstl0,
     cram_vddoffl0, cram_wl_enl0, cram_write_blbld, data_muxsel1_blbld,
     data_muxsel_blbld, en_8bconfig_b_blbld, j_rst_bl0, last_rsr3,
     row_testl1, smc_core_por_bottom1, smc_core_por_bottom2,
     smc_row_incl0, smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0,
     spi_ss_in_bbankd, tck_padl0, bl_bot, cm_banksel,
     cm_banksel_blbrd_2_, cm_clk_blbrd, cm_sdi_u0, cm_sdi_u1,
     cm_sdi_u2d, cm_sdo_u1d1, core_por_b0, core_por_bb, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     spi_ss_in_bbank, vddio_botbank, vddio_spi );
output  cm_banksel_blbld1_0_, cm_banksel_blbld_1_, cm_clk_blbld,
     core_por_b2, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, last_rsr3, row_testl1,
     smc_core_por_bottom1, smc_core_por_bottom2, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;


input  cm_banksel_blbrd_2_, cm_clk_blbrd, core_por_b0, core_por_bb,
     cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     vddio_botbank, vddio_spi;

output [1:0]  cm_sdo_u2d1;
output [4:0]  spi_ss_in_bbankd;
output [1:0]  cm_sdo_u0d1;
output [1:0]  cm_sdi_u1d;
output [1:0]  cm_sdo_u1d3;

inout [663:0]  bl_bot;

input [1:0]  cm_sdi_u0;
input [4:0]  spi_ss_in_bbank;
input [1:0]  cm_sdi_u2d;
input [1:0]  cm_sdi_u1;
input [1:0]  cm_sdo_u1d1;
input [1:0]  cm_banksel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1_buf;

wire  [0:1]  net233;

wire  [1:0]  cm_sdo_u0_buf;

wire  [0:1]  net297;

wire  [1:0]  dff_u2_d0;

wire  [1:0]  cm_sdi_u2d_buf;

wire  [0:1]  net321;

wire  [0:1]  net229;

wire  [0:1]  net317;

wire  [0:1]  net235;

wire  [0:1]  net234;

wire  [1:0]  cm_sdi_u0d1;

wire  [1:0]  cm_sdo_u2;

wire  [1:0]  dff_u0_d1;

wire  [1:0]  dff_u1_d1;

wire  [1:0]  cm_sdo_u0;



CHIP_route_bot_ice1f_blbank I_CHIP_route_bot_ice1f_blbank (
     .bl_bot(bl_bot[663:0]), .smc_writel0(smc_writel0),
     .smc_write(smc_write), .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_write(cram_write),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_pullup_b(cram_pullup_b), .cram_prec_blbld(cram_prec_blbld),
     .cram_prec(cram_prec), .core_por_bbl0(core_por_bbl0),
     .core_por_bb(core_por_bb), .cm_sdi_u2d(cm_sdi_u2d_buf[1:0]),
     .cm_sdi_u0d1(cm_sdi_u0d1[1:0]), .cm_clk_blbrd(cm_clk_blbrd),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1_0_),
     .cm_sdo_u0(cm_sdo_u0[1:0]), .cm_sdo_u2(cm_sdo_u2[1:0]));
tielo I561_1_ ( .tielo(net229[0]));
tielo I561_0_ ( .tielo(net229[1]));
tielo I562 ( .tielo(net230));
tielo I563 ( .tielo(net231));
tielo I564 ( .tielo(net232));
tielo I559_1_ ( .tielo(net233[0]));
tielo I559_0_ ( .tielo(net233[1]));
tielo I560_1_ ( .tielo(net234[0]));
tielo I560_0_ ( .tielo(net234[1]));
sg_bufx10_ice8p I532_1_ ( .in(net235[0]), .out(cm_sdi_u1d[1]));
sg_bufx10_ice8p I532_0_ ( .in(net235[1]), .out(cm_sdi_u1d[0]));
sg_bufx10_ice8p I484 ( .in(cram_pgateoff), .out(net327));
sg_bufx10_ice8p I482 ( .in(net239), .out(cram_pgateoffl0));
sg_bufx10_ice8p I516 ( .in(net241), .out(cm_banksel_blbld_1_));
sg_bufx10_ice8p I474 ( .in(net243), .out(net245));
sg_bufx10_ice8p I475 ( .in(net245), .out(smc_writel0));
sg_bufx10_ice8p I480 ( .in(net247), .out(net283));
sg_bufx10_ice8p I333 ( .in(j_rst_b), .out(j_rst_bl0));
sg_bufx10_ice8p I336 ( .in(core_por_bb), .out(net361));
sg_bufx10_ice8p I523 ( .in(smc_clk_mid), .out(cm_clk_blbld));
sg_bufx10_ice8p I478 ( .in(cram_vddoff), .out(net363));
sg_bufx10_ice8p I488 ( .in(predata_cram_pullup_b), .out(net295));
sg_bufx10_ice8p I473 ( .in(smc_write), .out(net243));
sg_bufx10_ice8p I496 ( .in(en_8bconfig_b_blbrd),
     .out(predata_en_8bconfig_b));
sg_bufx10_ice8p I527_1_ ( .in(cm_sdi_u0[1]), .out(net321[0]));
sg_bufx10_ice8p I527_0_ ( .in(cm_sdi_u0[0]), .out(net321[1]));
sg_bufx10_ice8p I459 ( .in(smc_row_inc), .out(net377));
sg_bufx10_ice8p I491 ( .in(cram_write), .out(predata_cram_write));
sg_bufx10_ice8p I568_4_ ( .in(spi_ss_in_bbank[4]),
     .out(spi_ss_in_bbankd[4]));
sg_bufx10_ice8p I568_3_ ( .in(spi_ss_in_bbank[3]),
     .out(spi_ss_in_bbankd[3]));
sg_bufx10_ice8p I568_2_ ( .in(spi_ss_in_bbank[2]),
     .out(spi_ss_in_bbankd[2]));
sg_bufx10_ice8p I568_1_ ( .in(spi_ss_in_bbank[1]),
     .out(spi_ss_in_bbankd[1]));
sg_bufx10_ice8p I568_0_ ( .in(spi_ss_in_bbank[0]),
     .out(spi_ss_in_bbankd[0]));
sg_bufx10_ice8p I467 ( .in(predata_muxsel1), .out(net291));
sg_bufx10_ice8p I505 ( .in(net273), .out(smc_rsr_rstl0));
sg_bufx10_ice8p I567 ( .in(core_por_b0), .out(core_por_b2));
sg_bufx10_ice8p I521 ( .in(net277), .out(cm_banksel_blbld1_0_));
sg_bufx10_ice8p I175 ( .in(net279), .out(data_muxsel_blbld));
sg_bufx10_ice8p I492 ( .in(net281), .out(cram_write_blbld));
sg_bufx10_ice8p I481 ( .in(net283), .out(cram_rstl0));
sg_bufx10_ice8p I439 ( .in(j_tck), .out(tck_padl0));
sg_bufx10_ice8p I495 ( .in(net287), .out(en_8bconfig_b_blbld));
sg_bufx10_ice8p I570 ( .in(net289), .out(core_por_bbl0));
sg_bufx10_ice8p I466 ( .in(net291), .out(data_muxsel1_blbld));
sg_bufx10_ice8p I486 ( .in(net293), .out(cram_prec_blbld));
sg_bufx10_ice8p I489 ( .in(net295), .out(cram_pullup_blbld));
sg_bufx10_ice8p I531_1_ ( .in(net297[0]), .out(net235[0]));
sg_bufx10_ice8p I531_0_ ( .in(net297[1]), .out(net235[1]));
sg_bufx10_ice8p I485 ( .in(cram_prec), .out(predata_cram_prec));
sg_bufx10_ice8p I533_1_ ( .in(cm_sdi_u1[1]), .out(net297[0]));
sg_bufx10_ice8p I533_0_ ( .in(cm_sdi_u1[0]), .out(net297[1]));
sg_bufx10_ice8p I520 ( .in(net303), .out(net277));
sg_bufx10_ice8p I517 ( .in(net305), .out(net241));
sg_bufx10_ice8p I493 ( .in(predata_cram_write), .out(net281));
sg_bufx10_ice8p I519 ( .in(cm_banksel[0]), .out(net303));
sg_bufx10_ice8p I509 ( .in(net311), .out(row_testl1));
sg_bufx10_ice8p I469 ( .in(net313), .out(smc_row_incl0));
sg_bufx10_ice8p I504 ( .in(smc_rsr_rst), .out(net331));
sg_bufx10_ice8p I529_1_ ( .in(net317[0]), .out(cm_sdi_u0d1[1]));
sg_bufx10_ice8p I529_0_ ( .in(net317[1]), .out(cm_sdi_u0d1[0]));
sg_bufx10_ice8p I476 ( .in(net319), .out(cram_vddoffl0));
sg_bufx10_ice8p I530_1_ ( .in(net321[0]), .out(net317[0]));
sg_bufx10_ice8p I530_0_ ( .in(net321[1]), .out(net317[1]));
sg_bufx10_ice8p I471 ( .in(net323), .out(net347));
sg_bufx10_ice8p I510 ( .in(net325), .out(net311));
sg_bufx10_ice8p I483 ( .in(net327), .out(net239));
sg_bufx10_ice8p I464 ( .in(predata_muxsel), .out(net279));
sg_bufx10_ice8p I503 ( .in(net331), .out(net273));
sg_bufx10_ice8p I494 ( .in(predata_en_8bconfig_b), .out(net287));
sg_bufx10_ice8p I490 ( .in(cram_pullup_b),
     .out(predata_cram_pullup_b));
sg_bufx10_ice8p I479 ( .in(cram_rst), .out(net247));
sg_bufx10_ice8p I465 ( .in(data_muxsel1_blbrd), .out(predata_muxsel1));
sg_bufx10_ice8p I525 ( .in(cm_clk_blbrd), .out(predata_smc_clk_out));
sg_bufx10_ice8p I518 ( .in(cm_banksel[1]), .out(net305));
sg_bufx10_ice8p I524 ( .in(predata_smc_clk_out), .out(smc_clk_mid));
sg_bufx10_ice8p I470 ( .in(net347), .out(cram_wl_enl0));
sg_bufx10_ice8p I511 ( .in(row_test0), .out(net325));
sg_bufx10_ice8p I293 ( .in(last_rsr1), .out(last_rsr2));
sg_bufx10_ice8p I541_1_ ( .in(dff_u0_d1[1]), .out(cm_sdo_u0d1[1]));
sg_bufx10_ice8p I541_0_ ( .in(dff_u0_d1[0]), .out(cm_sdo_u0d1[0]));
sg_bufx10_ice8p I539_1_ ( .in(cm_sdo_u1d1[1]), .out(cm_sdo_u1_buf[1]));
sg_bufx10_ice8p I539_0_ ( .in(cm_sdo_u1d1[0]), .out(cm_sdo_u1_buf[0]));
sg_bufx10_ice8p I455 ( .in(data_muxsel_blbrd), .out(predata_muxsel));
sg_bufx10_ice8p I526_1_ ( .in(cm_sdi_u2d[1]), .out(cm_sdi_u2d_buf[1]));
sg_bufx10_ice8p I526_0_ ( .in(cm_sdi_u2d[0]), .out(cm_sdi_u2d_buf[0]));
sg_bufx10_ice8p I569 ( .in(net361), .out(net289));
sg_bufx10_ice8p I477 ( .in(net363), .out(net319));
sg_bufx10_ice8p I566 ( .in(net387), .out(last_rsr3));
sg_bufx10_ice8p I540_1_ ( .in(dff_u1_d1[1]), .out(cm_sdo_u1d3[1]));
sg_bufx10_ice8p I540_0_ ( .in(dff_u1_d1[0]), .out(cm_sdo_u1d3[0]));
sg_bufx10_ice8p I497 ( .in(smc_wdis_dclk_blbrd),
     .out(predata_smc_wdis_dclk));
sg_bufx10_ice8p I487 ( .in(predata_cram_prec), .out(net293));
sg_bufx10_ice8p I498 ( .in(net373), .out(smc_wdis_dclk_blbld));
sg_bufx10_ice8p I499 ( .in(predata_smc_wdis_dclk), .out(net373));
sg_bufx10_ice8p I330 ( .in(net377), .out(net313));
sg_bufx10_ice8p I472 ( .in(cram_wl_en), .out(net323));
sg_dffbuf_modified I462_1_ ( .d(cm_sdo_u0_buf[1]), .clk(smc_clk_mid),
     .dffout(dff_u0_d1[1]), .r(net229[0]));
sg_dffbuf_modified I462_0_ ( .d(cm_sdo_u0_buf[0]), .clk(smc_clk_mid),
     .dffout(dff_u0_d1[0]), .r(net229[1]));
sg_dffbuf_modified I565 ( .d(last_rsr2), .clk(smc_clk_mid),
     .dffout(net387), .r(net232));
sg_dffbuf_modified I537_1_ ( .d(cm_sdo_u1_buf[1]), .clk(smc_clk_mid),
     .dffout(dff_u1_d1[1]), .r(net234[0]));
sg_dffbuf_modified I537_0_ ( .d(cm_sdo_u1_buf[0]), .clk(smc_clk_mid),
     .dffout(dff_u1_d1[0]), .r(net234[1]));
sg_dffbuf_modified I545_1_ ( .d(dff_u2_d0[1]),
     .clk(predata_smc_clk_out), .dffout(cm_sdo_u2d1[1]), .r(net231));
sg_dffbuf_modified I545_0_ ( .d(dff_u2_d0[0]),
     .clk(predata_smc_clk_out), .dffout(cm_sdo_u2d1[0]), .r(net231));
sg_dffbuf_modified I546_1_ ( .d(cm_sdo_u2[1]),
     .clk(predata_smc_clk_out), .dffout(dff_u2_d0[1]), .r(net230));
sg_dffbuf_modified I546_0_ ( .d(cm_sdo_u2[0]),
     .clk(predata_smc_clk_out), .dffout(dff_u2_d0[0]), .r(net230));
sg_dffbuf_modified I535_1_ ( .d(cm_sdo_u0[1]), .clk(cm_clk_blbld),
     .dffout(cm_sdo_u0_buf[1]), .r(net233[0]));
sg_dffbuf_modified I535_0_ ( .d(cm_sdo_u0[0]), .clk(cm_clk_blbld),
     .dffout(cm_sdo_u0_buf[0]), .r(net233[1]));
eh_io_pup_2_new_ice8p Ipor_spi ( .core_por_b(core_por_b0),
     .vdd_io(vddio_spi), .por_b(smc_core_por_bottom2));
eh_io_pup_2_new_ice8p Ipor_iob ( .core_por_b(core_por_b0),
     .vdd_io(vddio_botbank), .por_b(smc_core_por_bottom1));

endmodule
// Library - ice1chip, Cell - ring_route00_ice1f_june, View - schematic
// LAST TIME SAVED: Jun 29 09:50:50 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ring_route00_ice1f_june ( bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     end_of_startup, gint_hz, gsr, hiz_b0, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr,
     md_spi_b, mode0, mux_jtag_sel_b, pgate_l, pgate_r, reset_b_l,
     reset_b_r, sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_pad, update0, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r, bl_bot, bl_top, vppin, bm_sdo_o, cdone_in, creset_b_int,
     fabric_out_12_00, fabric_out_13_01, fabric_out_13_02, fromsdo,
     spi_ss_in_bbank, tck_pad, tdi_pad, tms_pad, trstb_pad,
     vddio_bottombank, vddio_spi );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     end_of_startup, gint_hz, gsr, hiz_b0, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, mux_jtag_sel_b, sdo_enable, shift0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, tdo_pad, update0;

inout  vppin;

input  cdone_in, creset_b_int, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fromsdo, tck_pad, tdi_pad, tms_pad, trstb_pad,
     vddio_bottombank, vddio_spi;

output [287:0]  wl_r;
output [287:0]  vdd_cntl_l;
output [287:0]  wl_l;
output [287:0]  pgate_l;
output [287:0]  reset_b_r;
output [3:0]  last_rsr;
output [287:0]  vdd_cntl_r;
output [7:0]  bm_sa_i;
output [3:0]  bm_sdi_i;
output [287:0]  reset_b_l;
output [3:0]  bm_banksel_i;
output [287:0]  pgate_r;

inout [663:0]  bl_top;
inout [663:0]  bl_bot;

input [3:0]  bm_sdo_o;
input [4:0]  spi_ss_in_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1d1;

wire  [1:0]  cm_sdi_u3d2;

wire  [1:0]  cm_sdi_u1d;

wire  [1:0]  cm_sdo_u1d3;

wire  [1:0]  cm_sdi_u1d3;

wire  [1:0]  cm_sdo_u2d1;

wire  [1:0]  cm_banksel;

wire  [1:0]  cm_sdo_u0d1;

wire  [1:0]  cm_sdo_u3;

wire  [3:3]  cm_banksel_bltrd1;

wire  [4:0]  spi_ss_in_bbankd;

wire  [1:0]  cm_sdi_u1;

wire  [1:1]  cm_banksel_bltld3;

wire  [1:0]  cm_sdo_u1;

wire  [1:0]  cm_sdi_u2d;

wire  [1:0]  cm_sdi_u0;



nvcm_ml_block_ice1f_june I_nvcm_ml_block_ice1f_june (
     .tgnd_fsm(tgnd_fsm), .tvdd_fsm(tvdd_fsm),
     .spi_ss_b(nvcm_spi_ss_b), .spi_sdi(nvcm_spi_sdi), .rst_b(rst_b),
     .nvcm_ce_b(cdone_in), .clk(spi_clk_out2fsm),
     .spi_sdo_oe_b(nvcm_spi_sdo_oe_b), .spi_sdo(nvcm_spi_sdo),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream),
     .fsm_tm_margin0_read(net398), .fsm_recall(net399), .bp0(bp0),
     .vpp(vppin), .nvcm_relextspi(nvcm_relextspi));
CHIP_route_lft2rgt_ice1f_june I_CHIP_route_rgt_ice1f (
     bm_banksel_i[3:0], bm_init_i, bm_rcapmux_en_i, bm_sa_i[7:0],
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i[3:0], bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bs_en0, cdone_out, ceb0, cm_banksel_blbrd_2_,
     cm_banksel[1:0], cm_banksel_bltrd1[3], cm_clk_blbrd,
     cm_clk_bltrd1, cm_sdi_u0[1:0], cm_sdi_u1[1:0], cm_sdi_u2d[1:0],
     cm_sdi_u3d2[1:0], core_por_b0, net228, core_por_b_rowu3,
     core_por_bb, cram_pgateoff, cram_prec, cram_prec_bltrd1,
     cram_pullup_b, cram_pullup_b_bltrd1, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, cram_write_bltrd1, data_muxsel1_blbrd,
     data_muxsel1_bltld3, data_muxsel_blbrd, data_muxsel_bltrd1,
     en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1, end_of_startup,
     gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     last_rsr[3:2], md_spi_b, mode0, mux_jtag_sel_b, nvcm_spi_sdi,
     nvcm_spi_ss_b, pgate_r[287:0], reset_b_r[287:0], row_test0, rst_b,
     sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rsr, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1, smc_write,
     smc_write_bltl1d1r, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_pad, update0, vdd_cntl_r[287:0], wl_r[287:0],
     bm_sdo_o[3:0], bp0, cdone_in, cm_sdo_u0d1[1:0], cm_sdo_u1d3[1:0],
     cm_sdo_u2d1[1:0], cm_sdo_u3[1:0], creset_b_int, fabric_out_12_00,
     fabric_out_13_01, fabric_out_13_02, fromsdo, {tgnd_fsm, tgnd_fsm,
     tgnd_fsm, tvdd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm, tvdd_fsm,
     tgnd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm,
     tgnd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm, tvdd_fsm},
     last_rsr3, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, smc_core_por_bottom1, smc_core_por_bottom2,
     spi_ss_in_bbankd[4:0], tck_pad, tdi_pad, tms_pad, trstb_pad,
     vddp_);
CHIP_route_top_ice1f I_CHIP_route_top_ice1f ( .bl_top(bl_top[663:0]),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltld1),
     .data_muxsel1_bltrd1(data_muxsel1_bltld3),
     .data_muxsel1_bltld3(data_muxsel1_bltld1),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_bltld3),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1),
     .core_por_b_rowu3(core_por_b_rowu3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .cm_prec_bltld3(cm_prec_bltld3), .cm_clk_bltrd1(cm_clk_bltrd1),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cm_banksel_bltrd1(cm_banksel_bltrd1[3]),
     .cm_banksel_bltld3(cm_banksel_bltld3[1]),
     .cm_sdo_u3(cm_sdo_u3[1:0]), .cm_sdo_u1(cm_sdo_u1[1:0]),
     .smc_write_bltld3(smc_write_bltld3),
     .smc_write_bltl1d1(smc_write_bltl1d1r));
CHIP_route_lft_ice1f I_CHIP_route_lft_ice1f ( .pgate_l(pgate_l[287:0]),
     .reset_l(reset_b_l[287:0]), .vdd_cntl_l(vdd_cntl_l[287:0]),
     .wl_l(wl_l[287:0]), .smc_write_bltld3(smc_write_bltld3),
     .tck_padl0(tck_padl0), .smc_writel0(smc_writel0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .smc_rsr_rstl0(smc_rsr_rstl0), .smc_row_incl0(smc_row_incl0),
     .row_testl1(row_testl1), .j_rst_bl0(j_rst_bl0),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_wl_enl0(cram_wl_enl0),
     .cram_vddoffl0(cram_vddoffl0), .cram_rstl0(cram_rstl0),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld),
     .cram_pgateoffl0(cram_pgateoffl0), .core_por_bbl0(core_por_bbl0),
     .cm_sdo_u1(cm_sdo_u1[1:0]), .cm_sdi_u1d(cm_sdi_u1d[1:0]),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbld(cm_banksel_blbld_1_),
     .cm_banksel_blbld1(cm_banksel_blbld1_0_),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3),
     .last_rsr(last_rsr[1:0]), .last_rsr0(last_rsr0),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel_bltld3(data_muxsel_bltld1),
     .data_muxsel1_bltld3(data_muxsel1_bltld1),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_bltld3),
     .cram_prec_bltld3(cm_prec_bltld3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdo_u1d1(cm_sdo_u1d1[1:0]), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cm_banksel_bltld3_1_(cm_banksel_bltld3[1]));
CHIP_route_bot_ice1f I_CHIP_route_bot_ice1f ( .bl_bot(bl_bot[663:0]),
     .core_por_b2(core_por_b2),
     .spi_ss_in_bbankd(spi_ss_in_bbankd[4:0]),
     .spi_ss_in_bbank(spi_ss_in_bbank[4:0]), .vddio_spi(vddio_spi),
     .vddio_botbank(vddio_bottombank), .smc_write(smc_write),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_rsr_rst(smc_rsr_rsr), .smc_row_inc(smc_row_inc),
     .row_test0(row_test0), .last_rsr1(last_rsr0), .j_tck(j_tck),
     .j_rst_b(j_rst_b), .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_blbrd(data_muxsel1_blbrd), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff),
     .core_por_bb(core_por_bb), .core_por_b0(core_por_b0),
     .cm_sdo_u1d1(cm_sdo_u1d1[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .cm_clk_blbrd(cm_clk_blbrd),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .cm_banksel(cm_banksel[1:0]), .tck_padl0(tck_padl0),
     .smc_writel0(smc_writel0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .smc_rsr_rstl0(smc_rsr_rstl0), .smc_row_incl0(smc_row_incl0),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .row_testl1(row_testl1), .last_rsr3(last_rsr3),
     .j_rst_bl0(j_rst_bl0), .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_wl_enl0(cram_wl_enl0),
     .cram_vddoffl0(cram_vddoffl0), .cram_rstl0(cram_rstl0),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld),
     .cram_pgateoffl0(cram_pgateoffl0), .core_por_bbl0(core_por_bbl0),
     .cm_sdo_u2d1(cm_sdo_u2d1[1:0]), .cm_sdo_u1d3(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0d1(cm_sdo_u0d1[1:0]), .cm_sdi_u1d(cm_sdi_u1d[1:0]),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbld_1_(cm_banksel_blbld_1_),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1_0_));
sg_bufx10_ice8p I_clkbuf ( .in(spi_clk_out), .out(spi_clk_out2fsm));

endmodule
// Library - ice1chip, Cell - LVDS_INBUFFER_ice1f, View - schematic
// LAST TIME SAVED: Apr 20 16:11:20 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module LVDS_INBUFFER_ice1f ( indiff, in_padn, in_padp, vddio, cbit[2],
     cbit[3], cbit[4] );
output  indiff;

inout  in_padn, in_padp, vddio;


input [2:4]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor3_hvt I56 ( .B(net0113), .Y(net0161), .A(cbit[3]), .C(cbit[2]));
nch_25od33  M10 ( .D(net1132), .B(gnd_), .G(net1138), .S(gnd_));
nch_25od33  M8 ( .D(net1138), .B(gnd_), .G(comp_out_25), .S(gnd_));
nch_25od33  M1 ( .D(lvdsen_b_25), .B(gnd_), .G(lvdsen_25), .S(gnd_));
pch_25od33  M9 ( .D(net1138), .B(vddio), .G(comp_out_25), .S(vddio));
pch_25od33  M0 ( .D(comp_out_25), .B(vddio), .G(lvdsen_25), .S(vddio));
pch_25od33  M11 ( .D(net1132), .B(vddio), .G(net1138), .S(vddio));
pch_25od33  M18 ( .D(comp_out_25), .B(vddio), .G(in_padp),
     .S(net1180));
pch_25od33  M13 ( .D(net1180), .B(vddio), .G(net1203), .S(net1184));
pch_25od33  M12 ( .D(net1184), .B(vddio), .G(lvdsen_b_25), .S(vddio));
pch_25od33  M19 ( .D(net1203), .B(vddio), .G(in_padn), .S(net1180));
pch_25od33  M2 ( .D(lvdsen_b_25), .B(vddio), .G(lvdsen_25), .S(vddio));
inv_hvt I129 ( .A(net0161), .Y(net1191));
inv_hvt I131 ( .A(indiff_b), .Y(indiff));
inv_hvt I55 ( .A(cbit[4]), .Y(net0113));
nch_25  x8 ( .D(indiff_b), .B(GND_), .G(net1138), .S(gnd_));
nch_25  M17 ( .D(net1204), .B(gnd_), .G(lvdsen_25), .S(gnd_));
nch_25  M16 ( .D(net1212), .B(gnd_), .G(net1203), .S(net1204));
nch_25  M23 ( .D(net0153), .B(GND_), .G(net1132), .S(gnd_));
nch_25  M21 ( .D(net1203), .B(GND_), .G(in_padn), .S(net1212));
nch_25  M20 ( .D(comp_out_25), .B(GND_), .G(in_padp), .S(net1212));
nch_25  x20 ( .D(lvdsen_25), .B(GND_), .G(net1191), .S(gnd_));
nch_25  x19 ( .D(net1149), .B(GND_), .G(net0161), .S(gnd_));
pch_25  x18 ( .D(net1149), .B(vddio), .G(lvdsen_25), .S(vddio));
pch_25  M5 ( .D(lvdsen_25), .B(vddio), .G(net1149), .S(vddio));
pch_hvt  x12 ( .D(indiff_b), .B(vdd_), .G(net0153), .S(vdd_));
pch_hvt  x13 ( .D(net0153), .B(vdd_), .G(indiff_b), .S(vdd_));

endmodule
// Library - ice1chip, Cell - PLVDS_pair_525M, View - schematic
// LAST TIME SAVED: Jun  6 15:28:18 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module PLVDS_pair_525M ( c_n, c_p, PAD_n, PAD_p, POC, cbit, i_n, i_p,
     oen_n, oen_p, tiegnd, vddio );
output  c_n, c_p;

inout  PAD_n, PAD_p;

input  POC, i_n, i_p, oen_n, oen_p, tiegnd, vddio;

input [4:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



PDUW08SDGZ_G_NOR I_ppart_0 ( .IE(cbit[3]), .POC(POC), .indiff(indiff),
     .PAD4LVDS(in_padp_0), .VDDIO(vddio), .REN(cbit[1]), .PAD(PAD_p),
     .C(c_p), .OEN(oen_p), .I(i_p));
PDUW08SDGZ_G_NOR I_npart_1 ( .IE(cbit[2]), .POC(POC), .indiff(tiegnd),
     .PAD4LVDS(in_padn_1), .VDDIO(vddio), .REN(cbit[0]), .PAD(PAD_n),
     .C(c_n), .OEN(oen_n), .I(i_n));
LVDS_INBUFFER_ice1f I_LVDS_INBUFFER ( indiff, in_padn_1, in_padp_0,
     vddio, cbit[3], cbit[2], cbit[4]);

endmodule
// Library - misc, Cell - ABIWTCZ4, View - schematic
// LAST TIME SAVED: Jun  8 08:11:43 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ABIWTCZ4 ( LOCK, PLLOUT, BYPASS, DIVF0, DIVF1, DIVF2, DIVF3,
     DIVF4, DIVF5, DIVF6, DIVQ0, DIVQ1, DIVQ2, DIVR0, DIVR1, DIVR2,
     DIVR3, FB, FSE, RANGE0, RANGE1, RANGE2, REF, RESET, VDDA );
output  LOCK, PLLOUT;

input  BYPASS, DIVF0, DIVF1, DIVF2, DIVF3, DIVF4, DIVF5, DIVF6, DIVQ0,
     DIVQ1, DIVQ2, DIVR0, DIVR1, DIVR2, DIVR3, FB, FSE, RANGE0, RANGE1,
     RANGE2, REF, RESET, VDDA;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD1DGZ_G, View - schematic
// LAST TIME SAVED: Sep  3 14:17:09 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module PVDD1DGZ_G ( VDD );
inout  VDD;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD2DGZ_G, View - schematic
// LAST TIME SAVED: Sep  3 14:16:20 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module PVDD2DGZ_G ( VDDPST );
inout  VDDPST;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD2POC_G, View - schematic
// LAST TIME SAVED: Sep  3 14:39:22 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module PVDD2POC_G ( POC, VDDPST );
output  POC;

inout  VDDPST;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - sbox1, View - schematic
// LAST TIME SAVED: Jun 22 18:19:36 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox1 ( b, l, r, t, c, cb, prog );
inout  b, l, r, t;

input  prog;

input [7:0]  c;
input [7:0]  cb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



sbox1m3to1_icc I232 ( .in2(r), .cb(cb[7:6]), .op(t), .in0(l), .in1(b),
     .c(c[7:6]), .prog(prog));
sbox1m3to1_icc I230 ( .in2(r), .cb(cb[3:2]), .op(l), .in0(b), .in1(t),
     .c(c[3:2]), .prog(prog));
sbox1m3to1_icc I226 ( .in2(r), .cb(cb[1:0]), .op(b), .in0(l), .in1(t),
     .c(c[1:0]), .prog(prog));
sbox1m3to1_icc I231 ( .in2(b), .cb(cb[5:4]), .op(r), .in0(l), .in1(t),
     .c(c[5:4]), .prog(prog));

endmodule
// Library - io, Cell - PVSS3DGZ_G, View - schematic
// LAST TIME SAVED: Sep 17 14:47:58 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module PVSS3DGZ_G ( VDDPST, VSS );
inout  VDDPST, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - ice1chip, Cell - IO_lft_bank_ice1f_v2, View - schematic
// LAST TIME SAVED: Jun  6 15:30:14 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module IO_lft_bank_ice1f_v2 ( in, pll_lock, pllout, pad, ien, lvds_en,
     oen, out, pll_bypass, pll_cbit, pll_fb, pll_fse, pll_ref,
     pll_reset, ren, vdda );
output  pll_lock, pllout;


input  pll_bypass, pll_fb, pll_fse, pll_ref, pll_reset, vdda;

output [23:0]  in;

inout [23:0]  pad;

input [23:0]  ien;
input [23:0]  oen;
input [23:0]  ren;
input [11:0]  lvds_en;
input [23:0]  out;
input [16:0]  pll_cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  ienb;



PLVDS_pair_525M plvds_1_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[2]), .oen_n(oen[3]),
     .PAD_n(pad[3]), .c_p(in[2]), .c_n(in[3]), .PAD_p(pad[2]),
     .i_n(out[3]), .i_p(out[2]), .cbit({lvds_en[1], ienb[2], ienb[3],
     ren[2], ren[3]}));
PLVDS_pair_525M plvds_0_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[0]), .oen_n(oen[1]),
     .PAD_n(pad[1]), .c_p(in[0]), .c_n(in[1]), .PAD_p(pad[0]),
     .i_n(out[1]), .i_p(out[0]), .cbit({lvds_en[0], ienb[0], ienb[1],
     ren[0], ren[1]}));
PLVDS_pair_525M plvds2 ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[4]), .oen_n(oen[5]),
     .PAD_n(pad[5]), .c_p(in[4]), .c_n(in[5]), .PAD_p(pad[4]),
     .i_n(out[5]), .i_p(out[4]), .cbit({lvds_en[2], ienb[4], ienb[5],
     ren[4], ren[5]}));
PLVDS_pair_525M plvds_5_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[10]), .oen_n(oen[11]),
     .PAD_n(pad[11]), .c_p(in[10]), .c_n(in[11]), .PAD_p(pad[10]),
     .i_n(out[11]), .i_p(out[10]), .cbit({lvds_en[5], ienb[10],
     ienb[11], ren[10], ren[11]}));
PLVDS_pair_525M plvds_4_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[8]), .oen_n(oen[9]),
     .PAD_n(pad[9]), .c_p(in[8]), .c_n(in[9]), .PAD_p(pad[8]),
     .i_n(out[9]), .i_p(out[8]), .cbit({lvds_en[4], ienb[8], ienb[9],
     ren[8], ren[9]}));
PLVDS_pair_525M plvds_3_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[6]), .oen_n(oen[7]),
     .PAD_n(pad[7]), .c_p(in[6]), .c_n(in[7]), .PAD_p(pad[6]),
     .i_n(out[7]), .i_p(out[6]), .cbit({lvds_en[3], ienb[6], ienb[7],
     ren[6], ren[7]}));
PLVDS_pair_525M plvds6 ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[12]), .oen_n(oen[13]),
     .PAD_n(pad[13]), .c_p(in[12]), .c_n(in[13]), .PAD_p(pad[12]),
     .i_n(out[13]), .i_p(out[12]), .cbit({lvds_en[6], ienb[12],
     ienb[13], ren[12], ren[13]}));
PLVDS_pair_525M plvds_9_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[18]), .oen_n(oen[19]),
     .PAD_n(pad[19]), .c_p(in[18]), .c_n(in[19]), .PAD_p(pad[18]),
     .i_n(out[19]), .i_p(out[18]), .cbit({lvds_en[9], ienb[18],
     ienb[19], ren[18], ren[19]}));
PLVDS_pair_525M plvds_8_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[16]), .oen_n(oen[17]),
     .PAD_n(pad[17]), .c_p(in[16]), .c_n(in[17]), .PAD_p(pad[16]),
     .i_n(out[17]), .i_p(out[16]), .cbit({lvds_en[8], ienb[16],
     ienb[17], ren[16], ren[17]}));
PLVDS_pair_525M plvds_7_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[14]), .oen_n(oen[15]),
     .PAD_n(pad[15]), .c_p(in[14]), .c_n(in[15]), .PAD_p(pad[14]),
     .i_n(out[15]), .i_p(out[14]), .cbit({lvds_en[7], ienb[14],
     ienb[15], ren[14], ren[15]}));
PLVDS_pair_525M plvds_11_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[22]), .oen_n(oen[23]),
     .PAD_n(pad[23]), .c_p(in[22]), .c_n(in[23]), .PAD_p(pad[22]),
     .i_n(out[23]), .i_p(out[22]), .cbit({lvds_en[11], ienb[22],
     ienb[23], ren[22], ren[23]}));
PLVDS_pair_525M plvds_10_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[20]), .oen_n(oen[21]),
     .PAD_n(pad[21]), .c_p(in[20]), .c_n(in[21]), .PAD_p(pad[20]),
     .i_n(out[21]), .i_p(out[20]), .cbit({lvds_en[10], ienb[20],
     ienb[21], ren[20], ren[21]}));
ABIWTCZ4 Ipll_bot ( .RESET(pll_reset), .REF(pll_ref),
     .RANGE2(pll_cbit[16]), .RANGE1(pll_cbit[15]),
     .RANGE0(pll_cbit[14]), .FSE(pll_fse), .FB(pll_fb),
     .DIVR3(pll_cbit[3]), .DIVR2(pll_cbit[2]), .DIVR1(pll_cbit[1]),
     .DIVR0(pll_cbit[0]), .DIVQ2(pll_cbit[13]), .DIVQ1(pll_cbit[12]),
     .DIVQ0(pll_cbit[11]), .DIVF5(pll_cbit[9]), .DIVF4(pll_cbit[8]),
     .DIVF3(pll_cbit[7]), .DIVF2(pll_cbit[6]), .DIVF1(pll_cbit[5]),
     .DIVF0(pll_cbit[4]), .BYPASS(pll_bypass), .PLLOUT(pllout),
     .LOCK(pll_lock), .VDDA(vdda), .DIVF6(pll_cbit[10]));
tielo4x I119 ( .tielo(tiegnd_lftpad));
inv_hvt I120_23_ ( .A(ien[23]), .Y(ienb[23]));
inv_hvt I120_22_ ( .A(ien[22]), .Y(ienb[22]));
inv_hvt I120_21_ ( .A(ien[21]), .Y(ienb[21]));
inv_hvt I120_20_ ( .A(ien[20]), .Y(ienb[20]));
inv_hvt I120_19_ ( .A(ien[19]), .Y(ienb[19]));
inv_hvt I120_18_ ( .A(ien[18]), .Y(ienb[18]));
inv_hvt I120_17_ ( .A(ien[17]), .Y(ienb[17]));
inv_hvt I120_16_ ( .A(ien[16]), .Y(ienb[16]));
inv_hvt I120_15_ ( .A(ien[15]), .Y(ienb[15]));
inv_hvt I120_14_ ( .A(ien[14]), .Y(ienb[14]));
inv_hvt I120_13_ ( .A(ien[13]), .Y(ienb[13]));
inv_hvt I120_12_ ( .A(ien[12]), .Y(ienb[12]));
inv_hvt I120_11_ ( .A(ien[11]), .Y(ienb[11]));
inv_hvt I120_10_ ( .A(ien[10]), .Y(ienb[10]));
inv_hvt I120_9_ ( .A(ien[9]), .Y(ienb[9]));
inv_hvt I120_8_ ( .A(ien[8]), .Y(ienb[8]));
inv_hvt I120_7_ ( .A(ien[7]), .Y(ienb[7]));
inv_hvt I120_6_ ( .A(ien[6]), .Y(ienb[6]));
inv_hvt I120_5_ ( .A(ien[5]), .Y(ienb[5]));
inv_hvt I120_4_ ( .A(ien[4]), .Y(ienb[4]));
inv_hvt I120_3_ ( .A(ien[3]), .Y(ienb[3]));
inv_hvt I120_2_ ( .A(ien[2]), .Y(ienb[2]));
inv_hvt I120_1_ ( .A(ien[1]), .Y(ienb[1]));
inv_hvt I120_0_ ( .A(ien[0]), .Y(ienb[0]));
PVDD1DGZ_G I129 ( .VDD(vdd_));
PVDD1DGZ_G I126_1_ ( .VDD(vdd_));
PVDD1DGZ_G I126_0_ ( .VDD(vdd_));
PVDD2DGZ_G I128 ( .VDDPST(vddio_leftbank));
PVDD2DGZ_G I121 ( .VDDPST(vddio_leftbank));
PVDD2DGZ_G I130 ( .VDDPST(vddio_leftbank));
PVDD2POC_G I122 ( .VDDPST(vddio_leftbank), .POC(poc_lft));
PVSS3DGZ_G gndummy12_1_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G gndummy12_0_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I123_1_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I123_0_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I127_1_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I127_0_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));

endmodule
// Library - misc, Cell - vpp_clamp_finger, View - schematic
// LAST TIME SAVED: Sep 17 15:01:43 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module vpp_clamp_finger ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .B(VSS), .D(net12), .G(VSS), .S(VSS));
nch_25  m1 ( .B(VSS), .D(VPP), .G(VDDIO), .S(net12));

endmodule
// Library - misc, Cell - vpp_clamp, View - schematic
// LAST TIME SAVED: Sep 17 14:58:48 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module vpp_clamp ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vpp_clamp_finger I0_3_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_2_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_1_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_0_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));

endmodule
// Library - io, Cell - pvpp, View - schematic
// LAST TIME SAVED: Oct  4 15:01:12 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module pvpp ( vpp, vppin );
inout  vpp, vppin;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I60_15_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_14_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_13_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_12_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_11_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_10_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_9_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_8_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_7_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_6_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_5_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_4_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_3_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_2_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_1_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_0_ ( .vddp_tieh(vddio_in));
rppolywo_m  R1 ( .MINUS(vpp), .PLUS(vppin), .BULK(gnd_));
vpp_clamp I59_15_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_14_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_13_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_12_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_11_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_10_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_9_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_8_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_7_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_6_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_5_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_4_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_3_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_2_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_1_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_0_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));

endmodule
// Library - ice1chip, Cell - IO_top_bank_ice1f, View - schematic
// LAST TIME SAVED: Jun  2 08:13:15 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module IO_top_bank_ice1f ( in, pad, vpp, vppin, ien, oen, out, ren );

inout  vpp, vppin;


output [23:0]  in;

inout [23:0]  pad;

input [23:0]  out;
input [23:0]  ren;
input [23:0]  oen;
input [23:0]  ien;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  n_ienb;

wire  [0:1]  net143;

wire  [0:3]  net223;

wire  [0:5]  net0166;

wire  [0:10]  net217;



tielo4x tielo4x_t ( .tielo(tiegnd_toppad));
pvpp vppfast_t ( .vppin(vppin), .vpp(vpp));
inv_hvt ien_inv_23_ ( .A(ien[23]), .Y(n_ienb[23]));
inv_hvt ien_inv_22_ ( .A(ien[22]), .Y(n_ienb[22]));
inv_hvt ien_inv_21_ ( .A(ien[21]), .Y(n_ienb[21]));
inv_hvt ien_inv_20_ ( .A(ien[20]), .Y(n_ienb[20]));
inv_hvt ien_inv_19_ ( .A(ien[19]), .Y(n_ienb[19]));
inv_hvt ien_inv_18_ ( .A(ien[18]), .Y(n_ienb[18]));
inv_hvt ien_inv_17_ ( .A(ien[17]), .Y(n_ienb[17]));
inv_hvt ien_inv_16_ ( .A(ien[16]), .Y(n_ienb[16]));
inv_hvt ien_inv_15_ ( .A(ien[15]), .Y(n_ienb[15]));
inv_hvt ien_inv_14_ ( .A(ien[14]), .Y(n_ienb[14]));
inv_hvt ien_inv_13_ ( .A(ien[13]), .Y(n_ienb[13]));
inv_hvt ien_inv_12_ ( .A(ien[12]), .Y(n_ienb[12]));
inv_hvt ien_inv_11_ ( .A(ien[11]), .Y(n_ienb[11]));
inv_hvt ien_inv_10_ ( .A(ien[10]), .Y(n_ienb[10]));
inv_hvt ien_inv_9_ ( .A(ien[9]), .Y(n_ienb[9]));
inv_hvt ien_inv_8_ ( .A(ien[8]), .Y(n_ienb[8]));
inv_hvt ien_inv_7_ ( .A(ien[7]), .Y(n_ienb[7]));
inv_hvt ien_inv_6_ ( .A(ien[6]), .Y(n_ienb[6]));
inv_hvt ien_inv_5_ ( .A(ien[5]), .Y(n_ienb[5]));
inv_hvt ien_inv_4_ ( .A(ien[4]), .Y(n_ienb[4]));
inv_hvt ien_inv_3_ ( .A(ien[3]), .Y(n_ienb[3]));
inv_hvt ien_inv_2_ ( .A(ien[2]), .Y(n_ienb[2]));
inv_hvt ien_inv_1_ ( .A(ien[1]), .Y(n_ienb[1]));
inv_hvt ien_inv_0_ ( .A(ien[0]), .Y(n_ienb[0]));
PVDD1DGZ_G vdd12_t_1_ ( .VDD(vdd_));
PVDD1DGZ_G vdd12_t_0_ ( .VDD(vdd_));
PVDD2POC_G vddio_poc2_t ( .VDDPST(vddio_topbank), .POC(poc_top));
PVDD2DGZ_G vcciodummy12_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vcciodummy12_0_ ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vddio1_t ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vddio34_t_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vddio34_t_0_ ( .VDDPST(vddio_topbank));
PVSS3DGZ_G gnddummy12_1_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnddummy12_0_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnddummy34_1_ ( .VSS(gnd_), .VDDPST(vddp_));
PVSS3DGZ_G gnddummy34_0_ ( .VSS(gnd_), .VDDPST(vddp_));
PVSS3DGZ_G gnd23_t_1_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnd23_t_0_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnd1_t ( .VSS(gnd_), .VDDPST(vddio_topbank));
PDUW08SDGZ_G_NOR pad_t_10_ ( .REN(ren[10]), .C(in[10]), .OEN(oen[10]),
     .IE(n_ienb[10]), .I(out[10]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net173), .VDDIO(vddio_topbank), .PAD(pad[10]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_12_ ( .REN(ren[12]), .C(in[12]), .OEN(oen[12]),
     .IE(n_ienb[12]), .I(out[12]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net143[0]), .VDDIO(vddio_topbank), .PAD(pad[12]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_11_ ( .REN(ren[11]), .C(in[11]), .OEN(oen[11]),
     .IE(n_ienb[11]), .I(out[11]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net143[1]), .VDDIO(vddio_topbank), .PAD(pad[11]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_23_ ( .REN(ren[23]), .C(in[23]), .OEN(oen[23]),
     .IE(n_ienb[23]), .I(out[23]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[0]), .VDDIO(vddio_topbank), .PAD(pad[23]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_22_ ( .REN(ren[22]), .C(in[22]), .OEN(oen[22]),
     .IE(n_ienb[22]), .I(out[22]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[1]), .VDDIO(vddio_topbank), .PAD(pad[22]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_21_ ( .REN(ren[21]), .C(in[21]), .OEN(oen[21]),
     .IE(n_ienb[21]), .I(out[21]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[2]), .VDDIO(vddio_topbank), .PAD(pad[21]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_20_ ( .REN(ren[20]), .C(in[20]), .OEN(oen[20]),
     .IE(n_ienb[20]), .I(out[20]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[3]), .VDDIO(vddio_topbank), .PAD(pad[20]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_19_ ( .REN(ren[19]), .C(in[19]), .OEN(oen[19]),
     .IE(n_ienb[19]), .I(out[19]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[4]), .VDDIO(vddio_topbank), .PAD(pad[19]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_18_ ( .REN(ren[18]), .C(in[18]), .OEN(oen[18]),
     .IE(n_ienb[18]), .I(out[18]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[5]), .VDDIO(vddio_topbank), .PAD(pad[18]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_17_ ( .REN(ren[17]), .C(in[17]), .OEN(oen[17]),
     .IE(n_ienb[17]), .I(out[17]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[6]), .VDDIO(vddio_topbank), .PAD(pad[17]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_16_ ( .REN(ren[16]), .C(in[16]), .OEN(oen[16]),
     .IE(n_ienb[16]), .I(out[16]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[7]), .VDDIO(vddio_topbank), .PAD(pad[16]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_15_ ( .REN(ren[15]), .C(in[15]), .OEN(oen[15]),
     .IE(n_ienb[15]), .I(out[15]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[8]), .VDDIO(vddio_topbank), .PAD(pad[15]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_14_ ( .REN(ren[14]), .C(in[14]), .OEN(oen[14]),
     .IE(n_ienb[14]), .I(out[14]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[9]), .VDDIO(vddio_topbank), .PAD(pad[14]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_13_ ( .REN(ren[13]), .C(in[13]), .OEN(oen[13]),
     .IE(n_ienb[13]), .I(out[13]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[10]), .VDDIO(vddio_topbank), .PAD(pad[13]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_3_ ( .REN(ren[3]), .C(in[3]), .OEN(oen[3]),
     .IE(n_ienb[3]), .I(out[3]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[0]), .VDDIO(vddio_topbank), .PAD(pad[3]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_2_ ( .REN(ren[2]), .C(in[2]), .OEN(oen[2]),
     .IE(n_ienb[2]), .I(out[2]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[1]), .VDDIO(vddio_topbank), .PAD(pad[2]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_1_ ( .REN(ren[1]), .C(in[1]), .OEN(oen[1]),
     .IE(n_ienb[1]), .I(out[1]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[2]), .VDDIO(vddio_topbank), .PAD(pad[1]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_0_ ( .REN(ren[0]), .C(in[0]), .OEN(oen[0]),
     .IE(n_ienb[0]), .I(out[0]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[3]), .VDDIO(vddio_topbank), .PAD(pad[0]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_9_ ( .REN(ren[9]), .C(in[9]), .OEN(oen[9]),
     .IE(n_ienb[9]), .I(out[9]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[0]), .VDDIO(vddio_topbank), .PAD(pad[9]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_8_ ( .REN(ren[8]), .C(in[8]), .OEN(oen[8]),
     .IE(n_ienb[8]), .I(out[8]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[1]), .VDDIO(vddio_topbank), .PAD(pad[8]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_7_ ( .REN(ren[7]), .C(in[7]), .OEN(oen[7]),
     .IE(n_ienb[7]), .I(out[7]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[2]), .VDDIO(vddio_topbank), .PAD(pad[7]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_6_ ( .REN(ren[6]), .C(in[6]), .OEN(oen[6]),
     .IE(n_ienb[6]), .I(out[6]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[3]), .VDDIO(vddio_topbank), .PAD(pad[6]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_5_ ( .REN(ren[5]), .C(in[5]), .OEN(oen[5]),
     .IE(n_ienb[5]), .I(out[5]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[4]), .VDDIO(vddio_topbank), .PAD(pad[5]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_4_ ( .REN(ren[4]), .C(in[4]), .OEN(oen[4]),
     .IE(n_ienb[4]), .I(out[4]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[5]), .VDDIO(vddio_topbank), .PAD(pad[4]),
     .POC(poc_top));

endmodule
// Library - TSMC_IO, Cell - PDDW08SDGZ_G, View - schematic
// LAST TIME SAVED: Oct  4 08:25:43 2010
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module PDDW08SDGZ_G ( C, PAD, I, OEN, POC, REN, VDDIO );
output  C;

inout  PAD;

input  I, OEN, POC, REN, VDDIO;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - ice1chip, Cell - IO_rgt_bank_ice1f, View - schematic
// LAST TIME SAVED: Jun  2 08:10:14 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module IO_rgt_bank_ice1f ( in, trstb_int, pad, TRSTb, ien, oen, out,
     ren );
output  trstb_int;


input  TRSTb;

output [24:0]  in;

inout [24:0]  pad;

input [24:0]  ien;
input [24:0]  out;
input [24:0]  oen;
input [25:0]  ren;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net117;

wire  [0:1]  net110;

wire  [24:0]  n_ienb;

wire  [0:1]  net184;

wire  [0:1]  net154;

wire  [0:4]  net144;

wire  [0:3]  net164;

wire  [0:3]  net134;

wire  [0:3]  net115;



tielo4x tielo4x_r ( .tielo(tiegnd_rgtpad));
tiehi4x tiehi4x_r ( .tiehi(tievdd_rgtpad));
inv_hvt I_ien_inv_24_ ( .A(ien[24]), .Y(n_ienb[24]));
inv_hvt I_ien_inv_23_ ( .A(ien[23]), .Y(n_ienb[23]));
inv_hvt I_ien_inv_22_ ( .A(ien[22]), .Y(n_ienb[22]));
inv_hvt I_ien_inv_21_ ( .A(ien[21]), .Y(n_ienb[21]));
inv_hvt I_ien_inv_20_ ( .A(ien[20]), .Y(n_ienb[20]));
inv_hvt I_ien_inv_19_ ( .A(ien[19]), .Y(n_ienb[19]));
inv_hvt I_ien_inv_18_ ( .A(ien[18]), .Y(n_ienb[18]));
inv_hvt I_ien_inv_17_ ( .A(ien[17]), .Y(n_ienb[17]));
inv_hvt I_ien_inv_16_ ( .A(ien[16]), .Y(n_ienb[16]));
inv_hvt I_ien_inv_15_ ( .A(ien[15]), .Y(n_ienb[15]));
inv_hvt I_ien_inv_14_ ( .A(ien[14]), .Y(n_ienb[14]));
inv_hvt I_ien_inv_13_ ( .A(ien[13]), .Y(n_ienb[13]));
inv_hvt I_ien_inv_12_ ( .A(ien[12]), .Y(n_ienb[12]));
inv_hvt I_ien_inv_11_ ( .A(ien[11]), .Y(n_ienb[11]));
inv_hvt I_ien_inv_10_ ( .A(ien[10]), .Y(n_ienb[10]));
inv_hvt I_ien_inv_9_ ( .A(ien[9]), .Y(n_ienb[9]));
inv_hvt I_ien_inv_8_ ( .A(ien[8]), .Y(n_ienb[8]));
inv_hvt I_ien_inv_7_ ( .A(ien[7]), .Y(n_ienb[7]));
inv_hvt I_ien_inv_6_ ( .A(ien[6]), .Y(n_ienb[6]));
inv_hvt I_ien_inv_5_ ( .A(ien[5]), .Y(n_ienb[5]));
inv_hvt I_ien_inv_4_ ( .A(ien[4]), .Y(n_ienb[4]));
inv_hvt I_ien_inv_3_ ( .A(ien[3]), .Y(n_ienb[3]));
inv_hvt I_ien_inv_2_ ( .A(ien[2]), .Y(n_ienb[2]));
inv_hvt I_ien_inv_1_ ( .A(ien[1]), .Y(n_ienb[1]));
inv_hvt I_ien_inv_0_ ( .A(ien[0]), .Y(n_ienb[0]));
PDDW08SDGZ_G trstb_r ( .REN(ren[25]), .C(trstb_int),
     .OEN(tievdd_rgtpad), .I(tiegnd_rgtpad), .VDDIO(vddio_rgtbank),
     .PAD(TRSTb), .POC(poc_rgt));
PVDD1DGZ_G vdd12_r_1_ ( .VDD(vdd_));
PVDD1DGZ_G vdd12_r_0_ ( .VDD(vdd_));
PDUW08SDGZ_G_NOR pad_r_13_ ( .REN(ren[13]), .C(in[13]), .OEN(oen[13]),
     .IE(n_ienb[13]), .I(out[13]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net154[0]), .VDDIO(vddio_rgtbank), .PAD(pad[13]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_12_ ( .REN(ren[12]), .C(in[12]), .OEN(oen[12]),
     .IE(n_ienb[12]), .I(out[12]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net154[1]), .VDDIO(vddio_rgtbank), .PAD(pad[12]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_7_ ( .REN(ren[7]), .C(in[7]), .OEN(oen[7]),
     .IE(n_ienb[7]), .I(out[7]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[0]), .VDDIO(vddio_rgtbank), .PAD(pad[7]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_6_ ( .REN(ren[6]), .C(in[6]), .OEN(oen[6]),
     .IE(n_ienb[6]), .I(out[6]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[1]), .VDDIO(vddio_rgtbank), .PAD(pad[6]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_5_ ( .REN(ren[5]), .C(in[5]), .OEN(oen[5]),
     .IE(n_ienb[5]), .I(out[5]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[2]), .VDDIO(vddio_rgtbank), .PAD(pad[5]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_4_ ( .REN(ren[4]), .C(in[4]), .OEN(oen[4]),
     .IE(n_ienb[4]), .I(out[4]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[3]), .VDDIO(vddio_rgtbank), .PAD(pad[4]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_3_ ( .REN(ren[3]), .C(in[3]), .OEN(oen[3]),
     .IE(n_ienb[3]), .I(out[3]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[0]), .VDDIO(vddio_rgtbank), .PAD(pad[3]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_2_ ( .REN(ren[2]), .C(in[2]), .OEN(oen[2]),
     .IE(n_ienb[2]), .I(out[2]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[1]), .VDDIO(vddio_rgtbank), .PAD(pad[2]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_1_ ( .REN(ren[1]), .C(in[1]), .OEN(oen[1]),
     .IE(n_ienb[1]), .I(out[1]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[2]), .VDDIO(vddio_rgtbank), .PAD(pad[1]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_0_ ( .REN(ren[0]), .C(in[0]), .OEN(oen[0]),
     .IE(n_ienb[0]), .I(out[0]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[3]), .VDDIO(vddio_rgtbank), .PAD(pad[0]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_9_ ( .REN(ren[9]), .C(in[9]), .OEN(oen[9]),
     .IE(n_ienb[9]), .I(out[9]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net184[0]), .VDDIO(vddio_rgtbank), .PAD(pad[9]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_8_ ( .REN(ren[8]), .C(in[8]), .OEN(oen[8]),
     .IE(n_ienb[8]), .I(out[8]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net184[1]), .VDDIO(vddio_rgtbank), .PAD(pad[8]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_11_ ( .REN(ren[11]), .C(in[11]), .OEN(oen[11]),
     .IE(n_ienb[11]), .I(out[11]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net117[0]), .VDDIO(vddio_rgtbank), .PAD(pad[11]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_10_ ( .REN(ren[10]), .C(in[10]), .OEN(oen[10]),
     .IE(n_ienb[10]), .I(out[10]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net117[1]), .VDDIO(vddio_rgtbank), .PAD(pad[10]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_24_ ( .REN(ren[24]), .C(in[24]), .OEN(oen[24]),
     .IE(n_ienb[24]), .I(out[24]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[0]), .VDDIO(vddio_rgtbank), .PAD(pad[24]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_23_ ( .REN(ren[23]), .C(in[23]), .OEN(oen[23]),
     .IE(n_ienb[23]), .I(out[23]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[1]), .VDDIO(vddio_rgtbank), .PAD(pad[23]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_22_ ( .REN(ren[22]), .C(in[22]), .OEN(oen[22]),
     .IE(n_ienb[22]), .I(out[22]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[2]), .VDDIO(vddio_rgtbank), .PAD(pad[22]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_21_ ( .REN(ren[21]), .C(in[21]), .OEN(oen[21]),
     .IE(n_ienb[21]), .I(out[21]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[3]), .VDDIO(vddio_rgtbank), .PAD(pad[21]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_18_ ( .REN(ren[18]), .C(in[18]), .OEN(oen[18]),
     .IE(n_ienb[18]), .I(out[18]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[0]), .VDDIO(vddio_rgtbank), .PAD(pad[18]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_17_ ( .REN(ren[17]), .C(in[17]), .OEN(oen[17]),
     .IE(n_ienb[17]), .I(out[17]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[1]), .VDDIO(vddio_rgtbank), .PAD(pad[17]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_16_ ( .REN(ren[16]), .C(in[16]), .OEN(oen[16]),
     .IE(n_ienb[16]), .I(out[16]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[2]), .VDDIO(vddio_rgtbank), .PAD(pad[16]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_15_ ( .REN(ren[15]), .C(in[15]), .OEN(oen[15]),
     .IE(n_ienb[15]), .I(out[15]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[3]), .VDDIO(vddio_rgtbank), .PAD(pad[15]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_14_ ( .REN(ren[14]), .C(in[14]), .OEN(oen[14]),
     .IE(n_ienb[14]), .I(out[14]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[4]), .VDDIO(vddio_rgtbank), .PAD(pad[14]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_20_ ( .REN(ren[20]), .C(in[20]), .OEN(oen[20]),
     .IE(n_ienb[20]), .I(out[20]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net110[0]), .VDDIO(vddio_rgtbank), .PAD(pad[20]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_19_ ( .REN(ren[19]), .C(in[19]), .OEN(oen[19]),
     .IE(n_ienb[19]), .I(out[19]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net110[1]), .VDDIO(vddio_rgtbank), .PAD(pad[19]),
     .POC(poc_rgt));
PVDD2DGZ_G vcciodummy2 ( .VDDPST(vddp_));
PVDD2DGZ_G vddio12_r_1_ ( .VDDPST(vddio_rgtbank));
PVDD2DGZ_G vddio12_r_0_ ( .VDDPST(vddio_rgtbank));
PVDD2DGZ_G vddio2_r ( .VDDPST(vddio_rgtbank));
PVDD2DGZ_G vcciodummy1 ( .VDDPST(vddio_rgtbank));
PVDD2POC_G vddpoc_r ( .VDDPST(vddio_rgtbank), .POC(poc_rgt));
PVDD2POC_G vppv25_r ( .VDDPST(vddp_), .POC(net0123));
PVSS3DGZ_G gnd23_r_1_ ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnd23_r_0_ ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnddummy2 ( .VSS(gnd_), .VDDPST(vddp_));
PVSS3DGZ_G gnddummy1 ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnd3_r ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnd1_r ( .VSS(gnd_), .VDDPST(vddio_rgtbank));

endmodule
// Library - ice1chip, Cell - IO_bot_bank_ice1f, View - schematic
// LAST TIME SAVED: Jun  2 08:14:10 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module IO_bot_bank_ice1f ( cdone_int, ctst_b_int, in, vddio_bottombank,
     vddio_spi, cdone, pad, cdone_out, ctst_b, ien, oen, out, ren );
output  cdone_int, ctst_b_int, vddio_bottombank, vddio_spi;

inout  cdone;

input  cdone_out, ctst_b;

output [23:0]  in;

inout [23:0]  pad;

input [23:0]  ien;
input [23:0]  ren;
input [23:0]  oen;
input [23:0]  out;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  n_ienb;

wire  [0:1]  net168;

wire  [0:4]  net228;

wire  [0:1]  net237;

wire  [0:1]  net236;

wire  [0:1]  net234;

wire  [0:1]  net188;

wire  [0:7]  net241;



tiehi4x tiehi4x ( .tiehi(tievdd_botpad));
tielo4x tielo4x ( .tielo(tiegnd_botpad));
inv_hvt I_ien_inv_23_ ( .A(ien[23]), .Y(n_ienb[23]));
inv_hvt I_ien_inv_22_ ( .A(ien[22]), .Y(n_ienb[22]));
inv_hvt I_ien_inv_21_ ( .A(ien[21]), .Y(n_ienb[21]));
inv_hvt I_ien_inv_20_ ( .A(ien[20]), .Y(n_ienb[20]));
inv_hvt I_ien_inv_19_ ( .A(ien[19]), .Y(n_ienb[19]));
inv_hvt I_ien_inv_18_ ( .A(ien[18]), .Y(n_ienb[18]));
inv_hvt I_ien_inv_17_ ( .A(ien[17]), .Y(n_ienb[17]));
inv_hvt I_ien_inv_16_ ( .A(ien[16]), .Y(n_ienb[16]));
inv_hvt I_ien_inv_15_ ( .A(ien[15]), .Y(n_ienb[15]));
inv_hvt I_ien_inv_14_ ( .A(ien[14]), .Y(n_ienb[14]));
inv_hvt I_ien_inv_13_ ( .A(ien[13]), .Y(n_ienb[13]));
inv_hvt I_ien_inv_12_ ( .A(ien[12]), .Y(n_ienb[12]));
inv_hvt I_ien_inv_11_ ( .A(ien[11]), .Y(n_ienb[11]));
inv_hvt I_ien_inv_10_ ( .A(ien[10]), .Y(n_ienb[10]));
inv_hvt I_ien_inv_9_ ( .A(ien[9]), .Y(n_ienb[9]));
inv_hvt I_ien_inv_8_ ( .A(ien[8]), .Y(n_ienb[8]));
inv_hvt I_ien_inv_7_ ( .A(ien[7]), .Y(n_ienb[7]));
inv_hvt I_ien_inv_6_ ( .A(ien[6]), .Y(n_ienb[6]));
inv_hvt I_ien_inv_5_ ( .A(ien[5]), .Y(n_ienb[5]));
inv_hvt I_ien_inv_4_ ( .A(ien[4]), .Y(n_ienb[4]));
inv_hvt I_ien_inv_3_ ( .A(ien[3]), .Y(n_ienb[3]));
inv_hvt I_ien_inv_2_ ( .A(ien[2]), .Y(n_ienb[2]));
inv_hvt I_ien_inv_1_ ( .A(ien[1]), .Y(n_ienb[1]));
inv_hvt I_ien_inv_0_ ( .A(ien[0]), .Y(n_ienb[0]));
PVDD1DGZ_G vdd12_b_1_ ( .VDD(vdd_));
PVDD1DGZ_G vdd12_b_0_ ( .VDD(vdd_));
PVDD2POC_G vddiopoc2_b ( .VDDPST(vddio_bottombank), .POC(poc_bot));
PVDD2POC_G pvdd2poc_g_spivcc ( .VDDPST(vddio_spi), .POC(poc_spi));
PVDD2DGZ_G vddio3_b ( .VDDPST(vddio_bottombank));
PVDD2DGZ_G vcciodummy1 ( .VDDPST(vddio_bottombank));
PVDD2DGZ_G vddio1_b ( .VDDPST(vddio_bottombank));
PVDD2DGZ_G vcciodummy2 ( .VDDPST(vddio_spi));
PVSS3DGZ_G gnddummy1 ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd34_b_1_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd34_b_0_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd12_b_1_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd12_b_0_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnddummy2 ( .VSS(gnd_), .VDDPST(vddio_spi));
PVSS3DGZ_G gnd5 ( .VSS(gnd_), .VDDPST(vddio_spi));
PDUW08SDGZ_G_NOR pad_b_21_ ( .REN(ren[21]), .C(in[21]), .OEN(oen[21]),
     .IE(n_ienb[21]), .I(out[21]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net234[0]), .VDDIO(vddio_spi), .PAD(pad[21]),
     .POC(poc_spi));
PDUW08SDGZ_G_NOR pad_b_20_ ( .REN(ren[20]), .C(in[20]), .OEN(oen[20]),
     .IE(n_ienb[20]), .I(out[20]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net234[1]), .VDDIO(vddio_spi), .PAD(pad[20]),
     .POC(poc_spi));
PDUW08SDGZ_G_NOR pad_b_11_ ( .REN(ren[11]), .C(in[11]), .OEN(oen[11]),
     .IE(n_ienb[11]), .I(out[11]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net237[0]), .VDDIO(vddio_bottombank), .PAD(pad[11]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_10_ ( .REN(ren[10]), .C(in[10]), .OEN(oen[10]),
     .IE(n_ienb[10]), .I(out[10]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net237[1]), .VDDIO(vddio_bottombank), .PAD(pad[10]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_13_ ( .REN(ren[13]), .C(in[13]), .OEN(oen[13]),
     .IE(n_ienb[13]), .I(out[13]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net188[0]), .VDDIO(vddio_bottombank), .PAD(pad[13]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_12_ ( .REN(ren[12]), .C(in[12]), .OEN(oen[12]),
     .IE(n_ienb[12]), .I(out[12]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net188[1]), .VDDIO(vddio_bottombank), .PAD(pad[12]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_14_ ( .REN(ren[14]), .C(in[14]), .OEN(oen[14]),
     .IE(n_ienb[14]), .I(out[14]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net198), .VDDIO(vddio_bottombank), .PAD(pad[14]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_7_ ( .REN(ren[7]), .C(in[7]), .OEN(oen[7]),
     .IE(n_ienb[7]), .I(out[7]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[0]), .VDDIO(vddio_bottombank), .PAD(pad[7]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_6_ ( .REN(ren[6]), .C(in[6]), .OEN(oen[6]),
     .IE(n_ienb[6]), .I(out[6]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[1]), .VDDIO(vddio_bottombank), .PAD(pad[6]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_5_ ( .REN(ren[5]), .C(in[5]), .OEN(oen[5]),
     .IE(n_ienb[5]), .I(out[5]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[2]), .VDDIO(vddio_bottombank), .PAD(pad[5]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_4_ ( .REN(ren[4]), .C(in[4]), .OEN(oen[4]),
     .IE(n_ienb[4]), .I(out[4]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[3]), .VDDIO(vddio_bottombank), .PAD(pad[4]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_3_ ( .REN(ren[3]), .C(in[3]), .OEN(oen[3]),
     .IE(n_ienb[3]), .I(out[3]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[4]), .VDDIO(vddio_bottombank), .PAD(pad[3]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_2_ ( .REN(ren[2]), .C(in[2]), .OEN(oen[2]),
     .IE(n_ienb[2]), .I(out[2]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[5]), .VDDIO(vddio_bottombank), .PAD(pad[2]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_1_ ( .REN(ren[1]), .C(in[1]), .OEN(oen[1]),
     .IE(n_ienb[1]), .I(out[1]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[6]), .VDDIO(vddio_bottombank), .PAD(pad[1]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_0_ ( .REN(ren[0]), .C(in[0]), .OEN(oen[0]),
     .IE(n_ienb[0]), .I(out[0]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[7]), .VDDIO(vddio_bottombank), .PAD(pad[0]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_9_ ( .REN(ren[9]), .C(in[9]), .OEN(oen[9]),
     .IE(n_ienb[9]), .I(out[9]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net236[0]), .VDDIO(vddio_bottombank), .PAD(pad[9]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_8_ ( .REN(ren[8]), .C(in[8]), .OEN(oen[8]),
     .IE(n_ienb[8]), .I(out[8]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net236[1]), .VDDIO(vddio_bottombank), .PAD(pad[8]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_19_ ( .REN(ren[19]), .C(in[19]), .OEN(oen[19]),
     .IE(n_ienb[19]), .I(out[19]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[0]), .VDDIO(vddio_bottombank), .PAD(pad[19]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_18_ ( .REN(ren[18]), .C(in[18]), .OEN(oen[18]),
     .IE(n_ienb[18]), .I(out[18]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[1]), .VDDIO(vddio_bottombank), .PAD(pad[18]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_17_ ( .REN(ren[17]), .C(in[17]), .OEN(oen[17]),
     .IE(n_ienb[17]), .I(out[17]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[2]), .VDDIO(vddio_bottombank), .PAD(pad[17]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_16_ ( .REN(ren[16]), .C(in[16]), .OEN(oen[16]),
     .IE(n_ienb[16]), .I(out[16]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[3]), .VDDIO(vddio_bottombank), .PAD(pad[16]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_15_ ( .REN(ren[15]), .C(in[15]), .OEN(oen[15]),
     .IE(n_ienb[15]), .I(out[15]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[4]), .VDDIO(vddio_bottombank), .PAD(pad[15]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR ctst_b_b ( .REN(tiegnd_botpad), .C(ctst_b_int),
     .OEN(tievdd_botpad), .IE(tievdd_botpad), .I(tiegnd_botpad),
     .indiff(tiegnd_botpad), .PAD4LVDS(net233),
     .VDDIO(vddio_bottombank), .PAD(ctst_b), .POC(poc_bot));
PDUW08SDGZ_G_NOR cdone_b ( .REN(tiegnd_botpad), .C(cdone_int),
     .OEN(cdone_out), .IE(tievdd_botpad), .I(tiegnd_botpad),
     .indiff(tiegnd_botpad), .PAD4LVDS(net148),
     .VDDIO(vddio_bottombank), .PAD(cdone), .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_23_ ( .REN(ren[23]), .C(in[23]), .OEN(oen[23]),
     .IE(n_ienb[23]), .I(out[23]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net168[0]), .VDDIO(vddio_spi), .PAD(pad[23]),
     .POC(poc_spi));
PDUW08SDGZ_G_NOR pad_b_22_ ( .REN(ren[22]), .C(in[22]), .OEN(oen[22]),
     .IE(n_ienb[22]), .I(out[22]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net168[1]), .VDDIO(vddio_spi), .PAD(pad[22]),
     .POC(poc_spi));

endmodule
// Library - ice1chip, Cell - padring_ice1f, View - schematic
// LAST TIME SAVED: Jun  2 08:15:39 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module padring_ice1f ( cdone_int, creset_b_int, in_bbank, in_lbank,
     in_rbank, in_tbank, pll_lock, pllout, trstb_int_pad,
     vddio_bottombank, vddio_spi, cdone, uio_bbank, uio_lbank,
     uio_rbank, uio_tbank, vpp, vppin, cdone_out, creset_b, ien,
     ien_bbank, ien_rbank, ien_tbank, lvds_en, oen_bbank, oen_lbank,
     oen_rbank, oen_tbank, out_bbank, out_lbank, out_rbank, out_tbank,
     pll_bypass, pll_cbit, pll_fb, pll_fse, pll_ref, pll_reset, ren,
     ren_bbank, ren_rbank, ren_tbank, trstb, vdda );
output  cdone_int, creset_b_int, pll_lock, pllout, trstb_int_pad,
     vddio_bottombank, vddio_spi;

inout  cdone, vpp, vppin;

input  cdone_out, creset_b, pll_bypass, pll_fb, pll_fse, pll_ref,
     pll_reset, trstb, vdda;

output [24:0]  in_rbank;
output [23:0]  in_tbank;
output [23:0]  in_bbank;
output [23:0]  in_lbank;

inout [23:0]  uio_tbank;
inout [24:0]  uio_rbank;
inout [23:0]  uio_bbank;
inout [23:0]  uio_lbank;

input [23:0]  out_tbank;
input [24:0]  out_rbank;
input [23:0]  out_bbank;
input [23:0]  ien_tbank;
input [24:0]  ien_rbank;
input [25:0]  ren_rbank;
input [16:0]  pll_cbit;
input [23:0]  ren_bbank;
input [23:0]  ren;
input [11:0]  lvds_en;
input [23:0]  ien_bbank;
input [23:0]  out_lbank;
input [23:0]  oen_tbank;
input [23:0]  ren_tbank;
input [23:0]  ien;
input [23:0]  oen_bbank;
input [24:0]  oen_rbank;
input [23:0]  oen_lbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



IO_lft_bank_ice1f_v2 iobank_l ( .ien(ien[23:0]),
     .lvds_en(lvds_en[11:0]), .ren(ren[23:0]), .pad(uio_lbank[23:0]),
     .in(in_lbank[23:0]), .oen(oen_lbank[23:0]), .out(out_lbank[23:0]),
     .vdda(vdda), .pll_ref(pll_ref), .pll_fse(pll_fse),
     .pll_cbit(pll_cbit[16:0]), .pll_fb(pll_fb),
     .pll_bypass(pll_bypass), .pll_lock(pll_lock), .pllout(pllout),
     .pll_reset(pll_reset));
IO_top_bank_ice1f iobank_t ( .vppin(vppin), .vpp(vpp),
     .ren(ren_tbank[23:0]), .out(out_tbank[23:0]),
     .oen(oen_tbank[23:0]), .ien(ien_tbank[23:0]), .in(in_tbank[23:0]),
     .pad(uio_tbank[23:0]));
IO_rgt_bank_ice1f iobank_r ( .ren(ren_rbank[25:0]),
     .ien(ien_rbank[24:0]), .oen(oen_rbank[24:0]), .in(in_rbank[24:0]),
     .pad(uio_rbank[24:0]), .out(out_rbank[24:0]), .TRSTb(trstb),
     .trstb_int(trstb_int_pad));
IO_bot_bank_ice1f iobank_b ( .vddio_bottombank(vddio_bottombank),
     .cdone_out(cdone_out), .ctst_b(creset_b), .ren(ren_bbank[23:0]),
     .out(out_bbank[23:0]), .oen(oen_bbank[23:0]),
     .ien(ien_bbank[23:0]), .in(in_bbank[23:0]), .pad(uio_bbank[23:0]),
     .vddio_spi(vddio_spi), .cdone(cdone), .cdone_int(cdone_int),
     .ctst_b_int(creset_b_int));

endmodule
// Library - xpmem, Cell - cram16x4, View - schematic
// LAST TIME SAVED: Jun 24 17:57:57 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module cram16x4 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [63:0]  q_b;
output [63:0]  q;

inout [3:0]  bl;

input [15:0]  r_gnd;
input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 I16_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[1:0]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[15:14]));
cram2x2 I16_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[1:0]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[13:12]));
cram2x2 I16_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[1:0]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[11:10]));
cram2x2 I16_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[1:0]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[9:8]));
cram2x2 I16_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[1:0]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[7:6]));
cram2x2 I16_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[1:0]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[5:4]));
cram2x2 I16_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[1:0]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[3:2]));
cram2x2 I16_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[3:2]), .q_b(q_b[63:60]),
     .q(q[63:60]), .wl(wl[15:14]));
cram2x2 Imstake_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[3:2]), .q_b(q_b[59:56]),
     .q(q[59:56]), .wl(wl[13:12]));
cram2x2 Imstake_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[3:2]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[11:10]));
cram2x2 Imstake_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[3:2]), .q_b(q_b[51:48]), .q(q[51:48]),
     .wl(wl[9:8]));
cram2x2 Imstake_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[3:2]), .q_b(q_b[47:44]), .q(q[47:44]),
     .wl(wl[7:6]));
cram2x2 Imstake_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[3:2]), .q_b(q_b[43:40]), .q(q[43:40]),
     .wl(wl[5:4]));
cram2x2 Imstake_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[3:2]), .q_b(q_b[39:36]), .q(q[39:36]),
     .wl(wl[3:2]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[35:32]), .q(q[35:32]),
     .wl(wl[1:0]));

endmodule
// Library - ice1chip, Cell - ring_route_ice1f, View - schematic
// LAST TIME SAVED: Jun 29 09:34:00 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module ring_route_ice1f ( bm_banksel_i, bm_init_i, bm_rcapmux_en_i,
     bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bs_en0, ceb0, end_of_startup, gint_hz, gsr,
     hiz_b0, in_bbank, in_lbank, in_rbank, in_tbank, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     .cdsNet0(last_rsr[1]), .cdsNet0(last_rsr[0]),
     .cdsNet0(last_rsr[3]), .cdsNet0(last_rsr[2]), md_spi_b, mode0,
     mux_jtag_sel_b, pgate_l, pgate_r, pll_lock, pllout, reset_l,
     reset_r, sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, trstb_pad, update0, vdd_cntl_l,
     vdd_cntl_r, wl_l, wl_r, bl_bot, bl_top, cdone, uio_bbank,
     uio_lbank, uio_rbank, uio_tbank, vpp, bm_sdo_o, creset_b,
     fabric_out_12_00, fabric_out_13_01, fabric_out_13_02, fromsdo,
     ien, ien_bbank, ien_rbank, ien_tbank, lvds_en, oen_bbank,
     oen_lbank, oen_rbank, oen_tbank, out_bbank, out_lbank, out_rbank,
     out_tbank, pll_bypass, pll_cbit, pll_fb, pll_fse, pll_ref,
     pll_reset, ren, ren_bbank, ren_rbank, ren_tbank, spi_ss_in_bbank,
     tck_pad, tdi_pad, tms_pad, trstb, vdda );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, ceb0, end_of_startup,
     gint_hz, gsr, hiz_b0, j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, md_spi_b, mode0, mux_jtag_sel_b,
     pll_lock, pllout, sdo_enable, shift0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, totdopad, trstb_pad, update0;

inout  cdone, vpp;

input  creset_b, fabric_out_12_00, fabric_out_13_01, fabric_out_13_02,
     fromsdo, pll_bypass, pll_fb, pll_fse, pll_ref, pll_reset, tck_pad,
     tdi_pad, tms_pad, trstb, vdda;

output [287:0]  vdd_cntl_r;
output [24:0]  in_rbank;
output [3:0]  bm_banksel_i;
output [3:0]  bm_sdi_i;
output [287:0]  pgate_l;
output [7:0]  bm_sa_i;
output [3:0]  last_rsr;
output [287:0]  pgate_r;
output [23:0]  in_bbank;
output [287:0]  reset_r;
output [287:0]  vdd_cntl_l;
output [287:0]  wl_l;
output [23:0]  in_lbank;
output [287:0]  wl_r;
output [287:0]  reset_l;
output [23:0]  in_tbank;

inout [663:0]  bl_top;
inout [23:0]  uio_tbank;
inout [663:0]  bl_bot;
inout [24:0]  uio_rbank;
inout [23:0]  uio_lbank;
inout [23:0]  uio_bbank;

input [24:0]  out_rbank;
input [3:0]  bm_sdo_o;
input [24:0]  ien_rbank;
input [24:0]  oen_rbank;
input [4:0]  spi_ss_in_bbank;
input [23:0]  out_tbank;
input [23:0]  oen_lbank;
input [23:0]  ien_bbank;
input [23:0]  out_lbank;
input [23:0]  ren;
input [23:0]  oen_tbank;
input [16:0]  pll_cbit;
input [25:0]  ren_rbank;
input [23:0]  out_bbank;
input [23:0]  oen_bbank;
input [11:0]  lvds_en;
input [23:0]  ien;
input [23:0]  ien_tbank;
input [23:0]  ren_tbank;
input [23:0]  ren_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ring_route00_ice1f_june I_ring_route00_ice1f (
     .spi_ss_in_bbank(spi_ss_in_bbank[4:0]),
     .fabric_out_12_00(fabric_out_12_00),
     .fabric_out_13_01(fabric_out_13_01),
     .fabric_out_13_02(fabric_out_13_02), .pgate_r(pgate_r[287:0]),
     .reset_b_r(reset_r[287:0]), .vdd_cntl_r(vdd_cntl_r[287:0]),
     .wl_r(wl_r[287:0]), .wl_l(wl_l[287:0]),
     .vdd_cntl_l(vdd_cntl_l[287:0]), .pgate_l(pgate_l[287:0]),
     .reset_b_l(reset_l[287:0]), .bl_top(bl_top[663:0]),
     .bl_bot(bl_bot[663:0]), .trstb_pad(trstb_pad), .tms_pad(tms_pad),
     .tdi_pad(tdi_pad), .tck_pad(tck_pad), .fromsdo(fromsdo),
     .creset_b_int(creset_b_int), .vddio_bottombank(vddio_bottombank),
     .vddio_spi(vddio_spi), .bm_sa_i(bm_sa_i[7:0]),
     .cdone_in(cdone_in), .bm_sdo_o(bm_sdo_o[3:0]), .vppin(vppin),
     .update0(update0), .tdo_pad(totdopad),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out), .shift0(shift0),
     .sdo_enable(sdo_enable), .mode0(mode0), .md_spi_b(md_spi_b),
     .last_rsr(last_rsr[3:0]),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .j_tdi(j_tdi), .j_tck(j_tck), .mux_jtag_sel_b(mux_jtag_sel_b),
     .hiz_b0(hiz_b0), .gsr(gsr), .gint_hz(gint_hz),
     .end_of_startup(end_of_startup), .ceb0(ceb0),
     .cdone_out(cdone_out), .bs_en0(bs_en0),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclk_i(bm_sclk_i),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bm_banksel_i(bm_banksel_i[3:0]));
padring_ice1f I_padring_ice1f ( .ien(ien[23:0]),
     .lvds_en(lvds_en[11:0]), .ren(ren[23:0]),
     .uio_lbank(uio_lbank[23:0]), .oen_lbank(oen_lbank[23:0]),
     .out_lbank(out_lbank[23:0]), .in_lbank(in_lbank[23:0]),
     .vdda(vdda), .pll_lock(pll_lock), .pllout(pllout),
     .pll_reset(pll_reset), .pll_bypass(pll_bypass), .pll_fb(pll_fb),
     .pll_cbit(pll_cbit[16:0]), .pll_fse(pll_fse), .pll_ref(pll_ref),
     .vddio_bottombank(vddio_bottombank), .uio_bbank(uio_bbank[23:0]),
     .uio_rbank(uio_rbank[24:0]), .uio_tbank(uio_tbank[23:0]),
     .in_bbank(in_bbank[23:0]), .in_rbank(in_rbank[24:0]),
     .in_tbank(in_tbank[23:0]), .ren_bbank(ren_bbank[23:0]),
     .oen_bbank(oen_bbank[23:0]), .oen_rbank(oen_rbank[24:0]),
     .oen_tbank(oen_tbank[23:0]), .out_bbank(out_bbank[23:0]),
     .out_rbank(out_rbank[24:0]), .out_tbank(out_tbank[23:0]),
     .ren_rbank(ren_rbank[25:0]), .ien_rbank(ien_rbank[24:0]),
     .ien_tbank(ien_tbank[23:0]), .ren_tbank(ren_tbank[23:0]),
     .ien_bbank(ien_bbank[23:0]), .vppin(vppin), .trstb(trstb),
     .creset_b(creset_b), .cdone_out(cdone_out),
     .creset_b_int(creset_b_int), .vpp(vpp), .cdone(cdone),
     .cdone_int(cdone_in), .trstb_int_pad(trstb_pad),
     .vddio_spi(vddio_spi));

endmodule
// Library - ice1chip, Cell - chip_ice1f, View - schematic
// LAST TIME SAVED: Jun  8 12:05:31 2011
// NETLIST TIME: Jun 29 10:32:28 2011
`timescale 1ns / 1ns 

module chip_ice1f ( cdone, uio_bbank, uio_lbank, uio_rbank, uio_tbank,
     vpp, creset_b, trstb, vdda );

inout  cdone, vpp;

input  creset_b, trstb, vdda;

inout [23:0]  uio_lbank;
inout [24:0]  uio_rbank;
inout [23:0]  uio_tbank;
inout [23:0]  uio_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [287:0]  wl_r;

wire  [3:0]  bm_sdo_o;

wire  [24:0]  out_rbank;

wire  [23:0]  oen_tbank;

wire  [287:0]  vdd_cntl_l;

wire  [287:0]  wl_l;

wire  [287:0]  pgate_r;

wire  [287:0]  reset_r;

wire  [287:0]  pgate_l;

wire  [287:0]  reset_l;

wire  [24:0]  oen_rbank;

wire  [23:0]  in_tbank;

wire  [24:0]  in_rbank;

wire  [23:0]  out_bbank;

wire  [4:0]  spi_ss_in_bbank;

wire  [23:0]  oen_bbank;

wire  [23:0]  out_lbank;

wire  [23:0]  out_tbank;

wire  [23:0]  oen_lbank;

wire  [1:0]  gclk_l2clktv_b;

wire  [23:0]  in_bbank;

wire  [383:0]  cf_rbank;

wire  [3:0]  bm_sdi_o;

wire  [7:0]  fo_dlyadj;

wire  [1:0]  gclk_r2clktv_b;

wire  [16:0]  pll_cbit;

wire  [287:0]  cf_tbank;

wire  [663:0]  bl_bot;

wire  [287:0]  cf_bbank;

wire  [23:0]  in_lbank;

wire  [3:0]  bm_banksel_i;

wire  [0:3]  last_rsr;

wire  [7:0]  bm_sa_i;

wire  [663:0]  bl_top;

wire  [383:0]  cf_lbank;

wire  [10:11]  in_bbank_pll;

wire  [287:0]  vdd_cntl_r;



pll_bufwrap_ice1f I_pll_sdo_buf ( .f_in(pll_sdo), .f_out(pll_sdod));
pll_wrapbuf_ice1f pll_wrap ( gclk_l2clktv_b[1:0], gclk_r2clktv_b[1:0],
     in_bbank_pll[10], in_bbank_pll[11], pll_bypass, pll_cbit[16:0],
     pll_fb, pll_fse, pll_lock_out, pll_ref, pll_reset, pll_sdo,
     cf_bbank[159], cf_bbank[135], cf_lbank[9:1], cf_lbank[33:25],
     cf_lbank[57:49], cf_lbank[81:73], cf_lbank[97], cf_lbank[99],
     cf_lbank[101], fabric_out_06_00, fabric_out_07_00, fo_bypass,
     fo_dlyadj[7:0], fo_fb, fo_ref, fo_reset, fo_sck, fp_sdi, icegate,
     in_bbank[10], in_bbank[11], pll_lock, pllout, gint_hz);
quad_x4_ice1 iquad_x4 ( bm_sdo_o[3:0], cf_bbank[287:0],
     cf_lbank[383:0], cf_rbank[383:0], cf_tbank[287:0], icegate,
     fabric_out_06_00, fabric_out_07_00, fabric_out_12_00_wb,
     fabric_out_13_01, fabric_out_13_02, fo_bypass, fo_dlyadj[7:0],
     fo_fb, fo_ref, fo_reset, fo_sck, fp_sdi, oen_bbank[23:0],
     oen_lbank[23:0], oen_rbank[24:0], oen_tbank[23:0],
     out_bbank[23:0], out_lbank[23:0], out_rbank[24:0],
     out_tbank[23:0], fromsdo, spi_ss_in_bbank[4:0], tck_pad, tdi_pad,
     tms_pad, bl_bot[663:0], bl_top[663:0], bm_banksel_i[3:0],
     bm_init_i, bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i,
     bm_sdi_o[3:0], bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0,
     ceb, end_of_startup, gclk_l2clktv_b[1:0], gclk_r2clktv_b[1:0],
     hiz_b0, jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[0],
     last_rsr[1], last_rsr[2], last_rsr[3], md_spi_b, mode0,
     mux_jtag_sel_b, {in_bbank[23:12], in_bbank_pll[11],
     in_bbank_pll[10], in_bbank[9:0]}, in_lbank[23:0], in_rbank[24:0],
     in_tbank[23:0], pgate_l[287:0], pgate_r[287:0], pll_lock_out,
     pll_sdod, gint_hz, gsr, gsr, reset_l[287:0], reset_r[287:0],
     j_tdi, sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, j_tck, totdopad, trstb_pad, update0,
     vdd_cntl_l[287:0], vdd_cntl_r[287:0], wl_l[287:0], wl_r[287:0]);
ring_route_ice1f I_ring_route1f ( bm_banksel_i[3:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i,
     bm_sdi_o[3:0], bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0,
     ceb, end_of_startup, gint_hz, gsr, hiz_b0, in_bbank[23:0],
     in_lbank[23:0], in_rbank[24:0], in_tbank[23:0], j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[1],
     last_rsr[0], last_rsr[3], last_rsr[2], md_spi_b, mode0,
     mux_jtag_sel_b, pgate_l[287:0], pgate_r[287:0], pll_lock, pllout,
     reset_l[287:0], reset_r[287:0], sdo_enable, shift0, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out, totdopad, trstb_pad, update0,
     vdd_cntl_l[287:0], vdd_cntl_r[287:0], wl_l[287:0], wl_r[287:0],
     bl_bot[663:0], bl_top[663:0], cdone, uio_bbank[23:0],
     uio_lbank[23:0], uio_rbank[24:0], uio_tbank[23:0], vpp,
     bm_sdo_o[3:0], creset_b, fabric_out_12_00_wb, fabric_out_13_01,
     fabric_out_13_02, fromsdo, {cf_lbank[324], cf_lbank[323],
     cf_lbank[300], cf_lbank[299], cf_lbank[276], cf_lbank[275],
     cf_lbank[252], cf_lbank[251], cf_lbank[228], cf_lbank[227],
     cf_lbank[204], cf_lbank[203], cf_lbank[180], cf_lbank[179],
     cf_lbank[132], cf_lbank[131], cf_lbank[108], cf_lbank[107],
     cf_lbank[84], cf_lbank[83], cf_lbank[60], cf_lbank[59],
     cf_lbank[36], cf_lbank[35]}, {cf_bbank[275], cf_bbank[276],
     cf_bbank[251], cf_bbank[252], cf_bbank[227], cf_bbank[228],
     cf_bbank[203], cf_bbank[204], cf_bbank[179], cf_bbank[180],
     cf_bbank[155], cf_bbank[156], cf_bbank[131], cf_bbank[132],
     cf_bbank[107], cf_bbank[108], cf_bbank[83], cf_bbank[84],
     cf_bbank[59], cf_bbank[60], cf_bbank[35], cf_bbank[36],
     cf_bbank[11], cf_bbank[12]}, {cf_rbank[347], cf_rbank[348],
     cf_rbank[323], cf_rbank[324], cf_rbank[299], cf_rbank[300],
     cf_rbank[251], cf_rbank[252], cf_rbank[227], cf_rbank[228],
     cf_rbank[203], cf_rbank[204], cf_rbank[179], cf_rbank[180],
     cf_rbank[155], cf_rbank[156], cf_rbank[131], cf_rbank[132],
     cf_rbank[83], cf_rbank[84], cf_rbank[59], cf_rbank[35],
     cf_rbank[36], cf_rbank[11], cf_rbank[12]}, {cf_tbank[275],
     cf_tbank[276], cf_tbank[251], cf_tbank[252], cf_tbank[227],
     cf_tbank[228], cf_tbank[203], cf_tbank[204], cf_tbank[179],
     cf_tbank[180], cf_tbank[155], cf_tbank[156], cf_tbank[131],
     cf_tbank[132], cf_tbank[107], cf_tbank[108], cf_tbank[83],
     cf_tbank[84], cf_tbank[59], cf_tbank[60], cf_tbank[35],
     cf_tbank[36], cf_tbank[11], cf_tbank[12]}, {cf_lbank[325],
     cf_lbank[301], cf_lbank[277], cf_lbank[253], cf_lbank[229],
     cf_lbank[205], cf_lbank[181], cf_lbank[133], cf_lbank[109],
     cf_lbank[85], cf_lbank[61], cf_lbank[37]}, oen_bbank[23:0],
     oen_lbank[23:0], oen_rbank[24:0], oen_tbank[23:0],
     out_bbank[23:0], out_lbank[23:0], out_rbank[24:0],
     out_tbank[23:0], pll_bypass, pll_cbit[16:0], pll_fb, pll_fse,
     pll_ref, pll_reset, {cf_lbank[322], cf_lbank[312], cf_lbank[298],
     cf_lbank[288], cf_lbank[274], cf_lbank[264], cf_lbank[250],
     cf_lbank[240], cf_lbank[226], cf_lbank[216], cf_lbank[202],
     cf_lbank[192], cf_lbank[178], cf_lbank[168], cf_lbank[130],
     cf_lbank[120], cf_lbank[106], cf_lbank[96], cf_lbank[82],
     cf_lbank[72], cf_lbank[58], cf_lbank[48], cf_lbank[34],
     cf_lbank[24]}, {cf_bbank[264], cf_bbank[274], cf_bbank[240],
     cf_bbank[250], cf_bbank[216], cf_bbank[226], cf_bbank[192],
     cf_bbank[202], cf_bbank[168], cf_bbank[178], cf_bbank[144],
     cf_bbank[154], cf_bbank[120], cf_bbank[130], cf_bbank[96],
     cf_bbank[106], cf_bbank[72], cf_bbank[82], cf_bbank[48],
     cf_bbank[58], cf_bbank[24], cf_bbank[34], cf_bbank[0],
     cf_bbank[10]}, {cf_rbank[38], cf_rbank[336], cf_rbank[346],
     cf_rbank[312], cf_rbank[322], cf_rbank[288], cf_rbank[298],
     cf_rbank[240], cf_rbank[250], cf_rbank[216], cf_rbank[226],
     cf_rbank[192], cf_rbank[202], cf_rbank[168], cf_rbank[178],
     cf_rbank[144], cf_rbank[154], cf_rbank[120], cf_rbank[130],
     cf_rbank[72], cf_rbank[82], cf_rbank[48], cf_rbank[24],
     cf_rbank[34], cf_rbank[0], cf_rbank[10]}, {cf_tbank[264],
     cf_tbank[274], cf_tbank[240], cf_tbank[250], cf_tbank[216],
     cf_tbank[226], cf_tbank[192], cf_tbank[202], cf_tbank[168],
     cf_tbank[178], cf_tbank[144], cf_tbank[154], cf_tbank[120],
     cf_tbank[130], cf_tbank[96], cf_tbank[106], cf_tbank[72],
     cf_tbank[82], cf_tbank[48], cf_tbank[58], cf_tbank[24],
     cf_tbank[34], cf_tbank[0], cf_tbank[10]}, spi_ss_in_bbank[4:0],
     tck_pad, tdi_pad, tms_pad, trstb, vdda);

endmodule
// Library - leafcell, Cell - misc_module4_ice1p, View - schematic
// LAST TIME SAVED: Jun  2 10:50:29 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module misc_module4_ice1p ( S_R, .cbit_colcntl({cbit[60], cbit[56],
     cbit[52], cbit[48], cbit[44], cbit[40], cbit[32], cbit[3]}), clk,
     clkb, glb2local, sp4, bl, b, glb_netwk, l, lc_trk_g0, lc_trk_g1,
     lc_trk_g2, lc_trk_g3, m, min0, min1, min2, min3, pgate, prog, r,
     reset_b, sp12, vdd_cntl, wl );
output  S_R, clk, clkb;


input  prog;

output [63:0]  cbit;
output [7:0]  sp4;
output [3:0]  glb2local;

inout [3:0]  bl;

input [5:0]  lc_trk_g2;
input [15:0]  reset_b;
input [1:0]  l;
input [7:0]  min1;
input [5:0]  lc_trk_g1;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [5:0]  lc_trk_g0;
input [7:0]  min3;
input [7:0]  min0;
input [7:0]  glb_netwk;
input [7:0]  sp12;
input [15:0]  wl;
input [1:0]  m;
input [7:0]  min2;
input [1:0]  b;
input [5:0]  lc_trk_g3;
input [1:0]  r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [63:0]  cbitb;

wire  [15:0]  r_vdd;



inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
pch_hvt  M0_15_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[15]), .S(r_vdd[15]));
pch_hvt  M0_14_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[14]), .S(r_vdd[14]));
pch_hvt  M0_13_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[13]), .S(r_vdd[13]));
pch_hvt  M0_12_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[12]), .S(r_vdd[12]));
pch_hvt  M0_11_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[11]), .S(r_vdd[11]));
pch_hvt  M0_10_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[10]), .S(r_vdd[10]));
pch_hvt  M0_9_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[9]), .S(r_vdd[9]));
pch_hvt  M0_8_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[8]), .S(r_vdd[8]));
pch_hvt  M0_7_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[7]), .S(r_vdd[7]));
pch_hvt  M0_6_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[6]), .S(r_vdd[6]));
pch_hvt  M0_5_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[5]), .S(r_vdd[5]));
pch_hvt  M0_4_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[4]), .S(r_vdd[4]));
pch_hvt  M0_3_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[3]), .S(r_vdd[3]));
pch_hvt  M0_2_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[2]), .S(r_vdd[2]));
pch_hvt  M0_1_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[1]), .S(r_vdd[1]));
pch_hvt  M0_0_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[0]), .S(r_vdd[0]));
clkmandcmuxrev0 I_clkmandcmuxrev0 ( .prog(progd),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]), .clk(clk),
     .clkb(clkb), .glb_netwk(glb_netwk[7:0]), .s_r(S_R),
     .glb2local(glb2local[3:0]), .cbit({cbit[2], cbit[1], cbit[0],
     cbit[27], cbit[25], cbit[26], cbit[24], cbit[23], cbit[21],
     cbit[22], cbit[20], cbit[19], cbit[17], cbit[18], cbit[16],
     cbit[15], cbit[13], cbit[14], cbit[12], cbit[31], cbit[29],
     cbit[30], cbit[28], cbit[11], cbit[9], cbit[10], cbit[8],
     cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}), .min2(min2[7:0]),
     .min1(min1[7:0]), .min0(min0[7:0]), .min3(min3[7:0]),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}));
sp12to4 I_sp12to4_7_ ( .prog(progd), .triout(sp4[7]),
     .cbitb(cbitb[62]), .drv(sp12[7]));
sp12to4 I_sp12to4_6_ ( .prog(progd), .triout(sp4[6]),
     .cbitb(cbitb[58]), .drv(sp12[6]));
sp12to4 I_sp12to4_5_ ( .prog(progd), .triout(sp4[5]),
     .cbitb(cbitb[54]), .drv(sp12[5]));
sp12to4 I_sp12to4_4_ ( .prog(progd), .triout(sp4[4]),
     .cbitb(cbitb[50]), .drv(sp12[4]));
sp12to4 I_sp12to4_3_ ( .prog(progd), .triout(sp4[3]),
     .cbitb(cbitb[46]), .drv(sp12[3]));
sp12to4 I_sp12to4_2_ ( .prog(progd), .triout(sp4[2]),
     .cbitb(cbitb[42]), .drv(sp12[2]));
sp12to4 I_sp12to4_1_ ( .prog(progd), .triout(sp4[1]), .cbitb(cbitb[5]),
     .drv(sp12[1]));
sp12to4 I_sp12to4_0_ ( .prog(progd), .triout(sp4[0]),
     .cbitb(cbitb[34]), .drv(sp12[0]));
sbox1 I_sbox1_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(progd));
sbox1 I_sbox1_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(progd));
cram16x4 I_cram16x4 ( .q(cbit[63:0]), .r_gnd(r_vdd[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));

endmodule
// Library - xpmem, Cell - cram2x2x5, View - schematic
// LAST TIME SAVED: May 11 15:38:01 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module cram2x2x5 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [19:0]  q_b;
output [19:0]  q;

inout [9:0]  bl;

input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  r_gnd;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - sbox11to9_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:53:05 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox11to9_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  b;
inout [9:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_l10 ( .prog(prog), .in6(t[4]), .in5(t[10]), .in4(r[2]),
     .in3(r[10]), .in2(r[7]), .in1(b[10]), .in0(b[5]), .out(l[10]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t10 ( .prog(prog), .in6(r[4]), .in5(r[10]), .in4(b[2]),
     .in3(b[10]), .in2(b[7]), .in1(l[10]), .in0(l[5]), .out(t[10]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t11 ( .prog(prog), .in6(r[5]), .in5(r[11]), .in4(b[3]),
     .in3(b[11]), .in2(b[8]), .in1(l[11]), .in0(l[6]), .out(t[11]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t9 ( .prog(prog), .in6(r[3]), .in5(r[9]), .in4(b[1]),
     .in3(b[9]), .in2(b[6]), .in1(l[9]), .in0(l[4]), .out(t[9]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l11 ( .prog(prog), .in6(t[5]), .in5(t[11]), .in4(r[3]),
     .in3(r[11]), .in2(r[8]), .in1(b[11]), .in0(b[6]), .out(l[11]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l9 ( .prog(prog), .in6(t[3]), .in5(t[9]), .in4(r[1]),
     .in3(r[9]), .in2(r[6]), .in1(b[9]), .in0(b[4]), .out(l[9]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox11to9_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:52:20 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox11to9_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  b;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r10 ( .prog(prog), .in6(b[4]), .in5(b[10]), .in4(l[2]),
     .in3(l[10]), .in2(l[7]), .in1(t[10]), .in0(t[5]), .out(r[10]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b10 ( .prog(prog), .in6(l[4]), .in5(l[10]), .in4(t[2]),
     .in3(t[10]), .in2(t[7]), .in1(r[10]), .in0(r[5]), .out(b[10]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b11 ( .prog(prog), .in6(l[5]), .in5(l[11]), .in4(t[3]),
     .in3(t[11]), .in2(t[8]), .in1(r[11]), .in0(r[6]), .out(b[11]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b9 ( .prog(prog), .in6(l[3]), .in5(l[9]), .in4(t[1]),
     .in3(t[9]), .in2(t[6]), .in1(r[9]), .in0(r[4]), .out(b[9]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r11 ( .prog(prog), .in6(b[5]), .in5(b[11]), .in4(l[3]),
     .in3(l[11]), .in2(l[8]), .in1(t[11]), .in0(t[6]), .out(r[11]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r9 ( .prog(prog), .in6(b[3]), .in5(b[9]), .in4(l[1]),
     .in3(l[9]), .in2(l[6]), .in1(t[9]), .in0(t[4]), .out(r[9]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox8to6_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:51:38 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox8to6_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  t;
inout [9:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  reset_b;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I554 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_l7 ( .prog(prog), .in6(t[1]), .in5(t[7]), .in4(r[11]),
     .in3(r[7]), .in2(r[4]), .in1(b[7]), .in0(b[2]), .out(l[7]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t7 ( .prog(prog), .in6(r[1]), .in5(r[7]), .in4(b[11]),
     .in3(b[7]), .in2(b[4]), .in1(l[7]), .in0(l[2]), .out(t[7]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t8 ( .prog(prog), .in6(r[2]), .in5(r[8]), .in4(b[0]),
     .in3(b[8]), .in2(b[5]), .in1(l[8]), .in0(l[3]), .out(t[8]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t6 ( .prog(prog), .in6(r[0]), .in5(r[6]), .in4(b[10]),
     .in3(b[6]), .in2(b[3]), .in1(l[6]), .in0(l[1]), .out(t[6]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l8 ( .prog(prog), .in6(t[2]), .in5(t[8]), .in4(r[0]),
     .in3(r[8]), .in2(r[5]), .in1(b[8]), .in0(b[3]), .out(l[8]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l6 ( .prog(prog), .in6(t[0]), .in5(t[6]), .in4(r[10]),
     .in3(r[6]), .in2(r[3]), .in1(b[6]), .in0(b[1]), .out(l[6]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - pll_ml_dff, View - schematic
// LAST TIME SAVED: Jun  9 15:25:37 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pll_ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - leafcell, Cell - sbox8to6_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:50:50 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox8to6_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r7 ( .prog(prog), .in6(b[1]), .in5(b[7]), .in4(l[11]),
     .in3(l[7]), .in2(l[4]), .in1(t[7]), .in0(t[2]), .out(r[7]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b7 ( .prog(prog), .in6(l[1]), .in5(l[7]), .in4(t[11]),
     .in3(t[7]), .in2(t[4]), .in1(r[7]), .in0(r[2]), .out(b[7]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b8 ( .prog(prog), .in6(l[2]), .in5(l[8]), .in4(t[0]),
     .in3(t[8]), .in2(t[5]), .in1(r[8]), .in0(r[3]), .out(b[8]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b6 ( .prog(prog), .in6(l[0]), .in5(l[6]), .in4(t[10]),
     .in3(t[6]), .in2(t[3]), .in1(r[6]), .in0(r[1]), .out(b[6]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r8 ( .prog(prog), .in6(b[2]), .in5(b[8]), .in4(l[0]),
     .in3(l[8]), .in2(l[5]), .in1(t[8]), .in0(t[3]), .out(r[8]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r6 ( .prog(prog), .in6(b[0]), .in5(b[6]), .in4(l[10]),
     .in3(l[6]), .in2(l[3]), .in1(t[6]), .in0(t[1]), .out(r[6]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox5to3_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:39:32 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox5to3_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  l;
inout [11:0]  t;
inout [11:0]  b;
inout [11:0]  r;
inout [9:0]  bl;

input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_l4 ( .prog(prog), .in6(t[10]), .in5(t[4]), .in4(r[8]),
     .in3(r[4]), .in2(r[1]), .in1(b[4]), .in0(b[11]), .out(l[4]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t4 ( .prog(prog), .in6(r[10]), .in5(r[4]), .in4(b[8]),
     .in3(b[4]), .in2(b[1]), .in1(l[4]), .in0(l[11]), .out(t[4]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t5 ( .prog(prog), .in6(r[11]), .in5(r[5]), .in4(b[9]),
     .in3(b[5]), .in2(b[2]), .in1(l[5]), .in0(l[0]), .out(t[5]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t3 ( .prog(prog), .in6(r[9]), .in5(r[3]), .in4(b[7]),
     .in3(b[3]), .in2(b[0]), .in1(l[3]), .in0(l[10]), .out(t[3]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l5 ( .prog(prog), .in6(t[11]), .in5(t[5]), .in4(r[9]),
     .in3(r[5]), .in2(r[2]), .in1(b[5]), .in0(b[0]), .out(l[5]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l3 ( .prog(prog), .in6(t[9]), .in5(t[3]), .in4(r[7]),
     .in3(r[3]), .in2(r[0]), .in1(b[3]), .in0(b[10]), .out(l[3]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox5to3_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:38:42 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox5to3_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  b;

input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r4 ( .prog(prog), .in6(b[10]), .in5(b[4]), .in4(l[8]),
     .in3(l[4]), .in2(l[1]), .in1(t[4]), .in0(t[11]), .out(r[4]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b4 ( .prog(prog), .in6(l[10]), .in5(l[4]), .in4(t[8]),
     .in3(t[4]), .in2(t[1]), .in1(r[4]), .in0(r[11]), .out(b[4]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b5 ( .prog(prog), .in6(l[11]), .in5(l[5]), .in4(t[9]),
     .in3(t[5]), .in2(t[2]), .in1(r[5]), .in0(r[0]), .out(b[5]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b3 ( .prog(prog), .in6(l[9]), .in5(l[3]), .in4(t[7]),
     .in3(t[3]), .in2(t[0]), .in1(r[3]), .in0(r[10]), .out(b[3]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r5 ( .prog(prog), .in6(b[11]), .in5(b[5]), .in4(l[9]),
     .in3(l[5]), .in2(l[2]), .in1(t[5]), .in0(t[0]), .out(r[5]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r3 ( .prog(prog), .in6(b[9]), .in5(b[3]), .in4(l[7]),
     .in3(l[3]), .in2(l[0]), .in1(t[3]), .in0(t[10]), .out(r[3]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox2to0_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:37:50 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox2to0_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbitb;
output [19:0]  cbit;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  b;
inout [11:0]  l;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_l1 ( .prog(prog), .in6(t[7]), .in5(t[1]), .in4(r[5]),
     .in3(r[1]), .in2(r[10]), .in1(b[1]), .in0(b[8]), .out(l[1]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_l0 ( .prog(prog), .in6(t[6]), .in5(t[0]), .in4(r[4]),
     .in3(r[0]), .in2(r[9]), .in1(b[0]), .in0(b[7]), .out(l[0]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));
sbox7to1_220 I_t1 ( .prog(prog), .in6(r[7]), .in5(r[1]), .in4(b[5]),
     .in3(b[1]), .in2(b[10]), .in1(l[1]), .in0(l[8]), .out(t[1]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_l2 ( .prog(prog), .in6(t[8]), .in5(t[2]), .in4(r[6]),
     .in3(r[2]), .in2(r[11]), .in1(b[2]), .in0(b[9]), .out(l[2]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_t2 ( .prog(prog), .in6(r[8]), .in5(r[2]), .in4(b[6]),
     .in3(b[2]), .in2(b[11]), .in1(l[2]), .in0(l[9]), .out(t[2]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t0 ( .prog(prog), .in6(r[6]), .in5(r[0]), .in4(b[4]),
     .in3(b[0]), .in2(b[9]), .in1(l[0]), .in0(l[7]), .out(t[0]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));

endmodule
// Library - leafcell, Cell - sbox2to0_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:53:10 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox2to0_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  b;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r1 ( .prog(prog), .in6(b[7]), .in5(b[1]), .in4(l[5]),
     .in3(l[1]), .in2(l[10]), .in1(t[1]), .in0(t[8]), .out(r[1]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_r0 ( .prog(prog), .in6(b[6]), .in5(b[0]), .in4(l[4]),
     .in3(l[0]), .in2(l[9]), .in1(t[0]), .in0(t[7]), .out(r[0]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));
sbox7to1_220 I_b1 ( .prog(prog), .in6(l[7]), .in5(l[1]), .in4(t[5]),
     .in3(t[1]), .in2(t[10]), .in1(r[1]), .in0(r[8]), .out(b[1]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_r2 ( .prog(prog), .in6(b[8]), .in5(b[2]), .in4(l[6]),
     .in3(l[2]), .in2(l[11]), .in1(t[2]), .in0(t[9]), .out(r[2]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_b2 ( .prog(prog), .in6(l[8]), .in5(l[2]), .in4(t[6]),
     .in3(t[2]), .in2(t[11]), .in1(r[2]), .in0(r[9]), .out(b[2]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b0 ( .prog(prog), .in6(l[6]), .in5(l[0]), .in4(t[4]),
     .in3(t[0]), .in2(t[9]), .in1(r[0]), .in0(r[7]), .out(b[0]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));

endmodule
// Library - leafcell, Cell - span4_switchandmem_v3, View - schematic
// LAST TIME SAVED: Oct 19 10:24:53 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module span4_switchandmem_v3 ( c, cc, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [7:0]  c;
output [15:8]  cc;

inout [11:0]  r;
inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  b;

input [15:0]  reset_b;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  n2;

wire  [0:19]  net0236;

wire  [19:0]  n1;

wire  [0:19]  net0248;

wire  [0:19]  net0245;

wire  [19:0]  n3;

wire  [0:19]  net0177;

wire  [0:19]  net0241;

wire  [19:0]  n6;

wire  [19:0]  n5;

wire  [19:0]  n0;

wire  [19:0]  n4;

wire  [0:19]  net0201;

wire  [19:0]  n7;

wire  [0:19]  net0189;

wire  [0:19]  net0250;



sbox11to9_p2_v2 I_sbox11to9_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb(net0241[0:19]), .cbit({n7[19:8], cc[15], n7[6], cc[14],
     n7[4:0]}), .wl(wl[15:14]), .vdd_cntl(vdd_cntl[15:14]),
     .reset_b(reset_b[15:14]), .pgate(pgate[15:14]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox11to9_p1_v2 I_sbox11to9_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb(net0236[0:19]), .cbit({n6[19:8], cc[13], n6[6], cc[12],
     n6[4:0]}), .wl(wl[13:12]), .vdd_cntl(vdd_cntl[13:12]),
     .reset_b(reset_b[13:12]), .pgate(pgate[13:12]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox8to6_p2_v2 I_sbox8to6_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb(net0248[0:19]), .cbit({n5[19:8], cc[11], n5[6], cc[10],
     n5[4:0]}), .wl(wl[11:10]), .vdd_cntl(vdd_cntl[11:10]),
     .reset_b(reset_b[11:10]), .pgate(pgate[11:10]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox8to6_p1_v2 I_sbox8to6_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb(net0177[0:19]), .cbit({n4[19:8], cc[9], n4[6], cc[8],
     n4[4:0]}), .wl(wl[9:8]), .vdd_cntl(vdd_cntl[9:8]),
     .reset_b(reset_b[9:8]), .pgate(pgate[9:8]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox5to3_p2_v2 I_sbox5to3_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb(net0189[0:19]), .cbit({n3[19:8], c[7], n3[6], c[6],
     n3[4:0]}), .wl(wl[7:6]), .vdd_cntl(vdd_cntl[7:6]),
     .reset_b(reset_b[7:6]), .pgate(pgate[7:6]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox5to3_p1_v2 I_sbox5to3_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb(net0201[0:19]), .cbit({n2[19:8], c[5], n2[6], c[4],
     n2[4:0]}), .wl(wl[5:4]), .vdd_cntl(vdd_cntl[5:4]),
     .reset_b(reset_b[5:4]), .pgate(pgate[5:4]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox2to0_p2_v2 I_sbox2to0_p2_v2 ( .b(b[11:0]), .cbitb(net0245[0:19]),
     .cbit({n1[19:8], c[3], n1[6], c[2], n1[4:0]}), .wl(wl[3:2]),
     .vdd_cntl(vdd_cntl[3:2]), .reset_b(reset_b[3:2]), .prog(prog),
     .pgate(pgate[3:2]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox2to0_p1_v2 I_sbox2to0_p1_v2 ( .cbitb(net0250[0:19]),
     .cbit({n0[19:8], c[1], n0[6], c[0], n0[4:0]}), .wl(wl[1:0]),
     .vdd_cntl(vdd_cntl[1:0]), .reset_b(reset_b[1:0]), .prog(prog),
     .pgate(pgate[1:0]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]), .b(b[11:0]));

endmodule
// Library - leafcell, Cell - span4_ice8p, View - schematic
// LAST TIME SAVED: Jan 12 15:03:31 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module span4_ice8p ( bram_cbit, ccntrl_cbit, bl, sp4_h_l, sp4_h_r,
     sp4_v_b, sp4_v_t, pgate, prog, reset_b, vdd_cntl, wl );


input  prog;

output [7:0]  bram_cbit;
output [7:0]  ccntrl_cbit;

inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_t;
inout [47:0]  sp4_h_r;
inout [9:0]  bl;

input [15:0]  vdd_cntl;
input [15:0]  reset_b;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  sp4_h_r_mid;

wire  [11:0]  sp4_v_b_mid;



rm7y  R0_47_ ( .MINUS(sp4_v_b[47]), .PLUS(sp4_v_t[34]));
rm7y  R0_46_ ( .MINUS(sp4_v_b[46]), .PLUS(sp4_v_t[35]));
rm7y  R0_45_ ( .MINUS(sp4_v_b[45]), .PLUS(sp4_v_t[32]));
rm7y  R0_44_ ( .MINUS(sp4_v_b[44]), .PLUS(sp4_v_t[33]));
rm7y  R0_43_ ( .MINUS(sp4_v_b[43]), .PLUS(sp4_v_t[30]));
rm7y  R0_42_ ( .MINUS(sp4_v_b[42]), .PLUS(sp4_v_t[31]));
rm7y  R0_41_ ( .MINUS(sp4_v_b[41]), .PLUS(sp4_v_t[28]));
rm7y  R0_40_ ( .MINUS(sp4_v_b[40]), .PLUS(sp4_v_t[29]));
rm7y  R0_39_ ( .MINUS(sp4_v_b[39]), .PLUS(sp4_v_t[26]));
rm7y  R0_38_ ( .MINUS(sp4_v_b[38]), .PLUS(sp4_v_t[27]));
rm7y  R0_37_ ( .MINUS(sp4_v_b[37]), .PLUS(sp4_v_t[24]));
rm7y  R0_36_ ( .MINUS(sp4_v_b[36]), .PLUS(sp4_v_t[25]));
rm7y  R0_35_ ( .MINUS(sp4_v_b[35]), .PLUS(sp4_v_t[22]));
rm7y  R0_34_ ( .MINUS(sp4_v_b[34]), .PLUS(sp4_v_t[23]));
rm7y  R0_33_ ( .MINUS(sp4_v_b[33]), .PLUS(sp4_v_t[20]));
rm7y  R0_32_ ( .MINUS(sp4_v_b[32]), .PLUS(sp4_v_t[21]));
rm7y  R0_31_ ( .MINUS(sp4_v_b[31]), .PLUS(sp4_v_t[18]));
rm7y  R0_30_ ( .MINUS(sp4_v_b[30]), .PLUS(sp4_v_t[19]));
rm7y  R0_29_ ( .MINUS(sp4_v_b[29]), .PLUS(sp4_v_t[16]));
rm7y  R0_28_ ( .MINUS(sp4_v_b[28]), .PLUS(sp4_v_t[17]));
rm7y  R0_27_ ( .MINUS(sp4_v_b[27]), .PLUS(sp4_v_t[14]));
rm7y  R0_26_ ( .MINUS(sp4_v_b[26]), .PLUS(sp4_v_t[15]));
rm7y  R0_25_ ( .MINUS(sp4_v_b[25]), .PLUS(sp4_v_t[12]));
rm7y  R0_24_ ( .MINUS(sp4_v_b[24]), .PLUS(sp4_v_t[13]));
rm7y  R0_23_ ( .MINUS(sp4_v_b[23]), .PLUS(sp4_v_t[10]));
rm7y  R0_22_ ( .MINUS(sp4_v_b[22]), .PLUS(sp4_v_t[11]));
rm7y  R0_21_ ( .MINUS(sp4_v_b[21]), .PLUS(sp4_v_t[8]));
rm7y  R0_20_ ( .MINUS(sp4_v_b[20]), .PLUS(sp4_v_t[9]));
rm7y  R0_19_ ( .MINUS(sp4_v_b[19]), .PLUS(sp4_v_t[6]));
rm7y  R0_18_ ( .MINUS(sp4_v_b[18]), .PLUS(sp4_v_t[7]));
rm7y  R0_17_ ( .MINUS(sp4_v_b[17]), .PLUS(sp4_v_t[4]));
rm7y  R0_16_ ( .MINUS(sp4_v_b[16]), .PLUS(sp4_v_t[5]));
rm7y  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[2]));
rm7y  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[3]));
rm7y  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[0]));
rm7y  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[1]));
rm7y  R0_11_ ( .MINUS(sp4_v_b_mid[11]), .PLUS(sp4_v_t[46]));
rm7y  R0_10_ ( .MINUS(sp4_v_b_mid[10]), .PLUS(sp4_v_t[47]));
rm7y  R0_9_ ( .MINUS(sp4_v_b_mid[9]), .PLUS(sp4_v_t[44]));
rm7y  R0_8_ ( .MINUS(sp4_v_b_mid[8]), .PLUS(sp4_v_t[45]));
rm7y  R0_7_ ( .MINUS(sp4_v_b_mid[7]), .PLUS(sp4_v_t[42]));
rm7y  R0_6_ ( .MINUS(sp4_v_b_mid[6]), .PLUS(sp4_v_t[43]));
rm7y  R0_5_ ( .MINUS(sp4_v_b_mid[5]), .PLUS(sp4_v_t[40]));
rm7y  R0_4_ ( .MINUS(sp4_v_b_mid[4]), .PLUS(sp4_v_t[41]));
rm7y  R0_3_ ( .MINUS(sp4_v_b_mid[3]), .PLUS(sp4_v_t[38]));
rm7y  R0_2_ ( .MINUS(sp4_v_b_mid[2]), .PLUS(sp4_v_t[39]));
rm7y  R0_1_ ( .MINUS(sp4_v_b_mid[1]), .PLUS(sp4_v_t[36]));
rm7y  R0_0_ ( .MINUS(sp4_v_b_mid[0]), .PLUS(sp4_v_t[37]));
span4_switchandmem_v3 I_span4_switchandmem_rev ( .cc(ccntrl_cbit[7:0]),
     .c(bram_cbit[7:0]), .wl(wl[15:0]), .vdd_cntl(vdd_cntl[15:0]),
     .reset_b(reset_b[15:0]), .prog(prog), .pgate(pgate[15:0]),
     .t(sp4_v_b_mid[11:0]), .r(sp4_h_r[11:0]), .l(sp4_h_r_mid[11:0]),
     .bl(bl[9:0]), .b(sp4_v_b[11:0]));
rm6w  R1_27_ ( .MINUS(sp4_h_r[47]), .PLUS(sp4_h_l[34]));
rm6w  R1_26_ ( .MINUS(sp4_h_r[46]), .PLUS(sp4_h_l[35]));
rm6w  R1_25_ ( .MINUS(sp4_h_r[45]), .PLUS(sp4_h_l[32]));
rm6w  R1_24_ ( .MINUS(sp4_h_r[44]), .PLUS(sp4_h_l[33]));
rm6w  R1_23_ ( .MINUS(sp4_h_r[43]), .PLUS(sp4_h_l[30]));
rm6w  R1_22_ ( .MINUS(sp4_h_r[42]), .PLUS(sp4_h_l[31]));
rm6w  R1_21_ ( .MINUS(sp4_h_r[41]), .PLUS(sp4_h_l[28]));
rm6w  R1_20_ ( .MINUS(sp4_h_r[40]), .PLUS(sp4_h_l[29]));
rm6w  R1_19_ ( .MINUS(sp4_h_r[39]), .PLUS(sp4_h_l[26]));
rm6w  R1_18_ ( .MINUS(sp4_h_r[38]), .PLUS(sp4_h_l[27]));
rm6w  R1_17_ ( .MINUS(sp4_h_r[37]), .PLUS(sp4_h_l[24]));
rm6w  R1_16_ ( .MINUS(sp4_h_r[36]), .PLUS(sp4_h_l[25]));
rm6w  R1_15_ ( .MINUS(sp4_h_r[35]), .PLUS(sp4_h_l[22]));
rm6w  R1_14_ ( .MINUS(sp4_h_r[34]), .PLUS(sp4_h_l[23]));
rm6w  R1_13_ ( .MINUS(sp4_h_r[23]), .PLUS(sp4_h_l[10]));
rm6w  R1_12_ ( .MINUS(sp4_h_r[22]), .PLUS(sp4_h_l[11]));
rm6w  R1_11_ ( .MINUS(sp4_h_r_mid[11]), .PLUS(sp4_h_l[46]));
rm6w  R1_10_ ( .MINUS(sp4_h_r_mid[10]), .PLUS(sp4_h_l[47]));
rm6w  R1_9_ ( .MINUS(sp4_h_r_mid[9]), .PLUS(sp4_h_l[44]));
rm6w  R1_8_ ( .MINUS(sp4_h_r_mid[8]), .PLUS(sp4_h_l[45]));
rm6w  R1_7_ ( .MINUS(sp4_h_r_mid[7]), .PLUS(sp4_h_l[42]));
rm6w  R1_6_ ( .MINUS(sp4_h_r_mid[6]), .PLUS(sp4_h_l[43]));
rm6w  R1_5_ ( .MINUS(sp4_h_r_mid[5]), .PLUS(sp4_h_l[40]));
rm6w  R1_4_ ( .MINUS(sp4_h_r_mid[4]), .PLUS(sp4_h_l[41]));
rm6w  R1_3_ ( .MINUS(sp4_h_r_mid[3]), .PLUS(sp4_h_l[38]));
rm6w  R1_2_ ( .MINUS(sp4_h_r_mid[2]), .PLUS(sp4_h_l[39]));
rm6w  R1_1_ ( .MINUS(sp4_h_r_mid[1]), .PLUS(sp4_h_l[36]));
rm6w  R1_0_ ( .MINUS(sp4_h_r_mid[0]), .PLUS(sp4_h_l[37]));
rm6w  R2_19_ ( .MINUS(sp4_h_r[33]), .PLUS(sp4_h_l[20]));
rm6w  R2_18_ ( .MINUS(sp4_h_r[32]), .PLUS(sp4_h_l[21]));
rm6w  R2_17_ ( .MINUS(sp4_h_r[31]), .PLUS(sp4_h_l[18]));
rm6w  R2_16_ ( .MINUS(sp4_h_r[30]), .PLUS(sp4_h_l[19]));
rm6w  R2_15_ ( .MINUS(sp4_h_r[29]), .PLUS(sp4_h_l[16]));
rm6w  R2_14_ ( .MINUS(sp4_h_r[28]), .PLUS(sp4_h_l[17]));
rm6w  R2_13_ ( .MINUS(sp4_h_r[27]), .PLUS(sp4_h_l[14]));
rm6w  R2_12_ ( .MINUS(sp4_h_r[26]), .PLUS(sp4_h_l[15]));
rm6w  R2_11_ ( .MINUS(sp4_h_r[25]), .PLUS(sp4_h_l[12]));
rm6w  R2_10_ ( .MINUS(sp4_h_r[24]), .PLUS(sp4_h_l[13]));
rm6w  R2_9_ ( .MINUS(sp4_h_r[21]), .PLUS(sp4_h_l[8]));
rm6w  R2_8_ ( .MINUS(sp4_h_r[20]), .PLUS(sp4_h_l[9]));
rm6w  R2_7_ ( .MINUS(sp4_h_r[19]), .PLUS(sp4_h_l[6]));
rm6w  R2_6_ ( .MINUS(sp4_h_r[18]), .PLUS(sp4_h_l[7]));
rm6w  R2_5_ ( .MINUS(sp4_h_r[17]), .PLUS(sp4_h_l[4]));
rm6w  R2_4_ ( .MINUS(sp4_h_r[16]), .PLUS(sp4_h_l[5]));
rm6w  R2_3_ ( .MINUS(sp4_h_r[15]), .PLUS(sp4_h_l[2]));
rm6w  R2_2_ ( .MINUS(sp4_h_r[14]), .PLUS(sp4_h_l[3]));
rm6w  R2_1_ ( .MINUS(sp4_h_r[13]), .PLUS(sp4_h_l[0]));
rm6w  R2_0_ ( .MINUS(sp4_h_r[12]), .PLUS(sp4_h_l[1]));

endmodule
// Library - xpmem, Cell - cram2x2x6, View - schematic
// LAST TIME SAVED: May 11 14:44:08 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module cram2x2x6 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [23:0]  q;
output [23:0]  q_b;

inout [11:0]  bl;

input [1:0]  r_gnd;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_5_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_base, View - schematic
// LAST TIME SAVED: Nov  5 15:41:50 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_base ( lc_trk_out, sp4_out, bl, min0, min1, min2,
     min3, pgate, prog, reset_b, sp12_in, vdd_cntl, wl );


input  prog;

output [1:0]  sp4_out;
output [3:0]  lc_trk_out;

inout [11:0]  bl;

input [1:0]  vdd_cntl;
input [15:0]  min3;
input [1:0]  sp12_in;
input [15:0]  min1;
input [1:0]  reset_b;
input [15:0]  min2;
input [1:0]  pgate;
input [1:0]  wl;
input [15:0]  min0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [23:0]  cbitb;

wire  [23:0]  cbit;



inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net60));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
g_mux I_mux2 ( .min(min2[15:0]), .prog(net60), .inmuxo(lc_trk_out[2]),
     .cbit({cbit[16], cbit[17], cbit[20], cbit[23], cbit[21]}),
     .cbitb({cbitb[16], cbitb[17], cbitb[20], cbitb[23], cbitb[21]}));
g_mux I_mux3 ( .min(min3[15:0]), .prog(net60), .inmuxo(lc_trk_out[3]),
     .cbit({cbit[18], cbit[19], cbit[22], cbit[15], cbit[13]}),
     .cbitb({cbitb[18], cbitb[19], cbitb[22], cbitb[15], cbitb[13]}));
g_mux I_mux1 ( .min(min1[15:0]), .prog(net60), .inmuxo(lc_trk_out[1]),
     .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}));
g_mux I_mux0 ( .min(min0[15:0]), .prog(net60), .inmuxo(lc_trk_out[0]),
     .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}));
cram2x2x6 I_mem2x2x6 ( .pgate(pgate[1:0]), .q(cbit[23:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[11:0]), .q_b(cbitb[23:0]));
sp12to4 I_sp12to4_1_ ( .triout(sp4_out[1]), .cbitb(cbitb[11]),
     .drv(sp12_in[1]), .prog(net60));
sp12to4 I_sp12to4_0_ ( .triout(sp4_out[0]), .cbitb(cbitb[9]),
     .drv(sp12_in[0]), .prog(net60));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0a, View - schematic
// LAST TIME SAVED: Jul 24 13:27:07 2007
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g0a ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g0;

inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;

input [7:0]  tnl_op;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[34], sp4_r_v_b[25]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[33], sp4_r_v_b[26]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[35], sp4_r_v_b[24]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[32], sp4_r_v_b[27]}),
     .sp4_out(sp4_v_b[13:12]), .sp12_in({sp12_v_b[3], sp12_v_b[1]}),
     .lc_trk_out(lc_trk_g0[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - pllcfg_sr26_40lp, View - schematic
// LAST TIME SAVED: Nov  2 13:15:11 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module pllcfg_sr26_40lp ( q, pll_sck, pll_sdi, reset );

input  pll_sck, pll_sdi, reset;

output [25:0]  q;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:25]  net16;



inv_hvt I472 ( .A(pll_sck), .Y(net11));
pll_ml_dff I4_25_ ( .R(reset), .D(q[24]), .CLK(net11), .QN(net16[0]),
     .Q(q[25]));
pll_ml_dff I4_24_ ( .R(reset), .D(q[23]), .CLK(net11), .QN(net16[1]),
     .Q(q[24]));
pll_ml_dff I4_23_ ( .R(reset), .D(q[22]), .CLK(net11), .QN(net16[2]),
     .Q(q[23]));
pll_ml_dff I4_22_ ( .R(reset), .D(q[21]), .CLK(net11), .QN(net16[3]),
     .Q(q[22]));
pll_ml_dff I4_21_ ( .R(reset), .D(q[20]), .CLK(net11), .QN(net16[4]),
     .Q(q[21]));
pll_ml_dff I4_20_ ( .R(reset), .D(q[19]), .CLK(net11), .QN(net16[5]),
     .Q(q[20]));
pll_ml_dff I4_19_ ( .R(reset), .D(q[18]), .CLK(net11), .QN(net16[6]),
     .Q(q[19]));
pll_ml_dff I4_18_ ( .R(reset), .D(q[17]), .CLK(net11), .QN(net16[7]),
     .Q(q[18]));
pll_ml_dff I4_17_ ( .R(reset), .D(q[16]), .CLK(net11), .QN(net16[8]),
     .Q(q[17]));
pll_ml_dff I4_16_ ( .R(reset), .D(q[15]), .CLK(net11), .QN(net16[9]),
     .Q(q[16]));
pll_ml_dff I4_15_ ( .R(reset), .D(q[14]), .CLK(net11), .QN(net16[10]),
     .Q(q[15]));
pll_ml_dff I4_14_ ( .R(reset), .D(q[13]), .CLK(net11), .QN(net16[11]),
     .Q(q[14]));
pll_ml_dff I4_13_ ( .R(reset), .D(q[12]), .CLK(net11), .QN(net16[12]),
     .Q(q[13]));
pll_ml_dff I4_12_ ( .R(reset), .D(q[11]), .CLK(net11), .QN(net16[13]),
     .Q(q[12]));
pll_ml_dff I4_11_ ( .R(reset), .D(q[10]), .CLK(net11), .QN(net16[14]),
     .Q(q[11]));
pll_ml_dff I4_10_ ( .R(reset), .D(q[9]), .CLK(net11), .QN(net16[15]),
     .Q(q[10]));
pll_ml_dff I4_9_ ( .R(reset), .D(q[8]), .CLK(net11), .QN(net16[16]),
     .Q(q[9]));
pll_ml_dff I4_8_ ( .R(reset), .D(q[7]), .CLK(net11), .QN(net16[17]),
     .Q(q[8]));
pll_ml_dff I4_7_ ( .R(reset), .D(q[6]), .CLK(net11), .QN(net16[18]),
     .Q(q[7]));
pll_ml_dff I4_6_ ( .R(reset), .D(q[5]), .CLK(net11), .QN(net16[19]),
     .Q(q[6]));
pll_ml_dff I4_5_ ( .R(reset), .D(q[4]), .CLK(net11), .QN(net16[20]),
     .Q(q[5]));
pll_ml_dff I4_4_ ( .R(reset), .D(q[3]), .CLK(net11), .QN(net16[21]),
     .Q(q[4]));
pll_ml_dff I4_3_ ( .R(reset), .D(q[2]), .CLK(net11), .QN(net16[22]),
     .Q(q[3]));
pll_ml_dff I4_2_ ( .R(reset), .D(q[1]), .CLK(net11), .QN(net16[23]),
     .Q(q[2]));
pll_ml_dff I4_1_ ( .R(reset), .D(q[0]), .CLK(net11), .QN(net16[24]),
     .Q(q[1]));
pll_ml_dff I4_0_ ( .R(reset), .D(pll_sdi), .CLK(net11), .QN(net16[25]),
     .Q(q[0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0b, View - schematic
// LAST TIME SAVED: Jul 24 13:26:14 2007
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g0b ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, glb2local, lft_op,
     pgate, prog, reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op,
     vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g0;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
input [3:0]  glb2local;
input [7:0]  bnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  top_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], glb2local[1]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], glb2local[2]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], glb2local[0]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], glb2local[3]}),
     .sp4_out(sp4_v_b[15:14]), .sp12_in({sp12_v_b[7], sp12_v_b[5]}),
     .lc_trk_out(lc_trk_g0[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1a, View - schematic
// LAST TIME SAVED: Jul 24 13:25:29 2007
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g1a ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [1:0]  wl;
input [7:0]  bnl_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[25], sp4_r_v_b[1]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[26], sp4_r_v_b[2]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[24], sp4_r_v_b[0]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[27], sp4_r_v_b[3]}),
     .sp4_out(sp4_v_b[17:16]), .sp12_in({sp12_v_b[11], sp12_v_b[9]}),
     .lc_trk_out(lc_trk_g1[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1b, View - schematic
// LAST TIME SAVED: Jul 24 13:24:39 2007
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g1b ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], sp4_r_v_b[5]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], sp4_r_v_b[6]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], sp4_r_v_b[4]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], sp4_r_v_b[7]}),
     .sp4_out(sp4_v_b[19:18]), .sp12_in({sp12_v_b[15], sp12_v_b[13]}),
     .lc_trk_out(lc_trk_g1[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2a, View - schematic
// LAST TIME SAVED: Jul 24 13:23:46 2007
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g2a ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g2;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;

input [7:0]  lft_op;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnl_op;
input [7:0]  slf_op;
input [1:0]  vdd_cntl;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  bnr_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[33], sp4_r_v_b[9]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[34], sp4_r_v_b[10]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[32], sp4_r_v_b[8]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[35], sp4_r_v_b[11]}),
     .sp4_out(sp4_v_b[21:20]), .sp12_in({sp12_v_b[19], sp12_v_b[17]}),
     .lc_trk_out(lc_trk_g2[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2b, View - schematic
// LAST TIME SAVED: Jul 24 13:22:58 2007
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g2b ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g2;

inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [7:0]  bnr_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[37], sp4_r_v_b[13]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[38], sp4_r_v_b[14]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[36], sp4_r_v_b[12]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[39], sp4_r_v_b[15]}),
     .sp4_out(sp4_v_b[23:22]), .sp12_in({sp12_v_b[23], sp12_v_b[21]}),
     .lc_trk_out(lc_trk_g2[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3a, View - schematic
// LAST TIME SAVED: May 11 14:44:38 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g3a ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g3;

inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  lft_op;
input [7:0]  bot_op;
input [7:0]  top_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
input [7:0]  tnr_op;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  bnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[41], sp4_r_v_b[17]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[42], sp4_r_v_b[18]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[40], sp4_r_v_b[16]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[43], sp4_r_v_b[19]}),
     .sp4_out(sp4_h_r[13:12]), .sp12_in({sp12_h_r[2], sp12_h_r[0]}),
     .lc_trk_out(lc_trk_g3[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3b, View - schematic
// LAST TIME SAVED: May 11 14:44:24 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g3b ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g3;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;

input [7:0]  top_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [7:0]  bot_op;
input [1:0]  wl;
input [7:0]  bnr_op;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [1:0]  vdd_cntl;
input [7:0]  slf_op;
input [7:0]  rgt_op;
input [7:0]  lft_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base I_gmux_12to4_g3b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[45], sp4_r_v_b[21]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[46], sp4_r_v_b[22]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[44], sp4_r_v_b[20]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[47], sp4_r_v_b[23]}),
     .sp4_out(sp4_h_r[15:14]), .sp12_in({sp12_h_r[6], sp12_h_r[4]}),
     .lc_trk_out(lc_trk_g3[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4, View - schematic
// LAST TIME SAVED: Jun  3 14:49:41 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module gmux_sp12to4 ( lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, bl,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bnl_op, bnr_op,
     bot_op, glb2local, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g3;

inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_r_v_b;

input [7:0]  rgt_op;
input [7:0]  top_op;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [7:0]  bnr_op;
input [3:0]  glb2local;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  tnr_op;
input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  tnl_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_g0a I_g0_30 ( .vdd_cntl(vdd_cntl[1:0]),
     .pgate(pgate[1:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp12_v_b(sp12_v_b[23:0]), .lc_trk_g0(lc_trk_g0[3:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g0b I_g0_74 ( .vdd_cntl(vdd_cntl[3:2]),
     .pgate(pgate[3:2]), .glb2local(glb2local[3:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .lc_trk_g0(lc_trk_g0[7:4]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[3:2]), .reset_b(reset_b[3:2]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g1a I_g1_30 ( .vdd_cntl(vdd_cntl[5:4]),
     .pgate(pgate[5:4]), .bl(bl[11:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]),
     .lft_op(lft_op[7:0]), .prog(prog), .rgt_op(rgt_op[7:0]),
     .reset_b(reset_b[5:4]), .slf_op(slf_op[7:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .wl(wl[5:4]), .lc_trk_g1(lc_trk_g1[3:0]));
gmux_sp12to4_g1b I_g1_74 ( .vdd_cntl(vdd_cntl[7:6]),
     .pgate(pgate[7:6]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g1(lc_trk_g1[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g2a I_g2_30 ( .vdd_cntl(vdd_cntl[9:8]), .wl(wl[9:8]),
     .reset_b(reset_b[9:8]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[3:0]), .pgate(pgate[9:8]));
gmux_sp12to4_g2b I_g2_74 ( .vdd_cntl(vdd_cntl[11:10]),
     .pgate(pgate[11:10]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[11:10]),
     .reset_b(reset_b[11:10]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g3a I_g3_30 ( .vdd_cntl(vdd_cntl[13:12]), .wl(wl[13:12]),
     .reset_b(reset_b[13:12]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .pgate(pgate[13:12]), .lc_trk_g3(lc_trk_g3[3:0]));
gmux_sp12to4_g3b I_g3_74 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g3(lc_trk_g3[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .prog(prog),
     .bl(bl[11:0]), .reset_b(reset_b[15:14]), .wl(wl[15:14]));

endmodule
// Library - leafcell, Cell - bram_routing_tracks4_ice1p, View -
//schematic
// LAST TIME SAVED: Jun  2 10:48:34 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_routing_tracks4_ice1p ( bram_cbit, clk, cntl_cbit,
     lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, s_r, bl, sp4_h_l,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r,
     sp12_v_b, sp12_v_t, bnl_op, bnr_op, bot_op, glb_netwk, lft_op,
     pgate, prog, reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op,
     vdd_cntl, wl );
output  clk, s_r;


input  prog;

output [7:0]  cntl_cbit;
output [7:0]  bram_cbit;
output [7:0]  lc_trk_g3;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g1;

inout [47:0]  sp4_v_t;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [23:0]  sp12_h_r;
inout [23:0]  sp12_v_t;
inout [25:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [7:0]  rgt_op;
input [7:0]  tnl_op;
input [15:0]  wl;
input [7:0]  top_op;
input [15:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  bot_op;
input [7:0]  bnl_op;
input [7:0]  tnr_op;
input [7:0]  glb_netwk;
input [15:0]  pgate;
input [7:0]  slf_op;
input [15:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net144;

wire  [1:0]  sp12_v_b_mid;

wire  [3:0]  net_glb2local;

wire  [1:0]  sp12_h_r_mid;



misc_module4_ice1p I_misc ( .cbit_colcntl(cntl_cbit[7:0]),
     .wl(wl[15:0]), .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18],
     sp12_h_r[16], sp12_h_r[14], sp12_h_r[12], sp12_h_r[10],
     sp12_h_r[8]}), .vdd_cntl(vdd_cntl[15:0]), .b(sp12_v_b[1:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .lc_trk_g1(lc_trk_g1[5:0]), .glb2local(net_glb2local[3:0]),
     .bl(bl[3:0]), .min3(glb_netwk[7:0]), .clk(clk),
     .min2(glb_netwk[7:0]), .reset_b(reset_b[15:0]), .prog(progd),
     .m(sp12_v_b_mid[1:0]), .r(sp12_h_r[1:0]), .S_R(s_r),
     .sp4(sp4_h_r[23:16]), .clkb(clkb), .lc_trk_g0(lc_trk_g0[5:0]),
     .glb_netwk(glb_netwk[7:0]), .min1(glb_netwk[7:0]),
     .min0(glb_netwk[7:0]), .l(sp12_h_r_mid[1:0]),
     .pgate(pgate[15:0]));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(progd));
rm8w  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm8w  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm8w  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm8w  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm8w  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm8w  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm8w  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm8w  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm8w  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm8w  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm8w  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm8w  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm8w  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm8w  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm8w  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm8w  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm8w  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm8w  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm8w  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm8w  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm8w  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm8w  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm8w  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm8w  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
span4_ice8p I_sp4_sw ( .ccntrl_cbit(net144[0:7]),
     .bram_cbit(bram_cbit[7:0]), .sp4_h_l(sp4_h_l[47:0]),
     .bl(bl[13:4]), .wl(wl[15:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_t(sp4_v_t[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .reset_b(reset_b[15:0]), .vdd_cntl(vdd_cntl[15:0]),
     .pgate(pgate[15:0]), .prog(progd));
rm7y  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7y  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7y  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7y  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7y  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7y  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7y  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7y  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7y  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7y  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7y  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7y  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7y  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7y  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7y  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7y  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7y  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7y  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7y  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7y  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7y  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7y  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7y  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7y  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
gmux_sp12to4 I_gmux_sp12to4 ( .reset_b(reset_b[15:0]),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .lft_op(lft_op[7:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .glb2local(net_glb2local[3:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .wl(wl[15:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .bl(bl[25:14]), .lc_trk_g3(lc_trk_g3[7:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .vdd_cntl(vdd_cntl[15:0]), .prog(progd));

endmodule
// Library - leafcell, Cell - tiehis, View - schematic
// LAST TIME SAVED: May 12 18:03:23 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module tiehis ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - tiehi, View - schematic
// LAST TIME SAVED: Aug 18 15:41:32 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module tiehi ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - odrv12_30, View - schematic
// LAST TIME SAVED: May 11 14:28:15 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module odrv12_30 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_h_r;

input  prog, slfop;

output [2:0]  sp4_h_r;
output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_r_v_b;

input [11:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



odrv12 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b[1]));
odrv12 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp12(sp12_v_b[0]));
odrv12 I70 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r));
odrv4 I69_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I71_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[2]));
odrv4 I71_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[1]));
odrv4 I71_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp4(sp4_v_b[0]));
odrv4 I73_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I73_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I73_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux3_0, View - schematic
// LAST TIME SAVED: Jun 24 10:59:05 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4k_inmux3_0 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_h_r;

input  op, prog;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min2;
input [15:0]  min1;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
input [15:0]  min3;
input [15:0]  bl;
input [15:0]  min0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [31:0]  cbit;

wire  [31:0]  cbitb;



in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12],
     cbit[13], cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12],
     cbitb[13], cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12_30 I_odrv74 ( .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));

endmodule
// Library - leafcell, Cell - odrv12_74, View - schematic
// LAST TIME SAVED: May 12 12:56:34 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module odrv12_74 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_v_b;

input  prog, slfop;

output [2:0]  sp4_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_h_r;
output [2:0]  sp4_r_v_b;

input [11:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



odrv12 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp12(sp12_h_r[1]));
odrv12 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r[0]));
odrv12 I71 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b));
odrv4 I68_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I68_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I68_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I70_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp4(sp4_v_b[2]));
odrv4 I70_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[1]));
odrv4 I70_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[0]));
odrv4 I72_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux7_4, View - schematic
// LAST TIME SAVED: Jun 24 10:56:58 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4k_inmux7_4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_v_b;

input  op, prog;

output [1:0]  sp12_h_r;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [2:0]  sp4_h_r;

input [1:0]  vdd_cntl;
input [15:0]  min0;
input [15:0]  bl;
input [15:0]  min1;
input [15:0]  min3;
input [1:0]  pgate;
input [1:0]  reset_b;
input [15:0]  min2;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [31:0]  cbit;

wire  [31:0]  cbitb;



in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12],
     cbit[13], cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12],
     cbitb[13], cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
odrv12_74 I_odrv74 ( .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux_8x4, View - schematic
// LAST TIME SAVED: May 12 18:08:28 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4k_inmux_8x4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, op, pgate, prog, reset_b, vdd_cntl, wl );

input  prog;

output [23:0]  sp4_h_r;
output [23:0]  sp4_r_v_b;
output [11:0]  sp12_v_b;
output [11:0]  sp12_h_r;
output [7:0]  in1;
output [7:0]  in2;
output [7:0]  in3;
output [7:0]  in0;
output [23:0]  sp4_v_b;

input [15:0]  bl;
input [7:0]  op;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g3;
input [7:0]  lc_trk_g2;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  reset_b;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I81 ( .A(prog), .Y(progb));
inv I82 ( .A(progb), .Y(progd));
tiehis I10 ( .tiehi(tiehi));
bram_4k_inmux3_0 I3 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[3]), .sp12_v_b(sp12_v_b[7:6]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(progd), .pgate(pgate[7:6]),
     .op(op[3]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[11:9]), .sp4_r_v_b(sp4_r_v_b[11:9]),
     .sp4_h_r(sp4_h_r[11:9]), .in3(in3[3]), .in2(in2[3]), .in1(in1[3]),
     .in0(in0[3]));
bram_4k_inmux3_0 I2 ( .vdd_cntl(vdd_cntl[5:4]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[2]), .sp12_v_b(sp12_v_b[5:4]), .wl(wl[5:4]),
     .reset_b(reset_b[5:4]), .prog(progd), .pgate(pgate[5:4]),
     .op(op[2]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[8:6]), .sp4_r_v_b(sp4_r_v_b[8:6]),
     .sp4_h_r(sp4_h_r[8:6]), .in3(in3[2]), .in2(in2[2]), .in1(in1[2]),
     .in0(in0[2]));
bram_4k_inmux3_0 I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[1]), .sp12_v_b(sp12_v_b[3:2]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(progd), .pgate(pgate[3:2]),
     .op(op[1]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[5:3]), .sp4_r_v_b(sp4_r_v_b[5:3]),
     .sp4_h_r(sp4_h_r[5:3]), .in3(in3[1]), .in2(in2[1]), .in1(in1[1]),
     .in0(in0[1]));
bram_4k_inmux3_0 I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[0]), .sp12_v_b(sp12_v_b[1:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(progd), .pgate(pgate[1:0]),
     .op(op[0]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .in3(in3[0]), .in2(in2[0]), .in1(in1[0]),
     .in0(in0[0]));
bram_4k_inmux7_4 I6 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[15:0]),
     .wl(wl[13:12]), .reset_b(reset_b[13:12]), .prog(progd),
     .pgate(pgate[13:12]), .op(op[6]), .min3({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp12_v_b(sp12_v_b[10]), .sp12_h_r(sp12_h_r[9:8]),
     .sp4_v_b(sp4_v_b[20:18]), .sp4_r_v_b(sp4_r_v_b[20:18]),
     .sp4_h_r(sp4_h_r[20:18]), .in3(in3[6]), .in2(in2[6]),
     .in1(in1[6]), .in0(in0[6]));
bram_4k_inmux7_4 I5 ( .vdd_cntl(vdd_cntl[11:10]), .bl(bl[15:0]),
     .wl(wl[11:10]), .reset_b(reset_b[11:10]), .prog(progd),
     .pgate(pgate[11:10]), .op(op[5]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[9]), .sp12_h_r(sp12_h_r[7:6]),
     .sp4_v_b(sp4_v_b[17:15]), .sp4_r_v_b(sp4_r_v_b[17:15]),
     .sp4_h_r(sp4_h_r[17:15]), .in3(in3[5]), .in2(in2[5]),
     .in1(in1[5]), .in0(in0[5]));
bram_4k_inmux7_4 I4 ( .vdd_cntl(vdd_cntl[9:8]), .bl(bl[15:0]),
     .wl(wl[9:8]), .reset_b(reset_b[9:8]), .prog(progd),
     .pgate(pgate[9:8]), .op(op[4]), .min3({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .sp12_v_b(sp12_v_b[8]),
     .sp12_h_r(sp12_h_r[5:4]), .sp4_v_b(sp4_v_b[14:12]),
     .sp4_r_v_b(sp4_r_v_b[14:12]), .sp4_h_r(sp4_h_r[14:12]),
     .in3(in3[4]), .in2(in2[4]), .in1(in1[4]), .in0(in0[4]));
bram_4k_inmux7_4 I7 ( .vdd_cntl(vdd_cntl[15:14]), .bl(bl[15:0]),
     .wl(wl[15:14]), .reset_b(reset_b[15:14]), .prog(progd),
     .pgate(pgate[15:14]), .op(op[7]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[11]), .sp12_h_r(sp12_h_r[11:10]),
     .sp4_v_b(sp4_v_b[23:21]), .sp4_r_v_b(sp4_r_v_b[23:21]),
     .sp4_h_r(sp4_h_r[23:21]), .in3(in3[7]), .in2(in2[7]),
     .in1(in1[7]), .in0(in0[7]));

endmodule
// Library - ice1chip, Cell - bram_4kprouting_left_ice1p, View -
//schematic
// LAST TIME SAVED: Jun  6 11:31:11 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4kprouting_left_ice1p ( bm_bweb, bm_clkr2rf_n40,
     bm_clkw2rf_n40, bm_d, bm_ren2rf_n40, bm_wen2rf_n40, bram_aa,
     bram_ab, bram_cbit_bot, bram_cbit_top, cntl_cbit_bot,
     cntl_cbit_top, bl, sp4_h_l_bot, sp4_h_l_top, sp4_h_r_bot,
     sp4_h_r_top, sp4_r_v_b_bot, sp4_r_v_b_top, sp4_v_b_bot,
     sp4_v_b_top, sp4_v_t_top, sp12_h_l_bot, sp12_h_l_top,
     sp12_h_r_bot, sp12_h_r_top, sp12_v_b_bot, sp12_v_t_top,
     bnl_op_bot, bnr_op_bot, bot_op_bot, glb_netwk, lft_op_bot,
     lft_op_top, pgate_bot, pgate_top, prog, reset_b_bot, reset_b_top,
     rgt_op_bot, rgt_op_top, slf_op_bot, slf_op_top, tnl_op_top,
     tnr_op_top, top_op_top, vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top
     );
output  bm_clkr2rf_n40, bm_clkw2rf_n40, bm_ren2rf_n40, bm_wen2rf_n40;


input  prog;

output [7:0]  cntl_cbit_bot;
output [7:0]  bram_cbit_top;
output [15:0]  bm_d;
output [7:0]  bram_cbit_bot;
output [10:0]  bram_ab;
output [7:0]  cntl_cbit_top;
output [10:0]  bram_aa;
output [15:0]  bm_bweb;

inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_v_t_top;
inout [41:0]  bl;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_h_r_bot;

input [7:0]  tnl_op_top;
input [7:0]  slf_op_top;
input [15:0]  wl_bot;
input [7:0]  top_op_top;
input [7:0]  rgt_op_bot;
input [15:0]  pgate_bot;
input [7:0]  lft_op_bot;
input [15:0]  reset_b_top;
input [7:0]  bnl_op_bot;
input [7:0]  lft_op_top;
input [7:0]  rgt_op_top;
input [7:0]  tnr_op_top;
input [15:0]  pgate_top;
input [7:0]  bnr_op_bot;
input [7:0]  bot_op_bot;
input [15:0]  reset_b_bot;
input [7:0]  glb_netwk;
input [15:0]  wl_top;
input [15:0]  vdd_cntl_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  slf_op_bot;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net226;

wire  [0:7]  net194;

wire  [0:7]  net195;

wire  [0:7]  net229;

wire  [0:7]  net228;

wire  [0:7]  net227;

wire  [0:7]  net193;

wire  [4:0]  in2_top;

wire  [4:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net196;



inv_hvt I3 ( .A(bram_cbit_bot0), .Y(bram_cbit_bot[0]));
bram_routing_tracks4_ice1p I_bram_routing_tracks4_ice1p_bot (
     .cntl_cbit(cntl_cbit_bot[7:0]), .bram_cbit({bram_cbit_bot[7:1],
     bram_cbit_bot0}), .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15],
     vdd_cntl_bot[12], vdd_cntl_bot[13], vdd_cntl_bot[10],
     vdd_cntl_bot[11], vdd_cntl_bot[8], vdd_cntl_bot[9],
     vdd_cntl_bot[6], vdd_cntl_bot[7], vdd_cntl_bot[4],
     vdd_cntl_bot[5], vdd_cntl_bot[2], vdd_cntl_bot[3],
     vdd_cntl_bot[0], vdd_cntl_bot[1]}), .s_r(bm_wen2rf_n40),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(rgt_op_top[7:0]),
     .tnl_op(lft_op_top[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3(net193[0:7]), .lc_trk_g2(net194[0:7]),
     .lc_trk_g1(net195[0:7]), .lc_trk_g0(net196[0:7]),
     .clk(bm_clkw2rf_n40), .sp12_v_t(sp12_v_b_top[23:0]),
     .sp12_v_b(sp12_v_b_bot[23:0]), .sp12_h_r(sp12_h_r_bot[23:0]),
     .sp12_h_l(sp12_h_l_bot[23:0]), .sp4_v_t(sp4_v_b_top[47:0]),
     .sp4_v_b(sp4_v_b_bot[47:0]), .sp4_r_v_b(sp4_r_v_b_bot[47:0]),
     .sp4_h_r(sp4_h_r_bot[47:0]), .sp4_h_l(sp4_h_l_bot[47:0]),
     .bl(bl[25:0]));
bram_routing_tracks4_ice1p I_bram_routing_tracks4_ice1p_top (
     .cntl_cbit(cntl_cbit_top[7:0]), .bram_cbit(bram_cbit_top[7:0]),
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .s_r(bm_ren2rf_n40), .wl({wl_top[14],
     wl_top[15], wl_top[12], wl_top[13], wl_top[10], wl_top[11],
     wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5],
     wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bot_op(slf_op_bot[7:0]),
     .bnr_op(rgt_op_bot[7:0]), .bnl_op(lft_op_bot[7:0]),
     .lc_trk_g3(net226[0:7]), .lc_trk_g2(net227[0:7]),
     .lc_trk_g1(net228[0:7]), .lc_trk_g0(net229[0:7]),
     .clk(bm_clkr2rf_n40), .sp12_v_t(sp12_v_t_top[23:0]),
     .sp12_v_b(sp12_v_b_top[23:0]), .sp12_h_r(sp12_h_r_top[23:0]),
     .sp12_h_l(sp12_h_l_top[23:0]), .sp4_v_t(sp4_v_t_top[47:0]),
     .sp4_v_b(sp4_v_b_top[47:0]), .sp4_r_v_b(sp4_r_v_b_top[47:0]),
     .sp4_h_r(sp4_h_r_top[47:0]), .sp4_h_l(sp4_h_l_top[47:0]),
     .bl(bl[25:0]));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_bot (
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .bl(bl[41:26]), .wl({wl_bot[14], wl_bot[15],
     wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8],
     wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2],
     wl_bot[3], wl_bot[0], wl_bot[1]}), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .op(slf_op_bot[7:0]), .lc_trk_g3(net193[0:7]),
     .lc_trk_g2(net194[0:7]), .lc_trk_g1(net195[0:7]),
     .lc_trk_g0(net196[0:7]), .sp12_h_r({sp12_h_r_bot[22],
     sp12_h_r_bot[6], sp12_h_r_bot[20], sp12_h_r_bot[4],
     sp12_h_r_bot[18], sp12_h_r_bot[2], sp12_h_r_bot[16],
     sp12_h_r_bot[0], sp12_h_r_bot[14], sp12_h_r_bot[12],
     sp12_h_r_bot[10], sp12_h_r_bot[8]}), .sp4_v_b({sp4_v_b_bot[46],
     sp4_v_b_bot[30], sp4_v_b_bot[14], sp4_v_b_bot[44],
     sp4_v_b_bot[28], sp4_v_b_bot[12], sp4_v_b_bot[42],
     sp4_v_b_bot[26], sp4_v_b_bot[10], sp4_v_b_bot[40],
     sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38], sp4_v_b_bot[22],
     sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20], sp4_v_b_bot[4],
     sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2], sp4_v_b_bot[32],
     sp4_v_b_bot[16], sp4_v_b_bot[0]}), .sp4_r_v_b({sp4_r_v_b_bot[47],
     sp4_r_v_b_bot[31], sp4_r_v_b_bot[15], sp4_r_v_b_bot[45],
     sp4_r_v_b_bot[29], sp4_r_v_b_bot[13], sp4_r_v_b_bot[43],
     sp4_r_v_b_bot[27], sp4_r_v_b_bot[11], sp4_r_v_b_bot[41],
     sp4_r_v_b_bot[25], sp4_r_v_b_bot[9], sp4_r_v_b_bot[39],
     sp4_r_v_b_bot[23], sp4_r_v_b_bot[7], sp4_r_v_b_bot[37],
     sp4_r_v_b_bot[21], sp4_r_v_b_bot[5], sp4_r_v_b_bot[35],
     sp4_r_v_b_bot[19], sp4_r_v_b_bot[3], sp4_r_v_b_bot[33],
     sp4_r_v_b_bot[17], sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46],
     sp4_h_r_bot[30], sp4_h_r_bot[14], sp4_h_r_bot[44],
     sp4_h_r_bot[28], sp4_h_r_bot[12], sp4_h_r_bot[42],
     sp4_h_r_bot[26], sp4_h_r_bot[10], sp4_h_r_bot[40],
     sp4_h_r_bot[24], sp4_h_r_bot[8], sp4_h_r_bot[38], sp4_h_r_bot[22],
     sp4_h_r_bot[6], sp4_h_r_bot[36], sp4_h_r_bot[20], sp4_h_r_bot[4],
     sp4_h_r_bot[34], sp4_h_r_bot[18], sp4_h_r_bot[2], sp4_h_r_bot[32],
     sp4_h_r_bot[16], sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]),
     .in2({in2_bot[4:0], bram_aa[10:8]}), .in1(bm_d[7:0]),
     .in0(bram_aa[7:0]), .sp12_v_b({sp12_v_b_bot[14], sp12_v_b_bot[12],
     sp12_v_b_bot[10], sp12_v_b_bot[8], sp12_v_b_bot[22],
     sp12_v_b_bot[6], sp12_v_b_bot[20], sp12_v_b_bot[4],
     sp12_v_b_bot[18], sp12_v_b_bot[2], sp12_v_b_bot[16],
     sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_top (
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .bl(bl[41:26]), .sp12_v_b({sp12_v_b_top[14],
     sp12_v_b_top[12], sp12_v_b_top[10], sp12_v_b_top[8],
     sp12_v_b_top[22], sp12_v_b_top[6], sp12_v_b_top[20],
     sp12_v_b_top[4], sp12_v_b_top[18], sp12_v_b_top[2],
     sp12_v_b_top[16], sp12_v_b_top[0]}), .wl({wl_top[14], wl_top[15],
     wl_top[12], wl_top[13], wl_top[10], wl_top[11], wl_top[8],
     wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2],
     wl_top[3], wl_top[0], wl_top[1]}), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .op(slf_op_top[7:0]), .lc_trk_g3(net226[0:7]),
     .lc_trk_g2(net227[0:7]), .lc_trk_g1(net228[0:7]),
     .lc_trk_g0(net229[0:7]), .sp12_h_r({sp12_h_r_top[22],
     sp12_h_r_top[6], sp12_h_r_top[20], sp12_h_r_top[4],
     sp12_h_r_top[18], sp12_h_r_top[2], sp12_h_r_top[16],
     sp12_h_r_top[0], sp12_h_r_top[14], sp12_h_r_top[12],
     sp12_h_r_top[10], sp12_h_r_top[8]}), .sp4_v_b({sp4_v_b_top[46],
     sp4_v_b_top[30], sp4_v_b_top[14], sp4_v_b_top[44],
     sp4_v_b_top[28], sp4_v_b_top[12], sp4_v_b_top[42],
     sp4_v_b_top[26], sp4_v_b_top[10], sp4_v_b_top[40],
     sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38], sp4_v_b_top[22],
     sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20], sp4_v_b_top[4],
     sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2], sp4_v_b_top[32],
     sp4_v_b_top[16], sp4_v_b_top[0]}), .sp4_r_v_b({sp4_r_v_b_top[47],
     sp4_r_v_b_top[31], sp4_r_v_b_top[15], sp4_r_v_b_top[45],
     sp4_r_v_b_top[29], sp4_r_v_b_top[13], sp4_r_v_b_top[43],
     sp4_r_v_b_top[27], sp4_r_v_b_top[11], sp4_r_v_b_top[41],
     sp4_r_v_b_top[25], sp4_r_v_b_top[9], sp4_r_v_b_top[39],
     sp4_r_v_b_top[23], sp4_r_v_b_top[7], sp4_r_v_b_top[37],
     sp4_r_v_b_top[21], sp4_r_v_b_top[5], sp4_r_v_b_top[35],
     sp4_r_v_b_top[19], sp4_r_v_b_top[3], sp4_r_v_b_top[33],
     sp4_r_v_b_top[17], sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46],
     sp4_h_r_top[30], sp4_h_r_top[14], sp4_h_r_top[44],
     sp4_h_r_top[28], sp4_h_r_top[12], sp4_h_r_top[42],
     sp4_h_r_top[26], sp4_h_r_top[10], sp4_h_r_top[40],
     sp4_h_r_top[24], sp4_h_r_top[8], sp4_h_r_top[38], sp4_h_r_top[22],
     sp4_h_r_top[6], sp4_h_r_top[36], sp4_h_r_top[20], sp4_h_r_top[4],
     sp4_h_r_top[34], sp4_h_r_top[18], sp4_h_r_top[2], sp4_h_r_top[32],
     sp4_h_r_top[16], sp4_h_r_top[0]}), .in3(bm_bweb[15:8]),
     .in2({in2_top[4:0], bram_ab[10:8]}), .in1(bm_d[15:8]),
     .in0(bram_ab[7:0]));

endmodule
// Library - leafcell, Cell - bram_2mux, View - schematic
// LAST TIME SAVED: Jun 24 10:40:59 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_2mux ( out, c, in0, in1 );
output  out;

input  c, in0, in1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate I14 ( .in(in1), .out(net52), .pp(net045), .nn(c));
txgate I33 ( .in(in0), .out(net52), .pp(c), .nn(net045));
inv I15 ( .A(net52), .Y(net029));
inv I0 ( .A(net029), .Y(out));
inv_hvt I1 ( .A(c), .Y(net045));

endmodule
// Library - leafcell, Cell - bram_cascade_addr, View - schematic
// LAST TIME SAVED: Jan  2 17:57:15 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_cascade_addr ( addr_2bot, addr_muxo, addr, addr_top, cbit,
     prog );

input  prog;

output [10:0]  addr_2bot;
output [10:0]  addr_muxo;

input [10:0]  addr_top;
input [10:0]  addr;
input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(cbit[1]), .Y(net71));
bram_bufferx4 I33 ( .in(cbit[0]), .out(net66));
nor2_hvt I65 ( .A(prog), .B(net71), .Y(net69));
spn4dbuf I_addr_2bot_10_ ( .T(net69), .A(addr_muxo[10]),
     .Y(addr_2bot[10]));
spn4dbuf I_addr_2bot_9_ ( .T(net69), .A(addr_muxo[9]),
     .Y(addr_2bot[9]));
spn4dbuf I_addr_2bot_8_ ( .T(net69), .A(addr_muxo[8]),
     .Y(addr_2bot[8]));
spn4dbuf I_addr_2bot_7_ ( .T(net69), .A(addr_muxo[7]),
     .Y(addr_2bot[7]));
spn4dbuf I_addr_2bot_6_ ( .T(net69), .A(addr_muxo[6]),
     .Y(addr_2bot[6]));
spn4dbuf I_addr_2bot_5_ ( .T(net69), .A(addr_muxo[5]),
     .Y(addr_2bot[5]));
spn4dbuf I_addr_2bot_4_ ( .T(net69), .A(addr_muxo[4]),
     .Y(addr_2bot[4]));
spn4dbuf I_addr_2bot_3_ ( .T(net69), .A(addr_muxo[3]),
     .Y(addr_2bot[3]));
spn4dbuf I_addr_2bot_2_ ( .T(net69), .A(addr_muxo[2]),
     .Y(addr_2bot[2]));
spn4dbuf I_addr_2bot_1_ ( .T(net69), .A(addr_muxo[1]),
     .Y(addr_2bot[1]));
spn4dbuf I_addr_2bot_0_ ( .T(net69), .A(addr_muxo[0]),
     .Y(addr_2bot[0]));
bram_2mux I_bram_2mux_10_ ( .c(net66), .out(addr_muxo[10]),
     .in0(addr[10]), .in1(addr_top[10]));
bram_2mux I_bram_2mux_9_ ( .c(net66), .out(addr_muxo[9]),
     .in0(addr[9]), .in1(addr_top[9]));
bram_2mux I_bram_2mux_8_ ( .c(net66), .out(addr_muxo[8]),
     .in0(addr[8]), .in1(addr_top[8]));
bram_2mux I_bram_2mux_7_ ( .c(net66), .out(addr_muxo[7]),
     .in0(addr[7]), .in1(addr_top[7]));
bram_2mux I_bram_2mux_6_ ( .c(net66), .out(addr_muxo[6]),
     .in0(addr[6]), .in1(addr_top[6]));
bram_2mux I_bram_2mux_5_ ( .c(net66), .out(addr_muxo[5]),
     .in0(addr[5]), .in1(addr_top[5]));
bram_2mux I_bram_2mux_4_ ( .c(net66), .out(addr_muxo[4]),
     .in0(addr[4]), .in1(addr_top[4]));
bram_2mux I_bram_2mux_3_ ( .c(net66), .out(addr_muxo[3]),
     .in0(addr[3]), .in1(addr_top[3]));
bram_2mux I_bram_2mux_2_ ( .c(net66), .out(addr_muxo[2]),
     .in0(addr[2]), .in1(addr_top[2]));
bram_2mux I_bram_2mux_1_ ( .c(net66), .out(addr_muxo[1]),
     .in0(addr[1]), .in1(addr_top[1]));
bram_2mux I_bram_2mux_0_ ( .c(net66), .out(addr_muxo[0]),
     .in0(addr[0]), .in1(addr_top[0]));

endmodule
// Library - leafcell, Cell - bram_2mux_lvt, View - schematic
// LAST TIME SAVED: Nov  8 18:34:36 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_2mux_lvt ( out, c, in0, in1 );
output  out;

input  c, in0, in1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I14 ( .in(in1), .out(net52), .pp(net045), .nn(c));
txgate_lvt I33 ( .in(in0), .out(net52), .pp(c), .nn(net045));
inv_lvt I15 ( .A(net52), .Y(net029));
inv_lvt I0 ( .A(net029), .Y(out));
inv_hvt I1 ( .A(c), .Y(net045));

endmodule
// Library - misc, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: May 13 14:45:34 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ml_mux2_hvt ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - tielo, View - schematic
// LAST TIME SAVED: Jul 23 17:02:44 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module tielo ( tielo );
output  tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M1 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));
nch_hvt  M2 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - leafcell, Cell - rf_4k_n40, View - schematic
// LAST TIME SAVED: Aug 16 16:53:19 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module rf_4k_n40 ( Q, AA, AB, AMA, AMB, BIST, BWEB, BWEBM, CLKR, CLKW,
     D, DM, PD, REB, REBM, WEB, WEBM );

input  BIST, CLKR, CLKW, PD, REB, REBM, WEB, WEBM;

output [15:0]  Q;

input [7:0]  AMA;
input [15:0]  DM;
input [7:0]  AA;
input [15:0]  D;
input [15:0]  BWEB;
input [15:0]  BWEBM;
input [7:0]  AB;
input [7:0]  AMB;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: May 12 17:56:32 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ml_mux2_hvt_schematic ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - bram_dff_mux, View - schematic
// LAST TIME SAVED: Oct  4 14:55:56 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_dff_mux ( q, bm_q, bm_sdi, ce, clk, rcapmux_en, rst );
output  q;

input  bm_q, bm_sdi, ce, clk, rcapmux_en, rst;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_mux2_hvt I5 ( .in1(net14), .in0(q), .out(net020), .sel(ce));
ml_dff I_ml_dff ( .R(rst), .D(net020), .CLK(clk), .QN(net10), .Q(q));
ml_mux2_hvt_schematic I1 ( .in1(bm_q), .in0(bm_sdi), .out(net14),
     .sel(rcapmux_en));

endmodule
// Library - leafcell, Cell - bram_4k_sr_v1, View - schematic
// LAST TIME SAVED: Oct 29 10:24:13 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4k_sr_v1 ( bm_dm, bm_sdo, bm_sweb, clk, rcapmux_en, rst,
     bm_q, bm_sdi, wdummymux_en );
output  bm_sdo;

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff I_dff15 ( .R(rst), .D(bm_dm[14]), .CLK(clk), .QN(net0258),
     .Q(rdummy_reg));
ml_dff I_dff0 ( .R(rst), .D(bm_sdi), .CLK(clk), .QN(net157),
     .Q(wdummy_reg));
bram_dff_mux I_dff_mux_15_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[14]),
     .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I_dff_mux_14_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[13]),
     .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I_dff_mux_13_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[12]),
     .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I_dff_mux_12_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[11]),
     .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I_dff_mux_11_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[10]),
     .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I_dff_mux_10_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[9]),
     .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I_dff_mux_9_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[8]),
     .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I_dff_mux_8_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[7]),
     .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I_dff_mux_7_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[6]),
     .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I_dff_mux_6_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[5]),
     .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I_dff_mux_5_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[4]),
     .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I_dff_mux_4_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[3]),
     .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I_dff_mux_3_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[2]),
     .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I_dff_mux_2_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[1]),
     .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I_dff_mux_1_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(net150),
     .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I_dff_mux_0_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[0]), .q(bm_dm[0]));
ml_mux2_hvt_schematic I_mux15 ( .in1(rdummy_reg), .in0(bm_dm[15]),
     .out(bm_sdo), .sel(rcapmux_en));
ml_mux2_hvt_schematic I_mux0 ( .in1(wdummy_reg), .in0(bm_dm[0]),
     .out(net150), .sel(wdummymux_en));

endmodule
// Library - leafcell, Cell - bram_4k_n40, View - schematic
// LAST TIME SAVED: Jan  2 17:48:30 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4k_n40 ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_pd, bm_rcapmux_en, bm_ren, bm_sa,
     bm_sclk, bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en,
     bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_pd, bm_rcapmux_en, bm_ren,
     bm_sclk, bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en,
     bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [7:0]  bm_sa;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [7:0]  bm_aa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  bm_dm;



bram_2mux_lvt I22 ( .c(bm_init), .out(net108), .in0(bm_clkr),
     .in1(bm_sclkrw));
bram_2mux_lvt I23 ( .c(bm_init), .out(net110), .in0(bm_clkw),
     .in1(bm_sclkrw));
inv_lvt I6 ( .A(bm_ren), .Y(reb));
inv_lvt I5 ( .A(bm_wen), .Y(web));
ml_mux2_hvt I20 ( .in1(net90), .in0(bm_pd), .out(net0118),
     .sel(bm_init));
bram_bufferx4 I19 ( .in(net0118), .out(net0111));
rf_4k_n40 I_rf_4k ( .PD(net0111), .DM(bm_dm[15:0]), .WEBM(bm_sweb),
     .WEB(web), .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]),
     .CLKW(net110), .CLKR(net108), .BWEBM({net0128, net0128, net0128,
     net0128, net0128, net0128, net0128, net0128, net0128, net0128,
     net0128, net0128, net0128, net0128, net0128, net0128}),
     .BWEB(bm_bweb[15:0]), .BIST(bm_init), .AMB(bm_sa[7:0]),
     .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]), .AA(bm_aa[7:0]),
     .Q(bm_q[15:0]));
bram_4k_sr_v1 I_bram_4k_sr ( .bm_sdo(bm_sdo), .bm_dm(bm_dm[15:0]),
     .rst(net90), .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
tielo I15 ( .tielo(net0128));
tielo I18 ( .tielo(net90));

endmodule
// Library - leafcell, Cell - o_mux_out_bram, View - schematic
// LAST TIME SAVED: Jun 24 10:30:25 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module o_mux_out_bram ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I181 ( .A(in), .Y(out));

endmodule
// Library - leafcell, Cell - bram_3muxinv, View - schematic
// LAST TIME SAVED: Jun 24 10:39:04 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_3muxinv ( out, c, .cdsNet0(in[0]), .cdsNet0(in[1]),
     .cdsNet0(in[2]) );
output  out;


input [2:0]  in;
input [1:0]  c;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  ci;

wire  [1:0]  cb;



txgate_lvt I21 ( .in(in[2]), .out(net52), .pp(cb[1]), .nn(ci[1]));
txgate_lvt I33 ( .in(in[0]), .out(net52), .pp(net048), .nn(net053));
txgate_lvt I20 ( .in(in[1]), .out(net52), .pp(net045), .nn(net051));
inv_lvt I0 ( .A(net52), .Y(out));
nand2_hvt I15 ( .A(ci[0]), .Y(net045), .B(cb[1]));
nand2_hvt I2 ( .A(cb[0]), .Y(net048), .B(cb[1]));
inv_hvt I19 ( .A(net045), .Y(net051));
inv_hvt I18 ( .A(net048), .Y(net053));
inv_hvt I14_1_ ( .A(c[1]), .Y(cb[1]));
inv_hvt I14_0_ ( .A(c[0]), .Y(cb[0]));
inv_hvt I1_1_ ( .A(cb[1]), .Y(ci[1]));
inv_hvt I1_0_ ( .A(cb[0]), .Y(ci[0]));

endmodule
// Library - leafcell, Cell - bram_2muxinv, View - schematic
// LAST TIME SAVED: Jun 24 10:38:19 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_2muxinv ( out, c, in0, in1 );
output  out;

input  c, in0, in1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I13 ( .in(in1), .out(net52), .pp(net045), .nn(c));
txgate_lvt I33 ( .in(in0), .out(net52), .pp(c), .nn(net045));
inv_lvt I0 ( .A(net52), .Y(out));
inv_hvt I1 ( .A(c), .Y(net045));

endmodule
// Library - leafcell, Cell - bram_rd_decoder0to7, View - schematic
// LAST TIME SAVED: Jun 24 10:39:29 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_rd_decoder0to7 ( rd, c, raq, rdi );


output [7:0]  rd;

input [1:0]  c;
input [7:0]  rdi;
input [10:8]  raq;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cb;

wire  [10:10]  raqb;

wire  [1:0]  cd;



nand2 I65 ( .A(mode16_b), .Y(raq8_b), .B(raq[8]));
inv I85 ( .A(raq[9]), .Y(net0245));
inv I68 ( .A(raq[10]), .Y(raqb[10]));
o_mux_out_bram I69 ( .in(net360), .out(rd[0]));
o_mux_out_bram I92 ( .out(rd[7]), .in(net378));
o_mux_out_bram I91 ( .out(rd[6]), .in(net333));
o_mux_out_bram I90 ( .out(rd[5]), .in(net372));
o_mux_out_bram I89 ( .out(rd[4]), .in(net362));
o_mux_out_bram I88 ( .out(rd[3]), .in(net390));
o_mux_out_bram I87 ( .out(rd[2]), .in(net329));
o_mux_out_bram I86 ( .out(rd[1]), .in(net384));
inv_lvt I104 ( .A(rdi[7]), .Y(net378));
nand2_hvt I106 ( .A(cd[1]), .Y(mode4_b), .B(cb[0]));
nand2_hvt I107 ( .A(cd[1]), .Y(mode2_b), .B(cd[0]));
nand2_hvt I105 ( .A(cb[1]), .Y(mode16_b), .B(cb[0]));
inv_hvt I22_1_ ( .A(cb[1]), .Y(cd[1]));
inv_hvt I22_0_ ( .A(cb[0]), .Y(cd[0]));
inv_hvt I53_1_ ( .A(c[1]), .Y(cb[1]));
inv_hvt I53_0_ ( .A(c[0]), .Y(cb[0]));
bram_3muxinv I3 ( net390, {mode2_b, raqb[10]}, net285, net357, rdi[3]);
bram_2muxinv I35 ( .in1(rdi[2]), .c(raq8_b), .out(net329),
     .in0(rdi[3]));
bram_2muxinv I36 ( .in1(rdi[4]), .c(raq8_b), .out(net362),
     .in0(rdi[5]));
bram_2muxinv I37 ( .in1(rdi[6]), .c(raq8_b), .out(net333),
     .in0(rdi[7]));
bram_2muxinv I34 ( .in1(rdi[0]), .c(raq8_b), .out(net360),
     .in0(rdi[1]));
bram_2muxinv I42 ( .in1(net360), .c(net0245), .out(net357),
     .in0(net329));
bram_2muxinv I43 ( .in1(net362), .c(net0245), .out(net285),
     .in0(net333));
bram_2muxinv I49 ( .in1(rdi[5]), .c(mode4_b), .out(net372),
     .in0(net285));
bram_2muxinv I50 ( .in1(rdi[1]), .c(mode4_b), .out(net384),
     .in0(net357));

endmodule
// Library - leafcell, Cell - bram_4muxinv, View - schematic
// LAST TIME SAVED: Jan  2 18:09:52 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4muxinv ( out, .cdsNet0(in[0]), .cdsNet0(in[1]),
     .cdsNet0(in[2]), .cdsNet0(in[3]), sel, selb );
output  out;


input [3:0]  selb;
input [3:0]  sel;
input [3:0]  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I0 ( .A(net47), .Y(out));
txgate_lvt I19 ( .in(in[3]), .out(net47), .pp(selb[3]), .nn(sel[3]));
txgate_lvt I17 ( .in(in[2]), .out(net47), .pp(selb[2]), .nn(sel[2]));
txgate_lvt I33 ( .in(in[0]), .out(net47), .pp(selb[0]), .nn(sel[0]));
txgate_lvt I16 ( .in(in[1]), .out(net47), .pp(selb[1]), .nn(sel[1]));

endmodule
// Library - leafcell, Cell - mux4plldly, View - schematic
// LAST TIME SAVED: Jun 28 10:07:29 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module mux4plldly ( mout, cbit, min );
output  mout;


input [1:0]  cbit;
input [3:0]  min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cbit_b;



txgate_hvt I11 ( .in(net_2_0), .out(net52), .pp(cbit[1]),
     .nn(cbit_b[1]));
txgate_hvt I8 ( .in(min[1]), .out(net_2_0), .pp(cbit_b[0]),
     .nn(cbit[0]));
txgate_hvt I9 ( .in(min[2]), .out(net_2_1), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I12 ( .in(net_2_1), .out(net52), .pp(cbit_b[1]),
     .nn(cbit[1]));
txgate_hvt Itg20 ( .in(min[0]), .out(net_2_0), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I10 ( .in(min[3]), .out(net_2_1), .pp(cbit_b[0]),
     .nn(cbit[0]));
inv_hvt I1_1_ ( .A(cbit[1]), .Y(cbit_b[1]));
inv_hvt I1_0_ ( .A(cbit[0]), .Y(cbit_b[0]));
inv_hvt I0 ( .A(net52), .Y(mout));

endmodule
// Library - leafcell, Cell - bram_wd_decoder0to7, View - schematic
// LAST TIME SAVED: Jun 24 10:50:20 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_wd_decoder0to7 ( wd, sel, wdi );


output [7:0]  wd;

input [3:0]  sel;
input [7:0]  wdi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  selb;

wire  [0:3]  net0202;

wire  [0:3]  net0210;



inv I74 ( .A(wdi[1]), .Y(net176));
inv I75 ( .A(wdi[2]), .Y(net162));
inv I76 ( .A(wdi[3]), .Y(net177));
inv I77 ( .A(wdi[3]), .Y(net159));
inv I78 ( .A(wdi[4]), .Y(net150));
inv I79 ( .A(wdi[5]), .Y(net152));
inv I80 ( .A(wdi[6]), .Y(net138));
inv I81 ( .A(wdi[7]), .Y(net132));
inv I22 ( .A(wdi[0]), .Y(net174));
bram_4muxinv I95 ( wd[5], net152, net150, net152, net159, net0202[0:3],
     selb[3:0]);
bram_4muxinv I96 ( wd[6], net138, net138, net152, net159, net0202[0:3],
     selb[3:0]);
bram_4muxinv I97 ( wd[7], net132, net138, net152, net159, net0202[0:3],
     selb[3:0]);
bram_4muxinv I91 ( wd[1], net176, net174, net176, net177, net0202[0:3],
     selb[3:0]);
bram_4muxinv I92 ( wd[2], net162, net162, net176, net177, net0202[0:3],
     selb[3:0]);
bram_4muxinv I93 ( wd[3], net177, net162, net176, net159, net0202[0:3],
     selb[3:0]);
bram_4muxinv I94 ( wd[4], net150, net150, net152, net159, net0202[0:3],
     selb[3:0]);
bram_4muxinv I3 ( wd[0], net174, net174, net176, net177, net0202[0:3],
     selb[3:0]);
inv_hvt I122_3_ ( .A(net0210[0]), .Y(net0202[0]));
inv_hvt I122_2_ ( .A(net0210[1]), .Y(net0202[1]));
inv_hvt I122_1_ ( .A(net0210[2]), .Y(net0202[2]));
inv_hvt I122_0_ ( .A(net0210[3]), .Y(net0202[3]));
inv_hvt I125_3_ ( .A(sel[3]), .Y(selb[3]));
inv_hvt I125_2_ ( .A(sel[2]), .Y(selb[2]));
inv_hvt I125_1_ ( .A(sel[1]), .Y(selb[1]));
inv_hvt I125_0_ ( .A(sel[0]), .Y(selb[0]));
inv_hvt I123_3_ ( .A(sel[3]), .Y(net0210[0]));
inv_hvt I123_2_ ( .A(sel[2]), .Y(net0210[1]));
inv_hvt I123_1_ ( .A(sel[1]), .Y(net0210[2]));
inv_hvt I123_0_ ( .A(sel[0]), .Y(net0210[3]));

endmodule
// Library - leafcell, Cell - bram_4mux, View - schematic
// LAST TIME SAVED: Jun 24 10:52:41 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4mux ( out, .cdsNet0(in[0]), .cdsNet0(in[1]),
     .cdsNet0(in[2]), .cdsNet0(in[3]), sel, selb );
output  out;


input [3:0]  sel;
input [3:0]  in;
input [3:0]  selb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I13 ( .A(net62), .Y(net48));
inv I14 ( .A(net48), .Y(out));
txgate_lvt I26 ( .in(in[3]), .out(net62), .pp(selb[3]), .nn(sel[3]));
txgate_lvt I33 ( .in(in[0]), .out(net62), .pp(selb[0]), .nn(sel[0]));
txgate_lvt I24 ( .in(in[1]), .out(net62), .pp(selb[1]), .nn(sel[1]));
txgate_lvt I25 ( .in(in[2]), .out(net62), .pp(selb[2]), .nn(sel[2]));

endmodule
// Library - leafcell, Cell - bram_wd_bweb, View - schematic
// LAST TIME SAVED: Jun 24 10:54:56 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_wd_bweb ( bweb, bwebi, sel, wai );


output [15:0]  bweb;

input [10:8]  wai;
input [3:0]  sel;
input [15:0]  bwebi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net0282;

wire  [3:0]  selb;

wire  [10:8]  wa_b;

wire  [0:2]  net168;

wire  [0:3]  net0226;

wire  [10:8]  wa;



nand2 I105 ( .A(wa[8]), .Y(nandwa89), .B(wa[9]));
nand2 I2 ( .A(wa_b[8]), .B(wa_b[9]), .Y(nandwa8b9b));
nand2 I104 ( .A(wa_b[8]), .Y(nandwa8b9), .B(wa[9]));
nand2 I103 ( .A(wa[8]), .Y(nandwa89b), .B(wa_b[9]));
nand3 I60 ( .C(wa_b[10]), .A(wa_b[8]), .Y(nandwa8b9b10b), .B(wa_b[9]));
nand3 I98 ( .Y(nandwa8910b), .B(wa[9]), .C(wa_b[10]), .A(wa[8]));
nand3 I97 ( .Y(nandwa8b910b), .B(wa[9]), .C(wa_b[10]), .A(wa_b[8]));
nand3 I96 ( .Y(nandwa89b10b), .B(wa_b[9]), .C(wa_b[10]), .A(wa[8]));
nand3 I99 ( .Y(nandwa8b9b10), .B(wa_b[9]), .C(wa[10]), .A(wa_b[8]));
nand3 I100 ( .Y(nandwa89b10), .B(wa_b[9]), .C(wa[10]), .A(wa[8]));
nand3 I101 ( .Y(nandwa8b910), .B(wa[9]), .C(wa[10]), .A(wa_b[8]));
nand3 I102 ( .Y(nandwa8910), .B(wa[9]), .C(wa[10]), .A(wa[8]));
inv I106 ( .A(wa_b[8]), .Y(wa8));
inv I71 ( .A(wa[8]), .Y(wa8b));
inv I82_2_ ( .A(wai[10]), .Y(net168[0]));
inv I82_1_ ( .A(wai[9]), .Y(net168[1]));
inv I82_0_ ( .A(wai[8]), .Y(net168[2]));
inv I95_2_ ( .A(wai[10]), .Y(wa_b[10]));
inv I95_1_ ( .A(wai[9]), .Y(wa_b[9]));
inv I95_0_ ( .A(wai[8]), .Y(wa_b[8]));
inv I83_2_ ( .A(net168[0]), .Y(wa[10]));
inv I83_1_ ( .A(net168[1]), .Y(wa[9]));
inv I83_0_ ( .A(net168[2]), .Y(wa[8]));
bram_4mux I107 ( bweb[1], bwebi[1], wa8b, nandwa89b, nandwa89b10b,
     net0226[0:3], selb[3:0]);
bram_4mux I108 ( bweb[2], bwebi[2], wa8, nandwa8b9, nandwa8b910b,
     net0226[0:3], selb[3:0]);
bram_4mux I109 ( bweb[3], bwebi[3], wa8b, nandwa89, nandwa8910b,
     net0226[0:3], selb[3:0]);
bram_4mux I110 ( bweb[4], bwebi[4], wa8, nandwa8b9b, nandwa8b9b10,
     net0226[0:3], selb[3:0]);
bram_4mux I111 ( bweb[5], bwebi[5], wa8b, nandwa89b, nandwa89b10,
     net0226[0:3], selb[3:0]);
bram_4mux I112 ( bweb[6], bwebi[6], wa8, nandwa8b9, nandwa8b910,
     net0226[0:3], selb[3:0]);
bram_4mux I113 ( bweb[7], bwebi[7], wa8b, nandwa89, nandwa8910,
     net0226[0:3], selb[3:0]);
bram_4mux I114 ( bweb[8], bwebi[8], wa8, nandwa8b9b, nandwa8b9b10b,
     net0226[0:3], selb[3:0]);
bram_4mux I115 ( bweb[9], bwebi[9], wa8b, nandwa89b, nandwa89b10b,
     net0226[0:3], selb[3:0]);
bram_4mux I116 ( bweb[10], bwebi[10], wa8, nandwa8b9, nandwa8b910b,
     net0226[0:3], selb[3:0]);
bram_4mux I117 ( bweb[11], bwebi[11], wa8b, nandwa89, nandwa8910b,
     net0226[0:3], selb[3:0]);
bram_4mux I118 ( bweb[12], bwebi[12], wa8, nandwa8b9b, nandwa8b9b10,
     net0226[0:3], selb[3:0]);
bram_4mux I119 ( bweb[13], bwebi[13], wa8b, nandwa89b, nandwa89b10,
     net0226[0:3], selb[3:0]);
bram_4mux I120 ( bweb[14], bwebi[14], wa8, nandwa8b9, nandwa8b910,
     net0226[0:3], selb[3:0]);
bram_4mux I121 ( bweb[15], bwebi[15], wa8b, nandwa89, nandwa8910,
     net0226[0:3], selb[3:0]);
bram_4mux I40 ( bweb[0], bwebi[0], wa8, nandwa8b9b, nandwa8b9b10b,
     net0226[0:3], selb[3:0]);
inv_hvt I122_3_ ( .A(net0282[0]), .Y(net0226[0]));
inv_hvt I122_2_ ( .A(net0282[1]), .Y(net0226[1]));
inv_hvt I122_1_ ( .A(net0282[2]), .Y(net0226[2]));
inv_hvt I122_0_ ( .A(net0282[3]), .Y(net0226[3]));
inv_hvt I123_3_ ( .A(sel[3]), .Y(net0282[0]));
inv_hvt I123_2_ ( .A(sel[2]), .Y(net0282[1]));
inv_hvt I123_1_ ( .A(sel[1]), .Y(net0282[2]));
inv_hvt I123_0_ ( .A(sel[0]), .Y(net0282[3]));
inv_hvt I125_3_ ( .A(sel[3]), .Y(selb[3]));
inv_hvt I125_2_ ( .A(sel[2]), .Y(selb[2]));
inv_hvt I125_1_ ( .A(sel[1]), .Y(selb[1]));
inv_hvt I125_0_ ( .A(sel[0]), .Y(selb[0]));

endmodule
// Library - leafcell, Cell - bram_bufferx6, View - schematic
// LAST TIME SAVED: Jan  2 18:54:54 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_bufferx6 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - bram_4k_buffer, View - schematic
// LAST TIME SAVED: Sep 30 18:29:20 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4k_buffer ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;

input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I14 ( .in(bm_sdo_i), .out(bm_sdo_o));
bram_bufferx6 I6 ( .in(bm_sdi_i), .out(bm_sdi_o));
bram_bufferx6 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx6 I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx6 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx6 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx6 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx6 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx6 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx6 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx6 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx6 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx6 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx6 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx6 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx6 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx6 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbank_pbuffer_v1, View -
//schematic
// LAST TIME SAVED: Jan  2 18:54:22 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_v1 ( bm_aa_2bot, bm_ab_2bot, bm_init_o,
     bm_q, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bm_aa,
     bm_aa_top, bm_ab, bm_ab_top, bm_bweb, bm_clkr, bm_clkw, bm_d,
     bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen, cbit, prog );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen, prog;

output [10:0]  bm_aa_2bot;
output [1:0]  bm_sclkrw_o;
output [10:0]  bm_ab_2bot;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [10:0]  bm_aa_top;
input [10:0]  bm_ab_top;
input [1:0]  bm_sweb_i;
input [1:0]  bm_sdo_i;
input [10:0]  bm_aa;
input [1:0]  bm_sdi_i;
input [10:0]  bm_ab;
input [7:0]  bm_sa_i;
input [8:0]  cbit;
input [1:0]  bm_sclkrw_i;
input [15:0]  bm_d;
input [15:0]  bm_bweb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  net231;

wire  [0:2]  net200;

wire  [0:2]  net232;

wire  [0:15]  net236;

wire  [15:0]  bm_q_fromip;

wire  [0:8]  cbitb;

wire  [10:0]  bm_ab_2ip;

wire  [1:0]  cbitd;

wire  [10:0]  bm_aa_2ip;

wire  [15:0]  bm_d_2ip;

wire  [3:0]  sel;



inv_hvt I41 ( .A(net178), .Y(sel[2]));
inv_hvt I55_1_ ( .A(cbitb[1]), .Y(cbitd[1]));
inv_hvt I55_0_ ( .A(cbitb[0]), .Y(cbitd[0]));
inv_hvt I43 ( .A(cbit[8]), .Y(cbitb[8]));
inv_hvt I54_1_ ( .A(cbit[1]), .Y(cbitb[1]));
inv_hvt I54_0_ ( .A(cbit[0]), .Y(cbitb[0]));
inv_hvt I56 ( .A(net172), .Y(sel[0]));
inv_hvt I42 ( .A(net175), .Y(sel[3]));
inv_hvt I40 ( .A(net181), .Y(sel[1]));
bram_cascade_addr I_cascade_addr4ra ( .prog(prog),
     .addr_2bot(bm_ab_2bot[10:0]), .cbit(cbit[7:6]),
     .addr_top(bm_ab_top[10:0]), .addr(bm_ab[10:0]),
     .addr_muxo(bm_ab_2ip[10:0]));
bram_cascade_addr I_cascade_addr4wa ( .prog(prog),
     .addr_2bot(bm_aa_2bot[10:0]), .cbit(cbit[5:4]),
     .addr_top(bm_aa_top[10:0]), .addr(bm_aa[10:0]),
     .addr_muxo(bm_aa_2ip[10:0]));
bram_4k_n40 I_bram_4k ( .bm_pd(cbitb[8]), .bm_ab(bm_ab_2ip[7:0]),
     .bm_aa(bm_aa_2ip[7:0]), .bm_q(bm_q_fromip[15:0]),
     .bm_sclk(bm_sclk_o), .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(net236[0:15]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d_2ip[15:0]), .bm_clkw(bm_clkw),
     .bm_sdo(net246));
bram_rd_decoder0to7 I_bram_rd_decoder8to15 ( .rd(bm_q[15:8]),
     .rdi(bm_q_fromip[15:8]), .c(cbit[3:2]), .raq(net200[0:2]));
bram_rd_decoder0to7 I_bram_rd_decoder0to7 ( .c(cbit[3:2]),
     .rd(bm_q[7:0]), .raq(net200[0:2]), .rdi(bm_q_fromip[7:0]));
bram_wd_decoder0to7 I_bram_wd_decoder8to15 ( .wd(bm_d_2ip[15:8]),
     .wdi(bm_d[15:8]), .sel(sel[3:0]));
bram_wd_decoder0to7 I_bram_wd_decoder0to7 ( .wd(bm_d_2ip[7:0]),
     .sel(sel[3:0]), .wdi(bm_d[7:0]));
nand2_hvt I92 ( .A(cbitb[0]), .Y(net172), .B(cbitb[1]));
nand2_hvt I39 ( .A(cbitd[0]), .Y(net175), .B(cbitd[1]));
nand2_hvt I38 ( .A(cbitb[0]), .Y(net178), .B(cbitd[1]));
nand2_hvt I37 ( .A(cbitd[0]), .Y(net181), .B(cbitb[1]));
inv I46_2_ ( .A(net231[0]), .Y(net200[0]));
inv I46_1_ ( .A(net231[1]), .Y(net200[1]));
inv I46_0_ ( .A(net231[2]), .Y(net200[2]));
ml_dff I_RAQ_2_ ( .R(prog), .D(bm_ab_2ip[10]), .CLK(bm_clkr),
     .QN(net231[0]), .Q(net232[0]));
ml_dff I_RAQ_1_ ( .R(prog), .D(bm_ab_2ip[9]), .CLK(bm_clkr),
     .QN(net231[1]), .Q(net232[1]));
ml_dff I_RAQ_0_ ( .R(prog), .D(bm_ab_2ip[8]), .CLK(bm_clkr),
     .QN(net231[2]), .Q(net232[2]));
bram_wd_bweb I_bram_wd_bweb ( .sel(sel[3:0]), .wai(bm_aa_2ip[10:8]),
     .bwebi(bm_bweb[15:0]), .bweb(net236[0:15]));
bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k_buffer I_bram_4k_buffer ( .bm_sdo_o(bm_sdo_o[0]),
     .bm_sdo_i(net246), .bm_sclkrw_i(bm_sclkrw_i[0]),
     .bm_sclkrw_o(bm_sclkrw_o[0]), .bm_sdi_o(bm_sdi_o[0]),
     .bm_sdi_i(bm_sdi_i[0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - ice1chip, Cell - bram_4kprouting_ice1p, View - schematic
// LAST TIME SAVED: Jun  6 10:11:51 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram_4kprouting_ice1p ( bm_aa_2bot, bm_ab_2bot, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, cntl_cbit_bot,
     cntl_cbit_top, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_aa_top, bm_ab_top, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_bot,
     bnr_op_bot, bot_op_bot, glb_netwk, lft_op_bot, lft_op_top,
     pgate_bot, pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot,
     rgt_op_top, tnl_op_top, tnr_op_top, top_op_top, vdd_cntl_bot,
     vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [1:0]  bm_sclkrw_o;
output [10:0]  bm_aa_2bot;
output [10:0]  bm_ab_2bot;
output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sweb_o;
output [7:0]  cntl_cbit_top;
output [7:0]  cntl_cbit_bot;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_h_r_bot;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_v_b_top;
inout [23:0]  sp12_h_r_top;
inout [41:0]  bl;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_v_b_bot;

input [7:0]  rgt_op_bot;
input [15:0]  reset_b_bot;
input [15:0]  pgate_bot;
input [15:0]  reset_b_top;
input [7:0]  lft_op_top;
input [15:0]  vdd_cntl_top;
input [7:0]  top_op_top;
input [7:0]  bnr_op_bot;
input [15:0]  wl_bot;
input [1:0]  bm_sdo_i;
input [7:0]  tnl_op_top;
input [7:0]  lft_op_bot;
input [10:0]  bm_ab_top;
input [7:0]  tnr_op_top;
input [7:0]  glb_netwk;
input [7:0]  rgt_op_top;
input [1:0]  bm_sdi_i;
input [15:0]  vdd_cntl_bot;
input [15:0]  wl_top;
input [1:0]  bm_sclkrw_i;
input [15:0]  pgate_top;
input [1:0]  bm_sweb_i;
input [7:0]  bnl_op_bot;
input [7:0]  bot_op_bot;
input [10:0]  bm_aa_top;
input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  bram_ab;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [10:0]  bram_aa;

wire  [7:0]  bram_cbit_bot;

wire  [7:0]  bram_cbit_top;



bram_4kprouting_left_ice1p I_bram_4kprouting_left_ice1p (
     .slf_op_top(slf_op_top[7:0]), .slf_op_bot(slf_op_bot[7:0]),
     .wl_bot(wl_bot[15:0]), .top_op_top(top_op_top[7:0]),
     .sp12_h_l_bot(sp12_h_l_bot[23:0]),
     .sp4_h_l_bot(sp4_h_l_bot[47:0]), .tnl_op_top(tnl_op_top[7:0]),
     .reset_b_top(reset_b_top[15:0]), .reset_b_bot(reset_b_bot[15:0]),
     .vdd_cntl_top(vdd_cntl_top[15:0]), .prog(prog),
     .pgate_top(pgate_top[15:0]), .pgate_bot(pgate_bot[15:0]),
     .lft_op_bot(lft_op_bot[7:0]), .bot_op_bot(bot_op_bot[7:0]),
     .rgt_op_bot(rgt_op_bot[7:0]), .bnl_op_bot(bnl_op_bot[7:0]),
     .sp4_h_r_top(sp4_h_r_top[47:0]),
     .sp12_v_t_top(sp12_v_t_top[23:0]),
     .sp12_v_b_bot(sp12_v_b_bot[23:0]),
     .sp4_h_r_bot(sp4_h_r_bot[47:0]),
     .sp12_h_r_bot(sp12_h_r_bot[23:0]),
     .sp4_v_t_top(sp4_v_t_top[47:0]), .sp4_v_b_bot(sp4_v_b_bot[47:0]),
     .sp12_h_r_top(sp12_h_r_top[23:0]), .bl(bl[41:0]),
     .sp4_h_l_top(sp4_h_l_top[47:0]), .lft_op_top(lft_op_top[7:0]),
     .wl_top(wl_top[15:0]), .sp12_h_l_top(sp12_h_l_top[23:0]),
     .sp4_v_b_top(sp4_v_b_top[47:0]), .rgt_op_top(rgt_op_top[7:0]),
     .vdd_cntl_bot(vdd_cntl_bot[15:0]), .bnr_op_bot(bnr_op_bot[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_bot[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_top[47:0]),
     .cntl_cbit_bot(cntl_cbit_bot[7:0]),
     .cntl_cbit_top(cntl_cbit_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bram_ab(bram_ab[10:0]), .bram_aa(bram_aa[10:0]),
     .bm_bweb(bm_bweb[15:0]), .bm_clkr2rf_n40(bm_clkr2rf_n40),
     .bm_clkw2rf_n40(bm_clkw2rf_n40), .bm_d(bm_d[15:0]),
     .bm_ren2rf_n40(bm_ren2rf_n40), .bm_wen2rf_n40(bm_wen2rf_n40),
     .bram_cbit_top(bram_cbit_top[7:0]),
     .bram_cbit_bot(bram_cbit_bot[7:0]), .tnr_op_top(tnr_op_top[7:0]));
bram_4kbank_pbuffer_v1 I_bram_4kbank_pbuffer ( .cbit({bram_cbit_bot[0],
     bram_cbit_top[7:0]}), .bm_aa(bram_aa[10:0]), .prog(prog),
     .bm_ab(bram_ab[10:0]), .bm_aa_2bot(bm_aa_2bot[10:0]),
     .bm_ab_2bot(bm_ab_2bot[10:0]), .bm_aa_top(bm_aa_top[10:0]),
     .bm_ab_top(bm_ab_top[10:0]), .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(bm_ren2rf_n40),
     .bm_wen(bm_wen2rf_n40), .bm_d(bm_d[15:0]),
     .bm_clkr(bm_clkr2rf_n40), .bm_clkw(bm_clkw2rf_n40),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));

endmodule
// Library - leafcell, Cell - clk_colbuf12k_icc, View - schematic
// LAST TIME SAVED: Jun 23 08:09:26 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module clk_colbuf12k_icc ( clko, cbit, clki );
output  clko;

input  cbit, clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_lvt I_nand2_lvt ( .A(clki), .Y(clkb), .B(cbit));
nch_lvt  M1 ( .D(clko), .B(gnd_), .G(clkb), .S(net7));
nch_lvt  M2 ( .D(net7), .B(gnd_), .G(cbit), .S(gnd_));
pch_lvt  M0 ( .D(clko), .B(vdd_), .G(clkb), .S(vdd_));

endmodule
// Library - ice8chip, Cell - clk_col_buf_x8_ice8p, View - schematic
// LAST TIME SAVED: Jun 23 08:10:00 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module clk_col_buf_x8_ice8p ( col_clk, clk_in, colbuf_cntl );


output [7:0]  col_clk;

input [7:0]  clk_in;
input [7:0]  colbuf_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_colbuf12k_icc I_colbuf12k_7_ ( .clki(clk_in[7]), .clko(col_clk[7]),
     .cbit(colbuf_cntl[7]));
clk_colbuf12k_icc I_colbuf12k_6_ ( .clki(clk_in[6]), .clko(col_clk[6]),
     .cbit(colbuf_cntl[6]));
clk_colbuf12k_icc I_colbuf12k_5_ ( .clki(clk_in[5]), .clko(col_clk[5]),
     .cbit(colbuf_cntl[5]));
clk_colbuf12k_icc I_colbuf12k_4_ ( .clki(clk_in[4]), .clko(col_clk[4]),
     .cbit(colbuf_cntl[4]));
clk_colbuf12k_icc I_colbuf12k_3_ ( .clki(clk_in[3]), .clko(col_clk[3]),
     .cbit(colbuf_cntl[3]));
clk_colbuf12k_icc I_colbuf12k_2_ ( .clki(clk_in[2]), .clko(col_clk[2]),
     .cbit(colbuf_cntl[2]));
clk_colbuf12k_icc I_colbuf12k_1_ ( .clki(clk_in[1]), .clko(col_clk[1]),
     .cbit(colbuf_cntl[1]));
clk_colbuf12k_icc I_colbuf12k_0_ ( .clki(clk_in[0]), .clko(col_clk[0]),
     .cbit(colbuf_cntl[0]));

endmodule
// Library - ice1chip, Cell - bram1x4_ice1f, View - schematic
// LAST TIME SAVED: Jun  6 10:13:33 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module bram1x4_ice1f ( bm_aa_2bot, bm_ab_2bot, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, glb_netwk_bot,
     glb_netwk_top, slf_op_01, slf_op_02, slf_op_03, slf_op_04,
     slf_op_05, slf_op_06, slf_op_07, slf_op_08, bl, pgate, reset_b,
     sp4_h_l_01, sp4_h_l_02, sp4_h_l_03, sp4_h_l_04, sp4_h_l_05,
     sp4_h_l_06, sp4_h_l_07, sp4_h_l_08, sp4_h_r_01, sp4_h_r_02,
     sp4_h_r_03, sp4_h_r_04, sp4_h_r_05, sp4_h_r_06, sp4_h_r_07,
     sp4_h_r_08, sp4_r_v_b_01, sp4_r_v_b_02, sp4_r_v_b_03,
     sp4_r_v_b_04, sp4_r_v_b_05, sp4_r_v_b_06, sp4_r_v_b_07,
     sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03, sp4_v_b_04,
     sp4_v_b_05, sp4_v_b_06, sp4_v_b_07, sp4_v_b_08, sp4_v_t_08,
     sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04, sp12_h_l_05,
     sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_r_01, sp12_h_r_02,
     sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06, sp12_h_r_07,
     sp12_h_r_08, sp12_v_b_01, sp12_v_t_08, vdd_cntl, wl, bm_aa_top,
     bm_ab_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_01, bnr_op_01, bot_op_01, glb_netwk_col,
     lft_op_01, lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06,
     lft_op_07, lft_op_08, prog, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, tnl_op_08,
     tnr_op_08, top_op_08 );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [7:0]  slf_op_06;
output [7:0]  slf_op_04;
output [1:0]  bm_sclkrw_o;
output [10:0]  bm_ab_2bot;
output [1:0]  bm_sdi_o;
output [10:0]  bm_aa_2bot;
output [1:0]  bm_sweb_o;
output [7:0]  glb_netwk_bot;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_08;
output [7:0]  slf_op_07;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_05;
output [7:0]  slf_op_03;
output [7:0]  glb_netwk_top;
output [7:0]  slf_op_02;
output [7:0]  slf_op_01;

inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_h_l_06;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_h_l_07;
inout [23:0]  sp12_h_l_05;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_h_r_08;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_r_v_b_01;
inout [23:0]  sp12_h_l_02;
inout [23:0]  sp12_h_r_01;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_v_b_05;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_h_r_07;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_v_t_08;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_r_v_b_04;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_r_08;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_v_t_08;
inout [47:0]  sp4_v_b_03;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_h_l_04;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_v_b_07;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_v_b_06;
inout [41:0]  bl;
inout [47:0]  sp4_r_v_b_05;
inout [23:0]  sp12_v_b_01;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_h_r_03;
inout [23:0]  sp12_h_l_04;
inout [143:16]  pgate;
inout [23:0]  sp12_h_r_07;
inout [143:16]  reset_b;
inout [23:0]  sp12_h_r_06;
inout [143:16]  vdd_cntl;
inout [143:16]  wl;
inout [23:0]  sp12_h_r_04;

input [7:0]  rgt_op_08;
input [7:0]  lft_op_08;
input [7:0]  rgt_op_06;
input [1:0]  bm_sweb_i;
input [7:0]  lft_op_06;
input [7:0]  rgt_op_04;
input [10:0]  bm_aa_top;
input [7:0]  glb_netwk_col;
input [10:0]  bm_ab_top;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_05;
input [7:0]  bnr_op_01;
input [1:0]  bm_sdo_i;
input [7:0]  bm_sa_i;
input [7:0]  lft_op_07;
input [7:0]  lft_op_02;
input [7:0]  lft_op_01;
input [7:0]  top_op_08;
input [7:0]  bot_op_01;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_01;
input [7:0]  lft_op_05;
input [7:0]  rgt_op_02;
input [1:0]  bm_sdi_i;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_03;
input [7:0]  tnl_op_08;
input [7:0]  lft_op_04;
input [1:0]  bm_sclkrw_i;
input [7:0]  bnl_op_01;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net985;

wire  [0:7]  net1049;

wire  [7:0]  colbuf_cntl_bot;

wire  [0:1]  net930;

wire  [0:23]  net1023;

wire  [0:7]  net928;

wire  [0:7]  net1177;

wire  [0:7]  net0666;

wire  [0:7]  net1119;

wire  [0:7]  net0501;

wire  [0:7]  net1120;

wire  [0:23]  net1151;

wire  [0:10]  net0807;

wire  [0:1]  net933;

wire  [0:7]  net863;

wire  [0:1]  net1121;

wire  [0:10]  net0806;

wire  [0:10]  net01011;

wire  [0:10]  net0874;

wire  [0:1]  net997;

wire  [0:1]  net993;

wire  [0:1]  net1127;

wire  [0:10]  net01010;

wire  [0:23]  net959;

wire  [0:1]  net999;

wire  [0:1]  net1125;

wire  [0:10]  net0875;

wire  [0:1]  net929;

wire  [0:1]  net935;

wire  [0:1]  net1122;

wire  [7:0]  colbuf_cntl_top;

wire  [0:1]  net994;



bram_4kprouting_ice1p I_bram_0825_08 ( .cntl_cbit_top(net0666[0:7]),
     .cntl_cbit_bot(net863[0:7]), .bm_aa_2bot(net0806[0:10]),
     .bm_ab_2bot(net0807[0:10]), .bm_aa_top(bm_aa_top[10:0]),
     .bm_ab_top(bm_ab_top[10:0]), .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sclkrw_i(net930[0:1]),
     .bm_sweb_i(net933[0:1]), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_sdi_i(net929[0:1]), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdo_o(net935[0:1]), .slf_op_top(slf_op_08[7:0]),
     .slf_op_bot(slf_op_07[7:0]), .wl_bot(wl[127:112]),
     .top_op_top(top_op_08[7:0]), .sp12_h_l_bot(sp12_h_l_07[23:0]),
     .sp4_h_l_bot(sp4_h_l_07[47:0]), .tnl_op_top(tnl_op_08[7:0]),
     .reset_b_top(reset_b[143:128]), .reset_b_bot(reset_b[127:112]),
     .vdd_cntl_top(vdd_cntl[143:128]), .prog(prog),
     .pgate_top(pgate[143:128]), .pgate_bot(pgate[127:112]),
     .lft_op_bot(lft_op_07[7:0]), .glb_netwk(glb_netwk_top[7:0]),
     .bm_wdummymux_en_i(net988), .bot_op_bot(slf_op_06[7:0]),
     .rgt_op_bot(rgt_op_07[7:0]), .bnl_op_bot(lft_op_06[7:0]),
     .sp4_h_r_top(sp4_h_r_08[47:0]), .sp12_v_t_top(sp12_v_t_08[23:0]),
     .sp12_v_b_bot(net959[0:23]), .bm_init_i(net984),
     .sp4_h_r_bot(sp4_h_r_07[47:0]), .sp12_h_r_bot(sp12_h_r_07[23:0]),
     .sp4_v_t_top(sp4_v_t_08[47:0]), .sp4_v_b_bot(sp4_v_b_07[47:0]),
     .sp12_h_r_top(sp12_h_r_08[23:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net983), .sp4_h_l_top(sp4_h_l_08[47:0]),
     .lft_op_top(lft_op_08[7:0]), .wl_top(wl[143:128]),
     .sp12_h_l_top(sp12_h_l_08[23:0]), .sp4_v_b_top(sp4_v_b_08[47:0]),
     .tnr_op_top(tnr_op_08[7:0]), .rgt_op_top(rgt_op_08[7:0]),
     .bm_sa_i(net985[0:7]), .bm_sclk_i(net986), .bm_sreb_i(net987),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .vdd_cntl_bot(vdd_cntl[127:112]), .bnr_op_bot(rgt_op_06[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_07[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_08[47:0]));
bram_4kprouting_ice1p I_bram_0825_06 ( .cntl_cbit_top(net928[0:7]),
     .cntl_cbit_bot(colbuf_cntl_top[7:0]), .bm_aa_2bot(net0874[0:10]),
     .bm_ab_2bot(net0875[0:10]), .bm_aa_top(net0806[0:10]),
     .bm_ab_top(net0807[0:10]), .bm_sdi_o(net929[0:1]),
     .bm_sclkrw_o(net930[0:1]), .bm_sclkrw_i(net994[0:1]),
     .bm_sweb_i(net997[0:1]), .bm_sweb_o(net933[0:1]),
     .bm_sdi_i(net993[0:1]), .bm_sdo_i(net935[0:1]),
     .bm_sdo_o(net999[0:1]), .slf_op_top(slf_op_06[7:0]),
     .slf_op_bot(slf_op_05[7:0]), .wl_top(wl[111:96]),
     .wl_bot(wl[95:80]), .top_op_top(slf_op_07[7:0]),
     .tnl_op_top(lft_op_07[7:0]), .reset_b_top(reset_b[111:96]),
     .reset_b_bot(reset_b[95:80]), .prog(prog),
     .pgate_top(pgate[111:96]), .pgate_bot(pgate[95:80]),
     .lft_op_top(lft_op_06[7:0]), .lft_op_bot(lft_op_05[7:0]),
     .glb_netwk(glb_netwk_top[7:0]), .bm_wdummymux_en_i(net1052),
     .bot_op_bot(slf_op_04[7:0]), .sp4_h_r_top(sp4_h_r_06[47:0]),
     .bnl_op_bot(lft_op_04[7:0]), .bnr_op_bot(rgt_op_04[7:0]),
     .sp4_h_r_bot(sp4_h_r_05[47:0]), .sp12_v_t_top(net959[0:23]),
     .sp12_v_b_bot(net1023[0:23]), .bm_init_i(net1048),
     .sp12_h_l_top(sp12_h_l_06[23:0]),
     .sp12_h_r_bot(sp12_h_r_05[23:0]),
     .sp12_h_l_bot(sp12_h_l_05[23:0]),
     .sp12_h_r_top(sp12_h_r_06[23:0]), .sp4_v_t_top(sp4_v_b_07[47:0]),
     .sp4_v_b_top(sp4_v_b_06[47:0]), .sp4_v_b_bot(sp4_v_b_05[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_05[47:0]),
     .sp4_h_l_top(sp4_h_l_06[47:0]), .tnr_op_top(rgt_op_07[7:0]),
     .sp4_h_l_bot(sp4_h_l_05[47:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net1047), .sp4_r_v_b_top(sp4_r_v_b_06[47:0]),
     .rgt_op_bot(rgt_op_05[7:0]), .rgt_op_top(rgt_op_06[7:0]),
     .bm_sa_i(net1049[0:7]), .bm_sclk_i(net1050), .bm_sreb_i(net1051),
     .bm_rcapmux_en_o(net983), .bm_init_o(net984),
     .bm_sa_o(net985[0:7]), .bm_sclk_o(net986), .bm_sreb_o(net987),
     .bm_wdummymux_en_o(net988), .vdd_cntl_top(vdd_cntl[111:96]),
     .vdd_cntl_bot(vdd_cntl[95:80]));
bram_4kprouting_ice1p I_bram_0825_04 ( .cntl_cbit_top(net0501[0:7]),
     .cntl_cbit_bot(colbuf_cntl_bot[7:0]), .bm_aa_2bot(net01010[0:10]),
     .bm_ab_2bot(net01011[0:10]), .bm_aa_top(net0874[0:10]),
     .bm_ab_top(net0875[0:10]), .bm_sdi_o(net993[0:1]),
     .bm_sclkrw_o(net994[0:1]), .bm_sclkrw_i(net1122[0:1]),
     .bm_sweb_i(net1125[0:1]), .bm_sweb_o(net997[0:1]),
     .bm_sdi_i(net1121[0:1]), .bm_sdo_i(net999[0:1]),
     .bm_sdo_o(net1127[0:1]), .slf_op_top(slf_op_04[7:0]),
     .slf_op_bot(slf_op_03[7:0]), .wl_top(wl[79:64]),
     .wl_bot(wl[63:48]), .top_op_top(slf_op_05[7:0]),
     .tnl_op_top(lft_op_05[7:0]), .reset_b_top(reset_b[79:64]),
     .reset_b_bot(reset_b[63:48]), .prog(prog),
     .pgate_top(pgate[79:64]), .pgate_bot(pgate[63:48]),
     .lft_op_top(lft_op_04[7:0]), .lft_op_bot(lft_op_03[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]), .bm_wdummymux_en_i(net1180),
     .bot_op_bot(slf_op_02[7:0]), .sp4_h_r_top(sp4_h_r_04[47:0]),
     .bnl_op_bot(lft_op_02[7:0]), .bnr_op_bot(rgt_op_02[7:0]),
     .sp4_h_r_bot(sp4_h_r_03[47:0]), .sp12_v_t_top(net1023[0:23]),
     .sp12_v_b_bot(net1151[0:23]), .bm_init_i(net1176),
     .sp12_h_l_top(sp12_h_l_04[23:0]),
     .sp12_h_r_bot(sp12_h_r_03[23:0]),
     .sp12_h_l_bot(sp12_h_l_03[23:0]),
     .sp12_h_r_top(sp12_h_r_04[23:0]), .sp4_v_t_top(sp4_v_b_05[47:0]),
     .sp4_v_b_top(sp4_v_b_04[47:0]), .sp4_v_b_bot(sp4_v_b_03[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_03[47:0]),
     .sp4_h_l_top(sp4_h_l_04[47:0]), .tnr_op_top(rgt_op_05[7:0]),
     .sp4_h_l_bot(sp4_h_l_03[47:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net1175), .sp4_r_v_b_top(sp4_r_v_b_04[47:0]),
     .rgt_op_bot(rgt_op_03[7:0]), .rgt_op_top(rgt_op_04[7:0]),
     .bm_sa_i(net1177[0:7]), .bm_sclk_i(net1178), .bm_sreb_i(net1179),
     .bm_rcapmux_en_o(net1047), .bm_init_o(net1048),
     .bm_sa_o(net1049[0:7]), .bm_sclk_o(net1050), .bm_sreb_o(net1051),
     .bm_wdummymux_en_o(net1052), .vdd_cntl_top(vdd_cntl[79:64]),
     .vdd_cntl_bot(vdd_cntl[63:48]));
bram_4kprouting_ice1p I_bram_0825_02 ( .cntl_cbit_top(net1120[0:7]),
     .cntl_cbit_bot(net1119[0:7]), .bm_aa_2bot(bm_aa_2bot[10:0]),
     .bm_ab_2bot(bm_ab_2bot[10:0]), .bm_aa_top(net01010[0:10]),
     .bm_ab_top(net01011[0:10]), .bm_sdi_o(net1121[0:1]),
     .bm_sclkrw_o(net1122[0:1]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sweb_o(net1125[0:1]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sdo_i(net1127[0:1]),
     .bm_sdo_o(bm_sdo_o[1:0]), .slf_op_top(slf_op_02[7:0]),
     .slf_op_bot(slf_op_01[7:0]), .wl_top(wl[47:32]),
     .wl_bot(wl[31:16]), .top_op_top(slf_op_03[7:0]),
     .tnl_op_top(lft_op_03[7:0]), .reset_b_top(reset_b[47:32]),
     .reset_b_bot(reset_b[31:16]), .prog(prog),
     .pgate_top(pgate[47:32]), .pgate_bot(pgate[31:16]),
     .lft_op_top(lft_op_02[7:0]), .lft_op_bot(lft_op_01[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_01[7:0]), .sp4_h_r_top(sp4_h_r_02[47:0]),
     .bnl_op_bot(bnl_op_01[7:0]), .bnr_op_bot(bnr_op_01[7:0]),
     .sp4_h_r_bot(sp4_h_r_01[47:0]), .sp12_v_t_top(net1151[0:23]),
     .sp12_v_b_bot(sp12_v_b_01[23:0]), .bm_init_i(bm_init_i),
     .sp12_h_l_top(sp12_h_l_02[23:0]),
     .sp12_h_r_bot(sp12_h_r_01[23:0]),
     .sp12_h_l_bot(sp12_h_l_01[23:0]),
     .sp12_h_r_top(sp12_h_r_02[23:0]), .sp4_v_t_top(sp4_v_b_03[47:0]),
     .sp4_v_b_top(sp4_v_b_02[47:0]), .sp4_v_b_bot(sp4_v_b_01[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_01[47:0]),
     .sp4_h_l_top(sp4_h_l_02[47:0]), .tnr_op_top(rgt_op_03[7:0]),
     .sp4_h_l_bot(sp4_h_l_01[47:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .sp4_r_v_b_top(sp4_r_v_b_02[47:0]), .rgt_op_bot(rgt_op_01[7:0]),
     .rgt_op_top(rgt_op_02[7:0]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(net1175), .bm_init_o(net1176),
     .bm_sa_o(net1177[0:7]), .bm_sclk_o(net1178), .bm_sreb_o(net1179),
     .bm_wdummymux_en_o(net1180), .vdd_cntl_top(vdd_cntl[47:32]),
     .vdd_cntl_bot(vdd_cntl[31:16]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_top (
     .colbuf_cntl(colbuf_cntl_top[7:0]), .col_clk(glb_netwk_top[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_bot (
     .colbuf_cntl(colbuf_cntl_bot[7:0]), .col_clk(glb_netwk_bot[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - delay150ps, View - schematic
// LAST TIME SAVED: Dec 21 17:50:49 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module delay150ps ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I4 ( .A(in), .Y(net12));
inv_hvt I0 ( .A(net013), .Y(out));
inv_hvt I6 ( .A(net12), .Y(net17));
inv_hvt I2 ( .A(net17), .Y(net013));

endmodule
// Library - io, Cell - ioin_mux_v3, View - schematic
// LAST TIME SAVED: Jun 24 11:14:10 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioin_mux_v3 ( inmuxo, cbit,
     cbitb, min[7:0], prog );
output  inmuxo;

input  prog;

input [3:0]  cbitb;
input [3:0]  cbit;
input [7:0]  min;
supply1 vdd_;
supply0 gnd_;
//////////wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_lvt I282 ( .A(prog), .Y(en), .B(cbitb[3]));
inv_lvt I281 ( .A(inmuxob), .Y(inmuxo));
nand2_lvt I_nand2 ( .A(st2), .Y(inmuxob), .B(en));
txgate_lvt I285 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I289 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I286 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I283 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_lvt I292 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I293 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I291 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I294 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I287 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I290 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I288 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I295 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I284 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc_v0, View - schematic
// LAST TIME SAVED: Dec  7 10:49:57 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc_v0 ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  spi;
output [1:0]  ti;

inout [5:0]  bl;

input [7:0]  min2;
input [7:0]  min1;
input [1:0]  vdd_cntl;
input [7:0]  min0;
input [1:0]  reset;
input [1:0]  padin;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



ioin_mux_v3 I_ioin_mux_bankcntl ( bankcntl, {cbit[11], cbit[8], cbit[9],
     cbit[10]}, {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0],
     prog);
ioin_mux_v3 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v3 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
inv_lvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_lvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
nor2_lvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_lvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nand2inv_v0, View - schematic
// LAST TIME SAVED: Dec  7 10:48:43 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioinmx2nand2inv_v0 ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  reset;
input [7:0]  min0;
input [7:0]  min1;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [7:0]  ce;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;

wire  [11:0]  cbit;



ioin_mux_v3 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v3 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
nand2_lvt I180 ( .A(update_b), .Y(updt), .B(bs_en));
inv_lvt I181 ( .A(update), .Y(update_b));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioin_mux_v2, View - schematic
// LAST TIME SAVED: Jun 24 11:10:53 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioin_mux_v2 ( inmuxo, cbit,
     cbitb, min[7:0], prog );
output  inmuxo;

input  prog;

input [3:0]  cbit;
input [7:0]  min;
input [3:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//////////wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_lvt I_nor2_lvt ( .A(prog), .Y(en), .B(cbitb[3]));
inv_lvt I281 ( .A(inmuxob), .Y(inmuxo));
nand2_lvt I_nand2 ( .A(st2), .Y(inmuxob), .B(en));
txgate_lvt I285 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I289 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I286 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I283 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_lvt I292 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I293 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I291 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I294 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I287 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I290 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I288 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I295 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I284 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));

endmodule
// Library - io, Cell - ioinmx1mux2_v1, View - schematic
// LAST TIME SAVED: Jun 24 11:09:14 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module ioinmx1mux2_v1 ( clk, ti, bl, ce, ceb, min, pgate, prog, reset,
     vdd_cntl, wl );
output  clk, ti;


input  ceb, prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [7:0]  min;
input [11:0]  ce;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;



clk_mux12to1_icc I_clk_mux12to1 ( .prog(prog), .min(ce[11:0]),
     .clk(clk), .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7],
     cbitb[10], cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7],
     cbit[10], cbit[6], cbit[4]}), .cenb(ceb));
ioin_mux_v2 I_ioin_mux ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1mem, View - schematic
// LAST TIME SAVED: Jun 24 11:12:19 2011
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox1mem ( b, bl, l, r, t, pgate, prog, reset, vdd_cntl, wl );
inout  b, l, r, t;

input  prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;



sbox1m3to1_icc I232 ( .in2(r), .cb({cbitb[3], cbitb[6]}), .op(t),
     .in0(l), .in1(b), .c({cbit[3], cbit[6]}), .prog(prog));
sbox1m3to1_icc I230 ( .in2(r), .cb({cbitb[1], cbitb[4]}), .op(l),
     .in0(b), .in1(t), .c({cbit[1], cbit[4]}), .prog(prog));
sbox1m3to1_icc I226 ( .in2(r), .cb({cbitb[8], cbitb[5]}), .op(b),
     .in0(l), .in1(t), .c({cbit[8], cbit[5]}), .prog(prog));
sbox1m3to1_icc I231 ( .in2(b), .cb({cbitb[10], cbitb[7]}), .op(r),
     .in0(l), .in1(t), .c({cbit[10], cbit[7]}), .prog(prog));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc_v4, View - schematic
// LAST TIME SAVED: Dec  7 10:50:25 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module sbox1_colbdlc_v4 ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [5:0]  ti;

inout [5:0]  bl;
inout [3:0]  r;
inout [3:0]  l;
inout [3:0]  sp4_v_b;
inout [3:0]  t_mid;

input [1:0]  oeb;
input [7:0]  min1;
input [1:0]  padin;
input [7:0]  min3;
input [7:0]  min4;
input [7:0]  min6;
input [11:0]  clk_in;
input [1:0]  out;
input [7:0]  min0;
input [11:0]  inclk_in;
input [1:0]  spioeb;
input [1:0]  spiout;
input [7:0]  ceb_in;
input [15:0]  reset;
input [7:0]  min2;
input [15:0]  vdd_cntl;
input [7:0]  min5;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spioob;

wire  [1:0]  spioo;

wire  [1:0]  oeboo;

wire  [1:0]  oeboob;



ioinmx2nor2invx2bdlc_v0 I5 ( .vdd_cntl(vdd_cntl[5:4]),
     .min2(min6[7:0]), .bankcntl(fabric_out), .bl(bl[5:0]),
     .prog(prog), .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx2nand2inv_v0 I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
ioinmx1mux2_v1 I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .ti(ti[2]), .min(min2[7:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]));
ioinmx1mux2_v1 I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .ti(ti[5]), .min(min5[7:0]), .wl(wl[15:14]), .reset(reset[15:14]),
     .pgate(pgate[15:14]));
inv_lvt I_inv_2_1_ ( .A(spioob[1]), .Y(pado[1]));
inv_lvt I_inv_2_0_ ( .A(spioob[0]), .Y(pado[0]));
inv_lvt I9_1_ ( .A(oeboo[1]), .Y(oeboob[1]));
inv_lvt I9_0_ ( .A(oeboo[0]), .Y(oeboob[0]));
inv_lvt I8_1_ ( .A(oeboob[1]), .Y(padeb[1]));
inv_lvt I8_0_ ( .A(oeboob[0]), .Y(padeb[0]));
inv_lvt inv_1_1_ ( .A(spioo[1]), .Y(spioob[1]));
inv_lvt inv_1_0_ ( .A(spioo[0]), .Y(spioob[0]));
mux2x1_hvt I10_1_ ( .in1(oeb[1]), .in0(spioeb[1]), .out(oeboo[1]),
     .sel(cdone_in));
mux2x1_hvt I10_0_ ( .in1(oeb[0]), .in0(spioeb[0]), .out(oeboo[0]),
     .sel(cdone_in));
mux2x1_hvt I_emux_1_ ( .in1(out[1]), .in0(spiout[1]), .out(spioo[1]),
     .sel(cdone_in));
mux2x1_hvt I_emux_0_ ( .in1(out[0]), .in0(spiout[0]), .out(spioo[0]),
     .sel(cdone_in));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - io, Cell - io_gmux_x2v3, View - schematic
// LAST TIME SAVED: Aug 25 13:36:12 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_gmux_x2v3 ( .cbit_colcntl({cbit[11], cbit[9]}), gout, bl,
     min0, min1, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [11:0]  cbit;
output [1:0]  gout;

inout [5:0]  bl;

input [15:0]  min1;
input [15:0]  min0;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux I_g_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux I_g_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare_v4, View - schematic
// LAST TIME SAVED: Aug 25 13:36:24 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module io_gmux_x16bare_v4 ( cbit_colcntl, lc_trk_g0, lc_trk_g1, bl,
     min0, min1, min2, min3, min4, min5, min6, min7, min8, min9, min10,
     min11, min12, min13, min14, min15, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [7:0]  cbit_colcntl;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g1;

inout [5:0]  bl;

input [15:0]  min9;
input [15:0]  min12;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min0;
input [15:0]  min7;
input [15:0]  min5;
input [15:0]  min3;
input [15:0]  min4;
input [15:0]  min10;
input [15:0]  min6;
input [15:0]  min8;
input [15:0]  min15;
input [15:0]  min14;
input [15:0]  min11;
input [15:0]  reset;
input [15:0]  min2;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net187;

wire  [0:1]  net114;

wire  [0:1]  net124;

wire  [0:1]  net188;



io_gmux_x2v3 I_io_gmux_x2_7 ( .cbit_colcntl(net114[0:1]),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[15:14]));
io_gmux_x2v3 I_io_gmux_x2_6 ( .cbit_colcntl(net124[0:1]),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[13:12]));
io_gmux_x2v3 I_io_gmux_x2_2 ( .cbit_colcntl(cbit_colcntl[5:4]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[5:4]));
io_gmux_x2v3 I_io_gmux_x2_0 ( .cbit_colcntl(cbit_colcntl[1:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[1:0]));
io_gmux_x2v3 _io_gmux_x2_1 ( .cbit_colcntl(cbit_colcntl[3:2]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[3:2]));
io_gmux_x2v3 I_io_gmux_x2_4 ( .cbit_colcntl(net187[0:1]),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[9:8]));
io_gmux_x2v3 I_io_gmux_x2_5 ( .cbit_colcntl(net188[0:1]),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[11:10]));
io_gmux_x2v3 I_io_gmux_x2_3 ( .cbit_colcntl(cbit_colcntl[7:6]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[7:6]));

endmodule
// Library - io, Cell - insel1_lvt_imp, View - schematic
// LAST TIME SAVED: Aug 12 13:25:22 2010
// NETLIST TIME: Jun 29 10:32:24 2011
`timescale 1ns / 1ns 

module insel1_lvt_imp ( out, in0, in1, in2, in3, sb, sel );
output  out;

input  in0, in1, in2, in3;

input [1:0]  sb;
input [1:0]  sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I39 ( .in(in3), .out(outd23), .pp(sb[0]), .nn(sel[0]));
txgate_lvt I40 ( .in(in2), .out(outd23), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I33 ( .in(outd01), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_lvt I_txgate1 ( .in(in1), .out(outd01), .pp(sb[0]),
     .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(outd01), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(outd23), .out(out), .pp(sb[1]), .nn(sel[1]));

endmodule
// Library - leafcell, Cell - oa4plldly_40lp, View - schematic
// LAST TIME SAVED: Jul 23 17:36:30 2010
// NETLIST TIME: Jun 29 10:32:23 2011
`timescale 1ns / 1ns 

module oa4plldly_40lp ( out, cbit, fda_en, in, prog );
output  out;

input  cbit, fda_en, in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I7 ( .A(net9), .Y(net6), .B(cbit));
anor21_hvt I1 ( .A(net031), .B(fda_en), .Y(out), .C(net6));
inv_hvt I3 ( .A(prog), .Y(net9));
inv_hvt I23 ( .A(in), .Y(net031));

endmodule
