// Library - ice384chip, Cell - nvcm_top_id_u40, View - schematic
// LAST TIME SAVED: Dec 13 15:09:51 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_top_id_u40 ( bp0, fsm_blkadd, fsm_blkadd_b, fsm_coladd,
     fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_redrow,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_recall,
     fsm_rowadd, fsm_sample, fsm_tm_allbank_sel, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_bgr_dis,
     fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_ref,
     fsm_tm_rprd, fsm_tm_tcol, fsm_tm_testdec, fsm_tm_testdec_wr,
     fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvpp, fsm_tm_xvpxa_int, fsm_trim_ipp,
     fsm_trim_multibl_read, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_trim_vbg, fsm_trim_vpgmwl, fsm_trim_vrdwl, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, idcode_msb20bits_out,
     nvcm_boot, nvcm_dis_idchk, nvcm_rdy, nvcm_relextspi, spi_sdo,
     spi_sdo_oe_b, status_wip, trim_spare, clk, idcode_msb20bits_in,
     nv_dataout, nvcm_ce_b, nvcm_max_coladd, nvcm_max_rowadd, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_redrow, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_recall, fsm_sample, fsm_tm_allbank_sel,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_bgr_dis, fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_tcol, fsm_tm_testdec, fsm_tm_testdec_wr,
     fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvpp, fsm_tm_xvpxa_int, fsm_trim_multibl_read, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot,
     nvcm_dis_idchk, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b,
     status_wip;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

output [3:0]  fsm_blkadd_b;
output [3:0]  fsm_trim_ipp;
output [19:0]  idcode_msb20bits_out;
output [8:0]  fsm_rowadd;
output [2:0]  fsm_trim_vpgmwl;
output [3:0]  trim_spare;
output [1:0]  fsm_tm_ref;
output [3:0]  fsm_blkadd;
output [2:0]  fsm_trim_rrefrd;
output [3:0]  fsm_trim_vbg;
output [2:0]  fsm_trim_vrdwl;
output [2:0]  fsm_trim_rrefpgm;
output [11:0]  fsm_coladd;

input [8:0]  nvcm_max_rowadd;
input [19:0]  idcode_msb20bits_in;
input [11:0]  nvcm_max_coladd;
input [8:0]  nv_dataout;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM_40nm, Cell - ml_bgr, View - schematic
// LAST TIME SAVED: Nov 28 11:56:25 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_bgr ( bgr, bgr_bias, sa_bias_25, en_25 );
inout  bgr, bgr_bias, sa_bias_25;

input  en_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



PNP_V45X45_LP  Q1 ( .C(GND_), .B(GND_), .E(in_pnpx1));
PNP_V45X45_LP  Q0 ( .C(GND_), .B(GND_), .E(net423));
RNPPO_LP_pcell2460 R4 ( .B(GND_), .MINUS(sa_bias_25), .PLUS(net0209));
RNPPO_LP_pcell2460 R3_0 ( .B(gnd_), .MINUS(net0278), .PLUS(bgr));
RNPPO_LP_pcell2460 R6_0 ( .B(gnd_), .MINUS(net0234), .PLUS(gnd_));
RNPPO_LP_pcell2460 R1_0 ( .B(gnd_), .MINUS(net0246), .PLUS(bgr));
RNPPO_LP_pcell2460 R10 ( .B(gnd_), .MINUS(gnd_), .PLUS(gnd_));
RNPPO_LP_pcell2460 R32 ( .B(gnd_), .MINUS(gnd_), .PLUS(net0261));
RNPPO_LP_pcell2460 R3_1 ( .B(gnd_), .MINUS(in_pnpx1), .PLUS(net0278));
RNPPO_LP_pcell2460 R1_1 ( .B(gnd_), .MINUS(in_pnpx8), .PLUS(net0246));
RNPPO_LP_pcell2460 R5_1 ( .B(gnd_), .MINUS(gnd_), .PLUS(net0243));
RNPPO_LP_pcell2460 R5_0 ( .B(gnd_), .MINUS(net0243), .PLUS(gnd_));
RNPPO_LP_pcell2460 R8_0 ( .B(gnd_), .MINUS(net0258), .PLUS(gnd_));
RNPPO_LP_pcell2460 R8_1 ( .B(gnd_), .MINUS(gnd_), .PLUS(net0258));
RNPPO_LP_pcell2460 R2 ( .B(gnd_), .MINUS(net423), .PLUS(in_pnpx8));
RNPPO_LP_pcell2460 R11 ( .B(gnd_), .MINUS(gnd_), .PLUS(gnd_));
RNPPO_LP_pcell2460 R0 ( .B(GND_), .MINUS(net0209), .PLUS(net0303));
RNPPO_LP_pcell2460 R7_1 ( .B(gnd_), .MINUS(gnd_), .PLUS(net0267));
RNPPO_LP_pcell2460 R7_0 ( .B(gnd_), .MINUS(net0267), .PLUS(gnd_));
RNPPO_LP_pcell2460 R6_1 ( .B(gnd_), .MINUS(gnd_), .PLUS(net0234));
RNPPO_LP_pcell2460 R35 ( .B(gnd_), .MINUS(net0255), .PLUS(gnd_));
RNPPO_LP_pcell2460 R34 ( .B(gnd_), .MINUS(gnd_), .PLUS(net0255));
RNPPO_LP_pcell2460 R33 ( .B(gnd_), .MINUS(net0261), .PLUS(gnd_));
P_25_LP  M22 ( .D(vddp_), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M62 ( .D(in_pnpx1), .B(vddp_), .G(net0224), .S(net0303));
P_25_LP  M83 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M98 ( .D(net0309), .B(vddp_), .G(net0309), .S(vddp_));
P_25_LP  M71 ( .D(sa_mirr_25), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
P_25_LP  M89 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M99 ( .D(net0323), .B(vddp_), .G(en_b_25), .S(vddp_));
P_25_LP  M74 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M40 ( .D(net0303), .B(vddp_), .G(en_b_25), .S(vddp_));
P_25_LP  M90 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M10 ( .D(sa_mirr_25), .B(vddp_), .G(en_25), .S(vddp_));
P_25_LP  M72 ( .D(net0224), .B(vddp_), .G(bgr_bias), .S(net0303));
P_25_LP  M80 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M73 ( .D(bgr), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M84 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M64 ( .D(bgr_bias), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
P_25_LP  M87 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M25 ( .D(bgr_bias), .B(vddp_), .G(en_25), .S(vddp_));
P_25_LP  M88 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
N_25_LP  M82 ( .D(sa_bias_25), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M58 ( .D(net0224), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M59 ( .D(net0224), .B(gnd_), .G(en_b_25), .S(GND_));
N_25_LP  M85 ( .D(sa_bias_25), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M100 ( .D(GND_), .B(gnd_), .G(tie_low), .S(GND_));
N_25_LP  M96 ( .D(net0224), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M86 ( .D(sa_bias_25), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M91 ( .D(GND_), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M94 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LP  M23 ( .D(bgr), .B(gnd_), .G(en_b_25), .S(GND_));
N_25_LP  M46 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LP  M27 ( .D(sa_bias_25), .B(gnd_), .G(en_b_25), .S(GND_));
N_25_LP  M92 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LP  M81 ( .D(sa_bias_25), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M95 ( .D(net0224), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LP  M97 ( .D(tie_low), .B(gnd_), .G(net0309), .S(GND_));
N_25_LP  M93 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LP  M3 ( .D(net436), .B(gnd_), .G(sa_bias_25), .S(GND_));
N_25_LPNVT  M60 ( .D(bgr_bias), .B(gnd_), .G(in_pnpx1), .S(net436));
N_25_LPNVT  M79 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LPNVT  M76 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LPNVT  M78 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LPNVT  M77 ( .D(gnd_), .B(gnd_), .G(tie_low), .S(gnd_));
N_25_LPNVT  M75 ( .D(sa_mirr_25), .B(gnd_), .G(in_pnpx8), .S(net436));
inv_25 I186 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_top, View - schematic
// LAST TIME SAVED: Sep 24 16:54:12 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_bgr_top ( bgr_int, fsm_bgr_dis_buf, fsm_nvcmen_buf,
     fsm_trim_vbg_buf );
inout  bgr_int;

input  fsm_bgr_dis_buf, fsm_nvcmen_buf;

input [3:0]  fsm_trim_vbg_buf;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net201;

wire  [3:0]  net200;

wire  [1:0]  net0169;

wire  [3:0]  net190;

wire  [3:0]  net192;

wire  [1:0]  net0170;

wire  [15:0]  bgr_dec_b_25;

wire  [3:0]  bgrtrim_b_25;

wire  [15:0]  vref;

wire  [3:0]  bgrtrim_25;



RNPPO_LP_pcell2460 R8 ( .B(gnd_), .MINUS(gnd_), .PLUS(vref[0]));
RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(vref[15]), .PLUS(net0147));
RNPPO_LP_pcell2460 R2 ( .B(gnd_), .MINUS(net0147), .PLUS(net124));
N_25_LPNVT  M8 ( .D(gnd_), .B(gnd_), .G(vref_reg), .S(gnd_));
N_25_LPNVT  M11 ( .D(gnd_), .B(gnd_), .G(bgr_int), .S(gnd_));
N_25_LPNVT  M60 ( .D(net124), .B(gnd_), .G(vref_reg), .S(net0155));
N_25_LPNVT  M0 ( .D(gnd_), .B(gnd_), .G(vref_reg), .S(gnd_));
N_25_LPNVT  M10 ( .D(gnd_), .B(gnd_), .G(vref_reg), .S(gnd_));
P_25_LP  M7_1_ ( .D(net0170[0]), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M7_0_ ( .D(net0170[1]), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M3 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M73 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M6_1_ ( .D(net0169[0]), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M6_0_ ( .D(net0169[1]), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M4 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M2 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M5 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
P_25_LP  M25 ( .D(net113), .B(vddp_), .G(bgr_en_b), .S(vddp_));
vdd_tiehigh I205 ( .vdd_tieh(net0167));
nand2_hvt I323 ( .B(fsm_nvcmen_buf), .A(net0281), .Y(net188));
ml_bgr_buf Iml_bgr_buf ( .sa_bias_25(sa_bias_25), .inp(bgr),
     .inn(vref[8]), .en_25(bgr_en_25), .sa_out(vref_reg));
nand4_25 I135_7_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[7]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_6_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[6]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_5_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[5]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_4_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[4]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_3_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[3]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_2_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[2]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_1_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[1]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_0_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[0]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_15_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[15]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_14_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[14]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_13_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[13]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_12_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[12]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_11_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[11]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_10_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[10]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_9_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[9]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_8_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[8]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
ml_vpp_ref_sw I169 ( .in(bgr_int), .out(net0238), .sel_b_25(bgr_en_b));
ml_vpp_ref_sw I170 ( .in(bgr_int), .out(vref_vdd),
     .sel_b_25(bgr_en_25));
ml_vpp_ref_sw ref_sw_7_ ( .in(net0238), .out(vref[7]),
     .sel_b_25(bgr_dec_b_25[7]));
ml_vpp_ref_sw ref_sw_6_ ( .in(net0238), .out(vref[6]),
     .sel_b_25(bgr_dec_b_25[6]));
ml_vpp_ref_sw ref_sw_5_ ( .in(net0238), .out(vref[5]),
     .sel_b_25(bgr_dec_b_25[5]));
ml_vpp_ref_sw ref_sw_4_ ( .in(net0238), .out(vref[4]),
     .sel_b_25(bgr_dec_b_25[4]));
ml_vpp_ref_sw ref_sw_3_ ( .in(net0238), .out(vref[3]),
     .sel_b_25(bgr_dec_b_25[3]));
ml_vpp_ref_sw ref_sw_2_ ( .in(net0238), .out(vref[2]),
     .sel_b_25(bgr_dec_b_25[2]));
ml_vpp_ref_sw ref_sw_1_ ( .in(net0238), .out(vref[1]),
     .sel_b_25(bgr_dec_b_25[1]));
ml_vpp_ref_sw ref_sw_0_ ( .in(net0238), .out(vref[0]),
     .sel_b_25(bgr_dec_b_25[0]));
ml_vpp_ref_sw ref_sw_15_ ( .in(net0238), .out(vref[15]),
     .sel_b_25(bgr_dec_b_25[15]));
ml_vpp_ref_sw ref_sw_14_ ( .in(net0238), .out(vref[14]),
     .sel_b_25(bgr_dec_b_25[14]));
ml_vpp_ref_sw ref_sw_13_ ( .in(net0238), .out(vref[13]),
     .sel_b_25(bgr_dec_b_25[13]));
ml_vpp_ref_sw ref_sw_12_ ( .in(net0238), .out(vref[12]),
     .sel_b_25(bgr_dec_b_25[12]));
ml_vpp_ref_sw ref_sw_11_ ( .in(net0238), .out(vref[11]),
     .sel_b_25(bgr_dec_b_25[11]));
ml_vpp_ref_sw ref_sw_10_ ( .in(net0238), .out(vref[10]),
     .sel_b_25(bgr_dec_b_25[10]));
ml_vpp_ref_sw ref_sw_9_ ( .in(net0238), .out(vref[9]),
     .sel_b_25(bgr_dec_b_25[9]));
ml_vpp_ref_sw ref_sw_8_ ( .in(net0238), .out(vref[8]),
     .sel_b_25(bgr_dec_b_25[8]));
ml_bgr_res_100_ohm I90 ( .t(vref[8]), .b(vref[7]));
ml_bgr_res_100_ohm I91 ( .t(vref[7]), .b(vref[6]));
ml_bgr_res_100_ohm I92 ( .t(vref[6]), .b(vref[5]));
ml_bgr_res_100_ohm I93 ( .t(vref[4]), .b(vref[3]));
ml_bgr_res_100_ohm I94 ( .t(vref[5]), .b(vref[4]));
ml_bgr_res_100_ohm I95 ( .t(vref[1]), .b(vref[0]));
ml_bgr_res_100_ohm I97 ( .t(vref[2]), .b(vref[1]));
ml_bgr_res_100_ohm I100 ( .t(vref[3]), .b(vref[2]));
ml_bgr_res_100_ohm I101 ( .t(vref[13]), .b(vref[14]));
ml_bgr_res_100_ohm I102 ( .t(vref[14]), .b(vref[15]));
ml_bgr_res_100_ohm I104 ( .t(vref[11]), .b(vref[12]));
ml_bgr_res_100_ohm I105 ( .t(vref[12]), .b(vref[13]));
ml_bgr_res_100_ohm I106 ( .t(vref[10]), .b(vref[11]));
ml_bgr_res_100_ohm I107 ( .t(vref[9]), .b(vref[10]));
ml_bgr_res_100_ohm I108 ( .t(vref[8]), .b(vref[9]));
ml_bgr Iml_bgr ( .bgr_bias(bgr_bias), .sa_bias_25(sa_bias_25),
     .en_25(bgr_en_25), .bgr(bgr));
inv_25 I186 ( .IN(net195), .OUT(bgr_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I139 ( .IN(net196), .OUT(bgr_en_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I198_3_ ( .IN(net201[0]), .OUT(bgrtrim_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_2_ ( .IN(net201[1]), .OUT(bgrtrim_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_1_ ( .IN(net201[2]), .OUT(bgrtrim_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_0_ ( .IN(net201[3]), .OUT(bgrtrim_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_3_ ( .IN(net200[0]), .OUT(bgrtrim_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_2_ ( .IN(net200[1]), .OUT(bgrtrim_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_1_ ( .IN(net200[2]), .OUT(bgrtrim_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_0_ ( .IN(net200[3]), .OUT(bgrtrim_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I192 ( .IN(net0313), .OUT(bgr2vdd_25_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I189 ( .IN(net0312), .OUT(bgr2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I88_3_ ( .A(fsm_trim_vbg_buf[3]), .Y(net190[0]));
inv_hvt I88_2_ ( .A(fsm_trim_vbg_buf[2]), .Y(net190[1]));
inv_hvt I88_1_ ( .A(fsm_trim_vbg_buf[1]), .Y(net190[2]));
inv_hvt I88_0_ ( .A(fsm_trim_vbg_buf[0]), .Y(net190[3]));
inv_hvt I167 ( .A(net188), .Y(net186));
inv_hvt I183 ( .A(net0167), .Y(net0326));
inv_hvt I168 ( .A(fsm_bgr_dis_buf), .Y(net0281));
inv_hvt I174 ( .A(net0326), .Y(vref_vdd));
inv_hvt I87_3_ ( .A(net190[0]), .Y(net192[0]));
inv_hvt I87_2_ ( .A(net190[1]), .Y(net192[1]));
inv_hvt I87_1_ ( .A(net190[2]), .Y(net192[2]));
inv_hvt I87_0_ ( .A(net190[3]), .Y(net192[3]));
ml_ls_vdd2vdd25 I80_3_ ( .in(net192[0]), .sup(vddp_),
     .out_vddio_b(net200[0]), .out_vddio(net201[0]), .in_b(net190[0]));
ml_ls_vdd2vdd25 I80_2_ ( .in(net192[1]), .sup(vddp_),
     .out_vddio_b(net200[1]), .out_vddio(net201[1]), .in_b(net190[1]));
ml_ls_vdd2vdd25 I80_1_ ( .in(net192[2]), .sup(vddp_),
     .out_vddio_b(net200[2]), .out_vddio(net201[2]), .in_b(net190[2]));
ml_ls_vdd2vdd25 I80_0_ ( .in(net192[3]), .sup(vddp_),
     .out_vddio_b(net200[3]), .out_vddio(net201[3]), .in_b(net190[3]));
ml_ls_vdd2vdd25 I177 ( .in(vref_vdd), .sup(vddp_),
     .out_vddio_b(net0312), .out_vddio(net0313), .in_b(net0326));
ml_ls_vdd2vdd25 I335 ( .in(net186), .sup(vddp_), .out_vddio_b(net195),
     .out_vddio(net196), .in_b(net188));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_buf, View - schematic
// LAST TIME SAVED: Aug  3 19:29:08 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_pump_vpxa_buf ( out, in );
output  out;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_25 I38 ( .IN(in), .OUT(net15), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
inv_25 I195 ( .IN(net15), .OUT(out), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_pump, View - schematic
// LAST TIME SAVED: Aug  3 19:29:12 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpp_pump ( pump_in, clkin_25, en_25 );
inout  pump_in;

input  clkin_25, en_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(net23), .B(vddp_), .G(net64), .S(vddp_));
N_25_LPNVT  M2 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
N_25_LPNVT  M3 ( .D(s_2), .B(GND_), .G(s_2), .S(s_3));
N_25_LPNVT  M22 ( .D(net23), .B(GND_), .G(net23), .S(s_0));
N_25_LPNVT  M4 ( .D(s_3), .B(GND_), .G(s_3), .S(pump_in));
N_25_LPNVT  M1 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
NCAP_25_LP  C0 ( .MINUS(clk_25), .PLUS(s_0));
NCAP_25_LP  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
NCAP_25_LP  C7 ( .MINUS(clk_25), .PLUS(s_2));
NCAP_25_LP  C1 ( .MINUS(clk_b_25), .PLUS(s_3));
inv_25 I230 ( .IN(clkin_25), .OUT(net0124), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I232 ( .IN(net088), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I233 ( .IN(net0100), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I234 ( .IN(net094), .OUT(net0106), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I235 ( .IN(net0106), .OUT(net0100), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I236 ( .IN(clkin_25), .OUT(net094), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I237 ( .IN(net0124), .OUT(net088), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I231 ( .IN(en_25), .OUT(net64), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd2vdd25_vpxa, View - schematic
// LAST TIME SAVED: Aug  3 19:29:06 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25_vpxa ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M1 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
P_25_LP  M2 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
P_25_LP  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));
P_25_LP  M0 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
N_25_LP  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
N_25_LP  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_hv2vddp_sw, View - schematic
// LAST TIME SAVED: Aug  3 19:29:03 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv2vddp_sw ( out_hv, hv2vddp, vddp_tieh, vpxa );
inout  out_hv;

input  hv2vddp, vddp_tieh, vpxa;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(net27), .B(vddp_), .G(sw_vddp_b), .S(vddp_));
P_25_LP  M1 ( .D(net27), .B(out_hv), .G(sw_vpp_b), .S(out_hv));
ml_ls_vdd2vdd25_vpxa I64 ( .in(net44), .sup(vddp_),
     .out_vddio_b(net060), .out_vddio(net37), .in_b(net46));
inv_25 I62 ( .IN(net37), .OUT(sw_vddp_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I71 ( .IN(net060), .OUT(net035), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I65 ( .A(hv2vddp), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(sw_vddp_b),
     .sel_25(net035), .out_b_hv(sw_vpp_b), .in_hv(out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ref, View - schematic
// LAST TIME SAVED: Nov  7 17:01:20 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpp_ref ( vref_25, bgr, pumpen_25, vppwl_25 );
inout  vref_25;

input  bgr, pumpen_25;

input [2:0]  vppwl_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_b_25;

wire  [7:0]  red_dec_25;



P_25_LP  M18 ( .D(net179), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
P_25_LP  M5 ( .D(ctrl_gate_25), .B(vddp_), .G(net0113), .S(net175));
P_25_LP  M6 ( .D(net0113), .B(vddp_), .G(net0113), .S(net175));
P_25_LP  M7 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
P_25_LP  M1 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(net175));
RNPPO_LP_pcell2460 R12 ( .B(GND_), .MINUS(net110), .PLUS(net113));
RNPPO_LP_pcell2460 R15 ( .B(GND_), .MINUS(net104), .PLUS(net0216));
RNPPO_LP_pcell2460 R18 ( .B(GND_), .MINUS(net0216), .PLUS(net139));
RNPPO_LP_pcell2460 R19 ( .B(GND_), .MINUS(net139), .PLUS(net0213));
RNPPO_LP_pcell2460 R22 ( .B(GND_), .MINUS(net0213), .PLUS(net98));
RNPPO_LP_pcell2460 R25 ( .B(GND_), .MINUS(net98),
     .PLUS(bgr_mirror_25));
RNPPO_LP_pcell2460 R24 ( .B(GND_), .MINUS(net98),
     .PLUS(bgr_mirror_25));
RNPPO_LP_pcell2460 R8 ( .B(GND_), .MINUS(gnd_), .PLUS(net0100));
RNPPO_LP_pcell2460 R14 ( .B(GND_), .MINUS(net113), .PLUS(net104));
RNPPO_LP_pcell2460 R1 ( .B(GND_), .MINUS(net0100), .PLUS(net0100));
RNPPO_LP_pcell2460 R2 ( .B(GND_), .MINUS(net0100), .PLUS(net0193));
RNPPO_LP_pcell2460 R10 ( .B(GND_), .MINUS(net0193), .PLUS(net110));
RNPPO_LP_pcell2460 R26 ( .B(GND_), .MINUS(bgr_mirror_25),
     .PLUS(net0129));
NCAP_25_LP  C2 ( .MINUS(gnd_), .PLUS(ctrl_gate_25));
NCAP_25_LP  C3 ( .MINUS(net0129), .PLUS(net0113));
N_25_LPNVT  M0 ( .D(net179), .B(GND_), .G(ctrl_gate_25),
     .S(bgr_mirror_25));
N_25_LP  M10 ( .D(net163), .B(GND_), .G(bgr), .S(gnd_));
N_25_LP  M14 ( .D(net0113), .B(GND_), .G(vppref_en_b_25), .S(gnd_));
N_25_LP  M15 ( .D(ctrl_gate_25), .B(GND_), .G(vppref_en_b_25),
     .S(gnd_));
N_25_LP  M8 ( .D(ctrl_gate_25), .B(GND_), .G(bgr_mirror_25),
     .S(net163));
N_25_LP  M13 ( .D(net0113), .B(GND_), .G(bgr), .S(net163));
nand3_25 I44_7_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[7]),
     .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_6_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[6]),
     .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_5_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[5]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_4_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[4]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_3_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[3]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_2_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[2]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_1_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[1]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_0_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[0]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
inv_25 I38 ( .IN(pumpen_25), .OUT(vppref_en_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_2_ ( .IN(vppwl_25[2]), .OUT(vppwl_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_1_ ( .IN(vppwl_25[1]), .OUT(vppwl_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_0_ ( .IN(vppwl_25[0]), .OUT(vppwl_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_vpp_ref_sw I281 ( .in(net0213), .out(vref_25),
     .sel_b_25(red_dec_25[6]));
ml_vpp_ref_sw I287 ( .in(net0216), .out(vref_25),
     .sel_b_25(red_dec_25[4]));
ml_vpp_ref_sw I283 ( .in(net98), .out(vref_25),
     .sel_b_25(red_dec_25[7]));
ml_vpp_ref_sw I290 ( .in(net0193), .out(vref_25),
     .sel_b_25(red_dec_25[0]));
ml_vpp_ref_sw I288 ( .in(net104), .out(vref_25),
     .sel_b_25(red_dec_25[3]));
ml_vpp_ref_sw I284 ( .in(net139), .out(vref_25),
     .sel_b_25(red_dec_25[5]));
ml_vpp_ref_sw I291 ( .in(net110), .out(vref_25),
     .sel_b_25(red_dec_25[1]));
ml_vpp_ref_sw I292 ( .in(net113), .out(vref_25),
     .sel_b_25(red_dec_25[2]));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ctrl, View - schematic
// LAST TIME SAVED: Aug  3 19:29:12 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpp_ctrl ( pumpen_25, vpint_en, vpp_2_vdd, vppdisc_vpxa,
     vppwl_25, vpxa, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_vpgmwl_buf, fsm_wgnden );
output  pumpen_25, vpint_en, vpp_2_vdd, vppdisc_vpxa;

inout  vpxa;

input  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint, fsm_wgnden;

output [2:0]  vppwl_25;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  net082;

wire  [2:0]  net068;

wire  [2:0]  net038;

wire  [2:0]  net092;



NCAP_25_LP  C7 ( .MINUS(GND_), .PLUS(net0122));
ml_ls_vdd2vdd25_vpxa I173 ( .in(fsm_pgmdisc_buf), .sup(vpxa),
     .out_vddio_b(net088), .out_vddio(net048), .in_b(net0106));
ml_dff_nvcm I77 ( .CLK(net084), .QN(vpp_pumpen_b), .R(pgm_dis),
     .D(vdd_tieh), .Q(vpp_pumpen));
inv_25 I95_2_ ( .IN(net068[0]), .OUT(vppwl_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_1_ ( .IN(net068[1]), .OUT(vppwl_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_0_ ( .IN(net068[2]), .OUT(vppwl_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I81 ( .IN(net073), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(net088), .OUT(vppdisc_vpxa), .P(vpxa), .Pb(vpxa),
     .G(gnd_), .Gb(gnd_));
nand3_hvt I79 ( .C(net086), .A(fsm_pgm_buf), .Y(pgm_dis),
     .B(fsm_nvcmen_buf));
nor2_hvt I111 ( .A(vpp_pumpen_b), .B(net080), .Y(net0133));
nor2_hvt I87 ( .A(vpp_pumpen), .Y(net036), .B(fsm_pgmdisc_buf));
nand4_hvt I75 ( .D(fsm_pgm_buf), .C(fsm_lshven_buf), .A(net0127),
     .Y(net046), .B(net0127));
inv_hvt I107 ( .A(net0122), .Y(net0124));
inv_hvt I109 ( .A(fsm_pgmvfy_buf), .Y(net0127));
inv_hvt I131 ( .A(net049), .Y(net080));
inv_hvt I110_2_ ( .A(net092[0]), .Y(net082[0]));
inv_hvt I110_1_ ( .A(net092[1]), .Y(net082[1]));
inv_hvt I110_0_ ( .A(net092[2]), .Y(net082[2]));
inv_hvt I76 ( .A(net046), .Y(net084));
inv_hvt I108 ( .A(fsm_pgmdisc_buf), .Y(net0122));
inv_hvt I78 ( .A(net0124), .Y(net086));
inv_hvt I113 ( .A(vpp_pumpen_b), .Y(vpint_en));
inv_hvt I91 ( .A(net036), .Y(net089));
inv_hvt I90 ( .A(net089), .Y(vpp_2_vdd));
inv_hvt I98_2_ ( .A(fsm_vpgmwl_buf[2]), .Y(net092[0]));
inv_hvt I98_1_ ( .A(fsm_vpgmwl_buf[1]), .Y(net092[1]));
inv_hvt I98_0_ ( .A(fsm_vpgmwl_buf[0]), .Y(net092[2]));
inv_hvt I112 ( .A(net0133), .Y(net0134));
inv_hvt I101 ( .A(fsm_pgmdisc_buf), .Y(net0106));
nand2_hvt I104 ( .A(fsm_tm_xforce), .Y(net049), .B(fsm_tm_xvppint));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_ls_vdd2vdd25 I96_2_ ( .in(net082[0]), .sup(vddp_),
     .out_vddio_b(net068[0]), .out_vddio(net038[0]), .in_b(net092[0]));
ml_ls_vdd2vdd25 I96_1_ ( .in(net082[1]), .sup(vddp_),
     .out_vddio_b(net068[1]), .out_vddio(net038[1]), .in_b(net092[1]));
ml_ls_vdd2vdd25 I96_0_ ( .in(net082[2]), .sup(vddp_),
     .out_vddio_b(net068[2]), .out_vddio(net038[2]), .in_b(net092[2]));
ml_ls_vdd2vdd25 I84 ( .in(net0133), .sup(vddp_), .out_vddio_b(net073),
     .out_vddio(net074), .in_b(net0134));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_reg, View - schematic
// LAST TIME SAVED: Nov  9 16:50:46 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpp_reg ( slow_25, bgr, pbias_25, pump_in, vpp_int, vpxa,
     pumpen_25, vppdisc_vpxa, vref_25 );
output  slow_25;

inout  bgr, pbias_25, pump_in, vpp_int, vpxa;

input  pumpen_25, vppdisc_vpxa, vref_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LPNVT  M22 ( .D(vpp_int), .B(GND_), .G(pump_gate), .S(pump_in));
N_25_LPNVT  M1 ( .D(GND_), .B(GND_), .G(pump_gate), .S(GND_));
N_25_LPNVT  M10 ( .D(net0203), .B(GND_), .G(net0208), .S(net0199));
N_25_LPNVT  M5 ( .D(pump_opamp_out), .B(GND_), .G(vpp_int),
     .S(pump_opamp_out));
N_25_LPNVT  M11 ( .D(net0199), .B(GND_), .G(vppdisc_vpxa),
     .S(net0271));
N_25_LP  M16 ( .D(net124), .B(GND_), .G(net124), .S(net155));
N_25_LP  M17 ( .D(net155), .B(GND_), .G(en_buf_25), .S(gnd_));
N_25_LP  M6 ( .D(vpp_int), .B(GND_), .G(en_buf_25), .S(net168));
N_25_LP  M3 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
N_25_LP  M20 ( .D(slow_25), .B(GND_), .G(pump_opamp_out), .S(gnd_));
N_25_LP  M7 ( .D(net168), .B(GND_), .G(pump_opamp_out), .S(gnd_));
N_25_LP  M4 ( .D(dis_pgate_25), .B(GND_), .G(net0208), .S(net0264));
N_25_LP  M41 ( .D(net0224), .B(GND_), .G(en_buf_25), .S(gnd_));
N_25_LP  M15 ( .D(pump_opamp_out), .B(GND_), .G(net124), .S(net155));
N_25_LP  M0 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net0175));
N_25_LP  M40 ( .D(net0264), .B(GND_), .G(vppdisc_vpxa), .S(gnd_));
P_25_LP  M2 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
P_25_LP  M9 ( .D(net0200), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
P_25_LP  M8_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
P_25_LP  M8_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
P_25_LP  M14 ( .D(pump_opamp_out), .B(net125), .G(vref_25),
     .S(net125));
P_25_LP  M18 ( .D(net122), .B(vpp_int), .G(net122), .S(vpp_int));
P_25_LP  M13 ( .D(net124), .B(net125), .G(vdiv), .S(net125));
P_25_LP  M32 ( .D(dis_pgate_25), .B(vpxa), .G(dis_pgate_25), .S(vpxa));
P_25_LP  M33 ( .D(dis_pgate_25), .B(vpxa), .G(vppdisc_vpxa), .S(vpxa));
P_25_LP  M12 ( .D(net125), .B(vddp_), .G(pbias_25), .S(vddp_));
P_25_LP  M19 ( .D(net134), .B(net122), .G(net134), .S(net122));
P_25_LP  M21 ( .D(net138), .B(net134), .G(net138), .S(net134));
P_25_LP  M23 ( .D(net142), .B(net138), .G(net142), .S(net138));
P_25_LP  M24 ( .D(vdiv), .B(net142), .G(vdiv), .S(net142));
P_25_LP  M25 ( .D(net0224), .B(vdiv), .G(net0224), .S(vdiv));
P_25_LP  M31 ( .D(net0203), .B(net0165), .G(dis_pgate_25),
     .S(net0165));
RNPPO_LP_pcell2460 R5 ( .B(GND_), .MINUS(net0165), .PLUS(vpp_int));
RNPPO_LP_pcell2460 R6 ( .B(GND_), .MINUS(gnd_), .PLUS(net0178));
RNPPO_LP_pcell2460 R14 ( .B(GND_), .MINUS(net0271), .PLUS(vdd_));
RNPPO_LP_pcell2460 R8 ( .B(GND_), .MINUS(gnd_), .PLUS(gnd_));
RNPPO_LP_pcell2460 R15 ( .B(GND_), .MINUS(net0271), .PLUS(vdd_));
RNPPO_LP_pcell2460 R16 ( .B(GND_), .MINUS(net0271), .PLUS(vdd_));
RNPPO_LP_pcell2460 R11 ( .B(GND_), .MINUS(vdd_), .PLUS(net0271));
RNPPO_LP_pcell2460 R12 ( .B(GND_), .MINUS(vdd_), .PLUS(net0271));
RNPPO_LP_pcell2460 R3 ( .B(GND_), .MINUS(pump_gate), .PLUS(pump_in));
RNPPO_LP_pcell2460 R7 ( .B(GND_), .MINUS(net0178), .PLUS(net0175));
RNPPO_LP_pcell2460 R13 ( .B(GND_), .MINUS(vdd_), .PLUS(net0271));
inv_25 I211 ( .IN(en_buf_b_25), .OUT(en_buf_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I212 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
vddp_tiehigh I261 ( .vddp_tieh(net0208));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_vco, View - schematic
// LAST TIME SAVED: Aug  3 19:29:13 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpp_vco ( clk_25_0, clk_25_1, pbias_25, slow_25, en_25,
     freq_25 );
output  clk_25_0, clk_25_1;

inout  pbias_25, slow_25;

input  en_25;

input [1:0]  freq_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:1]  freq_b_25;



P_25_LP  M10 ( .D(net236), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
P_25_LP  M9 ( .D(net248), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
P_25_LP  M3 ( .D(net189), .B(vddp_), .G(net173), .S(net248));
P_25_LP  M11 ( .D(net256), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
P_25_LP  M12 ( .D(net185), .B(vddp_), .G(net193), .S(net256));
P_25_LP  M19 ( .D(net193), .B(vddp_), .G(net195), .S(net260));
P_25_LP  M20 ( .D(net260), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
P_25_LP  M22 ( .D(pbias_osc_25), .B(vddp_), .G(en_b_25), .S(net228));
P_25_LP  M26_1_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25),
     .S(vddp_));
P_25_LP  M26_0_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25),
     .S(vddp_));
P_25_LP  M7 ( .D(net173), .B(vddp_), .G(net185), .S(net236));
P_25_LP  M27_1_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
P_25_LP  M27_0_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
P_25_LP  M28 ( .D(net212), .B(vddp_), .G(pbias_25), .S(vddp_));
P_25_LP  M29 ( .D(nbias_osc_25), .B(vddp_), .G(freq_25[0]),
     .S(net212));
P_25_LP  M30 ( .D(nbias_osc_25), .B(vddp_), .G(freq_b_25[1]),
     .S(net208));
P_25_LP  M21 ( .D(net228), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
N_25_LP  M6 ( .D(net177), .B(GND_), .G(nbias_osc_25), .S(GND_));
N_25_LP  M13 ( .D(net181), .B(GND_), .G(nbias_osc_25), .S(GND_));
N_25_LP  M14 ( .D(net185), .B(GND_), .G(net193), .S(net181));
N_25_LP  M8 ( .D(net189), .B(GND_), .G(net173), .S(net201));
N_25_LP  M17 ( .D(net193), .B(GND_), .G(net195), .S(net197));
N_25_LP  M18 ( .D(net197), .B(GND_), .G(nbias_osc_25), .S(GND_));
N_25_LP  M1 ( .D(net201), .B(GND_), .G(nbias_osc_25), .S(GND_));
N_25_LP  M23 ( .D(pbias_osc_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
N_25_LP  M5 ( .D(net173), .B(GND_), .G(net185), .S(net177));
N_25_LP  M24 ( .D(slow_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
N_25_LP  M25 ( .D(nbias_osc_25), .B(GND_), .G(en_25), .S(slow_25));
N_25_LPNVT  M15 ( .D(GND_), .B(GND_), .G(net185), .S(GND_));
N_25_LPNVT  M4 ( .D(GND_), .B(GND_), .G(net173), .S(GND_));
N_25_LPNVT  M16 ( .D(GND_), .B(GND_), .G(net193), .S(GND_));
N_25_LPNVT  M2 ( .D(GND_), .B(GND_), .G(net189), .S(GND_));
nand2_25 I96 ( .G(GND_), .Pb(vddp_), .A(net189), .Y(net195), .P(vddp_),
     .B(en_25), .Gb(GND_));
nand2_25 I205 ( .G(GND_), .Pb(vddp_), .A(net185), .Y(net0205),
     .P(vddp_), .B(en_25), .Gb(GND_));
inv_25 I201 ( .IN(net195), .OUT(clk_25_0), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(net0205), .OUT(clk_25_1), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I188 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I199 ( .IN(freq_25[1]), .OUT(freq_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));

endmodule
// Library - sbtlibn65lp, Cell - nor2_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:55 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nor2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(Y), .B(Pb), .G(B), .S(net15));
P_25_LP  M1 ( .D(net15), .B(Pb), .G(A), .S(P));
N_25_LP  M3 ( .D(Y), .B(Gb), .G(A), .S(G));
N_25_LP  M2 ( .D(Y), .B(Gb), .G(B), .S(G));

endmodule
// Library - NVCM_40nm, Cell - ml_vppint_top, View - schematic
// LAST TIME SAVED: Dec 15 15:09:50 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vppint_top ( vpint_en, vpp_int, vpxa, bgr, fsm_lshven_buf,
     fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf, fsm_pgmvfy_buf,
     fsm_tm_xforce, fsm_tm_xvppint, fsm_vpgmwl_buf, fsm_wgnden_buf );
output  vpint_en;

inout  vpp_int, vpxa;

input  bgr, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_wgnden_buf;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_25;

wire  [1:0]  freq_25;



ml_pump_vpxa_buf I95 ( .in(clkin_0_25), .out(net52));
ml_pump_vpxa_buf I81 ( .in(clkin_1_25), .out(net061));
ml_vpp_pump Ivpp_pump_0 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(clkin_1_25));
ml_vpp_pump Ivpp_pump_1 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net061));
ml_vpp_pump Ivpp_pump_2 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net52));
inv_25 I38 ( .IN(vddp_tieh), .OUT(freq_25[1]), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I91 ( .IN(vddp_tieh), .OUT(freq_25[0]), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_hv2vddp_sw Ivpxa_2vddp_sw ( .vpxa(vpxa), .hv2vddp(vpp_2_vdd),
     .vddp_tieh(vddp_tieh), .out_hv(vpp_int));
ml_vpp_ref Ivpp_ref ( .vref_25(vref_25), .vppwl_25(vppwl_25[2:0]),
     .pumpen_25(pumpen_25), .bgr(bgr));
ml_vpp_ctrl Ivpp_ctrl ( .vppdisc_vpxa(vppdisc_vpxa), .vpxa(vpxa),
     .vpint_en(vpint_en), .fsm_pgmvfy_buf(fsm_pgmvfy_buf),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .fsm_wgnden(fsm_wgnden_buf),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf), .vppwl_25(vppwl_25[2:0]),
     .vpp_2_vdd(vpp_2_vdd), .pumpen_25(pumpen_25));
ml_vpp_reg Ivpp_reg ( .vpxa(vpxa), .vppdisc_vpxa(vppdisc_vpxa),
     .bgr(bgr), .slow_25(slow_25), .pbias_25(pbias_25),
     .vref_25(vref_25), .pumpen_25(pumpen_25), .pump_in(pump_in),
     .vpp_int(vpp_int));
ml_vpp_vco Ivpp_vco ( .clk_25_1(clkin_1_25), .pbias_25(pbias_25),
     .slow_25(slow_25), .freq_25(freq_25[1:0]), .en_25(pumpen_25),
     .clk_25_0(clkin_0_25));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_3.3v, View - schematic
// LAST TIME SAVED: Aug  3 19:29:08 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_pump_vpxa_3_3v ( out, clkin_25, en_25 );
inout  out;

input  clkin_25, en_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M6 ( .D(net73), .B(vddp_), .G(net114), .S(vddp_));
N_25_LPNVT  M1 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
N_25_LPNVT  M2 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
N_25_LPNVT  M3 ( .D(s_2), .B(GND_), .G(s_2), .S(out));
N_25_LPNVT  M4 ( .D(net73), .B(GND_), .G(net73), .S(s_0));
NCAP_25_LP  C1 ( .MINUS(clk_25), .PLUS(s_0));
NCAP_25_LP  C2 ( .MINUS(clk_b_25), .PLUS(s_1));
NCAP_25_LP  C3 ( .MINUS(clk_25), .PLUS(s_2));
inv_25 I230 ( .IN(clkin_25), .OUT(net120), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I231 ( .IN(en_25), .OUT(net114), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I232 ( .IN(net78), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I233 ( .IN(net90), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I234 ( .IN(net84), .OUT(net96), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I235 ( .IN(net96), .OUT(net90), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I236 ( .IN(clkin_25), .OUT(net84), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I237 ( .IN(net120), .OUT(net78), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));

endmodule
// Library - sbtlibn65lp, Cell - ml_dlatch_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:55 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_dlatch_25 ( Q_25, D_25, EN_25, R_25 );
output  Q_25;

input  D_25, EN_25, R_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M8 ( .D(net31), .B(vddp_), .G(EN_25), .S(vddp_));
P_25_LP  M7 ( .D(net39), .B(vddp_), .G(EN_B_25), .S(vddp_));
P_25_LP  M3 ( .D(net52), .B(vddp_), .G(D_25), .S(net39));
P_25_LP  M2 ( .D(net52), .B(vddp_), .G(Q_25), .S(net31));
N_25_LP  M0 ( .D(net52), .B(GND_), .G(D_25), .S(net48));
N_25_LP  M1 ( .D(net48), .B(GND_), .G(EN_25), .S(GND_));
N_25_LP  M5 ( .D(net40), .B(GND_), .G(EN_B_25), .S(GND_));
N_25_LP  M6 ( .D(net52), .B(GND_), .G(Q_25), .S(net40));
nor2_25 I161 ( .A(net52), .Y(Q_25), .Gb(GND_), .G(GND_), .Pb(vddp_),
     .P(vddp_), .B(R_25));
inv_25 I156 ( .IN(EN_25), .OUT(EN_B_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_clk_reg, View - schematic
// LAST TIME SAVED: Aug  3 19:29:07 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_pump_clk_reg ( clk_out_25, clk_in_25, pump_chrg_25,
     pump_on_25 );
output  clk_out_25;

input  clk_in_25, pump_chrg_25, pump_on_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nand2_25 I78 ( .G(GND_), .Pb(vddp_), .A(pump_chrg_25), .Y(clk_freeze),
     .P(vddp_), .B(pump_on_25), .Gb(GND_));
inv_25 I72 ( .IN(net020), .OUT(clk_equal), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(vddp_tieh), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
exor2_25 I85 ( .A(clk_in_25), .Y(net020), .B(clk_out_25));
vddp_tiehigh I117 ( .vddp_tieh(vddp_tieh));
ml_dlatch_25 I63 ( .D_25(clk_in_25), .EN_25(clk_go), .R_25(net34),
     .Q_25(clk_out_25));
ml_dlatch_25 I64 ( .D_25(vddp_tieh), .EN_25(clk_equal),
     .R_25(clk_freeze), .Q_25(clk_go));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_x2, View - schematic
// LAST TIME SAVED: Aug  3 19:29:08 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_pump_vpxa_x2 ( vpxa_int, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, pumpen_25, vpxa_clk_25, vpxa_clk_b_25 );
inout  vpxa_int;

input  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25, pumpen_25,
     vpxa_clk_25, vpxa_clk_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_pump_vpxa_buf I80 ( .in(net43), .out(clkin_2_25));
ml_pump_vpxa_buf I79 ( .in(net47), .out(net22));
ml_pump_vpxa_buf I78 ( .in(net39), .out(clkin_0_25));
ml_pump_vpxa_buf I81 ( .in(net22), .out(clkin_1_25));
ml_pump_vpxa_3_3v Ivpxa_pump_0 ( .en_25(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_0_25));
ml_pump_vpxa_3_3v Ivpxa_pump_2 ( .en_25(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_2_25));
ml_pump_vpxa_3_3v Ivpxa_pump_1 ( .en_25(pumpen_25),
     .clkin_25(clkin_1_25), .out(vpxa_int));
ml_pump_clk_reg Iclk_reg_0 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_0_25), .pump_on_25(pumpen_25),
     .clk_out_25(net39));
ml_pump_clk_reg Iclk_reg_2 ( .clk_in_25(vpxa_clk_b_25),
     .pump_chrg_25(pump_chrg_2_25), .pump_on_25(pumpen_25),
     .clk_out_25(net43));
ml_pump_clk_reg Iclk_reg_1 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_1_25), .pump_on_25(pumpen_25),
     .clk_out_25(net47));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_osc, View - schematic
// LAST TIME SAVED: Sep 24 15:31:05 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpxa_osc ( vpxa_clk_25, bgr, freq_25, pumpen_25 );
output  vpxa_clk_25;

inout  bgr;

input  pumpen_25;

input [1:0]  freq_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  freq_buf_b_25;



N_25_LP  M11 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net044));
N_25_LP  M12 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
P_25_LP  M9 ( .D(net061), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
P_25_LP  M10 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
P_25_LP  M8_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
P_25_LP  M8_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
RNPPO_LP_pcell2460 R6 ( .B(GND_), .MINUS(gnd_), .PLUS(net043));
RNPPO_LP_pcell2460 R7 ( .B(GND_), .MINUS(net043), .PLUS(net044));
RNPPO_LP_pcell2460 R8 ( .B(GND_), .MINUS(gnd_), .PLUS(gnd_));
inv_25 I227 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I226 ( .IN(freq_25[0]), .OUT(freq_buf_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_vpp_vco Ivpx_vpp_vco ( .clk_25_1(net040), .pbias_25(pbias_25),
     .slow_25(net86), .freq_25({freq_25[1], freq_buf_b_25[0]}),
     .en_25(pumpen_25), .clk_25_0(vpxa_clk_25));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_ctrl, View - schematic
// LAST TIME SAVED: Aug  3 19:29:13 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpxa_ctrl ( pumpen, pumpen_25, vpxa_2_vdd, fsm_pumpen,
     fsm_tm_xforce, fsm_tm_xvpxaint );
output  pumpen, pumpen_25, vpxa_2_vdd;

input  fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I103 ( .A(vpxa_2_vdd), .B(net065), .Y(pumpen));
nand2_hvt I73 ( .A(fsm_tm_xvpxaint), .B(fsm_tm_xforce), .Y(net042));
inv_hvt I78 ( .A(pumpen), .Y(net075));
inv_hvt I77 ( .A(net042), .Y(net065));
inv_hvt I131 ( .A(fsm_pumpen), .Y(vpxa_2_vdd));
inv_25 I38 ( .IN(net045), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I173 ( .in(pumpen), .sup(vddp_), .out_vddio_b(net045),
     .out_vddio(net046), .in_b(net075));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:55 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_dff_25 ( Q_25, Q_B_25, CLK_25, D_25, R_25 );
output  Q_25, Q_B_25;

input  CLK_25, D_25, R_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_25 I96 ( .IN(Q_25), .OUT(Q_B_25), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I72 ( .IN(CLK_25), .OUT(net044), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I95 ( .IN(net044), .OUT(net038), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
ml_dlatch_25 Ilatch2 ( .D_25(net053), .EN_25(net038), .R_25(R_25),
     .Q_25(Q_25));
ml_dlatch_25 Ilatch1 ( .Q_25(net053), .EN_25(net044), .D_25(D_25),
     .R_25(R_25));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_n, View - schematic
// LAST TIME SAVED: Aug  3 19:28:59 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_core_sa_comp_n ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(out_div), .B(vddp_), .G(out_ref), .S(vddp_));
P_25_LP  M5 ( .D(out_div), .B(vddp_), .G(saen_25), .S(vddp_));
P_25_LP  M1 ( .D(out_ref), .B(vddp_), .G(saen_25), .S(vddp_));
P_25_LP  M7 ( .D(out_ref), .B(vddp_), .G(out_ref), .S(vddp_));
N_25_LP  M3 ( .D(out_div), .B(GND_), .G(in_div), .S(net049));
N_25_LP  M8 ( .D(out_ref), .B(GND_), .G(in_ref), .S(net049));
N_25_LP  M6_1_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
N_25_LP  M6_0_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_top_n, View - schematic
// LAST TIME SAVED: Aug  3 19:28:59 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_core_sa_comp_top_n ( pump_chrg_25, in_div, in_ref, sa_bias,
     saen_25 );
output  pump_chrg_25;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M6_1_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
N_25_LP  M6_0_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
nand2_25 I103 ( .G(gnd_), .Pb(vddp_), .A(saen_25), .Y(chrg_b_25),
     .P(vddp_), .B(net27), .Gb(gnd_));
inv_25 I102 ( .IN(chrg_b_25), .OUT(pump_chrg_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I104 ( .IN(out_div2), .OUT(net27), .P(vddp_), .Pb(vddp_),
     .G(net087), .Gb(gnd_));
ml_core_sa_comp_n Icore_sa_comp_n0 ( .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp_n Iml_core_sa_comp_n1 ( .out_div(out_div2),
     .out_ref(out_ref2), .in_div(in_div2), .in_ref(in_ref2),
     .sa_bias(sa_bias), .saen_25(saen_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd25_nor2, View - schematic
// LAST TIME SAVED: Aug  3 19:29:06 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ls_vdd25_nor2 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor2_25 I79 ( .A(in), .Y(out_vddio_b), .Gb(gnd_), .G(gnd_), .Pb(sup),
     .P(sup), .B(out_vddio));
nor2_25 I151 ( .A(out_vddio_b), .Y(out_vddio), .Gb(gnd_), .G(gnd_),
     .Pb(sup), .P(sup), .B(in_b));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_reg, View - schematic
// LAST TIME SAVED: Sep 24 15:38:09 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpxa_reg ( freq_25, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, vpxa_int, bgr, fsm_vrdwl, pumpen, vpxa_clk_25 );
output  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25;

inout  vpxa_int;

input  bgr, pumpen, vpxa_clk_25;

output [1:0]  freq_25;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vrdwl_b_vpxa;

wire  [2:0]  vrdwl_vpxa;

wire  [1:0]  freq_in_25;



P_25_LP  M11_1_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
P_25_LP  M11_0_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
P_25_LP  M37 ( .D(net226), .B(vpxa_int), .G(vrdwl_vpxa[2]),
     .S(net229));
P_25_LP  M1 ( .D(net223), .B(vddp_), .G(saen_b_25), .S(vddp_));
P_25_LP  M5 ( .D(net270), .B(vpxa_int), .G(vrdwl_vpxa[1]), .S(net226));
P_25_LP  M3 ( .D(net229), .B(vpxa_int), .G(saen_b_vpxa), .S(vpxa_int));
P_25_LP  M6 ( .D(net237), .B(vpxa_int), .G(vrdwl_vpxa[0]), .S(net270));
P_25_LP  M8_1_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
P_25_LP  M8_0_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
N_25_LP  M32 ( .D(net229), .B(GND_), .G(vrdwl_b_vpxa[2]), .S(net226));
N_25_LP  M0_3_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
N_25_LP  M0_2_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
N_25_LP  M0_1_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
N_25_LP  M0_0_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
N_25_LP  M7 ( .D(net270), .B(GND_), .G(vrdwl_b_vpxa[0]), .S(net237));
N_25_LP  M4 ( .D(net226), .B(GND_), .G(vrdwl_b_vpxa[1]), .S(net270));
N_25_LP  M2 ( .D(sa_bias), .B(GND_), .G(saen_b_25), .S(gnd_));
RNPPO_LP_pcell2460 R28 ( .B(GND_), .MINUS(in_div_2), .PLUS(in_div_1));
RNPPO_LP_pcell2460 R20 ( .B(GND_), .MINUS(in_div_2), .PLUS(in_div_1));
RNPPO_LP_pcell2460 R27 ( .B(GND_), .MINUS(in_div_2), .PLUS(in_div_1));
RNPPO_LP_pcell2460 R26 ( .B(GND_), .MINUS(in_div_0), .PLUS(net202));
RNPPO_LP_pcell2460 R29 ( .B(GND_), .MINUS(in_div_2), .PLUS(in_div_1));
RNPPO_LP_pcell2460 R17 ( .B(GND_), .MINUS(net232), .PLUS(net223));
RNPPO_LP_pcell2460 R2 ( .B(GND_), .MINUS(net270), .PLUS(net226));
RNPPO_LP_pcell2460 R18 ( .B(GND_), .MINUS(net226), .PLUS(net229));
RNPPO_LP_pcell2460 R0 ( .B(GND_), .MINUS(sa_bias), .PLUS(net232));
RNPPO_LP_pcell2460 R10 ( .B(GND_), .MINUS(net202), .PLUS(net237));
RNPPO_LP_pcell2460 R3 ( .B(GND_), .MINUS(net237), .PLUS(net270));
RNPPO_LP_pcell2460 R30 ( .B(GND_), .MINUS(in_div_1), .PLUS(in_div_0));
RNPPO_LP_pcell2460 R12 ( .B(GND_), .MINUS(gnd_), .PLUS(in_div_2));
RNPPO_LP_pcell2460 R31 ( .B(GND_), .MINUS(in_div_1), .PLUS(in_div_0));
ml_ls_vdd2vdd25_vpxa I191 ( .in(saen_25), .sup(vpxa_int),
     .out_vddio_b(saen_b_vpxa), .out_vddio(net0210), .in_b(saen_b_25));
ml_ls_vdd2vdd25_vpxa I87 ( .in(net171), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[2]), .out_vddio(vrdwl_b_vpxa[2]),
     .in_b(net175));
ml_ls_vdd2vdd25_vpxa I98 ( .in(net176), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[1]), .out_vddio(vrdwl_b_vpxa[1]),
     .in_b(net180));
ml_ls_vdd2vdd25_vpxa I99 ( .in(net181), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[0]), .out_vddio(vrdwl_b_vpxa[0]),
     .in_b(net185));
nand2_25 I194 ( .G(GND_), .Pb(vddp_), .A(net0179), .Y(freq_in_25[1]),
     .P(vddp_), .B(net0234), .Gb(GND_));
nand2_25 I145 ( .G(GND_), .Pb(vddp_), .A(net0171), .Y(freq_in_25[0]),
     .P(vddp_), .B(net0179), .Gb(GND_));
nand3_25 I193 ( .B(pump_chrg_1_b_25), .A(pump_chrg_2_25), .Y(net0171),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I192 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0179),
     .C(pump_chrg_0_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I159 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0234),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
inv_25 I196 ( .IN(net169), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I197 ( .IN(net168), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I195 ( .IN(pump_chrg_0_25), .OUT(pump_chrg_0_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
inv_25 I154 ( .IN(pump_chrg_1_25), .OUT(pump_chrg_1_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_dff_25 I125 ( .Q_B_25(net0187), .R_25(saen_b_25),
     .D_25(freq_in_25[1]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[1]));
ml_dff_25 I126 ( .Q_B_25(net0192), .R_25(saen_b_25),
     .D_25(freq_in_25[0]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[0]));
inv_hvt I85 ( .A(net171), .Y(net175));
inv_hvt I183 ( .A(fsm_vrdwl[2]), .Y(net171));
inv_hvt I83 ( .A(pumpen), .Y(net143));
inv_hvt I82 ( .A(net143), .Y(net145));
inv_hvt I184 ( .A(fsm_vrdwl[1]), .Y(net176));
inv_hvt I187 ( .A(fsm_vrdwl[0]), .Y(net181));
inv_hvt I186 ( .A(net181), .Y(net185));
inv_hvt I185 ( .A(net176), .Y(net180));
ml_ls_vdd2vdd25 I335 ( .in(net145), .sup(vddp_), .out_vddio_b(net168),
     .out_vddio(net169), .in_b(net143));
ml_core_sa_comp_top_n Icore_sa_comp_top_n2 (
     .pump_chrg_25(pump_chrg_2_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_2));
ml_core_sa_comp_top_n core_sa_comp_top_n0 (
     .pump_chrg_25(pump_chrg_0_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_0));
ml_core_sa_comp_top_n Icore_sa_comp_top_n1 (
     .pump_chrg_25(pump_chrg_1_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_1));

endmodule
// Library - NVCM_40nm, Cell - ml_hv2vdd_sw, View - schematic
// LAST TIME SAVED: Aug  3 19:29:03 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv2vdd_sw ( out_hv, hv2vdd, vddp_tieh );
inout  out_hv;

input  hv2vdd, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LPNVT  M2 ( .D(vdd_), .B(GND_), .G(hv2vdd_25), .S(net27));
N_25_LPNVT  M0 ( .D(net27), .B(GND_), .G(vddp_tieh), .S(out_hv));
inv_25 I62 ( .IN(net40), .OUT(hv2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I71 ( .A(net46), .Y(net44));
inv_hvt I72 ( .A(hv2vdd), .Y(net46));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net40),
     .out_vddio(net37), .in_b(net46));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_top, View - schematic
// LAST TIME SAVED: Dec 15 11:51:52 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpxa_top ( vpxa_int, bgr, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint, fsm_vrdwl );
inout  vpxa_int;

input  bgr, fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  freq_25;



inv_25 I73 ( .IN(vpxa_clk_25), .OUT(vpxa_clk_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_pump_vpxa_x2 Ipump_vpxa_x3 ( .vpxa_clk_b_25(vpxa_clk_b_25),
     .vpxa_clk_25(vpxa_clk_25), .pumpen_25(pumpen_25),
     .pump_chrg_2_25(pump_chrg_2_25), .pump_chrg_1_25(pump_chrg_1_25),
     .pump_chrg_0_25(pump_chrg_0_25), .vpxa_int(vpxa_int));
ml_vpxa_osc Ivpxa_osc ( .freq_25(freq_25[1:0]), .bgr(bgr),
     .pumpen_25(pumpen_25), .vpxa_clk_25(vpxa_clk_25));
ml_vpxa_ctrl Ivpxa_ctrl ( .fsm_pumpen(fsm_pumpen), .pumpen(pumpen),
     .pumpen_25(pumpen_25), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .vpxa_2_vdd(vpxa_2_vdd));
vddp_tiehigh I118 ( .vddp_tieh(vddp_tieh));
ml_vpxa_reg Ivpxa_reg ( .pump_chrg_0_25(pump_chrg_0_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_2_25(pump_chrg_2_25),
     .freq_25(freq_25[1:0]), .vpxa_clk_25(vpxa_clk_25),
     .pumpen(pumpen), .fsm_vrdwl(fsm_vrdwl[2:0]), .bgr(bgr),
     .vpxa_int(vpxa_int));
ml_hv2vdd_sw Ivpxa_2vdd_sw ( .vddp_tieh(vddp_tieh),
     .hv2vdd(vpxa_2_vdd), .out_hv(vpxa_int));

endmodule
// Library - NVCM_40nm, Cell - ml_rdhv_gen, View - schematic
// LAST TIME SAVED: Aug  3 19:29:08 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_rdhv_gen ( s_rdin_hv, srdsup_hv, s_rdin, vddp_tieh );
output  s_rdin_hv;

inout  srdsup_hv;

input  s_rdin, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_s_b_hv_sw Iml_s_b_25_sw ( .sbout_high_25(s_rdin_high_25),
     .sbout_gnd_25(net31), .sbout_hv(s_rdin_hv), .ssup_hv(srdsup_hv),
     .vddp_tieh(vddp_tieh));
ml_ls_vdd2vdd25 Iml_ls_vdd2vdd25 ( .in(s_rdin), .sup(vddp_),
     .out_vddio_b(net31), .out_vddio(s_rdin_high_25), .in_b(net35));
inv_hvt I439 ( .A(s_rdin), .Y(net35));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_top_ctrl, View - schematic
// LAST TIME SAVED: Aug  3 19:29:05 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hvmux_top_ctrl ( bgrext_en, bgrint_en, en_vblinhi,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp, fsm_lshven,
     fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en );
output  bgrext_en, bgrint_en, en_vblinhi, ngate_vddp, ngate_vpxa,
     sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint,
     vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint, vpxaint_ext,
     vtmode, ysup25_2vdd, ysup25_2vddp;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor4_hvt I186 ( .D(fsm_tm_rprd), .C(fsm_rd), .A(fsm_tm_rd_mode),
     .B(fsm_pgmvfy), .Y(net0349));
nand4_hvt I322 ( .D(fsm_lshven), .A(fsm_pgm), .C(fsm_lshven),
     .Y(pgmpulse_b), .B(net0236));
nand4_hvt I35 ( .D(fsm_lshven), .C(net0318), .A(fsm_pgm), .Y(net0196),
     .B(net0327));
anor21_hvt I245 ( .A(net0189), .B(net0193), .Y(vppint_ext),
     .C(net0190));
anor21_hvt I109 ( .A(net0201), .B(net0199), .Y(vpxa_ext), .C(net0190));
nand3_hvt I288 ( .Y(net0193), .B(pmprd), .C(pmprd),
     .A(fsm_tm_xvppint));
nand3_hvt I291 ( .Y(net0201), .B(vddp_rd_b), .C(gnd_tiel),
     .A(fsm_tm_xforce));
nand3_hvt I292 ( .Y(net0213), .B(net0321), .C(net0196), .A(net0321));
nand3_hvt I290 ( .Y(net0199), .B(pmprd), .C(pmprd), .A(gnd_tiel));
nand3_hvt I289 ( .Y(net0189), .B(vpint_en), .C(fsm_tm_xvppint),
     .A(fsm_tm_xforce));
nor3_hvt I286 ( .B(net0240), .Y(rd_vddp), .A(net0240),
     .C(fsm_nvcmen_b));
nor3_hvt I285 ( .B(tm_testdec), .Y(en_vblinhi), .A(fsm_nvcmen_b),
     .C(tm_allbl_l));
mux2_hvt I260 ( .in1(fsm_wgnden), .in0(fsm_wpen), .out(net0217),
     .sel(pgmpulse_b));
nor2_hvt I272 ( .A(net75), .B(net93), .Y(ysup25_2vdd));
nor2_hvt I279 ( .A(net0251), .B(net0266), .Y(sbhvsup_vppint));
nor2_hvt I283 ( .A(vddp_rd_b), .B(net0258), .Y(vpxa_vppd));
nor2_hvt I271 ( .A(net87), .B(net73), .Y(ysup25_2vddp));
nor2_hvt I273 ( .A(net0349), .B(net0240), .Y(vddp_rd));
nor2_hvt I281 ( .A(net0324), .B(fsm_nvcmen_b), .Y(net0251));
nor2_hvt I276 ( .A(net0272), .B(rd_vddp), .Y(ngate_vpxa));
nor2_hvt I280 ( .A(net0268), .B(net0213), .Y(sb25sup_vpxa));
nor2_hvt I275 ( .A(net0331), .B(net0270), .Y(ngate_vddp));
nor2_hvt I274 ( .A(fsm_tm_rprd), .B(gnd_tiel), .Y(net0240));
nor2_hvt I278 ( .A(net0264), .B(net0311), .Y(sbhvsup_vddp));
nor2_hvt I282 ( .A(net0256), .B(vddp_rd), .Y(vpxa_vpxaint));
nor2_hvt I277 ( .A(net0325), .B(net0260), .Y(sb25sup_vddp));
inv_hvt I294 ( .A(net77), .Y(vtmode));
inv_hvt I323 ( .A(fsm_pgmvfy), .Y(net0236));
inv_hvt I319 ( .A(ngate_vpxa), .Y(net0339));
inv_hvt I304 ( .A(net0251), .Y(net0311));
inv_hvt I315 ( .A(vddp_rd), .Y(vddp_rd_b));
inv_hvt I318 ( .A(ysup25_2vdd), .Y(ysup25_2vdd_b));
inv_hvt I314 ( .A(vpxa_vppd), .Y(net0297));
inv_hvt I309 ( .A(net0277), .Y(bgrext_en));
inv_hvt I317 ( .A(fsm_pgmvfy), .Y(net0327));
inv_hvt I316 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I297 ( .A(ysup25_2vddp), .Y(ysup25_2vddp_b));
inv_hvt I298 ( .A(rd_vddp), .Y(net0331));
inv_hvt I310 ( .A(fsm_pumpen), .Y(net0190));
inv_hvt I307 ( .A(sbhvsup_vddp), .Y(net0309));
inv_hvt I305 ( .A(sb25sup_vpxa), .Y(net0323));
inv_hvt I308 ( .A(sbhvsup_vppint), .Y(net0313));
inv_hvt I296 ( .A(net93), .Y(net87));
inv_hvt I295 ( .A(net80), .Y(net93));
inv_hvt I321 ( .A(fsm_tm_rprd), .Y(net0318));
inv_hvt I303 ( .A(pgmpulse_b), .Y(net0324));
inv_hvt I306 ( .A(pgmpulse_b), .Y(pgmpulse));
inv_hvt I300 ( .A(sb25sup_vddp), .Y(net0329));
inv_hvt I302 ( .A(rd_vddp), .Y(net0321));
inv_hvt I301 ( .A(net0213), .Y(net0325));
inv_hvt I311 ( .A(net0286), .Y(vpxaint_ext));
inv_hvt I312 ( .A(fsm_tm_xforce), .Y(pmprd));
inv_hvt I299 ( .A(ngate_vddp), .Y(net0335));
inv_hvt I313 ( .A(vpxa_vpxaint), .Y(net0319));
inv_hvt I233 ( .A(fsm_nvcmen_b), .Y(fsm_nvcmen_buf));
nand2_hvt I268 ( .A(fsm_nvcmen_buf), .Y(net0277), .B(fsm_tm_xvbg));
nand2_hvt I266 ( .A(fsm_nvcmen), .Y(net80), .B(net0217));
nand2_hvt I269 ( .A(bgrext_en), .Y(bgrint_en), .B(fsm_tm_xforce));
nand2_hvt I267 ( .A(fsm_pumpen), .Y(net0286), .B(fsm_tm_xvpxaint));
nand2_hvt I104 ( .A(fsm_nvcmen), .Y(net77), .B(tm_wleqbl));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
ml_pump_a_clkdly I219 ( .in(ysup25_2vddp_b), .out(net75));
ml_pump_a_clkdly I227 ( .in(net0297), .out(net0256));
ml_pump_a_clkdly I226 ( .in(net0319), .out(net0258));
ml_pump_a_clkdly I209 ( .in(net0323), .out(net0260));
ml_pump_a_clkdly I184 ( .in(ysup25_2vdd_b), .out(net73));
ml_pump_a_clkdly I217 ( .in(net0313), .out(net0264));
ml_pump_a_clkdly I216 ( .in(net0309), .out(net0266));
ml_pump_a_clkdly I208 ( .in(net0329), .out(net0268));
ml_pump_a_clkdly I198 ( .in(net0339), .out(net0270));
ml_pump_a_clkdly I197 ( .in(net0335), .out(net0272));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_ls25, View - schematic
// LAST TIME SAVED: Aug  3 19:29:05 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hvmux_ls25 ( bgrext_en_25, bgrint_en_25, ngate_vddp_25,
     ngate_vpxa_25, sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25, bgrext_en, bgrint_en,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp );
output  bgrext_en_25, bgrint_en_25, ngate_vddp_25, ngate_vpxa_25,
     sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25;

input  bgrext_en, bgrint_en, ngate_vddp, ngate_vpxa, sb25sup_vddp,
     sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint, vppint_ext, vpxa_ext,
     vpxa_vppd, vpxa_vpxaint, vpxaint_ext, vtmode, ysup25_2vdd,
     ysup25_2vddp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_25 I471 ( .IN(net0138), .OUT(bgrint_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I472 ( .IN(net0148), .OUT(bgrext_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I473 ( .IN(net0128), .OUT(vppint_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I474 ( .IN(net0123), .OUT(vpxa_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I475 ( .IN(net0158), .OUT(vpxaint_ext_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I476 ( .IN(net0133), .OUT(vpxa_vppd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I477 ( .IN(net0163), .OUT(vpxa_vpxaint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I406 ( .IN(net077), .OUT(ysup25_2vddp_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I463 ( .IN(net0168), .OUT(ysup25_2vdd_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I464 ( .IN(net0193), .OUT(vtmode_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I465 ( .IN(net0173), .OUT(ngate_vddp_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I466 ( .IN(net0183), .OUT(ngate_vpxa_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I467 ( .IN(net0188), .OUT(sb25sup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I468 ( .IN(net0153), .OUT(sb25sup_vpxa_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I469 ( .IN(net0203), .OUT(sbhvsup_vppint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I470 ( .IN(net0198), .OUT(sbhvsup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_hvt I457 ( .A(vpxa_vppd), .Y(net054));
inv_hvt I435 ( .A(vpxa_vpxaint), .Y(net0112));
inv_hvt I462 ( .A(bgrint_en), .Y(net058));
inv_hvt I461 ( .A(bgrext_en), .Y(net068));
inv_hvt I460 ( .A(vppint_ext), .Y(net066));
inv_hvt I455 ( .A(ysup25_2vddp), .Y(net0328));
inv_hvt I454 ( .A(ysup25_2vdd), .Y(net0312));
inv_hvt I447 ( .A(ngate_vpxa), .Y(net0318));
inv_hvt I439 ( .A(sbhvsup_vppint), .Y(net0326));
inv_hvt I446 ( .A(sb25sup_vddp), .Y(net0320));
inv_hvt I216 ( .A(ysup25_2vdd), .Y(net092));
inv_hvt I458 ( .A(vpxaint_ext), .Y(net060));
inv_hvt I442 ( .A(sbhvsup_vddp), .Y(net0324));
inv_hvt I443 ( .A(sb25sup_vpxa), .Y(net0322));
inv_hvt I450 ( .A(ngate_vddp), .Y(net0316));
inv_hvt I217 ( .A(net092), .Y(ysup25_2vdd_buf));
inv_hvt I451 ( .A(vtmode), .Y(net0314));
inv_hvt I459 ( .A(vpxa_ext), .Y(net082));
ml_ls_vdd2vdd25 I336 ( .in(vpxa_ext), .sup(vddp_),
     .out_vddio_b(net0123), .out_vddio(net0207), .in_b(net082));
ml_ls_vdd2vdd25 I337 ( .in(vppint_ext), .sup(vddp_),
     .out_vddio_b(net0128), .out_vddio(net0208), .in_b(net066));
ml_ls_vdd2vdd25 I338 ( .in(vpxa_vppd), .sup(vddp_),
     .out_vddio_b(net0133), .out_vddio(net0211), .in_b(net054));
ml_ls_vdd2vdd25 I339 ( .in(bgrint_en), .sup(vddp_),
     .out_vddio_b(net0138), .out_vddio(net0209), .in_b(net058));
ml_ls_vdd2vdd25 I332 ( .in(bgrext_en), .sup(vddp_),
     .out_vddio_b(net0148), .out_vddio(net0149), .in_b(net068));
ml_ls_vdd2vdd25 I238 ( .in(sb25sup_vpxa), .sup(vddp_),
     .out_vddio_b(net0153), .out_vddio(net0154), .in_b(net0322));
ml_ls_vdd2vdd25 I334 ( .in(vpxaint_ext), .sup(vddp_),
     .out_vddio_b(net0158), .out_vddio(net0214), .in_b(net060));
ml_ls_vdd2vdd25 I335 ( .in(vpxa_vpxaint), .sup(vddp_),
     .out_vddio_b(net0163), .out_vddio(net0206), .in_b(net0112));
ml_ls_vdd2vdd25 I212 ( .in(ysup25_2vdd), .sup(vddp_),
     .out_vddio_b(net0168), .out_vddio(net0169), .in_b(net0312));
ml_ls_vdd2vdd25 I226 ( .in(ngate_vddp), .sup(vddp_),
     .out_vddio_b(net0173), .out_vddio(net0174), .in_b(net0316));
ml_ls_vdd2vdd25 I203 ( .in(net0328), .sup(vddp_), .out_vddio_b(net077),
     .out_vddio(net078), .in_b(ysup25_2vddp));
ml_ls_vdd2vdd25 I221 ( .in(ngate_vpxa), .sup(vddp_),
     .out_vddio_b(net0183), .out_vddio(net0184), .in_b(net0318));
ml_ls_vdd2vdd25 I233 ( .in(sb25sup_vddp), .sup(vddp_),
     .out_vddio_b(net0188), .out_vddio(net0219), .in_b(net0320));
ml_ls_vdd2vdd25 I207 ( .in(vtmode), .sup(vddp_), .out_vddio_b(net0193),
     .out_vddio(net0194), .in_b(net0314));
ml_ls_vdd2vdd25 I260 ( .in(sbhvsup_vddp), .sup(vddp_),
     .out_vddio_b(net0198), .out_vddio(net0220), .in_b(net0324));
ml_ls_vdd2vdd25 I261 ( .in(sbhvsup_vppint), .sup(vddp_),
     .out_vddio_b(net0203), .out_vddio(net0204), .in_b(net0326));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_bgrxcvr, View - schematic
// LAST TIME SAVED: Aug  3 19:29:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_hvmux_bgrxcvr ( bgr, bgr_int, bgrint_en_25, vpp,
     bgrext_en_25, vddp_tieh );
inout  bgr, bgr_int, bgrint_en_25, vpp;

input  bgrext_en_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LPNVT  M0 ( .D(bgr), .B(GND_), .G(bgrint_en_25), .S(bgr_int));
N_25_LP  M2 ( .D(vpp), .B(GND_), .G(vddp_tieh), .S(net53));
N_25_LP  M1 ( .D(net53), .B(GND_), .G(bgrext_en_25), .S(bgr));

endmodule
// Library - NVCM_40nm, Cell - ml_ysup_25_switch, View - schematic
// LAST TIME SAVED: Aug  3 19:29:18 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_ysup_25_switch ( vdd, vddp, ysup_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25 );
inout  vdd, vddp, ysup_25;

input  ysup25_2vdd_25, ysup25_2vdd_buf, ysup25_2vddp_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(ysup_25), .B(ysup_25), .G(ysup25_2vdd_buf),
     .S(net73));
P_25_LP  M5 ( .D(net73), .B(vddp), .G(ysup25_2vddp_b_25), .S(vddp));
N_25_LPNVT  M13 ( .D(vdd), .B(GND_), .G(ysup25_2vdd_25), .S(ysup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_vblinhi, View - schematic
// LAST TIME SAVED: Aug  3 19:29:16 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_ymux_ctrl_vblinhi ( vblinhi, vpxa, en_vblinhi, vtmode,
     vtmode_25 );
inout  vblinhi, vpxa;

input  en_vblinhi, vtmode, vtmode_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M8 ( .D(vpxa), .B(GND_), .G(vtmode_25), .S(net035));
N_25_LP  M9 ( .D(net035), .B(GND_), .G(net035), .S(vblinhi));
P_11_LPHVT  M7_9_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_8_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_7_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_6_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_5_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_4_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_3_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_2_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_1_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
P_11_LPHVT  M7_0_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv),
     .S(vdd_));
N_11_LPHVT  M0_9_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_8_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_7_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_6_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_5_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_4_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_3_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_2_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_1_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
N_11_LPHVT  M0_0_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv),
     .S(gnd_));
nor2_hvt I191 ( .A(en_vblinhi), .B(vtmode_buf), .Y(ngate_inhi_lv));
inv_hvt I192 ( .A(net063), .Y(vtmode_buf));
inv_hvt I190 ( .A(vtmode), .Y(net063));
nand2_hvt I104 ( .A(net063), .Y(pgate_inhi_lv), .B(en_vblinhi));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_top, View - schematic
// LAST TIME SAVED: Aug  3 19:29:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_hvmux_top ( s_rdin_hv, bgr, bgr_int, ngate_25, sb25sup_25,
     sbhvsup_hv, srdsup_hv, vblinhi, vpp, vpp_int, vpxa, vpxa_int,
     ysup_25, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen,
     fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, s_rd,
     tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );

inout  bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv,
     vblinhi, vpp, vpp_int, vpxa, vpxa_int, ysup_25;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en;

output [3:0]  s_rdin_hv;

input [3:0]  s_rd;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_rdin;

wire  [3:0]  net294;



P_25_LP  M9 ( .D(vddp_tieh), .B(vddp_), .G(net299), .S(vddp_));
N_11_LPHVT  M1 ( .D(net299), .B(GND_), .G(net299), .S(gnd_));
inv_hvt I210_3_ ( .A(s_rd[3]), .Y(net294[0]));
inv_hvt I210_2_ ( .A(s_rd[2]), .Y(net294[1]));
inv_hvt I210_1_ ( .A(s_rd[1]), .Y(net294[2]));
inv_hvt I210_0_ ( .A(s_rd[0]), .Y(net294[3]));
inv_hvt I211_3_ ( .A(net294[0]), .Y(s_rdin[3]));
inv_hvt I211_2_ ( .A(net294[1]), .Y(s_rdin[2]));
inv_hvt I211_1_ ( .A(net294[2]), .Y(s_rdin[1]));
inv_hvt I211_0_ ( .A(net294[3]), .Y(s_rdin[0]));
ml_rdhv_gen Iml_rdhv_inv_3_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[3]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[3]));
ml_rdhv_gen Iml_rdhv_inv_2_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[2]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[2]));
ml_rdhv_gen Iml_rdhv_inv_1_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[1]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[1]));
ml_rdhv_gen Iml_rdhv_inv_0_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[0]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[0]));
ml_hv_hotswitch_enhance Ixcvr_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(vppint_ext_25), .hv_in_hv(vpp_int), .hv_out_hv(vpp));
ml_hvmux_top_ctrl Ihvmux_top_ctrl ( .fsm_tm_rprd(fsm_tm_rprd),
     .vpint_en(vpint_en), .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl),
     .tm_testdec(tm_testdec), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_lshven(fsm_lshven), .ysup25_2vddp(ysup25_2vddp),
     .ysup25_2vdd(ysup25_2vdd), .vtmode(vtmode),
     .vpxaint_ext(vpxaint_ext), .vpxa_vpxaint(vpxa_vpxaint),
     .vpxa_vppd(vpxa_vppd), .vpxa_ext(vpxa_ext),
     .vppint_ext(vppint_ext), .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .en_vblinhi(en_vblinhi),
     .bgrint_en(bgrint_en), .bgrext_en(bgrext_en));
ml_hvmux_ls25 Ihvmux_ls25 ( .ysup25_2vddp(ysup25_2vddp),
     .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vppint_25(sbhvsup_vppint_25), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en), .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vtmode_25(vtmode_25),
     .vpxaint_ext_25(vpxaint_ext_25),
     .vpxa_vpxaint_25(vpxa_vpxaint_25), .vpxa_vppd_25(vpxa_vppd_25),
     .vpxa_ext_25(net309), .vppint_ext_25(vppint_ext_25),
     .sbhvsup_vddp_25(sbhvsup_vddp_25),
     .sb25sup_vpxa_25(sb25sup_vpxa_25),
     .sb25sup_vddp_25(sb25sup_vddp_25), .ngate_vpxa_25(ngate_vpxa_25),
     .ngate_vddp_25(ngate_vddp_25), .bgrint_en_25(bgrint_en_25),
     .bgrext_en_25(bgrext_en_25));
ml_hvmux_bgrxcvr Ixcvr_bgr ( .vddp_tieh(vddp_tieh),
     .bgrext_en_25(bgrext_en_25), .vpp(vpp),
     .bgrint_en_25(bgrint_en_25), .bgr_int(bgr_int), .bgr(bgr));
ml_hv_hotswitch Ixcvr_vpxa_int ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa_int), .hv_out_hv(vpp));
ml_hvmux_hotswitch I212 ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(srdsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sbhvsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(sbhvsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sb25sup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sb25sup_vpxa_25), .sel_hv_a_25(sb25sup_vddp_25),
     .out_hv(sb25sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_ngate ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(ngate_vpxa_25), .sel_hv_a_25(ngate_vddp_25),
     .out_hv(ngate_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_1_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vddp_), .hvin_a_hv(vpxa_int));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_0_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vddp_), .hvin_a_hv(vpxa_int));
ml_ysup_25_switch Isw_ysup25_1_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ysup_25_switch Isw_ysup25_0_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_1_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_0_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yptest, View - schematic
// LAST TIME SAVED: Aug  3 19:29:17 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yptest ( yp_test_25, yp_test_b_25, yp_test,
     yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25, ysup_25 );
output  yp_test_25, yp_test_b_25;

input  yp_test, yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25,
     ysup_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I181 ( .A(yp_test), .Y(net40));
inv_25 I182 ( .IN(net028), .OUT(yp_test_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));
oai21x2_sup_25 I180 ( .A1(yp_test_b_low_ysup_25), .Y(yp_test_b_25),
     .A0(net37), .B0(yp_test_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(yp_test), .sup(ysup_25),
     .out_vddio_b(net028), .out_vddio(net37), .in_b(net40));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_hvsw_8f, View - schematic
// LAST TIME SAVED: Dec 15 15:10:09 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_chip_nvcm_hvsw_8f ( s_rdin_hv, bgr, ngate_25, sb25sup_25,
     sbhvsup_hv, srdsup_hv, vblinhi, vpp, vpp_int, vpxa, vpxa_int,
     ysup_25, fsm_bgr_dis, fsm_lshven, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_trim_vbg, fsm_vpgmwl,
     fsm_vrdwl, fsm_wgnden, fsm_wpen, s_rd, tm_allbl_l, tm_wleqbl );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi, vpp,
     vpp_int, vpxa, vpxa_int, ysup_25;

input  fsm_bgr_dis, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_wleqbl;

output [3:0]  s_rdin_hv;

input [2:0]  fsm_vpgmwl;
input [2:0]  fsm_vrdwl;
input [3:0]  s_rd;
input [3:0]  fsm_trim_vbg;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_bgr_top Ibgr_top ( .fsm_trim_vbg_buf(fsm_trim_vbg[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen), .fsm_bgr_dis_buf(fsm_bgr_dis),
     .bgr_int(bgr_int));
ml_vppint_top Ivppint_top ( .vpxa(vpxa),
     .fsm_vpgmwl_buf(fsm_vpgmwl[2:0]), .fsm_pgmdisc_buf(fsm_pgmdisc),
     .fsm_pgm_buf(fsm_pgm), .fsm_lshven_buf(fsm_lshven),
     .vpint_en(vpint_en), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmvfy_buf(fsm_pgmvfy), .fsm_wgnden_buf(fsm_wgnden),
     .fsm_nvcmen_buf(fsm_nvcmen), .bgr(bgr), .vpp_int(vpp_int),
     .fsm_tm_xvppint(fsm_tm_xvppint));
ml_vpxa_top Ivpxa_top ( .fsm_vrdwl(fsm_vrdwl[2:0]),
     .fsm_tm_xvpxaint(fsm_tm_xvpxaint), .fsm_tm_xforce(fsm_tm_xforce),
     .bgr(bgr), .vpxa_int(vpxa_int), .fsm_pumpen(fsm_pumpen));
ml_hvmux_top Ihvmux_top ( .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_lshven(fsm_lshven), .bgr(bgr), .bgr_int(bgr_int),
     .ngate_25(ngate_25), .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .vpp(vpp), .vpp_int(vpp_int),
     .vpxa(vpxa), .ysup_25(ysup_25), .vblinhi(vblinhi),
     .tm_testdec(fsm_tm_testdec), .srdsup_hv(srdsup_hv),
     .s_rd(s_rd[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rdin_hv(s_rdin_hv[3:0]), .vpint_en(vpint_en),
     .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl), .vpxa_int(vpxa_int));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_384, View - schematic
// LAST TIME SAVED: Dec 15 15:10:11 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_chip_nvcm_384 ( nv_dataout, vpp, vpp_int, vpxa_int,
     fsm_bgr_dis, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_multibl_read, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_pumpen,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxaint,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_trim_vbg,
     fsm_vpgmwl, fsm_vpxaset, fsm_vrdwl, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl
     );

inout  vpp, vpp_int, vpxa_int;

input  fsm_bgr_dis, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxaint,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl;

output [8:0]  nv_dataout;

input [2:0]  fsm_vpgmwl;
input [2:0]  fsm_trim_rrefpgm;
input [9:0]  fsm_coladd;
input [3:0]  fsm_trim_vbg;
input [2:0]  fsm_vrdwl;
input [1:0]  fsm_tm_ref;
input [7:0]  fsm_rowadd;
input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_rdin_hv;

wire  [3:0]  s_rd;



ml_chip_nvcm_core_384 Iml_chip_nvcm_core_384 (
     .fsm_tm_ref(fsm_tm_ref[1:0]), .fsm_wren(fsm_wren),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rdin_hv(s_rdin_hv[3:0]),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[8:0]),
     .fsm_pgmhv(fsm_pgmhv), .fsm_gwlbdis(fsm_gwlbdis),
     .vpp_int(vpp_int), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_pgm(fsm_pgm),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_din(fsm_din), .fsm_rd(fsm_rd), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_pgmdisc(fsm_pgmdisc),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ngate_25(ngate_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol), .bgr(bgr),
     .fsm_blkadd(fsm_blkadd[3:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi(vblinhi), .s_rd(s_rd[3:0]), .srdsup_hv(srdsup_hv),
     .ysup_25(ysup_25), .vpxa(vpxa));
ml_chip_nvcm_hvsw_8f Ihvsw ( .vpxa_int(vpxa_int), .bgr(bgr),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .vpp_int(vpp_int), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd), .fsm_wpen(fsm_wpen),
     .s_rdin_hv(s_rdin_hv[3:0]), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .srdsup_hv(srdsup_hv), .s_rd(s_rd[3:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .tm_allbl_l(tm_allbl_l),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_pumpen(fsm_pumpen), .sb25sup_25(sb25sup_25),
     .fsm_lshven(fsm_lshven), .sbhvsup_hv(sbhvsup_hv), .vpxa(vpxa),
     .ysup_25(ysup_25), .ngate_25(ngate_25), .fsm_wgnden(fsm_wgnden),
     .vblinhi(vblinhi), .tm_wleqbl(tm_wleqbl), .vpp(vpp),
     .fsm_vrdwl(fsm_vrdwl[2:0]), .fsm_bgr_dis(fsm_bgr_dis),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_vpgmwl(fsm_vpgmwl[2:0]), .fsm_tm_testdec(fsm_tm_testdec));

endmodule
// Library - leafcell, Cell - tiehi, View - schematic
// LAST TIME SAVED: Aug  3 19:21:04 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module tiehi ( tiehi );
output  tiehi;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));
N_11_LPHVT  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - leafcell, Cell - tielo, View - schematic
// LAST TIME SAVED: Aug  3 19:21:04 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module tielo ( tielo );
output  tielo;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_11_LPHVT  M2 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));
P_11_LPHVT  M1 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - ice8chip, Cell - sg_bufx10_ice8p, View - schematic
// LAST TIME SAVED: Jul 30 23:15:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module sg_bufx10_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - ice384chip, Cell - nvcm_ml_block_ice384_june, View -
//schematic
// LAST TIME SAVED: Jan 18 15:49:28 2012
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module nvcm_ml_block_ice384_june ( bp0, fsm_recall,
     fsm_tm_margin0_read, idcode_msb20bits_out, nvcm_boot,
     nvcm_dis_idchk, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b,
     tgnd_fsm, tvdd_fsm, vpp, vpp_int, vpxa_int, clk, nvcm_ce_b, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot,
     nvcm_dis_idchk, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b,
     tgnd_fsm, tvdd_fsm;

inout  vpp, vpp_int, vpxa_int;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

output [19:0]  idcode_msb20bits_out;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [8:0]  nv_dataout;

wire  [3:0]  fsm_blkadd;

wire  [3:0]  net178;

wire  [2:0]  fsm_trim_vrdwl;

wire  [2:0]  fsm_trim_vpgmwl;

wire  [3:0]  fsm_trim_vbg;

wire  [2:0]  fsm_trim_rrefrd;

wire  [2:0]  fsm_trim_rrefpgm;

wire  [3:0]  fsm_trim_ipp;

wire  [3:0]  fsm_blkadd_b;

wire  [1:0]  fsm_tm_ref_buf;

wire  [11:0]  fsm_coladd;

wire  [8:0]  fsm_rowadd;



nvcm_top_id_u40 I_nvcm_top_id_u40 ( .nvcm_dis_idchk(nvcm_dis_idchk),
     .idcode_msb20bits_out(idcode_msb20bits_out[19:0]),
     .idcode_msb20bits_in({tgnd_fsm, tgnd_fsm, tgnd_fsm, tvdd_fsm,
     tgnd_fsm, tgnd_fsm, tgnd_fsm, tvdd_fsm, tgnd_fsm, tgnd_fsm,
     tgnd_fsm, tvdd_fsm, tvdd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm,
     tgnd_fsm, tvdd_fsm, tgnd_fsm, tgnd_fsm}), .trim_spare({net178[0],
     net178[1], net178[2], net178[3]}), .fsm_tm_bgr_dis(fsm_bgr_dis),
     .fsm_tm_allbank_sel(fsm_tm_allbank_sel),
     .fsm_coladd(fsm_coladd[11:0]), .nvcm_max_coladd({tgnd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tgnd_fsm, tvdd_fsm, tgnd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm, tvdd_fsm}),
     .nvcm_max_rowadd({tgnd_fsm, tgnd_fsm, tgnd_fsm, tgnd_fsm,
     tvdd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm, tvdd_fsm}),
     .status_wip(net55), .fsm_tm_ref(fsm_tm_ref_buf[1:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .nvcm_boot(nvcm_boot),
     .spi_ss_b(spi_ss_b), .spi_sdi(spi_sdi),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_ce_b(nvcm_ce_b), .nv_dataout(nv_dataout[8:0]), .clk(clk),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .nvcm_relextspi(nvcm_relextspi), .nvcm_rdy(nvcm_rdy),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_trim_vrdwl(fsm_trim_vrdwl[2:0]),
     .fsm_trim_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_multibl_read(fsm_trim_multibl_read),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxa_int(fsm_tm_xvpxa_int), .fsm_tm_xvpp(fsm_tm_xvpp),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_vwleqbl(fsm_tm_vwleqbl),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_testdec_wr(fsm_tm_testdec_wr),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_tcol(fsm_tm_tcol),
     .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_margin0_read(fsm_tm_margin0_read),
     .fsm_tm_dma(fsm_tm_dma), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_sample(fsm_sample),
     .fsm_rowadd(fsm_rowadd[8:0]), .fsm_recall(fsm_recall),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_redrow(fsm_nv_redrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .bp0(bp0));
ml_chip_nvcm_384 I_ml_chip_nvcm_384 ( .vpp_int(vpp_int),
     .vpxa_int(vpxa_int), .fsm_tm_ref(fsm_tm_ref_buf[1:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .fsm_bgr_dis(fsm_bgr_dis),
     .tm_allbank_sel(fsm_tm_allbank_sel), .fsm_coladd(fsm_coladd[9:0]),
     .tm_wleqbl(fsm_tm_vwleqbl), .tm_testdec_wr(fsm_tm_testdec_wr),
     .tm_tcol(fsm_tm_tcol), .tm_dma(fsm_tm_dma),
     .tm_allwl_l(fsm_tm_allwl_l), .tm_allwl_h(fsm_tm_allwl_h),
     .tm_allbl_l(fsm_tm_allbl_l), .tm_allbl_h(fsm_tm_allbl_h),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vrdwl(fsm_trim_vrdwl[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxaint(fsm_tm_xvpxa_int), .fsm_tm_xvppint(fsm_tm_xvpp),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(rst_bd), .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rrow(fsm_nv_redrow), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_multibl_read(fsm_trim_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .nv_dataout(nv_dataout[8:0]), .vpp(vpp));
tiehi I442 ( .tiehi(tvdd_fsm));
tielo I369 ( .tielo(tgnd_fsm));
sg_bufx10_ice8p I541 ( .in(rst_b), .out(rst_bd));

endmodule
// Library - xpmem, Cell - ml_blsa_clk_buf, View - schematic
// LAST TIME SAVED: Jul 30 23:15:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_clk_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_powersurg_buf, View - schematic
// LAST TIME SAVED: Jul 30 23:15:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_powersurg_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I404 ( .A(net016), .Y(net012));
inv_hvt I405 ( .A(net012), .Y(o));
inv_hvt I391 ( .A(net77), .Y(net016));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jul 30 23:15:00 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_sch, View - schematic
// LAST TIME SAVED: Aug  3 19:22:00 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_sch ( dataout, bl, prec_sup, cram_prec, cram_pullup_b,
     cram_write, data_muxsel, datain, latch_clock, latch_reset,
     prec_hold_b, smc_wdic_clk );
output  dataout;

inout  bl, prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, datain,
     latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_11_LPHVT  MN8 ( .D(sa_out), .B(gnd_), .G(cram_pullup_b), .S(gnd_));
N_11_LPHVT  M1 ( .D(net0166), .B(gnd_), .G(n_gate), .S(gnd_));
N_11_LPHVT  MN3 ( .D(sa_out), .B(gnd_), .G(bl), .S(gnd_));
N_11_LPHVT  MN6 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
N_11_LPHVT  MN12 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
P_11_LPHVT  MP9 ( .D(bl), .B(vdd_), .G(net084), .S(net0148));
P_11_LPHVT  M0 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
P_11_LPHVT  M3 ( .D(net0110), .B(vdd_), .G(cram_write), .S(prec_sup));
P_11_LPHVT  MP8 ( .D(net0148), .B(vdd_), .G(dataout), .S(vdd_));
P_11_LPHVT  MP12 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
P_11_LPHVT  M2 ( .D(bl), .B(vdd_), .G(prec_hold_b), .S(net0110));
P_11_LPHVT  MP4 ( .D(net0143), .B(vdd_), .G(cram_pullup_b), .S(vdd_));
P_11_LPHVT  MP5 ( .D(sa_out), .B(vdd_), .G(bl), .S(net0143));
ml_dff Idff ( .R(latch_reset), .D(dff_in), .CLK(latch_clock),
     .QN(write_data_b), .Q(dff_data));
nor2_hvt I223 ( .A(net084), .B(write_data_b), .Y(n_gate));
inv_hvt I163 ( .A(write_data_b), .Y(dataout));
inv_hvt I159 ( .A(cram_prec), .Y(net0161));
inv_hvt I160 ( .A(cram_write), .Y(net084));
mux2_hvt I161 ( .in1(sa_out), .in0(datain), .out(latch_in),
     .sel(data_muxsel));
mux2_hvt I164 ( .in1(dff_data), .in0(latch_in), .out(dff_in),
     .sel(smc_wdic_clk));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_yp3_sup_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:56 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module oai21x2_yp3_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M6 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));
P_25_LP  M5 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));
P_25_LP  M4 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
N_25_LP  M12 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
N_25_LP  M1 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
N_25_LP  M0 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));

endmodule
// Library - xpmem, Cell - ml_blsa_tile, View - schematic
// LAST TIME SAVED: Jan  7 13:26:29 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_tile ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [53:0]  bl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [53:0]  dataout;

wire  [13:0]  ck;



inv_hvt I172 ( .A(net48), .Y(data_out));
inv_hvt I171 ( .A(dataout[53]), .Y(net48));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_powersurg_buf I161 ( .in(cram_write), .o(net53));
ml_powersurg_buf I165 ( .in(net57), .o(net55));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net57));
ml_powersurg_buf I163 ( .in(net55), .o(net59));
ml_powersurg_buf I162 ( .in(net65), .o(net61));
ml_powersurg_buf I169 ( .in(net61), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net53), .o(net65));
ml_powersurg_buf I168 ( .in(net59), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_47_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[47]),
     .dataout(dataout[47]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_46_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[46]),
     .dataout(dataout[46]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_45_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[45]),
     .dataout(dataout[45]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_44_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[44]),
     .dataout(dataout[44]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_43_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[43]),
     .dataout(dataout[43]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_42_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[42]),
     .dataout(dataout[42]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net55));
ml_blsa_sch I170_53_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[53]), .dataout(dataout[53]),
     .cram_prec(net57));
ml_blsa_sch I170_52_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[52]), .dataout(dataout[52]),
     .cram_prec(net57));
ml_blsa_sch I170_51_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[51]), .dataout(dataout[51]),
     .cram_prec(net57));
ml_blsa_sch I170_50_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[50]), .dataout(dataout[50]),
     .cram_prec(net57));
ml_blsa_sch I170_49_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[49]), .dataout(dataout[49]),
     .cram_prec(net57));
ml_blsa_sch I170_48_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[48]), .dataout(dataout[48]),
     .cram_prec(net57));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net59));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_1st, View - schematic
// LAST TIME SAVED: Jul 30 23:15:06 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_tile_1st ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [55:0]  bl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:1]  data_dummy_in;

wire  [5:1]  data_in;

wire  [55:0]  dataout;

wire  [14:0]  ck;



ml_dff I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net132), .Q(net154));
ml_dff I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net137), .Q(data_dummy_in[4]));
ml_dff I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net142), .Q(data_dummy_in[2]));
ml_dff I179 ( .R(latch_reset), .D(datain), .CLK(ck[14]), .QN(net147),
     .Q(data_dummy_in[1]));
ml_dff I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net152), .Q(data_dummy_in[3]));
inv_hvt I171 ( .A(dataout[55]), .Y(net121));
inv_hvt I172 ( .A(net121), .Y(data_out));
inv_hvt I224 ( .A(net0130), .Y(ck[14]));
inv_hvt I225 ( .A(net0129), .Y(net0130));
inv_hvt I226 ( .A(net0126), .Y(net0129));
inv_hvt I229 ( .A(latch_clock), .Y(net0122));
inv_hvt I227 ( .A(net0124), .Y(net0126));
inv_hvt I228 ( .A(net0122), .Y(net0124));
mux2_hvt I197 ( .in1(net154), .in0(dataout[4]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I232 ( .in1(data_dummy_in[2]), .in0(dataout[1]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I230 ( .in1(data_dummy_in[4]), .in0(dataout[3]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I233 ( .in1(data_dummy_in[1]), .in0(dataout[0]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I231 ( .in1(data_dummy_in[3]), .in0(dataout[2]),
     .out(data_in[3]), .sel(data_muxsel1));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[14]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[13]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[12]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[11]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[10]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[9]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[8]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[7]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[6]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[4]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[3]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[2]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[1]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(datain), .cram_prec(cram_prec_out),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_47_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[47]),
     .dataout(dataout[47]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_46_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[46]),
     .dataout(dataout[46]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_45_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[45]),
     .dataout(dataout[45]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_44_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[44]),
     .dataout(dataout[44]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_43_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[43]),
     .dataout(dataout[43]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_42_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[42]),
     .dataout(dataout[42]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[41]),
     .dataout(dataout[41]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[40]),
     .dataout(dataout[40]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[39]),
     .dataout(dataout[39]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[38]),
     .dataout(dataout[38]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[37]),
     .dataout(dataout[37]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[36]),
     .dataout(dataout[36]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[35]),
     .dataout(dataout[35]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[34]),
     .dataout(dataout[34]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[33]),
     .dataout(dataout[33]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[32]),
     .dataout(dataout[32]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_55_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[54]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[55]),
     .dataout(dataout[55]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_54_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[53]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[54]),
     .dataout(dataout[54]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_53_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[53]),
     .dataout(dataout[53]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_52_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[52]),
     .dataout(dataout[52]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_51_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[51]),
     .dataout(dataout[51]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_50_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[50]),
     .dataout(dataout[50]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_49_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[49]),
     .dataout(dataout[49]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_48_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[48]),
     .dataout(dataout[48]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[31]),
     .dataout(dataout[31]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[30]),
     .dataout(dataout[30]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[29]),
     .dataout(dataout[29]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[28]),
     .dataout(dataout[28]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[27]),
     .dataout(dataout[27]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[26]),
     .dataout(dataout[26]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[25]),
     .dataout(dataout[25]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[24]),
     .dataout(dataout[24]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[23]),
     .dataout(dataout[23]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[22]),
     .dataout(dataout[22]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[21]),
     .dataout(dataout[21]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[20]),
     .dataout(dataout[20]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[19]),
     .dataout(dataout[19]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[18]),
     .dataout(dataout[18]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[17]),
     .dataout(dataout[17]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[16]),
     .dataout(dataout[16]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_powersurg_buf I161 ( .in(cram_write), .o(net104));
ml_powersurg_buf I165 ( .in(net108), .o(net106));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net108));
ml_powersurg_buf I163 ( .in(net106), .o(net110));
ml_powersurg_buf I162 ( .in(net116), .o(net112));
ml_powersurg_buf I169 ( .in(net112), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net104), .o(net116));
ml_powersurg_buf I168 ( .in(net110), .o(cram_prec_out));

endmodule
// Library - xpmem, Cell - ml_blprecwrt_en, View - schematic
// LAST TIME SAVED: Jul 30 23:15:06 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blprecwrt_en ( data_out, action, clkin, data_in, rst );
output  data_out;

input  action, clkin, data_in, rst;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor3_hvt I105 ( .B(net86), .Y(net94), .A(net98), .C(rst));
nor2_hvt I103 ( .A(net88), .B(net94), .Y(net98));
inv_hvt I66 ( .A(net89), .Y(net88));
inv_hvt I168 ( .A(action), .Y(net86));
inv_hvt I165 ( .A(net98), .Y(data_out));
nand3_hvt I160 ( .Y(net89), .B(data_in), .C(action), .A(clkin));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_1st_ice1f, View - schematic
// LAST TIME SAVED: Aug  3 19:22:01 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_tilex2_1st_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [109:0]  bl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M3 ( .D(prec_sup), .B(vdd_), .G(net106), .S(vdd_));
ml_blsa_tile Iml_blsa_tile_1 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_wdic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[109:56]));
ml_blsa_tile_1st Iml_blsa_tile_1st_0 ( .prec_sup(prec_sup),
     .prec_hold_b(prec_hold_b), .bl(bl[55:0]),
     .cram_pullup_b(cram_pullup_buf), .latch_clock(latch_clock_out),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .datain(datain), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_mid),
     .cram_prec(prec_en_mid), .data_out(data_tile),
     .cram_write_out(wrt_out), .cram_prec_out(prec_en_last));
nor2_hvt I385 ( .A(latch_reset), .B(net86), .Y(net117));
tiehi I284 ( .tiehi(prec_hold_b));
inv_hvt I190 ( .A(net095), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net095));
inv_hvt I202 ( .A(latch_reset), .Y(net0113));
inv_hvt I203 ( .A(net0113), .Y(latch_reset_buf));
inv_hvt I196 ( .A(cram_pullup_b), .Y(net0109));
inv_hvt I204 ( .A(net0105), .Y(smc_wdic_clk_buf));
inv_hvt I200 ( .A(prec_hold_b), .Y(net106));
inv_hvt I205 ( .A(smc_wdic_clk), .Y(net0105));
inv_hvt I221 ( .A(net138), .Y(net110));
inv_hvt I197 ( .A(net0109), .Y(cram_pullup_buf));
inv_hvt I198 ( .A(net099), .Y(latch_clock_out));
inv_hvt I199 ( .A(latch_clock_in), .Y(net099));
inv_hvt I201 ( .A(net117), .Y(net118));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net118), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net138));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net86));

endmodule
// Library - leafcell, Cell - tiehis, View - schematic
// LAST TIME SAVED: Aug  3 19:21:04 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module tiehis ( tiehi );
output  tiehi;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPRVT  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));
N_11_LPRVT  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - xpmem, Cell - ml_buf_ice5, View - schematic
// LAST TIME SAVED: Jul 30 23:15:06 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_buf_ice5 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_last, View - schematic
// LAST TIME SAVED: Jul 30 23:15:06 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_tile_last ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [17:0]  bl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:0]  ck;

wire  [17:0]  dataout;



ml_dff Idff ( .R(latch_reset), .D(dataout[16]), .CLK(ck[0]),
     .QN(net50), .Q(net45));
ml_dff I179 ( .R(latch_reset), .D(net58), .CLK(ck[0]), .QN(net49),
     .Q(net61));
mux2_hvt I174 ( .in1(net45), .in0(dataout[17]), .out(net58),
     .sel(data_muxsel));
tiehis I185 ( .tiehi(net040));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_buf_ice5 I205 ( .in(net61), .o(data_out), .sel(net040));
ml_powersurg_buf I169 ( .in(cram_write), .o(cram_write_out));
ml_powersurg_buf I168 ( .in(cram_prec), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[16]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[17]), .dataout(dataout[17]));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[15]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[16]), .dataout(dataout[16]));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex1_last_ice1f, View - schematic
// LAST TIME SAVED: Nov  3 11:49:01 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_tilex1_last_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [71:0]  bl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M0 ( .D(prec_sup), .B(vdd_), .G(net0122), .S(vdd_));
nor2_hvt I385 ( .A(net0111), .B(latch_reset), .Y(net0121));
ml_blsa_tile_last Iml_blsa_tile_last ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .bl(bl[71:54]),
     .latch_reset(latch_reset_buf), .datain(datain_io),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_1st), .cram_prec_out(prec_en_1st),
     .latch_clock(latch_clock_out), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blsa_tile Iml_blsa_tile_0 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_dic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_1st), .cram_prec(prec_en_1st),
     .data_out(datain_io), .cram_write_out(wrt_out),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
tiehi I284 ( .tiehi(prec_hold_b));
inv_hvt I197 ( .A(prec_hold_b), .Y(net0122));
inv_hvt I194 ( .A(smc_wdic_clk), .Y(net0125));
inv_hvt I196 ( .A(net0124), .Y(net066));
inv_hvt I187 ( .A(net0121), .Y(net068));
inv_hvt I193 ( .A(latch_reset), .Y(net0127));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net0133));
inv_hvt I204 ( .A(net0137), .Y(latch_clock_out));
inv_hvt I208 ( .A(net0125), .Y(smc_dic_clk_buf));
inv_hvt I192 ( .A(latch_clock_in), .Y(net0137));
inv_hvt I190 ( .A(net0139), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net0139));
inv_hvt I203 ( .A(net0133), .Y(cram_pullup_b_buf));
inv_hvt I207 ( .A(net0127), .Y(latch_reset_buf));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net068), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net0124));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net0111));

endmodule
// Library - xpmem, Cell - ml_buf_ice1f, View - schematic
// LAST TIME SAVED: Jan  7 14:21:36 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_buf_ice1f ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_dff_bl, View - schematic
// LAST TIME SAVED: Jul 30 23:15:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_dff_bl ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yp3, View - schematic
// LAST TIME SAVED: Aug  3 19:29:16 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp3 ( yp3_25, yp3_b_25, yp3_b_high_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, ysup_25 );
output  yp3_25, yp3_b_25;

input  yp3_b_high_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, ysup_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



oai21x2_yp3_sup_25 I209 ( .A1(yp3_b_low_ysup_25), .Y(yp3_b_25),
     .A0(net069), .B0(yp3_b_high_b_ysup_25), .ysup_25(ysup_25));
inv_hvt I201 ( .A(yp3_sel), .Y(net075));
inv_hvt I101 ( .A(net075), .Y(net070));
inv_25 I204 ( .IN(yp3_25_b), .OUT(yp3_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd25_nor2 I192 ( .in(net070), .sup(ysup_25),
     .out_vddio_b(yp3_25_b), .out_vddio(net069), .in_b(net075));

endmodule
// Library - xpmem, Cell - ml_blsa_bank_ice384, View - schematic
// LAST TIME SAVED: Dec 16 17:07:19 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_blsa_bank_ice384 ( cm_sdo_u, bl, banksel, cm_sdi_u,
     cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk,
     smc_write );


input  banksel, cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk,
     smc_write;

output [1:0]  cm_sdo_u;

inout [181:0]  bl;

input [1:0]  cm_sdi_u;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tilex2_1st_ice1f I_lt_01 ( .wrt_in(wrt_out_1),
     .prec_in(prec_out_1), .latch_reset(latch_reset_buf),
     .datain(sdi0_buf), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .bl(bl[109:0]), .cram_prec(cram_prec_buf), .wrt_out(wrt_out_0),
     .prec_out(prec_out_0), .data_out(data_out_0),
     .latch_clock_in(net0137), .smc_write(smc_write_buf),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_out(net440),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf_b_ret));
ml_blsa_tilex1_last_ice1f I_lt_2 ( .smc_write(smc_write_buf),
     .bl(bl[181:110]), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(smc_clk), .latch_clock_out(net0137),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf),
     .wrt_in(cram_write_buf), .prec_in(net377),
     .latch_reset(latch_reset_buf), .datain(data_out_0),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_1), .prec_out(prec_out_1),
     .data_out(cm_sdo_u[1]));
ml_buf_ice1f I247 ( .in(cm_sdi_u[1]), .o(net0237), .sel(net527));
ml_buf_ice1f I249 ( .in(net519), .o(cor_en_8bpcfg_buf), .sel(net527));
ml_buf_ice1f I265 ( .in(net527), .o(cm_sdo_u[0]), .sel(net451));
ml_buf_ice1f I257 ( .in(smc_wdic_clk), .o(smc_wdic_clk_buf),
     .sel(banksel));
ml_buf_ice1f I203 ( .in(data_muxsel1), .o(data_muxsel1_buf),
     .sel(banksel));
ml_buf_ice1f I205 ( .in(latch_reset), .o(latch_reset_buf),
     .sel(net529));
ml_buf_ice1f I207 ( .in(cram_write), .o(cram_write_buf),
     .sel(banksel));
ml_buf_ice1f I208 ( .in(cram_pullup_logic_b), .o(cram_pullup_b_buf),
     .sel(cram_pullup_logic_b));
ml_buf_ice1f I201 ( .in(cram_prec), .o(cram_prec_buf), .sel(banksel));
ml_buf_ice1f I294b ( .in(banksel), .o(smc_write_buf), .sel(smc_write));
ml_buf_ice1f I216 ( .in(net528), .o(net474), .sel(net528));
ml_buf_ice1f I245 ( .in(cm_sdi_u[0]), .o(sdi0_buf), .sel(net527));
ml_buf_ice1f I187 ( .in(smc_clk), .o(smc_clk_buf), .sel(smc_clk));
ml_buf_ice1f I188 ( .in(net525), .o(smc_clk_buf_b_ret), .sel(net525));
ml_buf_ice1f I204 ( .in(data_muxsel), .o(data_muxsel_buf),
     .sel(banksel));
ml_buf_ice1f I227 ( .in(net532), .o(net489), .sel(net532));
nor3_hvt I217 ( .B(net531), .Y(net492), .A(net531), .C(net531));
nor3_hvt I220 ( .B(net500), .Y(net496), .A(net500), .C(net500));
nor3_hvt I218 ( .B(net492), .Y(net500), .A(net492), .C(net492));
nand3_hvt I231 ( .Y(net503), .B(net507), .C(net507), .A(net507));
nand3_hvt I230 ( .Y(net507), .B(net511), .C(net511), .A(net511));
nand3_hvt I224 ( .Y(net511), .B(net526), .C(net526), .A(net526));
nor2_hvt I254 ( .B(net515), .Y(net522), .A(cram_pullup_b));
inv_hvt I253 ( .A(cor_en_8bpcfg_b), .Y(net519));
inv_hvt I256 ( .A(banksel), .Y(net515));
inv_hvt I255 ( .A(net522), .Y(cram_pullup_logic_b));
inv_hvt I189 ( .A(smc_clk), .Y(net525));
tiehi I268 ( .tiehi(net526));
tiehi I272 ( .tiehi(net527));
tiehi I271 ( .tiehi(net528));
tiehi I273 ( .tiehi(net529));
tiehi I267 ( .tiehi(net377));
tiehi I270 ( .tiehi(net531));
tiehi I269 ( .tiehi(net532));
ml_dff_bl I_ml_dff_bl ( .R(latch_reset_buf), .D(net527), .CLK(smc_clk),
     .QN(net536), .Q(net451));

endmodule
// Library - ice384chip, Cell - CHIP_route_top_ice384, View - schematic
// LAST TIME SAVED: Nov  4 18:18:36 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module CHIP_route_top_ice384 ( cm_sdo_u1, cm_sdo_u3, bl_top,
     cm_banksel_bltld3, cm_banksel_bltrd1, cm_clk_bltld3,
     cm_clk_bltrd1, cm_prec_bltld3, cm_sdi_u1d3, cm_sdi_u3d2,
     core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1r,
     smc_write_bltl1d1, smc_write_bltld3 );


input  cm_clk_bltld3, cm_clk_bltrd1, cm_prec_bltld3, core_por_b_rowu1,
     core_por_b_rowu3, cram_prec_bltrd1, cram_pullup_b_bltrd1,
     cram_pullup_bltld3, cram_write_bltld3, cram_write_bltrd1,
     data_muxsel1_bltld3, data_muxsel1_bltrd1, data_muxsel_bltld3,
     data_muxsel_bltrd1, en_8bconfig_b_bltld3, en_8bconfig_b_bltrd1,
     smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1r, smc_write_bltl1d1,
     smc_write_bltld3;

output [1:0]  cm_sdo_u3;
output [1:0]  cm_sdo_u1;

inout [363:0]  bl_top;

input [1:0]  cm_sdi_u1d3;
input [1:1]  cm_banksel_bltld3;
input [3:3]  cm_banksel_bltrd1;
input [1:0]  cm_sdi_u3d2;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_bank_ice384 I_bltr ( .bl(bl_top[363:182]),
     .smc_write(smc_write_bltl1d1),
     .smc_wdic_clk(smc_wdis_dclk_bltrd1r), .smc_clk(cm_clk_bltrd1),
     .cm_sdi_u(cm_sdi_u3d2[1:0]), .latch_reset(core_por_b_rowu3),
     .cm_sdo_u(cm_sdo_u3[1:0]), .data_muxsel1(data_muxsel1_bltrd1),
     .data_muxsel(data_muxsel_bltrd1), .cram_write(cram_write_bltrd1),
     .cram_prec(cram_prec_bltrd1),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltrd1),
     .cram_pullup_b(cram_pullup_b_bltrd1),
     .banksel(cm_banksel_bltrd1[3]));
ml_blsa_bank_ice384 I_bltlu1 ( .bl({bl_top[0], bl_top[1], bl_top[2],
     bl_top[3], bl_top[4], bl_top[5], bl_top[6], bl_top[7], bl_top[8],
     bl_top[9], bl_top[10], bl_top[11], bl_top[12], bl_top[13],
     bl_top[14], bl_top[15], bl_top[16], bl_top[17], bl_top[18],
     bl_top[19], bl_top[20], bl_top[21], bl_top[22], bl_top[23],
     bl_top[24], bl_top[25], bl_top[26], bl_top[27], bl_top[28],
     bl_top[29], bl_top[30], bl_top[31], bl_top[32], bl_top[33],
     bl_top[34], bl_top[35], bl_top[36], bl_top[37], bl_top[38],
     bl_top[39], bl_top[40], bl_top[41], bl_top[42], bl_top[43],
     bl_top[44], bl_top[45], bl_top[46], bl_top[47], bl_top[48],
     bl_top[49], bl_top[50], bl_top[51], bl_top[52], bl_top[53],
     bl_top[54], bl_top[55], bl_top[56], bl_top[57], bl_top[58],
     bl_top[59], bl_top[60], bl_top[61], bl_top[62], bl_top[63],
     bl_top[64], bl_top[65], bl_top[66], bl_top[67], bl_top[68],
     bl_top[69], bl_top[70], bl_top[71], bl_top[72], bl_top[73],
     bl_top[74], bl_top[75], bl_top[76], bl_top[77], bl_top[78],
     bl_top[79], bl_top[80], bl_top[81], bl_top[82], bl_top[83],
     bl_top[84], bl_top[85], bl_top[86], bl_top[87], bl_top[88],
     bl_top[89], bl_top[90], bl_top[91], bl_top[92], bl_top[93],
     bl_top[94], bl_top[95], bl_top[96], bl_top[97], bl_top[98],
     bl_top[99], bl_top[100], bl_top[101], bl_top[102], bl_top[103],
     bl_top[104], bl_top[105], bl_top[106], bl_top[107], bl_top[108],
     bl_top[109], bl_top[110], bl_top[111], bl_top[112], bl_top[113],
     bl_top[114], bl_top[115], bl_top[116], bl_top[117], bl_top[118],
     bl_top[119], bl_top[120], bl_top[121], bl_top[122], bl_top[123],
     bl_top[124], bl_top[125], bl_top[126], bl_top[127], bl_top[128],
     bl_top[129], bl_top[130], bl_top[131], bl_top[132], bl_top[133],
     bl_top[134], bl_top[135], bl_top[136], bl_top[137], bl_top[138],
     bl_top[139], bl_top[140], bl_top[141], bl_top[142], bl_top[143],
     bl_top[144], bl_top[145], bl_top[146], bl_top[147], bl_top[148],
     bl_top[149], bl_top[150], bl_top[151], bl_top[152], bl_top[153],
     bl_top[154], bl_top[155], bl_top[156], bl_top[157], bl_top[158],
     bl_top[159], bl_top[160], bl_top[161], bl_top[162], bl_top[163],
     bl_top[164], bl_top[165], bl_top[166], bl_top[167], bl_top[168],
     bl_top[169], bl_top[170], bl_top[171], bl_top[172], bl_top[173],
     bl_top[174], bl_top[175], bl_top[176], bl_top[177], bl_top[178],
     bl_top[179], bl_top[180], bl_top[181]}),
     .smc_write(smc_write_bltld3), .smc_wdic_clk(smc_wdis_dclk_bltld3),
     .smc_clk(cm_clk_bltld3), .cm_sdi_u(cm_sdi_u1d3[1:0]),
     .latch_reset(core_por_b_rowu1), .cm_sdo_u(cm_sdo_u1[1:0]),
     .data_muxsel1(data_muxsel1_bltld3),
     .data_muxsel(data_muxsel_bltld3), .cram_write(cram_write_bltld3),
     .cram_prec(cm_prec_bltld3),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltld3),
     .cram_pullup_b(cram_pullup_bltld3),
     .banksel(cm_banksel_bltld3[1]));

endmodule
// Library - ice384chip, Cell - CHIP_route_bot_ice384_blbank, View -
//schematic
// LAST TIME SAVED: Nov  4 18:25:54 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module CHIP_route_bot_ice384_blbank ( cm_sdo_u0, cm_sdo_u2, bl_bot,
     cm_banksel_blbld1_0_, cm_banksel_blbrd_2_, cm_clk_blbld,
     cm_clk_blbrd, cm_sdi_u0d1, cm_sdi_u2d, core_por_bb, core_por_bbl0,
     cram_prec, cram_prec_blbld, cram_pullup_b, cram_pullup_blbld,
     cram_write, cram_write_blbld, data_muxsel1_blbld,
     data_muxsel1_blbrd, data_muxsel_blbld, data_muxsel_blbrd,
     en_8bconfig_b_blbld, en_8bconfig_b_blbrd, smc_wdis_dclk_blbld,
     smc_wdis_dclk_blbrd, smc_write, smc_writel0 );


input  cm_banksel_blbld1_0_, cm_banksel_blbrd_2_, cm_clk_blbld,
     cm_clk_blbrd, core_por_bb, core_por_bbl0, cram_prec,
     cram_prec_blbld, cram_pullup_b, cram_pullup_blbld, cram_write,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel1_blbrd,
     data_muxsel_blbld, data_muxsel_blbrd, en_8bconfig_b_blbld,
     en_8bconfig_b_blbrd, smc_wdis_dclk_blbld, smc_wdis_dclk_blbrd,
     smc_write, smc_writel0;

output [1:0]  cm_sdo_u0;
output [1:0]  cm_sdo_u2;

inout [363:0]  bl_bot;

input [1:0]  cm_sdi_u2d;
input [1:0]  cm_sdi_u0d1;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



CHIP_route_top_ice384 I_CHIP_route_top_ice384 ( .bl_top(bl_bot[363:0]),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_blbld),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_blbrd),
     .en_8bconfig_b_bltld3(en_8bconfig_b_blbld),
     .data_muxsel_bltrd1(data_muxsel_blbrd),
     .data_muxsel_bltld3(data_muxsel_blbld),
     .data_muxsel1_bltrd1(data_muxsel1_blbrd),
     .data_muxsel1_bltld3(data_muxsel1_blbld),
     .cram_write_bltrd1(cram_write),
     .cram_write_bltld3(cram_write_blbld),
     .cram_pullup_bltld3(cram_pullup_blbld),
     .cram_pullup_b_bltrd1(cram_pullup_b),
     .cram_prec_bltrd1(cram_prec), .core_por_b_rowu3(core_por_bb),
     .core_por_b_rowu1(core_por_bbl0), .cm_sdi_u3d2(cm_sdi_u2d[1:0]),
     .cm_sdi_u1d3(cm_sdi_u0d1[1:0]), .cm_prec_bltld3(cram_prec_blbld),
     .cm_clk_bltrd1(cm_clk_blbrd), .cm_clk_bltld3(cm_clk_blbld),
     .cm_banksel_bltrd1(cm_banksel_blbrd_2_),
     .cm_banksel_bltld3(cm_banksel_blbld1_0_),
     .cm_sdo_u3(cm_sdo_u2[1:0]), .cm_sdo_u1(cm_sdo_u0[1:0]),
     .smc_write_bltld3(smc_writel0), .smc_write_bltl1d1(smc_write));

endmodule
// Library - ice8chip, Cell - sg_dffbuf_modified, View - schematic
// LAST TIME SAVED: Aug 19 09:09:59 2010
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module sg_dffbuf_modified ( dffout, clk, d, r );
output  dffout;

input  clk, d, r;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_dff I0 ( .R(r), .D(d), .CLK(clk), .QN(net9), .Q(net10));
sg_bufx10_ice8p I5 ( .in(net10), .out(dffout));

endmodule
// Library - ice8chip, Cell - eh_io_pup_2_new_ice8p, View - schematic
// LAST TIME SAVED: Oct  3 11:29:53 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module eh_io_pup_2_new_ice8p ( por_b, core_por_b, vdd_io );
output  por_b;

input  core_por_b, vdd_io;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M5 ( .D(net0221), .B(vdd_io), .G(net0221), .S(vdd_io));
P_25_LP  M3 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
P_25_LP  M7 ( .D(v_in), .B(vdd_io), .G(net145), .S(net0221));
P_25_LP  M6 ( .D(net0221), .B(vdd_io), .G(net0221), .S(vdd_io));
P_25_LP  M4 ( .D(net0221), .B(vdd_io), .G(net0221), .S(vdd_io));
P_25_LP  M11 ( .D(net104), .B(vdd_), .G(v_in), .S(vdd_));
P_25_LP  M1 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
P_11_LPHVT  M0 ( .D(net84), .B(vdd_), .G(net104), .S(vdd_));
P_11_LPHVT  MP8 ( .D(net104), .B(vdd_), .G(core_por_b), .S(vdd_));
N_11_LPHVT  M2 ( .D(net84), .B(gnd_), .G(net104), .S(gnd_));
N_11_LPHVT  MN1 ( .D(net0196), .B(gnd_), .G(core_por_b), .S(gnd_));
N_25_LP  M8 ( .D(net104), .B(gnd_), .G(v_in), .S(net104));
N_25_LP  M23 ( .D(net104), .B(gnd_), .G(v_in), .S(net0196));
N_25_LP  M22 ( .D(net104), .B(gnd_), .G(v_in), .S(net104));
N_25_LP  MN6 ( .D(v_in), .B(gnd_), .G(net145), .S(gnd_));
N_25_LP  M10 ( .D(net0175), .B(gnd_), .G(net147), .S(net158));
N_25_LP  M28 ( .D(gnd_), .B(gnd_), .G(core_por_b), .S(gnd_));
N_25_LP  M14 ( .D(v_in), .B(gnd_), .G(net147), .S(net0224));
RNPPO_LP_pcell2460 R66 ( .B(gnd_), .MINUS(gnd_), .PLUS(net145));
N_25_LPNVT  M27 ( .D(net0224), .B(gnd_), .G(net0224), .S(net0132));
N_25_LPNVT  M24 ( .D(net0132), .B(gnd_), .G(net0132), .S(net0220));
N_25_LPNVT  M25 ( .D(net0220), .B(gnd_), .G(net0220), .S(net0216));
N_25_LPNVT  M9 ( .D(net158), .B(gnd_), .G(net158), .S(net154));
N_25_LPNVT  M13 ( .D(net150), .B(gnd_), .G(net150), .S(net162));
N_25_LPNVT  M16 ( .D(v_in), .B(gnd_), .G(net147), .S(v_in));
N_25_LPNVT  M20 ( .D(net162), .B(gnd_), .G(net162), .S(net0112));
N_25_LPNVT  M12 ( .D(net154), .B(gnd_), .G(net154), .S(net150));
N_25_LPNVT  M26 ( .D(net0216), .B(gnd_), .G(net0216), .S(gnd_));
N_25_LPNVT  M21 ( .D(net0112), .B(gnd_), .G(net0112), .S(gnd_));
sg_bufx10_ice8p I_clkbuf ( .in(net84), .out(por_b));
vdd_tiehigh I96 ( .vdd_tieh(net147));

endmodule
// Library - ice384chip, Cell - CHIP_route_bot_ice384, View - schematic
// LAST TIME SAVED: Dec 28 13:28:46 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module CHIP_route_bot_ice384 ( cm_banksel_blbld1_0_,
     cm_banksel_blbld_1_, cm_clk_blbld, cm_sdi_u1d, cm_sdo_u0d1,
     cm_sdo_u1d3, cm_sdo_u2d1, core_por_bbl0, cram_pgateoffl0,
     cram_prec_blbld, cram_pullup_blbld, cram_rstl0, cram_vddoffl0,
     cram_wl_enl0, cram_write_blbld, data_muxsel1_blbld,
     data_muxsel_blbld, en_8bconfig_b_blbld, j_rst_bl0, last_rsr3,
     row_testl1, smc_core_por_bottom1, smc_core_por_bottom2,
     smc_row_incl0, smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0,
     spi_ss_in_bbankd, tck_padl0, bl_bot, cm_banksel,
     cm_banksel_blbrd_2_, cm_clk_blbrd, cm_sdi_u0, cm_sdi_u1,
     cm_sdi_u2d, cm_sdo_u1d1, core_por_b0, core_por_bb, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     spi_ss_in_bbank, vddio_botbank, vddio_spi );
output  cm_banksel_blbld1_0_, cm_banksel_blbld_1_, cm_clk_blbld,
     core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, last_rsr3, row_testl1,
     smc_core_por_bottom1, smc_core_por_bottom2, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;


input  cm_banksel_blbrd_2_, cm_clk_blbrd, core_por_b0, core_por_bb,
     cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     vddio_botbank, vddio_spi;

output [1:0]  cm_sdo_u0d1;
output [1:0]  cm_sdi_u1d;
output [4:0]  spi_ss_in_bbankd;
output [1:0]  cm_sdo_u1d3;
output [1:0]  cm_sdo_u2d1;

inout [363:0]  bl_bot;

input [1:0]  cm_sdi_u0;
input [1:0]  cm_sdi_u2d;
input [4:0]  spi_ss_in_bbank;
input [1:0]  cm_banksel;
input [1:0]  cm_sdi_u1;
input [1:0]  cm_sdo_u1d1;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net231;

wire  [1:0]  dff_u1_d1;

wire  [1:0]  cm_sdo_u0_buf;

wire  [1:0]  cm_sdo_u1_buf;

wire  [1:0]  dff_u2_d0;

wire  [1:0]  net227;

wire  [1:0]  cm_sdo_u2;

wire  [1:0]  cm_sdi_u0d1;

wire  [1:0]  cm_sdo_u0;

wire  [1:0]  dff_u0_d1;

wire  [1:0]  net232;



CHIP_route_bot_ice384_blbank I_CHIP_route_bot_ice384_blbank (
     .bl_bot(bl_bot[363:0]), .smc_writel0(smc_writel0),
     .smc_write(smc_write), .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_write(cram_write),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_pullup_b(cram_pullup_b), .cram_prec_blbld(cram_prec_blbld),
     .cram_prec(cram_prec), .core_por_bbl0(core_por_bbl0),
     .core_por_bb(core_por_bb), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u0d1(cm_sdi_u0d1[1:0]), .cm_clk_blbrd(cm_clk_blbrd),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1_0_),
     .cm_sdo_u0(cm_sdo_u0[1:0]), .cm_sdo_u2(cm_sdo_u2[1:0]));
tielo I561_1_ ( .tielo(net227[0]));
tielo I561_0_ ( .tielo(net227[1]));
tielo I562 ( .tielo(net228));
tielo I563 ( .tielo(net229));
tielo I564 ( .tielo(net230));
tielo I559_1_ ( .tielo(net231[0]));
tielo I559_0_ ( .tielo(net231[1]));
tielo I560_1_ ( .tielo(net232[0]));
tielo I560_0_ ( .tielo(net232[1]));
sg_bufx10_ice8p I484 ( .in(cram_pgateoff), .out(cram_pgateoffl0));
sg_bufx10_ice8p I333 ( .in(j_rst_b), .out(j_rst_bl0));
sg_bufx10_ice8p I336 ( .in(core_por_bb), .out(core_por_bbl0));
sg_bufx10_ice8p I523 ( .in(smc_clk_mid), .out(cm_clk_blbld));
sg_bufx10_ice8p I478 ( .in(cram_vddoff), .out(cram_vddoffl0));
sg_bufx10_ice8p I473 ( .in(smc_write), .out(smc_writel0));
sg_bufx10_ice8p I496 ( .in(en_8bconfig_b_blbrd),
     .out(en_8bconfig_b_blbld));
sg_bufx10_ice8p I527_1_ ( .in(cm_sdi_u0[1]), .out(cm_sdi_u0d1[1]));
sg_bufx10_ice8p I527_0_ ( .in(cm_sdi_u0[0]), .out(cm_sdi_u0d1[0]));
sg_bufx10_ice8p I459 ( .in(smc_row_inc), .out(smc_row_incl0));
sg_bufx10_ice8p I491 ( .in(cram_write), .out(cram_write_blbld));
sg_bufx10_ice8p I568_4_ ( .in(spi_ss_in_bbank[4]),
     .out(spi_ss_in_bbankd[4]));
sg_bufx10_ice8p I568_3_ ( .in(spi_ss_in_bbank[3]),
     .out(spi_ss_in_bbankd[3]));
sg_bufx10_ice8p I568_2_ ( .in(spi_ss_in_bbank[2]),
     .out(spi_ss_in_bbankd[2]));
sg_bufx10_ice8p I568_1_ ( .in(spi_ss_in_bbank[1]),
     .out(spi_ss_in_bbankd[1]));
sg_bufx10_ice8p I568_0_ ( .in(spi_ss_in_bbank[0]),
     .out(spi_ss_in_bbankd[0]));
sg_bufx10_ice8p I439 ( .in(j_tck), .out(tck_padl0));
sg_bufx10_ice8p I485 ( .in(cram_prec), .out(cram_prec_blbld));
sg_bufx10_ice8p I533_1_ ( .in(cm_sdi_u1[1]), .out(cm_sdi_u1d[1]));
sg_bufx10_ice8p I533_0_ ( .in(cm_sdi_u1[0]), .out(cm_sdi_u1d[0]));
sg_bufx10_ice8p I519 ( .in(cm_banksel[0]), .out(cm_banksel_blbld1_0_));
sg_bufx10_ice8p I504 ( .in(smc_rsr_rst), .out(smc_rsr_rstl0));
sg_bufx10_ice8p I490 ( .in(cram_pullup_b), .out(cram_pullup_blbld));
sg_bufx10_ice8p I479 ( .in(cram_rst), .out(cram_rstl0));
sg_bufx10_ice8p I465 ( .in(data_muxsel1_blbrd),
     .out(data_muxsel1_blbld));
sg_bufx10_ice8p I525 ( .in(cm_clk_blbrd), .out(predata_smc_clk_out));
sg_bufx10_ice8p I518 ( .in(cm_banksel[1]), .out(cm_banksel_blbld_1_));
sg_bufx10_ice8p I524 ( .in(predata_smc_clk_out), .out(smc_clk_mid));
sg_bufx10_ice8p I511 ( .in(row_test0), .out(row_testl1));
sg_bufx10_ice8p I293 ( .in(last_rsr1), .out(last_rsr2));
sg_bufx10_ice8p I541_1_ ( .in(dff_u0_d1[1]), .out(cm_sdo_u0d1[1]));
sg_bufx10_ice8p I541_0_ ( .in(dff_u0_d1[0]), .out(cm_sdo_u0d1[0]));
sg_bufx10_ice8p I539_1_ ( .in(cm_sdo_u1d1[1]), .out(cm_sdo_u1_buf[1]));
sg_bufx10_ice8p I539_0_ ( .in(cm_sdo_u1d1[0]), .out(cm_sdo_u1_buf[0]));
sg_bufx10_ice8p I455 ( .in(data_muxsel_blbrd),
     .out(data_muxsel_blbld));
sg_bufx10_ice8p I566 ( .in(net385), .out(last_rsr3));
sg_bufx10_ice8p I540_1_ ( .in(dff_u1_d1[1]), .out(cm_sdo_u1d3[1]));
sg_bufx10_ice8p I540_0_ ( .in(dff_u1_d1[0]), .out(cm_sdo_u1d3[0]));
sg_bufx10_ice8p I497 ( .in(smc_wdis_dclk_blbrd),
     .out(smc_wdis_dclk_blbld));
sg_bufx10_ice8p I472 ( .in(cram_wl_en), .out(cram_wl_enl0));
sg_dffbuf_modified I462_1_ ( .d(cm_sdo_u0_buf[1]), .clk(smc_clk_mid),
     .dffout(dff_u0_d1[1]), .r(net227[0]));
sg_dffbuf_modified I462_0_ ( .d(cm_sdo_u0_buf[0]), .clk(smc_clk_mid),
     .dffout(dff_u0_d1[0]), .r(net227[1]));
sg_dffbuf_modified I565 ( .d(last_rsr2), .clk(smc_clk_mid),
     .dffout(net385), .r(net230));
sg_dffbuf_modified I537_1_ ( .d(cm_sdo_u1_buf[1]), .clk(smc_clk_mid),
     .dffout(dff_u1_d1[1]), .r(net232[0]));
sg_dffbuf_modified I537_0_ ( .d(cm_sdo_u1_buf[0]), .clk(smc_clk_mid),
     .dffout(dff_u1_d1[0]), .r(net232[1]));
sg_dffbuf_modified I545_1_ ( .d(dff_u2_d0[1]),
     .clk(predata_smc_clk_out), .dffout(cm_sdo_u2d1[1]), .r(net229));
sg_dffbuf_modified I545_0_ ( .d(dff_u2_d0[0]),
     .clk(predata_smc_clk_out), .dffout(cm_sdo_u2d1[0]), .r(net229));
sg_dffbuf_modified I546_1_ ( .d(cm_sdo_u2[1]),
     .clk(predata_smc_clk_out), .dffout(dff_u2_d0[1]), .r(net228));
sg_dffbuf_modified I546_0_ ( .d(cm_sdo_u2[0]),
     .clk(predata_smc_clk_out), .dffout(dff_u2_d0[0]), .r(net228));
sg_dffbuf_modified I535_1_ ( .d(cm_sdo_u0[1]), .clk(cm_clk_blbld),
     .dffout(cm_sdo_u0_buf[1]), .r(net231[0]));
sg_dffbuf_modified I535_0_ ( .d(cm_sdo_u0[0]), .clk(cm_clk_blbld),
     .dffout(cm_sdo_u0_buf[0]), .r(net231[1]));
eh_io_pup_2_new_ice8p Ipor_spi ( .core_por_b(core_por_b0),
     .vdd_io(vddio_spi), .por_b(smc_core_por_bottom2));
eh_io_pup_2_new_ice8p Ipor_iob ( .core_por_b(core_por_b0),
     .vdd_io(vddio_botbank), .por_b(smc_core_por_bottom1));

endmodule
// Library - ice384chip, Cell - smc_and_jtag_id_u40, View - schematic
// LAST TIME SAVED: Dec 13 13:46:03 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module smc_and_jtag_id_u40 ( bm_bank_sdi, bm_banksel, bm_clk, bm_init,
     bm_rcapmux_en, bm_sa, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_banksel, cm_clk, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2, cm_sdi_u3, data_muxsel, data_muxsel1,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0, j_hiz_b,
     j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck, j_tdi,
     j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, psdo, rst_b,
     smc_load_nvcm_bstream, smc_osc_fsel, smc_oscoff_b, smc_podt_off,
     smc_podt_rst, smc_read, smc_row_inc, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rsr_rst, smc_rwl_en, smc_seq_rst,
     smc_wcram_rst, smc_wdis_dclk, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, tdo_oe_pad, tdo_pad,
     bm_bank_sdo, boot, bp0, bschain_sdo, cdone_in, cm_last_rsr,
     cm_monitor_cell, cm_sdo_u0, cm_sdo_u1, cm_sdo_u2, cm_sdo_u3,
     cnt_podt_out, coldboot_sel, creset_b, idcode_msb20bits, nvcm_boot,
     nvcm_dis_idchk, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, osc_clk, por_b, psdi, spi_clk_in, spi_sdi,
     spi_ss_in_b, tck_pad, tdi_pad, tms_pad, trst_pad, warmboot_sel );
output  bm_clk, bm_init, bm_rcapmux_en, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_clk, data_muxsel,
     data_muxsel1, en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0,
     j_hiz_b, j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck,
     j_tdi, j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, rst_b,
     smc_load_nvcm_bstream, smc_oscoff_b, smc_podt_off, smc_podt_rst,
     smc_read, smc_row_inc, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rsr_rst, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_wdis_dclk, smc_write, smc_wset_prec, smc_wset_precgnd,
     smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_oe_pad, tdo_pad;

input  boot, bp0, bschain_sdo, cdone_in, cm_last_rsr, cnt_podt_out,
     creset_b, nvcm_boot, nvcm_dis_idchk, nvcm_rdy, nvcm_relextspi,
     nvcm_spi_sdo, nvcm_spi_sdo_oe_b, osc_clk, por_b, spi_clk_in,
     spi_sdi, spi_ss_in_b, tck_pad, tdi_pad, tms_pad, trst_pad;

output [1:0]  smc_osc_fsel;
output [3:0]  cm_banksel;
output [1:0]  cm_sdi_u3;
output [3:0]  bm_banksel;
output [3:0]  bm_bank_sdi;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_sdi_u0;
output [10:0]  bm_sa;
output [1:0]  cm_sdi_u2;
output [7:1]  psdo;

input [1:0]  warmboot_sel;
input [3:0]  bm_bank_sdo;
input [3:0]  cm_monitor_cell;
input [1:0]  coldboot_sel;
input [19:0]  idcode_msb20bits;
input [1:0]  cm_sdo_u0;
input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdo_u3;
input [7:1]  psdi;
input [1:0]  cm_sdo_u2;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - xpmem, Cell - ml_buf_ice5_2, View - schematic
// LAST TIME SAVED: Jun 14 11:22:45 2010
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_buf_ice5_2 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_rowdrv2_last, View - schematic
// LAST TIME SAVED: Aug  3 19:22:03 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_rowdrv2_last ( pgate, reset, smc_rsr_out, vddctrl, wl,
     wl_rd_sup, wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write
     );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_11_LPHVT  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
N_11_LPHVT  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
P_11_LPHVT  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));
N_11_LPRVT  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
P_11_LPRVT  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
ml_dff I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));

endmodule
// Library - xpmem, Cell - ml_rowdrvsup2, View - schematic
// LAST TIME SAVED: Aug  3 19:22:04 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_rowdrvsup2 ( wl_rd_sup, wl_rden_b );
inout  wl_rd_sup, wl_rden_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  MP15 ( .D(net045), .B(vdd_), .G(act_rd_b), .S(vdd_));
P_11_LPHVT  MP13 ( .D(wl_rden_b), .B(vdd_), .G(net059), .S(vdd_));
N_11_LPHVT  MN14 ( .D(net0158), .B(gnd_), .G(act_rd), .S(gnd_));
N_11_LPHVT  MN16 ( .D(wl_rd_sup), .B(gnd_), .G(act_rd_b), .S(gnd_));
RNPPO_LP_pcell2460 R17 ( .B(gnd_), .MINUS(net0104), .PLUS(net0110));
RNPPO_LP_pcell2460 R2 ( .B(gnd_), .MINUS(net089), .PLUS(net095));
RNPPO_LP_pcell2460 R1 ( .B(gnd_), .MINUS(net095), .PLUS(net0158));
RNPPO_LP_pcell2460 R18 ( .B(gnd_), .MINUS(wl_rd_sup), .PLUS(net0104));
RNPPO_LP_pcell2460 R7 ( .B(gnd_), .MINUS(net080), .PLUS(net092));
RNPPO_LP_pcell2460 R3 ( .B(gnd_), .MINUS(net092), .PLUS(net089));
RNPPO_LP_pcell2460 R9 ( .B(gnd_), .MINUS(net083), .PLUS(net086));
RNPPO_LP_pcell2460 R8 ( .B(gnd_), .MINUS(net086), .PLUS(net080));
RNPPO_LP_pcell2460 R10 ( .B(gnd_), .MINUS(net077), .PLUS(net083));
RNPPO_LP_pcell2460 R13 ( .B(gnd_), .MINUS(net0108), .PLUS(net0107));
RNPPO_LP_pcell2460 R11 ( .B(gnd_), .MINUS(net071), .PLUS(net077));
RNPPO_LP_pcell2460 R12 ( .B(gnd_), .MINUS(net0108), .PLUS(net071));
RNPPO_LP_pcell2460 R15 ( .B(gnd_), .MINUS(net0113), .PLUS(wl_rd_sup));
RNPPO_LP_pcell2460 R16 ( .B(gnd_), .MINUS(net0110), .PLUS(net045));
RNPPO_LP_pcell2460 R14 ( .B(gnd_), .MINUS(net0107), .PLUS(net0113));
inv_hvt I217 ( .A(wl_rden_b), .Y(net0142));
inv_hvt I220 ( .A(net0142), .Y(act_rd_b));
inv_hvt I180 ( .A(act_rd_b), .Y(act_rd));
tielo I223 ( .tielo(net059));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yp21, View - schematic
// LAST TIME SAVED: Aug  3 19:29:16 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp21 ( yp21, yp21_b_25, yp21_b_low_b, yp21_sel,
     ysup_25 );
output  yp21, yp21_b_25;

input  yp21_b_low_b, yp21_sel, ysup_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_25 I213 ( .IN(yp21_b_25_b), .OUT(yp21_b_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
nand2_hvt I206 ( .A(yp21_sel_b), .Y(net50), .B(yp21_b_low_b));
inv_hvt I207 ( .A(net50), .Y(net68));
inv_hvt I208 ( .A(yp21_sel), .Y(yp21_sel_b));
inv_hvt I209 ( .A(yp21_sel_b), .Y(yp21));
ml_ls_vdd25_nor2 I194 ( .in(net68), .sup(ysup_25),
     .out_vddio_b(yp21_b_25_b), .out_vddio(net72), .in_b(net50));

endmodule
// Library - xpmem, Cell - ml_rowdrv2, View - schematic
// LAST TIME SAVED: Aug  3 19:22:02 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_rowdrv2 ( pgate, reset, smc_rsr_out, vddctrl, wl, wl_rd_sup,
     wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_11_LPHVT  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
N_11_LPHVT  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
P_11_LPHVT  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));
N_11_LPRVT  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
P_11_LPRVT  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
ml_dff I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile_last, View - schematic
// LAST TIME SAVED: Jan 24 11:25:01 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_rowdrv_tile_last ( pgate, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  reset;
output [15:0]  wl;
output [15:0]  vddctrl;
output [15:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



nor2_hvt I211 ( .A(smc_rsr_out[15]), .Y(net049), .B(smc_rsr_inc_out));
inv_hvt I215 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I216 ( .A(net041), .Y(por_rst_buf));
inv_hvt I217 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I391 ( .A(net049), .Y(smc_rsr_inc_last));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I213 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net079));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I214 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I212 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I190 ( .A(net079), .Y(smc_rsr_1st_out));
ml_rowdrv2_last Iml_rowdrv2_last ( .smc_rsr_inc(smc_rsr_inc_last),
     .smc_rsr_in(smc_rsr_out[14]), .rsr_rst(rsr_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_rst(cram_rst_buf),
     .smc_rsr_out(smc_rsr_out[15]), .reset(reset[15]), .wl(wl[15]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile, View - schematic
// LAST TIME SAVED: Jul 30 23:15:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_rowdrv_tile ( pgate, por_rst_out, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  por_rst_out, smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  pgate;
output [15:0]  reset;
output [15:0]  wl;
output [15:0]  vddctrl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



inv_hvt I223 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I216 ( .A(cram_rst), .Y(net057));
inv_hvt I218 ( .A(net069), .Y(smc_write_buf));
inv_hvt I215 ( .A(cram_vddoff), .Y(net061));
inv_hvt I219 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I220 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I214 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I213 ( .A(smc_write), .Y(net069));
inv_hvt I221 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I212 ( .A(cram_wl_en), .Y(net055));
inv_hvt I217 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I190 ( .A(net037), .Y(smc_rsr_1st_out));
inv_hvt I211 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net037));
inv_hvt I210 ( .A(rsr_rst), .Y(net047));
inv_hvt I192 ( .A(por_rst), .Y(net041));
inv_hvt I222 ( .A(net041), .Y(por_rst_out));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I224 ( .A(net055), .Y(cram_wl_en_buf));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_15_ ( .reset(reset[15]), .wl(wl[15]),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[14]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[15]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_bank_384, View - schematic
// LAST TIME SAVED: Nov 10 15:44:55 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_rowdrv_bank_384 ( jtag_rowtest_mode_b, last_rsr, pgate,
     reset, vddctrl, wl, banksel, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst,
     smc_rsr_inc, smc_write, trst_b );
output  jtag_rowtest_mode_b, last_rsr;

input  banksel, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst, smc_rsr_inc,
     smc_write, trst_b;

output [79:0]  pgate;
output [79:0]  reset;
output [79:0]  wl;
output [79:0]  vddctrl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  smc_rsr_1st_out_buf;

wire  [3:0]  smc_rsr_inc_out;

wire  [3:0]  smc_rsr_1st_out;

wire  [4:0]  smc_rsr_out;

wire  [3:0]  por_rst_out;



tielo I252 ( .tielo(net308));
nand3_hvt I231 ( .Y(net252), .B(net256), .C(net256), .A(net256));
nand3_hvt I230 ( .Y(net256), .B(net261), .C(net261), .A(net261));
nand3_hvt I224 ( .B(net392), .Y(net261), .A(net392), .C(net392));
nand2_hvt I233 ( .A(smc_rsr_inc), .B(banksel), .Y(net269));
mux2_hvt I161 ( .in1(jtag_clk), .in0(net373), .out(net276),
     .sel(net366));
nor3_hvt I238 ( .B(por_rst), .Y(net336), .A(net304), .C(trst));
nor3_hvt I232 ( .C(rsr_rst), .A(jtag_rowtest_rst), .B(net308),
     .Y(net309));
nor3_hvt I218 ( .B(net321), .Y(net311), .A(net321), .C(net321));
nor3_hvt I220 ( .B(net311), .Y(net315), .A(net311), .C(net311));
nor3_hvt I217 ( .C(net392), .A(net392), .B(net392), .Y(net321));
nor3_hvt I244 ( .B(por_rst), .Y(net323), .A(net386),
     .C(smc_rsr_1st_out_buf[0]));
nor2_hvt I239 ( .A(jtag_rowtest_rst), .B(net336), .Y(net304));
nor2_hvt I193 ( .A(por_rst), .B(rsr_set_1st), .Y(net340));
nor2_hvt I245 ( .A(rsr_set_1st), .B(net323), .Y(net386));
inv_hvt I247 ( .A(net366), .Y(jtag_rowtest_mode_b));
inv_hvt I241 ( .A(net304), .Y(net366));
inv_hvt I192 ( .A(net309), .Y(rsr_set_1st));
inv_hvt I234 ( .A(net269), .Y(net373));
inv_hvt I35 ( .A(net374), .Y(smc_rsr_1st_out_buf[0]));
inv_hvt I240 ( .A(trst_b), .Y(trst));
inv_hvt I210 ( .A(net378), .Y(last_rsr));
inv_hvt I391 ( .A(net340), .Y(rst_row_reg));
inv_hvt I36 ( .A(smc_rsr_1st_out[0]), .Y(net374));
inv_hvt I209 ( .A(smc_rsr_out[4]), .Y(net378));
inv_hvt I205 ( .A(net386), .Y(smc_rsr_in_1st));
tiehi I269 ( .tiehi(net453));
tiehi I249 ( .tiehi(net392));
tiehi I250 ( .tiehi(net393));
ml_buf_ice5_2 I227 ( .in(net392), .o(net425), .sel(net392));
ml_buf_ice5_2 I216 ( .in(net392), .o(net428), .sel(net392));
ml_buf_ice5_2 I198 ( .sel(banksel), .in(cram_wl_en),
     .o(cram_wl_en_buf));
ml_buf_ice5_2 I196 ( .sel(banksel), .in(cram_rst), .o(cram_rst_buf));
ml_buf_ice5_2 I199 ( .sel(net393), .in(por_rst), .o(por_rst_buf));
ml_buf_ice5_2 I197 ( .sel(banksel), .in(cram_vddoff),
     .o(cram_vddoff_buf));
ml_buf_ice5_2 I195 ( .sel(banksel), .in(cram_pgateoff),
     .o(cram_pgateoff_buf));
ml_buf_ice5_2 I201 ( .sel(banksel), .in(smc_write), .o(smc_write_buf));
ml_buf_ice5_2 I203 ( .sel(net276), .in(net276), .o(smc_rsr_inc_buf));
ml_buf_ice5_2 I213 ( .in(net453), .o(net452), .sel(net453));
ml_rowdrv_tile_last I_ml_rowdrv_tile_last (
     .smc_rsr_inc_out(smc_rsr_inc_out_last), .pgate(pgate[79:64]),
     .wl(wl[79:64]), .vddctrl(vddctrl[79:64]), .reset(reset[79:64]),
     .smc_rsr_1st_out(net475), .smcc_rsr_out(smc_rsr_out[4]),
     .smc_write(smc_write_buf), .smc_rsr_inc(smc_rsr_inc_buf),
     .smc_rsr_in(smc_rsr_out[3]), .rsr_rst(rst_row_reg),
     .por_rst(por_rst_out[3]), .cram_wl_en(cram_wl_en_buf),
     .cram_vddoff(cram_vddoff_buf), .cram_rst(cram_rst_buf),
     .cram_pgateoff(cram_pgateoff_buf));
ml_rowdrv_tile I_ml_rowdrv_tile_3_ ( .por_rst_out(por_rst_out[3]),
     .smc_rsr_inc_out(smc_rsr_inc_out[3]),
     .smcc_rsr_out(smc_rsr_out[3]),
     .smc_rsr_1st_out(smc_rsr_1st_out[3]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out_last), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[2]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[63:48]), .vddctrl(vddctrl[63:48]), .reset(reset[63:48]),
     .pgate(pgate[63:48]));
ml_rowdrv_tile I_ml_rowdrv_tile_2_ ( .por_rst_out(por_rst_out[2]),
     .smc_rsr_inc_out(smc_rsr_inc_out[2]),
     .smcc_rsr_out(smc_rsr_out[2]),
     .smc_rsr_1st_out(smc_rsr_1st_out[2]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[3]), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[1]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[47:32]), .vddctrl(vddctrl[47:32]), .reset(reset[47:32]),
     .pgate(pgate[47:32]));
ml_rowdrv_tile I_ml_rowdrv_tile_1_ ( .por_rst_out(por_rst_out[1]),
     .smc_rsr_inc_out(smc_rsr_inc_out[1]),
     .smcc_rsr_out(smc_rsr_out[1]),
     .smc_rsr_1st_out(smc_rsr_1st_out[1]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[2]), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[0]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[31:16]), .vddctrl(vddctrl[31:16]), .reset(reset[31:16]),
     .pgate(pgate[31:16]));
ml_rowdrv_tile I_ml_rowdrv_tile_0_ ( .por_rst_out(por_rst_out[0]),
     .smc_rsr_inc_out(smc_rsr_inc_out[0]),
     .smcc_rsr_out(smc_rsr_out[0]),
     .smc_rsr_1st_out(smc_rsr_1st_out[0]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[1]), .smc_rsr_in(smc_rsr_in_1st),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[15:0]), .vddctrl(vddctrl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]));

endmodule
// Library - ice384chip, Cell - CHIP_route_lft_ice384, View - schematic
// LAST TIME SAVED: Nov 16 16:14:00 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module CHIP_route_lft_ice384 ( cm_banksel_bltld3_1_, cm_clk_bltld3,
     cm_sdi_u1d3, cm_sdo_u1d1, core_por_b_rowu1, cram_prec_bltld3,
     cram_pullup_bltld3, cram_write_bltld3, data_muxsel1_bltld3,
     data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     last_rsr, pgate_l, reset_l, smc_wdis_dclk_bltld3,
     smc_write_bltld3, vdd_cntl_l, wl_l, cm_banksel_blbld1,
     cm_banksel_blbld, cm_clk_blbld, cm_sdi_u1d, cm_sdo_u1,
     core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0 );
output  cm_banksel_bltld3_1_, cm_clk_bltld3, core_por_b_rowu1,
     cram_prec_bltld3, cram_pullup_bltld3, cram_write_bltld3,
     data_muxsel1_bltld3, data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     smc_wdis_dclk_bltld3, smc_write_bltld3;

input  cm_clk_blbld, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;

output [1:0]  cm_sdo_u1d1;
output [159:0]  pgate_l;
output [159:0]  wl_l;
output [1:0]  last_rsr;
output [159:0]  reset_l;
output [159:0]  vdd_cntl_l;
output [1:0]  cm_sdi_u1d3;

input [0:0]  cm_banksel_blbld1;
input [1:0]  cm_sdi_u1d;
input [1:0]  cm_sdo_u1;
input [1:1]  cm_banksel_blbld;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1d0;

wire  [1:1]  cm_banksel_bltld;

wire  [1:0]  cm_sdi_u1d0;

wire  [1:0]  dff_out;

wire  [1:0]  net299;



ml_rowdrv_bank_384 I_ml_rowdrv_bank384_bot ( .wl(wl_l[79:0]),
     .pgate(pgate_l[79:0]), .reset(reset_l[79:0]),
     .vddctrl(vdd_cntl_l[79:0]), .trst_b(j_rst_bl0),
     .smc_write(smc_writel0),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu0_b),
     .last_rsr(last_rsr[0]), .banksel(cm_banksel_blbld1[0]),
     .cram_pgateoff(cram_pgateoffl0), .cram_rst(cram_rstl0),
     .cram_vddoff(cram_vddoffl0), .cram_wl_en(cram_wl_enl0),
     .jtag_clk(tck_padl0), .jtag_rowtest_rst(row_testl1),
     .por_rst(core_por_bbl0), .rsr_rst(smc_rsr_rstl0),
     .smc_rsr_inc(smc_row_incl0));
ml_rowdrv_bank_384 I_ml_rowdrv_bank384_top ( .wl({wl_l[80], wl_l[81],
     wl_l[82], wl_l[83], wl_l[84], wl_l[85], wl_l[86], wl_l[87],
     wl_l[88], wl_l[89], wl_l[90], wl_l[91], wl_l[92], wl_l[93],
     wl_l[94], wl_l[95], wl_l[96], wl_l[97], wl_l[98], wl_l[99],
     wl_l[100], wl_l[101], wl_l[102], wl_l[103], wl_l[104], wl_l[105],
     wl_l[106], wl_l[107], wl_l[108], wl_l[109], wl_l[110], wl_l[111],
     wl_l[112], wl_l[113], wl_l[114], wl_l[115], wl_l[116], wl_l[117],
     wl_l[118], wl_l[119], wl_l[120], wl_l[121], wl_l[122], wl_l[123],
     wl_l[124], wl_l[125], wl_l[126], wl_l[127], wl_l[128], wl_l[129],
     wl_l[130], wl_l[131], wl_l[132], wl_l[133], wl_l[134], wl_l[135],
     wl_l[136], wl_l[137], wl_l[138], wl_l[139], wl_l[140], wl_l[141],
     wl_l[142], wl_l[143], wl_l[144], wl_l[145], wl_l[146], wl_l[147],
     wl_l[148], wl_l[149], wl_l[150], wl_l[151], wl_l[152], wl_l[153],
     wl_l[154], wl_l[155], wl_l[156], wl_l[157], wl_l[158],
     wl_l[159]}), .pgate({pgate_l[80], pgate_l[81], pgate_l[82],
     pgate_l[83], pgate_l[84], pgate_l[85], pgate_l[86], pgate_l[87],
     pgate_l[88], pgate_l[89], pgate_l[90], pgate_l[91], pgate_l[92],
     pgate_l[93], pgate_l[94], pgate_l[95], pgate_l[96], pgate_l[97],
     pgate_l[98], pgate_l[99], pgate_l[100], pgate_l[101],
     pgate_l[102], pgate_l[103], pgate_l[104], pgate_l[105],
     pgate_l[106], pgate_l[107], pgate_l[108], pgate_l[109],
     pgate_l[110], pgate_l[111], pgate_l[112], pgate_l[113],
     pgate_l[114], pgate_l[115], pgate_l[116], pgate_l[117],
     pgate_l[118], pgate_l[119], pgate_l[120], pgate_l[121],
     pgate_l[122], pgate_l[123], pgate_l[124], pgate_l[125],
     pgate_l[126], pgate_l[127], pgate_l[128], pgate_l[129],
     pgate_l[130], pgate_l[131], pgate_l[132], pgate_l[133],
     pgate_l[134], pgate_l[135], pgate_l[136], pgate_l[137],
     pgate_l[138], pgate_l[139], pgate_l[140], pgate_l[141],
     pgate_l[142], pgate_l[143], pgate_l[144], pgate_l[145],
     pgate_l[146], pgate_l[147], pgate_l[148], pgate_l[149],
     pgate_l[150], pgate_l[151], pgate_l[152], pgate_l[153],
     pgate_l[154], pgate_l[155], pgate_l[156], pgate_l[157],
     pgate_l[158], pgate_l[159]}), .reset({reset_l[80], reset_l[81],
     reset_l[82], reset_l[83], reset_l[84], reset_l[85], reset_l[86],
     reset_l[87], reset_l[88], reset_l[89], reset_l[90], reset_l[91],
     reset_l[92], reset_l[93], reset_l[94], reset_l[95], reset_l[96],
     reset_l[97], reset_l[98], reset_l[99], reset_l[100], reset_l[101],
     reset_l[102], reset_l[103], reset_l[104], reset_l[105],
     reset_l[106], reset_l[107], reset_l[108], reset_l[109],
     reset_l[110], reset_l[111], reset_l[112], reset_l[113],
     reset_l[114], reset_l[115], reset_l[116], reset_l[117],
     reset_l[118], reset_l[119], reset_l[120], reset_l[121],
     reset_l[122], reset_l[123], reset_l[124], reset_l[125],
     reset_l[126], reset_l[127], reset_l[128], reset_l[129],
     reset_l[130], reset_l[131], reset_l[132], reset_l[133],
     reset_l[134], reset_l[135], reset_l[136], reset_l[137],
     reset_l[138], reset_l[139], reset_l[140], reset_l[141],
     reset_l[142], reset_l[143], reset_l[144], reset_l[145],
     reset_l[146], reset_l[147], reset_l[148], reset_l[149],
     reset_l[150], reset_l[151], reset_l[152], reset_l[153],
     reset_l[154], reset_l[155], reset_l[156], reset_l[157],
     reset_l[158], reset_l[159]}), .vddctrl({vdd_cntl_l[80],
     vdd_cntl_l[81], vdd_cntl_l[82], vdd_cntl_l[83], vdd_cntl_l[84],
     vdd_cntl_l[85], vdd_cntl_l[86], vdd_cntl_l[87], vdd_cntl_l[88],
     vdd_cntl_l[89], vdd_cntl_l[90], vdd_cntl_l[91], vdd_cntl_l[92],
     vdd_cntl_l[93], vdd_cntl_l[94], vdd_cntl_l[95], vdd_cntl_l[96],
     vdd_cntl_l[97], vdd_cntl_l[98], vdd_cntl_l[99], vdd_cntl_l[100],
     vdd_cntl_l[101], vdd_cntl_l[102], vdd_cntl_l[103],
     vdd_cntl_l[104], vdd_cntl_l[105], vdd_cntl_l[106],
     vdd_cntl_l[107], vdd_cntl_l[108], vdd_cntl_l[109],
     vdd_cntl_l[110], vdd_cntl_l[111], vdd_cntl_l[112],
     vdd_cntl_l[113], vdd_cntl_l[114], vdd_cntl_l[115],
     vdd_cntl_l[116], vdd_cntl_l[117], vdd_cntl_l[118],
     vdd_cntl_l[119], vdd_cntl_l[120], vdd_cntl_l[121],
     vdd_cntl_l[122], vdd_cntl_l[123], vdd_cntl_l[124],
     vdd_cntl_l[125], vdd_cntl_l[126], vdd_cntl_l[127],
     vdd_cntl_l[128], vdd_cntl_l[129], vdd_cntl_l[130],
     vdd_cntl_l[131], vdd_cntl_l[132], vdd_cntl_l[133],
     vdd_cntl_l[134], vdd_cntl_l[135], vdd_cntl_l[136],
     vdd_cntl_l[137], vdd_cntl_l[138], vdd_cntl_l[139],
     vdd_cntl_l[140], vdd_cntl_l[141], vdd_cntl_l[142],
     vdd_cntl_l[143], vdd_cntl_l[144], vdd_cntl_l[145],
     vdd_cntl_l[146], vdd_cntl_l[147], vdd_cntl_l[148],
     vdd_cntl_l[149], vdd_cntl_l[150], vdd_cntl_l[151],
     vdd_cntl_l[152], vdd_cntl_l[153], vdd_cntl_l[154],
     vdd_cntl_l[155], vdd_cntl_l[156], vdd_cntl_l[157],
     vdd_cntl_l[158], vdd_cntl_l[159]}), .smc_write(smc_write_bltld3),
     .smc_rsr_inc(net303), .rsr_rst(net289),
     .por_rst(core_por_b_rowu1), .jtag_rowtest_rst(net345),
     .jtag_clk(net305), .cram_wl_en(net273), .cram_vddoff(net335),
     .cram_rst(net319), .cram_pgateoff(net295),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu1_b),
     .last_rsr(last_rsr[1]), .banksel(net231), .trst_b(net311));
tielo I74 ( .tielo(net219));
sg_bufx10_ice8p I28 ( .in(smc_writel0), .out(net221));
sg_bufx10_ice8p I35 ( .in(net291), .out(net223));
sg_bufx10_ice8p I45 ( .in(row_testl1), .out(net225));
sg_bufx10_ice8p I44 ( .in(net225), .out(net227));
sg_bufx10_ice8p I2 ( .in(cram_write_bltld), .out(net229));
sg_bufx10_ice8p I67 ( .in(cm_banksel_bltld[1]), .out(net231));
sg_bufx10_ice8p I39 ( .in(net237), .out(net233));
sg_bufx10_ice8p I4 ( .in(data_muxsel1_blbld),
     .out(data_muxsel1_bltld));
sg_bufx10_ice8p I40 ( .in(cram_wl_enl0), .out(net237));
sg_bufx10_ice8p I37 ( .in(cram_vddoffl0), .out(net239));
sg_bufx10_ice8p I22 ( .in(core_por_bbl0), .out(net241));
sg_bufx10_ice8p I5 ( .in(data_muxsel1_bltld), .out(net243));
sg_bufx10_ice8p I527 ( .in(net327), .out(en_8bconfig_b_bltld3));
sg_bufx10_ice8p I523 ( .in(net283), .out(data_muxsel_bltld3));
sg_bufx10_ice8p I524 ( .in(net243), .out(data_muxsel1_bltld3));
sg_bufx10_ice8p I526 ( .in(net343), .out(cram_prec_bltld3));
sg_bufx10_ice8p I33 ( .in(cram_rstl0), .out(net253));
sg_bufx10_ice8p I70_1_ ( .in(cm_sdo_u1[1]), .out(cm_sdo_u1d0[1]));
sg_bufx10_ice8p I70_0_ ( .in(cm_sdo_u1[0]), .out(cm_sdo_u1d0[0]));
sg_bufx10_ice8p I528 ( .in(net337), .out(smc_wdis_dclk_bltld3));
sg_bufx10_ice8p I18 ( .in(smc_rsr_rstl0), .out(net259));
sg_bufx10_ice8p I529 ( .in(net293), .out(cram_pullup_bltld3));
sg_bufx10_ice8p I3 ( .in(cram_write_blbld), .out(cram_write_bltld));
sg_bufx10_ice8p I532 ( .in(net363), .out(cm_clk_bltld3));
sg_bufx10_ice8p I79 ( .in(cm_clk_blbld), .out(cm_clk_bltld));
sg_bufx10_ice8p I8 ( .in(cram_pullup_blbld), .out(cram_pullup_bltld));
sg_bufx10_ice8p I7 ( .in(data_muxsel_blbld), .out(data_muxsel_bltld));
sg_bufx10_ice8p I554 ( .in(net233), .out(net273));
sg_bufx10_ice8p I27 ( .in(net221), .out(net275));
sg_bufx10_ice8p I25 ( .in(smc_row_incl0), .out(net277));
sg_bufx10_ice8p I47 ( .in(net357), .out(net279));
sg_bufx10_ice8p I68_1_ ( .in(cm_sdi_u1d[1]), .out(cm_sdi_u1d0[1]));
sg_bufx10_ice8p I68_0_ ( .in(cm_sdi_u1d[0]), .out(cm_sdi_u1d0[0]));
sg_bufx10_ice8p I6 ( .in(data_muxsel_bltld), .out(net283));
sg_bufx10_ice8p I38 ( .in(net239), .out(net285));
sg_bufx10_ice8p I19 ( .in(net259), .out(net287));
sg_bufx10_ice8p I546 ( .in(net287), .out(net289));
sg_bufx10_ice8p I36 ( .in(cram_pgateoffl0), .out(net291));
sg_bufx10_ice8p I9 ( .in(cram_pullup_bltld), .out(net293));
sg_bufx10_ice8p I547 ( .in(net223), .out(net295));
sg_bufx10_ice8p I552 ( .in(net275), .out(smc_write_bltld3));
sg_bufx10_ice8p I69_1_ ( .in(cm_sdi_u1d0[1]), .out(net299[0]));
sg_bufx10_ice8p I69_0_ ( .in(cm_sdi_u1d0[0]), .out(net299[1]));
sg_bufx10_ice8p I549 ( .in(net349), .out(net303));
sg_bufx10_ice8p I544 ( .in(net279), .out(net305));
sg_bufx10_ice8p I530_1_ ( .in(net299[0]), .out(cm_sdi_u1d3[1]));
sg_bufx10_ice8p I530_0_ ( .in(net299[1]), .out(cm_sdi_u1d3[0]));
sg_bufx10_ice8p I545 ( .in(net353), .out(net311));
sg_bufx10_ice8p I531 ( .in(net231), .out(cm_banksel_bltld3_1_));
sg_bufx10_ice8p I551 ( .in(net331), .out(net319));
sg_bufx10_ice8p I553 ( .in(net355), .out(core_por_b_rowu1));
sg_bufx10_ice8p I81 ( .in(cm_clk_bltld), .out(net363));
sg_bufx10_ice8p I15 ( .in(en_8bconfig_b_blbld),
     .out(en_8bconfig_b_bltld));
sg_bufx10_ice8p I14 ( .in(en_8bconfig_b_bltld), .out(net327));
sg_bufx10_ice8p I0 ( .in(cram_prec_blbld), .out(cram_prec_bltld));
sg_bufx10_ice8p I34 ( .in(net253), .out(net331));
sg_bufx10_ice8p I49 ( .in(j_rst_bl0), .out(net333));
sg_bufx10_ice8p I550 ( .in(net285), .out(net335));
sg_bufx10_ice8p I13 ( .in(smc_wdis_dclk_bltld), .out(net337));
sg_bufx10_ice8p I66 ( .in(cm_banksel_blbld[1]),
     .out(cm_banksel_bltld[1]));
sg_bufx10_ice8p I80_1_ ( .in(dff_out[1]), .out(cm_sdo_u1d1[1]));
sg_bufx10_ice8p I80_0_ ( .in(dff_out[0]), .out(cm_sdo_u1d1[0]));
sg_bufx10_ice8p I1 ( .in(cram_prec_bltld), .out(net343));
sg_bufx10_ice8p I548 ( .in(net227), .out(net345));
sg_bufx10_ice8p I525 ( .in(net229), .out(cram_write_bltld3));
sg_bufx10_ice8p I26 ( .in(net277), .out(net349));
sg_bufx10_ice8p I12 ( .in(smc_wdis_dclk_blbld),
     .out(smc_wdis_dclk_bltld));
sg_bufx10_ice8p I48 ( .in(net333), .out(net353));
sg_bufx10_ice8p I21 ( .in(net241), .out(net355));
sg_bufx10_ice8p I46 ( .in(tck_padl0), .out(net357));
sg_dffbuf_modified I73_1_ ( .d(cm_sdo_u1d0[1]), .clk(net363),
     .dffout(dff_out[1]), .r(net219));
sg_dffbuf_modified I73_0_ ( .d(cm_sdo_u1d0[0]), .clk(net363),
     .dffout(dff_out[0]), .r(net219));
sg_dffbuf_modified I77 ( .d(last_rsr[0]), .clk(net363),
     .dffout(last_rsr0), .r(net219));

endmodule
// Library - leafcell, Cell - bram_bufferx4, View - schematic
// LAST TIME SAVED: Aug 12 09:08:27 2010
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module bram_bufferx4 ( out, in );
output  out;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - creset_filter, View - schematic
// LAST TIME SAVED: Nov 18 18:04:19 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module creset_filter ( out, in );
output  out;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M2 ( .D(net13), .B(vdd_), .G(pbias), .S(vdd_));
P_11_LPHVT  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(vdd_));
P_11_LPHVT  M3 ( .D(net13), .B(vdd_), .G(net042), .S(vdd_));
P_11_LPHVT  M1 ( .D(vdd_), .B(vdd_), .G(net13), .S(vdd_));
P_11_LPHVT  MP41 ( .D(pbias), .B(vdd_), .G(net9), .S(vdd_));
RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(net17), .PLUS(pbias));
N_11_LPHVT  M0 ( .D(net13), .B(gnd_), .G(in), .S(gnd_));
N_11_LPHVT  MN31 ( .D(net17), .B(gnd_), .G(net9), .S(gnd_));
bram_bufferx4 I11 ( .in(net042), .out(out));
inv_hvt I6 ( .A(net13), .Y(net042));
inv_hvt I4 ( .A(in), .Y(net9));

endmodule
// Library - ice8chip, Cell - eh_core_pup_2, View - schematic
// LAST TIME SAVED: Jan  7 13:56:08 2012
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module eh_core_pup_2 ( por_b );
output  por_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



RNPPO_LP_pcell2460 RR16 ( .B(gnd_), .MINUS(vdd_), .PLUS(net0108));
RNPPO_LP_pcell2460 R12 ( .B(gnd_), .MINUS(net154), .PLUS(net157));
RNPPO_LP_pcell2460 R6 ( .B(gnd_), .MINUS(out_1), .PLUS(net124));
RNPPO_LP_pcell2460 R9 ( .B(gnd_), .MINUS(net118), .PLUS(net130));
RNPPO_LP_pcell2460 R15 ( .B(gnd_), .MINUS(net166), .PLUS(div_1));
RNPPO_LP_pcell2460 R13 ( .B(gnd_), .MINUS(net157), .PLUS(net145));
RNPPO_LP_pcell2460 R1 ( .B(gnd_), .MINUS(net068), .PLUS(net048));
RNPPO_LP_pcell2460 R2 ( .B(gnd_), .MINUS(net0145), .PLUS(net068));
RNPPO_LP_pcell2460 R4 ( .B(gnd_), .MINUS(net142), .PLUS(net079));
RNPPO_LP_pcell2460 R5 ( .B(gnd_), .MINUS(div_1), .PLUS(net142));
RNPPO_LP_pcell2460 R41 ( .B(gnd_), .MINUS(net039), .PLUS(net042));
RNPPO_LP_pcell2460 R40 ( .B(gnd_), .MINUS(net042), .PLUS(vdd_));
RNPPO_LP_pcell2460 R11 ( .B(gnd_), .MINUS(net109), .PLUS(net154));
RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(net048), .PLUS(net039));
RNPPO_LP_pcell2460 R10 ( .B(gnd_), .MINUS(net130), .PLUS(net109));
RNPPO_LP_pcell2460 R8 ( .B(gnd_), .MINUS(net127), .PLUS(net118));
RNPPO_LP_pcell2460 R14 ( .B(gnd_), .MINUS(net145), .PLUS(net166));
RNPPO_LP_pcell2460 R3 ( .B(gnd_), .MINUS(net079), .PLUS(net0145));
RNPPO_LP_pcell2460 R7 ( .B(gnd_), .MINUS(net124), .PLUS(net127));
N_11_LPHVT  M7 ( .D(net049), .B(gnd_), .G(net157), .S(gnd_));
N_11_LPHVT  M0 ( .D(net057), .B(gnd_), .G(net157), .S(gnd_));
N_11_LPHVT  M6 ( .D(net053), .B(gnd_), .G(net157), .S(gnd_));
N_11_LPHVT  M3 ( .D(gnd_), .B(gnd_), .G(out_2), .S(gnd_));
N_11_LPHVT  M1 ( .D(out_1), .B(gnd_), .G(out_2), .S(gnd_));
N_25_LP  M22 ( .D(out_1), .B(gnd_), .G(net048), .S(gnd_));
inv_hvt I7 ( .A(out_1), .Y(out_2));
inv_hvt I9 ( .A(out_2), .Y(out_3));
inv_hvt I11 ( .A(out_3), .Y(por_b));

endmodule
// Library - ice8chip, Cell - SMC_CORE_POR_right_ice8p, View -
//schematic
// LAST TIME SAVED: Sep 29 09:25:02 2010
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module SMC_CORE_POR_right_ice8p ( core_por_b0, core_por_bb, smc_por_b,
     creset_b, smc_core_por_bottom1, smc_core_por_bottom2,
     vddio_rightbank );
output  core_por_b0, core_por_bb, smc_por_b;

input  creset_b, smc_core_por_bottom1, smc_core_por_bottom2,
     vddio_rightbank;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



sg_bufx10_ice8p I500 ( .in(net032), .out(core_por_bb));
eh_io_pup_2_new_ice8p Ieh_io_pup_2_new_ice8p ( .core_por_b(net026),
     .vdd_io(vddio_rightbank), .por_b(net3));
eh_core_pup_2 Ieh_core_pup_2 ( .por_b(net026));
nand2_hvt I6 ( .A(net026), .Y(net021), .B(creset_b));
inv_hvt I11 ( .A(net04), .Y(smc_por_b));
inv_hvt I701 ( .A(core_por_b0), .Y(net032));
inv_hvt I7 ( .A(net021), .Y(core_por_b0));
nand4_hvt I2 ( .D(core_por_b0), .C(smc_core_por_bottom2), .A(net3),
     .Y(net04), .B(smc_core_por_bottom1));

endmodule
// Library - ice8chip, Cell - ml_cram_logic_ice8p, View - schematic
// LAST TIME SAVED: Aug  3 19:20:07 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_cram_logic_ice8p ( cram_pgateoff, cram_prec, cram_pullup_b,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, smc_clk_out, por,
     smc_clk, smc_read, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rwl_en, smc_seq_rst, smc_wcram_rst, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en );
output  cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, smc_clk_out;

input  por, smc_clk, smc_read, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_write, smc_wset_prec, smc_wset_precgnd, smc_wwlwrt_dis,
     smc_wwlwrt_en;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



NCAP_25_LP  C2 ( .MINUS(GND_), .PLUS(net326));
NCAP_25_LP  C1 ( .MINUS(GND_), .PLUS(net306));
NCAP_25_LP  C0 ( .MINUS(GND_), .PLUS(net314));
tielo I480 ( .tielo(net235));
sg_bufx10_ice8p I461 ( .in(net321), .out(cram_pullup_b));
sg_bufx10_ice8p I446 ( .in(net245), .out(cram_prec));
sg_bufx10_ice8p I457 ( .in(net234), .out(cram_wl_en));
sg_bufx10_ice8p I467 ( .in(net226), .out(cram_pgateoff));
sg_bufx10_ice8p I447 ( .in(cram_write_int), .out(cram_write));
sg_bufx10_ice8p I526 ( .in(net295), .out(cram_vddoff));
nand2_hvt I213 ( .A(net285), .Y(net222), .B(net311));
mux2_hvt I430 ( .in1(net407), .in0(net254), .out(net226),
     .sel(net235));
mux2_hvt I428 ( .in1(cram_write_int), .in0(net319), .out(net230),
     .sel(net285));
mux2_hvt I429 ( .in1(net254), .in0(net230), .out(net234),
     .sel(net235));
mux2_hvt I295 ( .in1(net255), .in0(net293), .out(net238),
     .sel(net285));
nor2_hvt I402 ( .A(net240), .B(smc_wset_precgnd), .Y(net242));
nor2_hvt I329 ( .A(net287), .B(smc_seq_rst), .Y(net245));
nor2_hvt I398 ( .A(smc_rpull_b), .B(net247), .Y(net248));
nor2_hvt I393 ( .A(set_wl_write), .B(reset_logic), .Y(net251));
nor2_hvt I364 ( .A(net426), .B(smc_seq_rst), .Y(net254));
nor2_hvt I400 ( .A(net255), .B(smc_wset_prec), .Y(net257));
nor2_hvt I366 ( .A(reset_logic), .B(net417), .Y(net260));
nor2_hvt I223 ( .A(net359), .B(por), .Y(net263));
nor2_hvt I390 ( .A(smc_write), .B(smc_seq_rst), .Y(net266));
nor2_hvt I392 ( .A(net240), .B(cram_rst), .Y(net269));
nor2_hvt I389 ( .A(net442), .B(reset_logic), .Y(net272));
nor2_hvt I385 ( .A(smc_rprec), .B(net274), .Y(net368));
nor2_hvt I414 ( .A(net276), .B(smc_wwlwrt_en), .Y(net278));
nor2_hvt I391 ( .A(cram_rst), .B(reset_logic), .Y(net281));
inv_hvt I458 ( .A(net272), .Y(rst_rpull_rwl));
inv_hvt I452 ( .A(net266), .Y(net285));
inv_hvt I451 ( .A(net238), .Y(net287));
inv_hvt I459 ( .A(smc_rwl_en), .Y(net289));
inv_hvt I373 ( .A(set_wl_write), .Y(net314));
inv_hvt I346 ( .A(net368), .Y(net293));
inv_hvt I464 ( .A(net222), .Y(net295));
inv_hvt I468 ( .A(net456), .Y(net297));
inv_hvt I454 ( .A(net260), .Y(dis_pgatewrt));
inv_hvt I403 ( .A(net242), .Y(net444));
inv_hvt I450 ( .A(net257), .Y(net303));
inv_hvt I448 ( .A(net281), .Y(net443));
inv_hvt I442 ( .A(net306), .Y(net307));
inv_hvt I444 ( .A(net315), .Y(net306));
inv_hvt I453 ( .A(net269), .Y(net311));
inv_hvt I445 ( .A(net307), .Y(net326));
inv_hvt I435 ( .A(net314), .Y(net315));
inv_hvt I4 ( .A(sm_clk_b), .Y(smc_clk_out));
inv_hvt I421 ( .A(net421), .Y(net319));
inv_hvt I462 ( .A(net247), .Y(net321));
inv_hvt I3 ( .A(smc_clk), .Y(sm_clk_b));
inv_hvt I449 ( .A(net251), .Y(net325));
inv_hvt I443 ( .A(net326), .Y(cram_write_int));
inv_hvt I465 ( .A(cram_rst_int_b), .Y(cram_rst));
inv_hvt I456 ( .A(net263), .Y(reset_logic));
inv_hvt I463 ( .A(net451), .Y(net247));
inv_hvt I460 ( .A(net248), .Y(net335));
inv_hvt I466 ( .A(net297), .Y(cram_rst_int_b));
inv_hvt I256 ( .A(net436), .Y(set_wl_write));
inv_hvt I455 ( .A(net278), .Y(net341));
nor3_hvt I472 ( .B(net347), .Y(net343), .A(net347), .C(net347));
nor3_hvt I471 ( .B(net351), .Y(net347), .A(net351), .C(net351));
nor3_hvt I470 ( .B(net363), .Y(net351), .A(net363), .C(net363));
nor3_hvt I217 ( .B(vdd_tieh), .Y(net355), .A(vdd_tieh), .C(vdd_tieh));
nor3_hvt I386 ( .B(smc_seq_rst), .Y(net359), .A(smc_write),
     .C(smc_read));
nor3_hvt I469 ( .B(net355), .Y(net363), .A(net355), .C(net355));
nor3_hvt I387 ( .B(smc_rwl_en), .Y(net274), .A(net368),
     .C(reset_logic));
nand3_hvt I476 ( .Y(net370), .B(net386), .C(net386), .A(net386));
nand3_hvt I477 ( .Y(net374), .B(net370), .C(net370), .A(net370));
nand3_hvt I478 ( .Y(net378), .B(net374), .C(net374), .A(net374));
nand3_hvt I479 ( .Y(net382), .B(net378), .C(net378), .A(net378));
nand3_hvt I426 ( .Y(net386), .B(vdd_tieh), .C(vdd_tieh), .A(vdd_tieh));
ml_dff I432 ( .R(dis_pgatewrt), .D(net412), .CLK(smc_clk_out),
     .QN(net406), .Q(net407));
ml_dff I431 ( .R(dis_pgatewrt), .D(net254), .CLK(sm_clk_b),
     .QN(net411), .Q(net412));
ml_dff I411 ( .R(reset_logic), .D(smc_wwlwrt_dis), .CLK(smc_clk),
     .QN(net416), .Q(net417));
ml_dff I408 ( .R(rst_rpull_rwl), .D(vdd_tieh), .CLK(net289),
     .QN(net421), .Q(net400));
ml_dff I405 ( .R(dis_pgatewrt), .D(vdd_tieh), .CLK(set_wl_write),
     .QN(net426), .Q(net399));
ml_dff I412 ( .R(net325), .D(net303), .CLK(smc_clk_out), .QN(net394),
     .Q(net255));
ml_dff I410 ( .R(dis_pgatewrt), .D(net341), .CLK(smc_clk_out),
     .QN(net436), .Q(net276));
ml_dff I108 ( .R(reset_logic), .D(smc_rrst_pullwlen),
     .CLK(smc_clk_out), .QN(net402), .Q(net442));
ml_dff I413 ( .R(net443), .D(net444), .CLK(smc_clk_out), .QN(net446),
     .Q(net240));
ml_dff I407 ( .R(rst_rpull_rwl), .D(net335), .CLK(smc_clk_out),
     .QN(net451), .Q(net397));
ml_dff I406 ( .R(reset_logic), .D(smc_wcram_rst), .CLK(smc_clk_out),
     .QN(net456), .Q(net457));
tiehi I427 ( .tiehi(vdd_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_vblinhi_pgm_drv, View -
//schematic
// LAST TIME SAVED: Aug  3 19:29:17 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_vblinhi_pgm_drv ( vblinhi_pgm_25, ysup_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25 );
inout  vblinhi_pgm_25, ysup_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(net10), .B(vblinhi_pgm_25), .G(en_blinhi_pgm_b),
     .S(vblinhi_pgm_25));
P_25_LP  M5 ( .D(net10), .B(ysup_25), .G(en_blinhi_pgm_b_ysup_25),
     .S(ysup_25));
N_25_LPNVT  M13 ( .D(vdd_), .B(GND_), .G(en_blinhi_pgm_b_ysup_25),
     .S(vblinhi_pgm_25));

endmodule
// Library - xpmem, Cell - ml_dff_osc, View - schematic
// LAST TIME SAVED: Jul 30 23:15:05 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_dff_osc ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - misc, Cell - ml_mux3_hvt, View - schematic
// LAST TIME SAVED: Aug  3 19:21:11 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_mux3_hvt ( out, in0, in1, in2, sel );
output  out;

input  in0, in1, in2;

input [3:0]  sel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_11_LPHVT  MN19 ( .D(out), .B(gnd_), .G(sel[3]), .S(gnd_));
inv_hvt I21 ( .A(sel[0]), .Y(net30));
inv_hvt I24 ( .A(sel[1]), .Y(net28));
inv_hvt I25 ( .A(sel[2]), .Y(net26));
txgate_hvt I23 ( .in(in1), .out(out), .pp(net28), .nn(sel[1]));
txgate_hvt I20 ( .in(in0), .out(out), .pp(net30), .nn(sel[0]));
txgate_hvt I26 ( .in(in2), .out(out), .pp(net26), .nn(sel[2]));

endmodule
// Library - misc, Cell - ml_osc_stage, View - schematic
// LAST TIME SAVED: Aug  3 19:21:12 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_osc_stage ( out, clkin, oscen_b, pbias, sel_trim );
output  out;

input  clkin, oscen_b, pbias;

input [3:0]  sel_trim;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M2 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net452));
P_11_LPHVT  MP30 ( .D(net452), .B(vdd_), .G(oscen_b), .S(vdd_));
P_11_LPHVT  MP72 ( .D(net456), .B(vdd_), .G(sel_trim[2]), .S(net452));
P_11_LPHVT  MP33 ( .D(out), .B(vdd_), .G(in_bot), .S(vdd_));
P_11_LPHVT  M3 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net456));
N_11_LPHVT  MN41 ( .D(loadbot_0), .B(gnd_), .G(net419), .S(gnd_));
N_11_LPHVT  MN39 ( .D(loadbot_2), .B(gnd_), .G(net419), .S(gnd_));
N_11_LPHVT  MN29 ( .D(out), .B(gnd_), .G(in_bot), .S(gnd_));
N_11_LPHVT  MN42 ( .D(loadbot_1), .B(gnd_), .G(net419), .S(gnd_));
NCAP_25_LP  C5 ( .MINUS(gnd_), .PLUS(loadbot_0));
NCAP_25_LP  C6 ( .MINUS(gnd_), .PLUS(loadbot_1));
NCAP_25_LP  C4 ( .MINUS(gnd_), .PLUS(loadbot_2));
inv_hvt I229 ( .A(net403), .Y(net419));
nor2_hvt I228 ( .A(clkin), .B(oscen_b), .Y(net403));
ml_mux3_hvt Iml_mux3_hvt_bot ( .in1(loadbot_1), .in0(loadbot_0),
     .out(in_bot), .sel(sel_trim[3:0]), .in2(loadbot_2));

endmodule
// Library - misc, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_mux2_hvt ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - misc, Cell - ml_osc_logic, View - schematic
// LAST TIME SAVED: Oct  7 11:48:52 2010
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_osc_logic ( sel_trim, clkin, smc_osc_fsel, smc_oscen );

input  clkin, smc_oscen;

output [3:0]  sel_trim;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:1]  in_sel;



ml_dff_osc I174 ( .R(reset_ff), .D(net050), .CLK(clkin_buf_b),
     .QN(net150), .Q(net172));
ml_dff_osc I238 ( .R(reset_ff), .D(net050), .CLK(clkin_buf),
     .QN(net154), .Q(net177));
ml_dff_osc I244 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf),
     .QN(net155), .Q(net182));
ml_dff_osc I245 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf_b),
     .QN(net153), .Q(net187));
ml_dff_osc I242 ( .R(reset_ff), .D(net048), .CLK(clkin_buf_b),
     .QN(net191), .Q(net192));
ml_dff_osc I243 ( .R(reset_ff), .D(net048), .CLK(clkin_buf),
     .QN(net152), .Q(net197));
nor2_hvt I256 ( .A(smc_osc_fsel[1]), .B(smc_osc_fsel[0]),
     .Y(in_sel[2]));
inv_hvt I293 ( .A(net197), .Y(net052));
inv_hvt I263 ( .A(clkin_buf), .Y(net065));
inv_hvt I283 ( .A(clkin_buf_b), .Y(clkin_buf));
inv_hvt I284 ( .A(smc_oscen), .Y(reset_ff));
inv_hvt I282 ( .A(clkin), .Y(clkin_buf_b));
inv_hvt I255 ( .A(smc_osc_fsel[1]), .Y(in_sel[1]));
inv_hvt I294 ( .A(net192), .Y(net054));
inv_hvt I295 ( .A(net177), .Y(net057));
inv_hvt I296 ( .A(net172), .Y(net061));
inv_hvt I261 ( .A(in_sel[2]), .Y(net050));
inv_hvt I262 ( .A(in_sel[1]), .Y(net048));
inv_hvt I299 ( .A(net059), .Y(net0143));
inv_hvt I297 ( .A(net065), .Y(net063));
inv_hvt I302 ( .A(net094), .Y(net096));
inv_hvt I298 ( .A(net063), .Y(net059));
inv_hvt I304 ( .A(net0143), .Y(net092));
inv_hvt I303 ( .A(net092), .Y(net094));
inv_hvt I301 ( .A(net096), .Y(clkin_buf_delay));
inv_hvt I285 ( .A(net058), .Y(sel_trim[3]));
tiehis I281 ( .tiehi(net058));
ml_mux2_hvt I279 ( .in1(net182), .in0(net187), .out(sel_trim[0]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I277 ( .in1(net057), .in0(net061), .out(sel_trim[2]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I278 ( .in1(net052), .in0(net054), .out(sel_trim[1]),
     .sel(clkin_buf_delay));

endmodule
// Library - misc, Cell - ml_osc, View - schematic
// LAST TIME SAVED: Sep 24 14:35:17 2011
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_osc ( clk_out, smc_osc_fsel, smc_oscen );
output  clk_out;

input  smc_oscen;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sel_trim;



P_11_LPHVT  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(net0101));
P_11_LPHVT  MP41 ( .D(pbias), .B(vdd_), .G(smc_oscen), .S(vdd_));
P_11_LPHVT  M0 ( .D(net0101), .B(vdd_), .G(oscen_b), .S(vdd_));
N_11_LPHVT  MN31 ( .D(net437), .B(gnd_), .G(smc_oscen), .S(gnd_));
RNPPO_LP_pcell2460 R1 ( .B(gnd_), .MINUS(net437), .PLUS(net383));
RNPPO_LP_pcell2460 R18 ( .B(gnd_), .MINUS(net437), .PLUS(net437));
RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(net437), .PLUS(net437));
RNPPO_LP_pcell2460 R3 ( .B(gnd_), .MINUS(net366), .PLUS(net076));
RNPPO_LP_pcell2460 R2 ( .B(gnd_), .MINUS(net383), .PLUS(net366));
RNPPO_LP_pcell2460 R5 ( .B(gnd_), .MINUS(net070), .PLUS(pbias));
RNPPO_LP_pcell2460 R4 ( .B(gnd_), .MINUS(net076), .PLUS(net070));
ml_dff_osc I174 ( .R(oscen_b), .D(clkby2_b), .CLK(clk_dffin),
     .QN(clkby2_b), .Q(clkby2));
ml_dff_osc I279 ( .R(oscen_b), .D(net063), .CLK(net0115), .QN(net063),
     .Q(net066));
nand2_hvt I175 ( .A(out_bot), .Y(clk_dffin), .B(out_top));
inv_hvt I280 ( .A(clkby2), .Y(net0115));
inv_hvt I222 ( .A(clkby2), .Y(clkby2_b_buf));
inv_hvt I220 ( .A(clkby2_b), .Y(clkby2_buf));
inv_hvt I176 ( .A(net063), .Y(clk_out));
inv_hvt I198 ( .A(smc_oscen), .Y(oscen_b));
ml_osc_stage Istage_bot ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_b_buf), .out(out_bot), .sel_trim(sel_trim[3:0]));
ml_osc_stage Istage_top ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_buf), .out(out_top), .sel_trim(sel_trim[3:0]));
ml_osc_logic Iosc_logic ( .sel_trim(sel_trim[3:0]),
     .smc_oscen(smc_oscen), .smc_osc_fsel(smc_osc_fsel[1:0]),
     .clkin(clk_out));

endmodule
// Library - misc, Cell - ml_osc_top, View - schematic
// LAST TIME SAVED: Oct 13 10:43:19 2010
// NETLIST TIME: Jan 18 18:48:18 2012
`timescale 1ns / 1ns 

module ml_osc_top ( cnt_podt_out, smc_clk, crst_b, por_b, smc_osc_fsel,
     smc_oscoff_b, smc_podt_off, smc_podt_rst );
output  cnt_podt_out, smc_clk;

input  crst_b, por_b, smc_oscoff_b, smc_podt_off, smc_podt_rst;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  q_b;

wire  [10:0]  q;



ml_dff_osc I230 ( .R(cnt_rst), .D(net076), .CLK(q_b[10]), .QN(net067),
     .Q(net063));
ml_dff_osc I243 ( .R(rst_off_latch), .D(net0174), .CLK(clk_out_b),
     .QN(smc_off_b), .Q(net0152));
ml_dff_osc I228_10_ ( .R(cnt_rst), .D(q_b[10]), .CLK(q[9]),
     .QN(q_b[10]), .Q(q[10]));
ml_dff_osc I228_9_ ( .R(cnt_rst), .D(q_b[9]), .CLK(q[8]), .QN(q_b[9]),
     .Q(q[9]));
ml_dff_osc I228_8_ ( .R(cnt_rst), .D(q_b[8]), .CLK(q[7]), .QN(q_b[8]),
     .Q(q[8]));
ml_dff_osc I228_7_ ( .R(cnt_rst), .D(q_b[7]), .CLK(q[6]), .QN(q_b[7]),
     .Q(q[7]));
ml_dff_osc I228_6_ ( .R(cnt_rst), .D(q_b[6]), .CLK(q[5]), .QN(q_b[6]),
     .Q(q[6]));
ml_dff_osc I228_5_ ( .R(cnt_rst), .D(q_b[5]), .CLK(q[4]), .QN(q_b[5]),
     .Q(q[5]));
ml_dff_osc I228_4_ ( .R(cnt_rst), .D(q_b[4]), .CLK(q[3]), .QN(q_b[4]),
     .Q(q[4]));
ml_dff_osc I228_3_ ( .R(cnt_rst), .D(q_b[3]), .CLK(q[2]), .QN(q_b[3]),
     .Q(q[3]));
ml_dff_osc I228_2_ ( .R(cnt_rst), .D(q_b[2]), .CLK(q[1]), .QN(q_b[2]),
     .Q(q[2]));
ml_dff_osc I228_1_ ( .R(cnt_rst), .D(q_b[1]), .CLK(q[0]), .QN(q_b[1]),
     .Q(q[1]));
ml_dff_osc I228_0_ ( .R(cnt_rst), .D(q_b[0]), .CLK(clk_in),
     .QN(q_b[0]), .Q(q[0]));
nand2_hvt I227 ( .A(smc_off_b), .B(rst_osc_b), .Y(disable_osc));
nand2_hvt I270 ( .A(crst_b), .Y(net064), .B(por_b));
inv_hvt I233 ( .A(clk_out), .Y(clk_out_b));
inv_hvt I271 ( .A(net064), .Y(rst_osc_b));
inv_hvt I267 ( .A(net078), .Y(clk_in));
inv_hvt I262 ( .A(net067), .Y(cnt_podt_out));
inv_hvt I275 ( .A(smc_oscoff_b), .Y(net0174));
inv_hvt I277 ( .A(net054), .Y(cnt_rst));
inv_hvt I229 ( .A(rst_osc_b), .Y(net090));
inv_hvt I253 ( .A(net0124), .Y(rst_off_latch));
inv_hvt I232 ( .A(clk_out_b), .Y(smc_clk));
nor2_hvt I272 ( .A(net066), .B(disable_osc), .Y(smc_oscen));
nor2_hvt I266 ( .A(clk_out), .B(smc_podt_off), .Y(net078));
nor2_hvt I273 ( .A(smc_oscoff_b), .B(rst_osc_b), .Y(net066));
nor2_hvt I276 ( .A(net090), .B(smc_podt_rst), .Y(net054));
nor2_hvt I274 ( .A(smc_oscoff_b), .B(cnt_rst), .Y(net0124));
tiehis I179 ( .tiehi(net076));
ml_osc Iml_osc ( .smc_osc_fsel(smc_osc_fsel[1:0]), .clk_out(clk_out),
     .smc_oscen(smc_oscen));

endmodule
// Library - ice384chip, Cell - CHIP_route_lft2rgt_ice384, View -
//schematic
// LAST TIME SAVED: Dec 23 16:05:28 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module CHIP_route_lft2rgt_ice384 ( bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bldld, cm_banksel_bltrd1_3_,
     cm_clk_blbrd, cm_clk_bltrd1, cm_sdi_u0, cm_sdi_u1, cm_sdi_u2d,
     cm_sdi_u3d2, core_por_b0, core_por_b_rowu3, core_por_bb,
     cram_pgateoff, cram_prec, cram_prec_bltrd1, cram_pullup_b,
     cram_pullup_b_bltrd1, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, cram_write_bltrd1, data_muxsel1_blbrd,
     data_muxsel1_bltrd1, data_muxsel_blbrd, data_muxsel_bltrd1,
     en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1, end_of_startup,
     gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr,
     md_spi_b, mode0, mux_jtag_sel, nvcm_spi_sdi, nvcm_spi_ss_b,
     pgate_r, reset_b_r, row_test0, rst_b, sdo_enable, shift0,
     smc_load_nvcm_bstream, smc_row_inc, smc_rsr_rst,
     smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1, smc_write0,
     smc_write_bltl1d1, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, update0, vdd_cntl_r, wl_r, bp0, cdone_in,
     cm_sdo_u0d1, cm_sdo_u1d3, cm_sdo_u2d1, cm_sdo_u3, creset_b_int,
     fromsdo, idcode_msb20bits, last_rsr3, nvcm_boot, nvcm_dis_idchk,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, spi_ss_in_bbank,
     tck_pad, tdi_pad, tms_pad, trstb_pad, vddio_rightbank );
output  bs_en0, cdone_out, ceb0, cm_banksel_blbrd_2_,
     cm_banksel_bltrd1_3_, cm_clk_blbrd, cm_clk_bltrd1, core_por_b0,
     core_por_b_rowu3, core_por_bb, cram_pgateoff, cram_prec,
     cram_prec_bltrd1, cram_pullup_b, cram_pullup_b_bltrd1, cram_rst,
     cram_vddoff, cram_wl_en, cram_write, cram_write_bltrd1,
     data_muxsel1_blbrd, data_muxsel1_bltrd1, data_muxsel_blbrd,
     data_muxsel_bltrd1, en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1,
     end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, mux_jtag_sel, nvcm_spi_sdi, nvcm_spi_ss_b, row_test0,
     rst_b, sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1,
     smc_write0, smc_write_bltl1d1, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, update0;

input  bp0, cdone_in, creset_b_int, fromsdo, last_rsr3, nvcm_boot,
     nvcm_dis_idchk, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, smc_core_por_bottom1, smc_core_por_bottom2,
     tck_pad, tdi_pad, tms_pad, trstb_pad, vddio_rightbank;

output [1:0]  last_rsr;
output [1:0]  cm_sdi_u0;
output [159:0]  vdd_cntl_r;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_sdi_u3d2;
output [159:0]  pgate_r;
output [159:0]  wl_r;
output [1:0]  cm_sdi_u2d;
output [1:0]  cm_banksel_bldld;
output [159:0]  reset_b_r;

input [1:0]  cm_sdo_u0d1;
input [1:0]  cm_sdo_u2d1;
input [1:0]  cm_sdo_u1d3;
input [19:0]  idcode_msb20bits;
input [1:0]  cm_sdo_u3;
input [4:0]  spi_ss_in_bbank;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  smc_osco_fsel;

wire  [3:0]  net0388;

wire  [3:0]  net0387;

wire  [10:0]  net0462;

wire  [3:0]  cm_banksel;

wire  [1:0]  cdsbus0;

wire  [1:0]  dff_out_top;

wire  [6:0]  net0409;



smc_and_jtag_id_u40 I_smc_and_jtag_id_u40 (
     .nvcm_dis_idchk(nvcm_dis_idchk), .bm_sa({net0462[0], net0462[1],
     net0462[2], net0462[3], net0462[4], net0462[5], net0462[6],
     net0462[7], net0462[8], net0462[9], net0462[10]}),
     .warmboot_sel({net497, net497}), .trst_pad(trstb_pad),
     .tms_pad(tms_pad), .tdi_pad(tdi_pad), .tck_pad(tck_pad),
     .spi_ss_in_b(spi_ss_in_bbank[4]), .cdone_in(cdone_in),
     .spi_sdi(spi_ss_in_bbank[2]), .spi_clk_in(spi_ss_in_bbank[3]),
     .psdi({net497, net497, net497, net497, net497, net497, net497}),
     .por_b(smc_por_b0), .osc_clk(osc_clk),
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .idcode_msb20bits(idcode_msb20bits[19:0]),
     .creset_b(crst_filterout), .coldboot_sel(spi_ss_in_bbank[1:0]),
     .cnt_podt_out(cnt_podt_out), .cm_sdo_u3(dff_out_top[1:0]),
     .cm_sdo_u2(cm_sdo_u2d1[1:0]), .cm_sdo_u1(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0(cm_sdo_u0d1[1:0]), .cm_monitor_cell({net497, net497,
     net497, net497}), .cm_last_rsr(last_rsr3), .bschain_sdo(fromsdo),
     .bp0(bp0), .boot(net497), .bm_bank_sdo({net497, net497, net497,
     net497}), .tdo_pad(totdopad), .tdo_oe_pad(sdo_enable),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out),
     .smc_wwlwrt_en(smc_wwlwrt_en), .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wdis_dclk(smc_wdis_dclk_blbrd),
     .smc_wcram_rst(smc_wcram_rst), .smc_seq_rst(smc_seq_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rsr_rst(smc_rsr_rst),
     .smc_rrst_pullwlen(smc_rrst_pullwlen), .smc_rpull_b(smc_rpull_b),
     .smc_rprec(smc_rprec), .smc_row_inc(smc_row_inc),
     .smc_read(smc_read), .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .psdo({net0409[0], net0409[1], net0409[2], net0409[3], net0409[4],
     net0409[5], net0409[6]}), .nvcm_spi_ss_b(nvcm_spi_ss_b),
     .nvcm_spi_sdi(nvcm_spi_sdi), .md_spi_b(md_spi_b),
     .j_upd_dr(update0), .j_tdi(j_tdi), .j_tck(j_tck),
     .j_shift0(shift0), .j_sft_dr(shiftromsmc), .j_rst_b(j_rst_b),
     .j_row_test(row_test0), .j_mode(mode0), .j_hiz_b(hiz_b0),
     .j_ceb0(ceb0), .gsr(net439), .gint_hz(net440),
     .end_of_startup(net441), .en_8bconfig_b(en_8bconfig_b_blbrd),
     .data_muxsel1(data_muxsel1_blbrd),
     .data_muxsel(data_muxsel_blbrd), .cm_sdi_u3(cdsbus0[1:0]),
     .cm_sdi_u2(cm_sdi_u2d[1:0]), .cm_sdi_u1(cm_sdi_u1[1:0]),
     .cm_sdi_u0(cm_sdi_u0[1:0]), .cm_clk(cm_clk),
     .cm_banksel(cm_banksel[3:0]), .cdone_out(cdone_out),
     .bs_en(bs_en0), .bm_wdummymux_en(net0458), .bm_sweb(net0381),
     .bm_sreb(net0382), .bm_sclkrw(net0383), .bm_rcapmux_en(net0384),
     .bm_init(net0385), .bm_clk(net0386), .bm_banksel({net0387[0],
     net0387[1], net0387[2], net0387[3]}), .bm_bank_sdi({net0388[0],
     net0388[1], net0388[2], net0388[3]}));
CHIP_route_lft_ice384 I_chip_route_lft2rgt_ice384 ( .wl_l(wl_r[159:0]),
     .vdd_cntl_l(vdd_cntl_r[159:0]), .reset_l(reset_b_r[159:0]),
     .pgate_l(pgate_r[159:0]), .tck_padl0(j_tck),
     .smc_writel0(smc_write0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbrd),
     .smc_rsr_rstl0(smc_rsr_rst), .smc_row_incl0(smc_row_inc),
     .row_testl1(row_test0), .j_rst_bl0(j_rst_b),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbrd),
     .data_muxsel_blbld(data_muxsel_blbrd),
     .data_muxsel1_blbld(data_muxsel1_blbrd),
     .cram_write_blbld(cram_write), .cram_wl_enl0(cram_wl_en),
     .cram_vddoffl0(cram_vddoff), .cram_rstl0(cram_rst),
     .cram_pullup_blbld(cram_pullup_b), .cram_prec_blbld(cram_prec),
     .cram_pgateoffl0(cram_pgateoff), .core_por_bbl0(core_por_bb),
     .cm_sdo_u1(cm_sdo_u3[1:0]), .cm_sdi_u1d(cdsbus0[1:0]),
     .cm_clk_blbld(cm_clk_blbrd), .cm_banksel_blbld(cm_banksel[3]),
     .cm_banksel_blbld1(cm_banksel_blbrd_2_),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltrd1),
     .last_rsr(last_rsr[1:0]), .last_rsr0(net485),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu2_b),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltrd1),
     .data_muxsel1_bltld3(data_muxsel1_bltrd1),
     .cram_write_bltld3(cram_write_bltrd1),
     .cram_pullup_bltld3(cram_pullup_b_bltrd1),
     .cram_prec_bltld3(cram_prec_bltrd1),
     .core_por_b_rowu1(core_por_b_rowu3),
     .smc_write_bltld3(smc_write_bltl1d1),
     .cm_sdo_u1d1(dff_out_top[1:0]), .cm_sdi_u1d3(cm_sdi_u3d2[1:0]),
     .cm_clk_bltld3(cm_clk_bltrd1),
     .cm_banksel_bltld3_1_(cm_banksel_bltrd1_3_));
creset_filter I561 ( .in(creset_b_int), .out(crst_filterout));
sg_bufx10_ice8p I558 ( .in(net441), .out(end_of_startup));
sg_bufx10_ice8p I559 ( .in(net439), .out(gsr));
sg_bufx10_ice8p I560 ( .in(net440), .out(gint_hz));
sg_bufx10_ice8p I551 ( .in(en_8bconfig_b_blbrd), .out(net0327));
sg_bufx10_ice8p I683_1_ ( .in(cm_banksel[1]),
     .out(cm_banksel_bldld[1]));
sg_bufx10_ice8p I683_0_ ( .in(cm_banksel[0]),
     .out(cm_banksel_bldld[0]));
sg_bufx10_ice8p I681 ( .in(cm_banksel[2]), .out(cm_banksel_blbrd_2_));
SMC_CORE_POR_right_ice8p I_SMC_CORE_POR_right (
     .core_por_b0(core_por_b0), .core_por_bb(core_por_bb),
     .vddio_rightbank(vddio_rightbank), .smc_por_b(smc_por_b0),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .creset_b(crst_filterout));
ml_cram_logic_ice8p ml_cram_logic_ice8p_1f (
     .smc_wwlwrt_en(smc_wwlwrt_en), .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wcram_rst(smc_wcram_rst), .smc_seq_rst(smc_seq_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rrst_pullwlen(smc_rrst_pullwlen),
     .smc_rpull_b(smc_rpull_b), .smc_rprec(smc_rprec),
     .smc_read(smc_read), .smc_clk(cm_clk), .por(core_por_bb),
     .smc_clk_out(cm_clk_blbrd), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff));
inv_hvt Imux4jtag_sel ( .A(trstb_pad), .Y(mux_jtag_sel));
ml_osc_top I_ml_osc_top ( .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]), .por_b(core_por_b0),
     .crst_b(crst_filterout), .smc_clk(osc_clk),
     .cnt_podt_out(cnt_podt_out));
tielo I553 ( .tielo(net497));

endmodule
// Library - ice384chip, Cell - ring_route00_ice384, View - schematic
// LAST TIME SAVED: Jan 12 15:26:11 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module ring_route00_ice384 ( bs_en0, cdone_out, ceb0, end_of_startup,
     gint_hz, gsr, hiz_b0, j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr, md_spi_b, mode0,
     mux_jtag_sel_b, pgate_l, pgate_r, reset_b_l, reset_b_r,
     sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_pad, update0, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r, bl_bot, bl_top, vppin, cdone_in, creset_b_int, fromsdo,
     spi_ss_in_bbank, tck_pad, tdi_pad, tms_pad, trstb_pad,
     vddio_bottombank, vddio_spi );
output  bs_en0, cdone_out, ceb0, end_of_startup, gint_hz, gsr, hiz_b0,
     j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, md_spi_b, mode0, mux_jtag_sel_b,
     sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_pad, update0;

inout  vppin;

input  cdone_in, creset_b_int, fromsdo, tck_pad, tdi_pad, tms_pad,
     trstb_pad, vddio_bottombank, vddio_spi;

output [159:0]  vdd_cntl_r;
output [159:0]  pgate_r;
output [159:0]  wl_r;
output [159:0]  wl_l;
output [159:0]  reset_b_l;
output [159:0]  vdd_cntl_l;
output [159:0]  pgate_l;
output [3:0]  last_rsr;
output [159:0]  reset_b_r;

inout [363:0]  bl_top;
inout [363:0]  bl_bot;

input [4:0]  spi_ss_in_bbank;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdi_u2d;

wire  [1:1]  cm_banksel_bltld3;

wire  [1:0]  cm_banksel;

wire  [1:0]  cm_sdi_u3d2;

wire  [1:0]  cm_sdo_u3;

wire  [1:0]  cm_sdo_u1;

wire  [1:0]  cm_sdo_u1d1;

wire  [1:0]  cm_sdo_u2d1;

wire  [1:0]  cm_sdi_u1d3;

wire  [1:0]  cm_sdi_u1;

wire  [3:3]  cm_banksel_bltrd1;

wire  [19:0]  idcode_msb20bits;

wire  [1:0]  cm_sdi_u0;

wire  [4:0]  spi_ss_in_bbankd;

wire  [1:0]  cm_sdo_u0d1;

wire  [1:0]  cm_sdi_u1d;

wire  [1:0]  cm_sdo_u1d3;



NCAP_25_LP  C7 ( .MINUS(gnd_), .PLUS(vpxa_int));
NCAP_25_LP  C3 ( .MINUS(gnd_), .PLUS(vdd_));
NCAP_25_LP  C1 ( .MINUS(gnd_), .PLUS(vpp_int));
nvcm_ml_block_ice384_june I_nvcm_ml_block_ice384_june (
     .vpp_int(vpp_int), .vpxa_int(vpxa_int),
     .nvcm_dis_idchk(nvcm_dis_idchk),
     .idcode_msb20bits_out(idcode_msb20bits[19:0]), .tvdd_fsm(net373),
     .tgnd_fsm(net374), .spi_ss_b(nvcm_spi_ss_b),
     .spi_sdi(nvcm_spi_sdi), .rst_b(rst_b), .nvcm_ce_b(cdone_in),
     .clk(spi_clk_out2fsm), .spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .spi_sdo(nvcm_spi_sdo), .nvcm_rdy(nvcm_rdy),
     .nvcm_boot(nvcm_boot),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream),
     .fsm_tm_margin0_read(net385), .fsm_recall(net386), .bp0(bp0),
     .vpp(vppin), .nvcm_relextspi(nvcm_relextspi));
CHIP_route_bot_ice384 I_CHIP_route_bot_ice384 ( .bl_bot(bl_bot[363:0]),
     .smc_write(smc_write), .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_rsr_rst(smc_rsr_rsr), .smc_row_inc(smc_row_inc),
     .row_test0(row_test0),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1_0_), .j_tck(j_tck),
     .j_rst_b(j_rst_b), .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .cram_wl_enl0(cram_wl_enl0),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_blbrd(data_muxsel1_blbrd), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff),
     .core_por_bb(core_por_bb),
     .cm_banksel_blbld_1_(cm_banksel_blbld_1_),
     .core_por_b0(core_por_b0), .cm_sdo_u1d1(cm_sdo_u1d1[1:0]),
     .cm_sdi_u2d(cm_sdi_u2d[1:0]), .cm_sdi_u1(cm_sdi_u1[1:0]),
     .cm_sdi_u0(cm_sdi_u0[1:0]), .cm_clk_blbrd(cm_clk_blbrd),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .cm_banksel(cm_banksel[1:0]), .smc_writel0(smc_writel0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .smc_rsr_rstl0(smc_rsr_rstl0), .smc_row_incl0(smc_row_incl0),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .row_testl1(row_testl1), .last_rsr3(last_rsr3),
     .j_rst_bl0(j_rst_bl0), .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbld(data_muxsel1_blbld), .last_rsr1(last_rsr0),
     .cram_write_blbld(cram_write_blbld),
     .cram_vddoffl0(cram_vddoffl0), .cram_rstl0(cram_rstl0),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld),
     .cram_pgateoffl0(cram_pgateoffl0), .core_por_bbl0(core_por_bbl0),
     .cm_sdo_u2d1(cm_sdo_u2d1[1:0]), .cm_sdo_u1d3(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0d1(cm_sdo_u0d1[1:0]), .tck_padl0(tck_padl0),
     .cm_clk_blbld(cm_clk_blbld), .cm_sdi_u1d(cm_sdi_u1d[1:0]),
     .spi_ss_in_bbank(spi_ss_in_bbank[4:0]),
     .spi_ss_in_bbankd(spi_ss_in_bbankd[4:0]), .vddio_spi(vddio_spi),
     .vddio_botbank(vddio_bottombank));
CHIP_route_lft2rgt_ice384 I_CHIP_route_rgt_ice384 (
     .nvcm_dis_idchk(nvcm_dis_idchk), .vdd_cntl_r(vdd_cntl_r[159:0]),
     .reset_b_r(reset_b_r[159:0]), .pgate_r(pgate_r[159:0]),
     .wl_r(wl_r[159:0]), .vddio_rightbank(vddp_), .tms_pad(tms_pad),
     .tdi_pad(tdi_pad), .tck_pad(tck_pad),
     .spi_ss_in_bbank(spi_ss_in_bbankd[4:0]),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot), .last_rsr3(last_rsr3),
     .fromsdo(fromsdo), .cm_sdo_u3(cm_sdo_u3[1:0]),
     .cm_sdo_u2d1(cm_sdo_u2d1[1:0]), .cm_sdo_u1d3(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0d1(cm_sdo_u0d1[1:0]), .cdone_in(cdone_in), .bp0(bp0),
     .update0(update0), .totdopad(tdo_pad),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out),
     .smc_write0(smc_write),
     .smc_wdis_dclk_bltrd1(smc_wdis_dclk_bltrd1),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_rsr_rst(smc_rsr_rsr), .smc_row_inc(smc_row_inc),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .shift0(shift0),
     .sdo_enable(sdo_enable), .rst_b(rst_b), .row_test0(row_test0),
     .nvcm_spi_ss_b(nvcm_spi_ss_b), .nvcm_spi_sdi(nvcm_spi_sdi),
     .mode0(mode0), .md_spi_b(md_spi_b), .last_rsr(last_rsr[3:2]),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .j_tdi(j_tdi), .j_tck(j_tck), .j_rst_b(j_rst_b), .hiz_b0(hiz_b0),
     .gsr(gsr), .gint_hz(gint_hz), .end_of_startup(end_of_startup),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_bltrd1(data_muxsel1_bltld3),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .cram_write_bltrd1(cram_write_bltrd1), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_pullup_b(cram_pullup_b),
     .cram_prec_bltrd1(cram_prec_bltrd1), .cram_prec(cram_prec),
     .cram_pgateoff(cram_pgateoff), .core_por_bb(core_por_bb),
     .core_por_b_rowu3(core_por_b_rowu3),
     .smc_write_bltl1d1(smc_write_bltl1d1r), .core_por_b0(core_por_b0),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .cm_clk_bltrd1(cm_clk_bltrd1), .cm_clk_blbrd(cm_clk_blbrd),
     .cm_banksel_bltrd1_3_(cm_banksel_bltrd1[3]),
     .cm_banksel_bldld(cm_banksel[1:0]),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_), .ceb0(ceb0),
     .cdone_out(cdone_out), .bs_en0(bs_en0),
     .creset_b_int(creset_b_int), .mux_jtag_sel(mux_jtag_sel_b),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .idcode_msb20bits(idcode_msb20bits[19:0]), .trstb_pad(trstb_pad));
CHIP_route_lft_ice384 I_CHIP_route_lft_ice384 ( .wl_l(wl_l[159:0]),
     .vdd_cntl_l(vdd_cntl_l[159:0]), .reset_l(reset_b_l[159:0]),
     .pgate_l(pgate_l[159:0]), .smc_writel0(smc_writel0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .smc_rsr_rstl0(smc_rsr_rstl0), .smc_row_incl0(smc_row_incl0),
     .row_testl1(row_testl1), .j_rst_bl0(j_rst_bl0),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_wl_enl0(cram_wl_enl0),
     .cram_vddoffl0(cram_vddoffl0), .cram_rstl0(cram_rstl0),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld),
     .cram_pgateoffl0(cram_pgateoffl0), .core_por_bbl0(core_por_bbl0),
     .cm_sdo_u1(cm_sdo_u1[1:0]), .cm_sdi_u1d(cm_sdi_u1d[1:0]),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbld(cm_banksel_blbld_1_),
     .cm_banksel_blbld1(cm_banksel_blbld1_0_),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel1_bltld3(data_muxsel1_bltld1),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_bltld3),
     .cram_prec_bltld3(cm_prec_bltld3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .cm_sdo_u1d1(cm_sdo_u1d1[1:0]), .last_rsr(last_rsr[1:0]),
     .last_rsr0(last_rsr0), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3),
     .data_muxsel_bltld3(data_muxsel_bltld1),
     .cm_banksel_bltld3_1_(cm_banksel_bltld3[1]),
     .smc_write_bltld3(smc_write_bltld3), .tck_padl0(tck_padl0));
CHIP_route_top_ice384 I_CHIP_route_top_ice384 ( .bl_top(bl_top[363:0]),
     .smc_write_bltld3(smc_write_bltld3),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltld1),
     .data_muxsel1_bltrd1(data_muxsel1_bltld3),
     .data_muxsel1_bltld3(data_muxsel1_bltld1),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_bltld3),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1),
     .core_por_b_rowu3(core_por_b_rowu3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .cm_prec_bltld3(cm_prec_bltld3), .cm_clk_bltrd1(cm_clk_bltrd1),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cm_banksel_bltrd1(cm_banksel_bltrd1[3]),
     .cm_banksel_bltld3(cm_banksel_bltld3[1]),
     .cm_sdo_u3(cm_sdo_u3[1:0]), .cm_sdo_u1(cm_sdo_u1[1:0]),
     .smc_write_bltl1d1(smc_write_bltl1d1r));
sg_bufx10_ice8p I_clkbuf ( .in(spi_clk_out), .out(spi_clk_out2fsm));

endmodule
// Library - umc40lp, Cell - RNPPO_LP, View - schematic
// LAST TIME SAVED: Jan 18 18:48:13 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module RNPPO_LP_pcell2461 ( MINUS, PLUS, B );
inout  MINUS, PLUS;

input  B;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



primRes3  R9 ( .MINUS(MINUS), .PLUS(n9), .B(B));
primRes3  R8 ( .MINUS(n9), .PLUS(n8), .B(B));
primRes3  R7 ( .MINUS(n8), .PLUS(n7), .B(B));
primRes3  R6 ( .MINUS(n7), .PLUS(n6), .B(B));
primRes3  R5 ( .MINUS(n6), .PLUS(n5), .B(B));
primRes3  R4 ( .MINUS(n5), .PLUS(n4), .B(B));
primRes3  R3 ( .MINUS(n4), .PLUS(n3), .B(B));
primRes3  R2 ( .MINUS(n3), .PLUS(n2), .B(B));
primRes3  R1 ( .MINUS(n2), .PLUS(n1), .B(B));
primRes3  R0 ( .MINUS(n1), .PLUS(PLUS), .B(B));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_1f, View - schematic
// LAST TIME SAVED: Aug  3 19:29:15 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_ctrl_1f ( yp1, yp1_b_25, yp2, yp2_b_25, yp3_25,
     yp3_b_25, yp_test_25, yp_test_b_25, vblinhi_pgm_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b, yp1_sel,
     yp2_b_low_b, yp2_sel, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, yp_test,
     ysup_25 );

inout  vblinhi_pgm_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b,
     yp2_b_low_b, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, ysup_25;

output [1:0]  yp_test_b_25;
output [7:0]  yp3_25;
output [5:0]  yp1;
output [7:0]  yp3_b_25;
output [7:0]  yp2_b_25;
output [7:0]  yp2;
output [1:0]  yp_test_25;
output [5:0]  yp1_b_25;

input [5:0]  yp1_sel;
input [7:0]  yp2_sel;
input [1:0]  yp_test;
input [7:0]  yp3_sel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_1_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1]), .yp_test(yp_test[1]),
     .yp_test_25(yp_test_25[1]));
ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_0_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[0]), .yp_test(yp_test[0]),
     .yp_test_25(yp_test_25[0]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_7_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[7]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[7]), .yp3_25(yp3_25[7]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_6_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[6]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[6]), .yp3_25(yp3_25[6]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_5_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[5]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[5]), .yp3_25(yp3_25[5]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_4_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[4]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[4]), .yp3_25(yp3_25[4]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_3_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[3]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[3]), .yp3_25(yp3_25[3]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_2_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[2]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[2]), .yp3_25(yp3_25[2]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_1_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[1]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[1]), .yp3_25(yp3_25[1]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_0_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[0]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[0]), .yp3_25(yp3_25[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_7_ ( .yp21_sel(yp2_sel[7]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[7]), .yp21(yp2[7]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_6_ ( .yp21_sel(yp2_sel[6]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[6]), .yp21(yp2[6]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_5_ ( .yp21_sel(yp2_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[5]), .yp21(yp2[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_4_ ( .yp21_sel(yp2_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[4]), .yp21(yp2[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_3_ ( .yp21_sel(yp2_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[3]), .yp21(yp2[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_2_ ( .yp21_sel(yp2_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[2]), .yp21(yp2[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_1_ ( .yp21_sel(yp2_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[1]), .yp21(yp2[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_0_ ( .yp21_sel(yp2_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[0]), .yp21(yp2[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_5_ ( .yp21_sel(yp1_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[5]), .yp21(yp1[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_4_ ( .yp21_sel(yp1_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[4]), .yp21(yp1[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_3_ ( .yp21_sel(yp1_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[3]), .yp21(yp1[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_2_ ( .yp21_sel(yp1_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[2]), .yp21(yp1[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_1_ ( .yp21_sel(yp1_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[1]), .yp21(yp1[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_0_ ( .yp21_sel(yp1_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[0]), .yp21(yp1[0]));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_1_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_0_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - umc40lp, Cell - RNPPO_LP, View - schematic
// LAST TIME SAVED: Jan 18 18:48:13 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module RNPPO_LP_pcell2462 ( MINUS, PLUS, B );
inout  MINUS, PLUS;

input  B;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



primRes3  R99 ( .MINUS(MINUS), .PLUS(n99), .B(B));
primRes3  R98 ( .MINUS(n99), .PLUS(n98), .B(B));
primRes3  R97 ( .MINUS(n98), .PLUS(n97), .B(B));
primRes3  R96 ( .MINUS(n97), .PLUS(n96), .B(B));
primRes3  R95 ( .MINUS(n96), .PLUS(n95), .B(B));
primRes3  R94 ( .MINUS(n95), .PLUS(n94), .B(B));
primRes3  R93 ( .MINUS(n94), .PLUS(n93), .B(B));
primRes3  R92 ( .MINUS(n93), .PLUS(n92), .B(B));
primRes3  R91 ( .MINUS(n92), .PLUS(n91), .B(B));
primRes3  R90 ( .MINUS(n91), .PLUS(n90), .B(B));
primRes3  R89 ( .MINUS(n90), .PLUS(n89), .B(B));
primRes3  R88 ( .MINUS(n89), .PLUS(n88), .B(B));
primRes3  R87 ( .MINUS(n88), .PLUS(n87), .B(B));
primRes3  R86 ( .MINUS(n87), .PLUS(n86), .B(B));
primRes3  R85 ( .MINUS(n86), .PLUS(n85), .B(B));
primRes3  R84 ( .MINUS(n85), .PLUS(n84), .B(B));
primRes3  R83 ( .MINUS(n84), .PLUS(n83), .B(B));
primRes3  R82 ( .MINUS(n83), .PLUS(n82), .B(B));
primRes3  R81 ( .MINUS(n82), .PLUS(n81), .B(B));
primRes3  R80 ( .MINUS(n81), .PLUS(n80), .B(B));
primRes3  R79 ( .MINUS(n80), .PLUS(n79), .B(B));
primRes3  R78 ( .MINUS(n79), .PLUS(n78), .B(B));
primRes3  R77 ( .MINUS(n78), .PLUS(n77), .B(B));
primRes3  R76 ( .MINUS(n77), .PLUS(n76), .B(B));
primRes3  R75 ( .MINUS(n76), .PLUS(n75), .B(B));
primRes3  R74 ( .MINUS(n75), .PLUS(n74), .B(B));
primRes3  R73 ( .MINUS(n74), .PLUS(n73), .B(B));
primRes3  R72 ( .MINUS(n73), .PLUS(n72), .B(B));
primRes3  R71 ( .MINUS(n72), .PLUS(n71), .B(B));
primRes3  R70 ( .MINUS(n71), .PLUS(n70), .B(B));
primRes3  R69 ( .MINUS(n70), .PLUS(n69), .B(B));
primRes3  R68 ( .MINUS(n69), .PLUS(n68), .B(B));
primRes3  R67 ( .MINUS(n68), .PLUS(n67), .B(B));
primRes3  R66 ( .MINUS(n67), .PLUS(n66), .B(B));
primRes3  R65 ( .MINUS(n66), .PLUS(n65), .B(B));
primRes3  R64 ( .MINUS(n65), .PLUS(n64), .B(B));
primRes3  R63 ( .MINUS(n64), .PLUS(n63), .B(B));
primRes3  R62 ( .MINUS(n63), .PLUS(n62), .B(B));
primRes3  R61 ( .MINUS(n62), .PLUS(n61), .B(B));
primRes3  R60 ( .MINUS(n61), .PLUS(n60), .B(B));
primRes3  R59 ( .MINUS(n60), .PLUS(n59), .B(B));
primRes3  R58 ( .MINUS(n59), .PLUS(n58), .B(B));
primRes3  R57 ( .MINUS(n58), .PLUS(n57), .B(B));
primRes3  R56 ( .MINUS(n57), .PLUS(n56), .B(B));
primRes3  R55 ( .MINUS(n56), .PLUS(n55), .B(B));
primRes3  R54 ( .MINUS(n55), .PLUS(n54), .B(B));
primRes3  R53 ( .MINUS(n54), .PLUS(n53), .B(B));
primRes3  R52 ( .MINUS(n53), .PLUS(n52), .B(B));
primRes3  R51 ( .MINUS(n52), .PLUS(n51), .B(B));
primRes3  R50 ( .MINUS(n51), .PLUS(n50), .B(B));
primRes3  R49 ( .MINUS(n50), .PLUS(n49), .B(B));
primRes3  R48 ( .MINUS(n49), .PLUS(n48), .B(B));
primRes3  R47 ( .MINUS(n48), .PLUS(n47), .B(B));
primRes3  R46 ( .MINUS(n47), .PLUS(n46), .B(B));
primRes3  R45 ( .MINUS(n46), .PLUS(n45), .B(B));
primRes3  R44 ( .MINUS(n45), .PLUS(n44), .B(B));
primRes3  R43 ( .MINUS(n44), .PLUS(n43), .B(B));
primRes3  R42 ( .MINUS(n43), .PLUS(n42), .B(B));
primRes3  R41 ( .MINUS(n42), .PLUS(n41), .B(B));
primRes3  R40 ( .MINUS(n41), .PLUS(n40), .B(B));
primRes3  R39 ( .MINUS(n40), .PLUS(n39), .B(B));
primRes3  R38 ( .MINUS(n39), .PLUS(n38), .B(B));
primRes3  R37 ( .MINUS(n38), .PLUS(n37), .B(B));
primRes3  R36 ( .MINUS(n37), .PLUS(n36), .B(B));
primRes3  R35 ( .MINUS(n36), .PLUS(n35), .B(B));
primRes3  R34 ( .MINUS(n35), .PLUS(n34), .B(B));
primRes3  R33 ( .MINUS(n34), .PLUS(n33), .B(B));
primRes3  R32 ( .MINUS(n33), .PLUS(n32), .B(B));
primRes3  R31 ( .MINUS(n32), .PLUS(n31), .B(B));
primRes3  R30 ( .MINUS(n31), .PLUS(n30), .B(B));
primRes3  R29 ( .MINUS(n30), .PLUS(n29), .B(B));
primRes3  R28 ( .MINUS(n29), .PLUS(n28), .B(B));
primRes3  R27 ( .MINUS(n28), .PLUS(n27), .B(B));
primRes3  R26 ( .MINUS(n27), .PLUS(n26), .B(B));
primRes3  R25 ( .MINUS(n26), .PLUS(n25), .B(B));
primRes3  R24 ( .MINUS(n25), .PLUS(n24), .B(B));
primRes3  R23 ( .MINUS(n24), .PLUS(n23), .B(B));
primRes3  R22 ( .MINUS(n23), .PLUS(n22), .B(B));
primRes3  R21 ( .MINUS(n22), .PLUS(n21), .B(B));
primRes3  R20 ( .MINUS(n21), .PLUS(n20), .B(B));
primRes3  R19 ( .MINUS(n20), .PLUS(n19), .B(B));
primRes3  R18 ( .MINUS(n19), .PLUS(n18), .B(B));
primRes3  R17 ( .MINUS(n18), .PLUS(n17), .B(B));
primRes3  R16 ( .MINUS(n17), .PLUS(n16), .B(B));
primRes3  R15 ( .MINUS(n16), .PLUS(n15), .B(B));
primRes3  R14 ( .MINUS(n15), .PLUS(n14), .B(B));
primRes3  R13 ( .MINUS(n14), .PLUS(n13), .B(B));
primRes3  R12 ( .MINUS(n13), .PLUS(n12), .B(B));
primRes3  R11 ( .MINUS(n12), .PLUS(n11), .B(B));
primRes3  R10 ( .MINUS(n11), .PLUS(n10), .B(B));
primRes3  R9 ( .MINUS(n10), .PLUS(n9), .B(B));
primRes3  R8 ( .MINUS(n9), .PLUS(n8), .B(B));
primRes3  R7 ( .MINUS(n8), .PLUS(n7), .B(B));
primRes3  R6 ( .MINUS(n7), .PLUS(n6), .B(B));
primRes3  R5 ( .MINUS(n6), .PLUS(n5), .B(B));
primRes3  R4 ( .MINUS(n5), .PLUS(n4), .B(B));
primRes3  R3 ( .MINUS(n4), .PLUS(n3), .B(B));
primRes3  R2 ( .MINUS(n3), .PLUS(n2), .B(B));
primRes3  R1 ( .MINUS(n2), .PLUS(n1), .B(B));
primRes3  R0 ( .MINUS(n1), .PLUS(PLUS), .B(B));

endmodule
// Library - umc40nm_io, Cell - SDDIOBREAK_sbt_a, View - schematic
// LAST TIME SAVED: Jan 17 18:29:00 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module SDDIOBREAK_sbt_a ( VDDIO );
input  VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



DIOP_25_LP  D1 ( .PLUS(gnd_), .MINUS(VDDIO));
N_25OD33_LP  NM4 ( .D(VDDIO), .B(gnd_), .G(net_1260), .S(gnd_));
N_25OD33_LP  NM0 ( .D(gnd_), .B(gnd_), .G(net_1259), .S(gnd_));
N_25OD33_LP  NM1 ( .D(net_1260), .B(gnd_), .G(net_1259), .S(gnd_));
P_25OD33_LP  PM3 ( .D(net_1260), .B(VDDIO), .G(net_1259), .S(VDDIO));
RNPPO_LP_pcell2461 R0 ( .B(vdd_), .MINUS(net39), .PLUS(VDDIO));
RNPPO_LP_pcell2462 R2 ( .B(gnd_), .MINUS(net36), .PLUS(net39));
RNPPO_LP_pcell2462 R3 ( .B(VDDIO), .MINUS(net_1259), .PLUS(net36));

endmodule
// Library - misc, Cell - vpp_clamp_finger, View - schematic
// LAST TIME SAVED: Jan  6 16:00:42 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module vpp_clamp_finger ( VDDIO, VPP );
input  VDDIO, VPP;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M0 ( .D(net12), .B(gnd_), .G(gnd_), .S(gnd_));
N_25_LP  m1 ( .D(VPP), .B(gnd_), .G(VDDIO), .S(net12));

endmodule
// Library - misc, Cell - vpp_clamp, View - schematic
// LAST TIME SAVED: Jan  6 16:00:44 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module vpp_clamp ( VDDIO, VPP );
input  VDDIO, VPP;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



vpp_clamp_finger I0_3_ ( .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_2_ ( .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_1_ ( .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_0_ ( .VDDIO(VDDIO), .VPP(VPP));

endmodule
// Library - io, Cell - pvpp, View - schematic
// LAST TIME SAVED: Jan  6 16:00:48 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module pvpp ( vpp, vppin );
inout  vpp, vppin;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



RNPPO_LP_pcell2460 R1 ( .B(gnd_), .MINUS(vpp), .PLUS(vppin));
vddp_tiehigh I60_15_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_14_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_13_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_12_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_11_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_10_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_9_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_8_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_7_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_6_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_5_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_4_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_3_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_2_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_1_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_0_ ( .vddp_tieh(vddio_in));
vpp_clamp I59_15_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_14_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_13_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_12_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_11_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_10_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_9_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_8_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_7_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_6_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_5_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_4_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_3_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_2_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_1_ ( .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_0_ ( .VDDIO(vddio_in), .VPP(vpp));

endmodule
// Library - umc40nm_io, Cell - SVSS_sbt_a, View - schematic
// LAST TIME SAVED: Jan 17 18:27:29 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module SVSS_sbt_a ( VDDIO );
input  VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



DIOP_25_LP  D1 ( .PLUS(gnd_), .MINUS(VDDIO));
P_25OD33_LP  PM3 ( .D(net_1260), .B(VDDIO), .G(net_1259), .S(VDDIO));
N_25OD33_LP  NM2 ( .D(VDDIO), .B(gnd_), .G(net_1260), .S(gnd_));
N_25OD33_LP  NM0 ( .D(gnd_), .B(gnd_), .G(net_1259), .S(gnd_));
N_25OD33_LP  NM1 ( .D(net_1260), .B(gnd_), .G(net_1259), .S(gnd_));
RNPPO_LP_pcell2462 R3 ( .B(VDDIO), .MINUS(net_1259), .PLUS(net36));
RNPPO_LP_pcell2461 R0 ( .B(vdd_), .MINUS(net39), .PLUS(VDDIO));
RNPPO_LP_pcell2462 R2 ( .B(gnd_), .MINUS(net36), .PLUS(net39));

endmodule
// Library - umc40nm_io, Cell - SVDDIO_sbt_a, View - schematic
// LAST TIME SAVED: Jan 17 18:24:45 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module SVDDIO_sbt_a ( VDDIO );
inout  VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



DIOP_25_LP  D1 ( .PLUS(gnd_), .MINUS(VDDIO));
RNPPO_LP_pcell2461 R0 ( .B(vdd_), .MINUS(net25), .PLUS(VDDIO));
RNPPO_LP_pcell2462 R2 ( .B(gnd_), .MINUS(net22), .PLUS(net25));
RNPPO_LP_pcell2462 R3 ( .B(VDDIO), .MINUS(net_1259), .PLUS(net22));
N_25OD33_LP  NM2 ( .D(VDDIO), .B(gnd_), .G(net_1260), .S(gnd_));
N_25OD33_LP  NM0 ( .D(gnd_), .B(gnd_), .G(net_1259), .S(gnd_));
N_25OD33_LP  NM1 ( .D(net_1260), .B(gnd_), .G(net_1259), .S(gnd_));
P_25OD33_LP  PM3 ( .D(net_1260), .B(VDDIO), .G(net_1259), .S(VDDIO));

endmodule
// Library - umc40lp, Cell - RNPPO_LP, View - schematic
// LAST TIME SAVED: Jan 18 18:48:13 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module RNPPO_LP_pcell2463 ( MINUS, PLUS, B );
inout  MINUS, PLUS;

input  B;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



primRes3  R19 ( .MINUS(MINUS), .PLUS(n19), .B(B));
primRes3  R18 ( .MINUS(n19), .PLUS(n18), .B(B));
primRes3  R17 ( .MINUS(n18), .PLUS(n17), .B(B));
primRes3  R16 ( .MINUS(n17), .PLUS(n16), .B(B));
primRes3  R15 ( .MINUS(n16), .PLUS(n15), .B(B));
primRes3  R14 ( .MINUS(n15), .PLUS(n14), .B(B));
primRes3  R13 ( .MINUS(n14), .PLUS(n13), .B(B));
primRes3  R12 ( .MINUS(n13), .PLUS(n12), .B(B));
primRes3  R11 ( .MINUS(n12), .PLUS(n11), .B(B));
primRes3  R10 ( .MINUS(n11), .PLUS(n10), .B(B));
primRes3  R9 ( .MINUS(n10), .PLUS(n9), .B(B));
primRes3  R8 ( .MINUS(n9), .PLUS(n8), .B(B));
primRes3  R7 ( .MINUS(n8), .PLUS(n7), .B(B));
primRes3  R6 ( .MINUS(n7), .PLUS(n6), .B(B));
primRes3  R5 ( .MINUS(n6), .PLUS(n5), .B(B));
primRes3  R4 ( .MINUS(n5), .PLUS(n4), .B(B));
primRes3  R3 ( .MINUS(n4), .PLUS(n3), .B(B));
primRes3  R2 ( .MINUS(n3), .PLUS(n2), .B(B));
primRes3  R1 ( .MINUS(n2), .PLUS(n1), .B(B));
primRes3  R0 ( .MINUS(n1), .PLUS(PLUS), .B(B));

endmodule
// Library - umc40nm_io, Cell - SVDD_sbt_a, View - schematic
// LAST TIME SAVED: Jan 18 10:36:12 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module SVDD_sbt_a (  );supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25OD33_LP  M3 ( .D(net_1254), .B(vdd_), .G(net_1255), .S(vdd_));
DION_25_LP  D0 ( .PLUS(gnd_), .MINUS(vdd_));
N_11_LPHVT  NM0 ( .D(vdd_), .B(gnd_), .G(net_1254), .S(gnd_));
N_25OD33_LP  M1 ( .D(net_1254), .B(gnd_), .G(net_1255), .S(gnd_));
N_25OD33_LP  M0 ( .D(gnd_), .B(gnd_), .G(net_1255), .S(gnd_));
RNPPO_LP_pcell2463 R0 ( .B(vdd_), .MINUS(net_1255), .PLUS(vdd_));

endmodule
// Library - leafcell, Cell - tielo4x, View - schematic
// LAST TIME SAVED: Aug  3 19:21:04 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module tielo4x ( tielo );
output  tielo;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M0 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));
N_11_LPHVT  M1 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_a_clkdly, View - schematic
// LAST TIME SAVED: Aug  3 19:29:07 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_pump_a_clkdly ( out, in );
output  out;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M80 ( .D(vdd_), .B(vdd_), .G(net66), .S(vdd_));
inv_hvt I206 ( .A(in), .Y(net66));
inv_hvt I205 ( .A(net66), .Y(net70));
inv_hvt I207 ( .A(net70), .Y(out));

endmodule
// Library - umc40nm_io, Cell - LS21, View - schematic
// LAST TIME SAVED: Aug 23 17:58:20 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module LS21 ( AO, A, VDDIO );
output  AO;

input  A, VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25OD33_LP  POFF1 ( .D(net59), .B(VDDIO), .G(A), .S(net52));
P_25OD33_LP  PL1 ( .D(net52), .B(VDDIO), .G(AO), .S(VDDIO));
P_25OD33_LP  PL ( .D(net56), .B(VDDIO), .G(net59), .S(VDDIO));
P_25OD33_LP  POFF ( .D(AO), .B(VDDIO), .G(net067), .S(net56));
N_25OD33_LP  N1 ( .D(net59), .B(gnd_), .G(A), .S(gnd_));
N_25OD33_LP  N0 ( .D(AO), .B(gnd_), .G(net067), .S(gnd_));
inv IIV0 ( .A(A), .Y(net067));

endmodule
// Library - umc40nm_io, Cell - LS41, View - schematic
// LAST TIME SAVED: Aug 22 16:50:05 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module LS41 ( AOB, DV2, net044, A, VDDIO, nor_in );
output  AOB, DV2, net044;

input  A, VDDIO, nor_in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nor2 I8 ( .B(DV2), .A(nor_in), .Y(net096));
P_11_LPRVT  PM0 ( .D(DV2), .B(vdd_), .G(net055), .S(vdd_));
P_11_LPRVT  PM1 ( .D(net055), .B(vdd_), .G(DV2), .S(vdd_));
N_25OD33_LP  N1 ( .D(DV2), .B(gnd_), .G(net040), .S(gnd_));
N_25OD33_LP  N0 ( .D(net055), .B(gnd_), .G(net044), .S(gnd_));
inv I9 ( .A(net096), .Y(AOB));
not IVT0 ( net044, A);
not IVT1 ( net040, net044);

endmodule
// Library - umc40nm_io, Cell - LS1, View - schematic
// LAST TIME SAVED: Aug 11 16:04:31 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module LS1 ( AO, AOB, A, VDDIO );
output  AO, AOB;

input  A, VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25OD33_LP  POFF1 ( .D(AOB), .B(VDDIO), .G(net63), .S(net42));
P_25OD33_LP  PL1 ( .D(net42), .B(VDDIO), .G(AO), .S(VDDIO));
P_25OD33_LP  PL ( .D(net46), .B(VDDIO), .G(AOB), .S(VDDIO));
P_25OD33_LP  POFF ( .D(AO), .B(VDDIO), .G(net063), .S(net46));
N_25OD33_LP  NM0 ( .D(AO), .B(gnd_), .G(AOB), .S(gnd_));
N_25OD33_LP  N1 ( .D(AOB), .B(gnd_), .G(net63), .S(gnd_));
N_25OD33_LP  N0 ( .D(AO), .B(gnd_), .G(net063), .S(gnd_));
inv IIV1 ( .A(net063), .Y(net63));
inv II15 ( .A(A), .Y(net063));

endmodule
// Library - umc40nm_io, Cell - NAND2_25OD33, View - schematic
// LAST TIME SAVED: Aug  9 18:13:12 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module NAND2_25OD33 ( Y, A, B, VDDIO );
output  Y;

input  A, B, VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25OD33_LP  M1 ( .D(Y), .B(gnd_), .G(A), .S(net025));
N_25OD33_LP  M3 ( .D(net025), .B(gnd_), .G(B), .S(gnd_));
P_25OD33_LP  M0 ( .D(Y), .B(VDDIO), .G(A), .S(VDDIO));
P_25OD33_LP  M2 ( .D(Y), .B(VDDIO), .G(B), .S(VDDIO));

endmodule
// Library - umc40nm_io, Cell - LS3U, View - schematic
// LAST TIME SAVED: Aug 26 17:07:37 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module LS3U ( AOB, A, VDDIO );
output  AOB;

input  A, VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25OD33_LP  POFF1 ( .D(AOB), .B(VDDIO), .G(net49), .S(net035));
P_25OD33_LP  PL1 ( .D(net035), .B(VDDIO), .G(net68), .S(VDDIO));
P_25OD33_LP  PL ( .D(net55), .B(VDDIO), .G(AOB), .S(VDDIO));
P_25OD33_LP  POFF ( .D(net68), .B(VDDIO), .G(net45), .S(net55));
N_25OD33_LP  N1 ( .D(AOB), .B(gnd_), .G(net49), .S(gnd_));
N_25OD33_LP  N0 ( .D(net68), .B(gnd_), .G(net45), .S(gnd_));
inv IIV1 ( .A(net45), .Y(net49));
inv I15 ( .A(A), .Y(net45));

endmodule
// Library - umc40nm_io, Cell - SUMB_sbt_HX, View - schematic
// LAST TIME SAVED: Nov 23 09:48:09 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module SUMB_sbt_HX ( DI, PGATE, PAD, DO, IE, OEN, REN, VDDIO, nor_in );
output  DI, PGATE;

inout  PAD;

input  DO, IE, OEN, REN, VDDIO, nor_in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



LS21 I489 ( .A(DO), .AO(DO1), .VDDIO(VDDIO));
LS41 I580 ( .A(DV), .DV2(net_107), .AOB(DI), .VDDIO(VDDIO),
     .net044(net_181), .nor_in(nor_in));
LS1 I493 ( .A(IE), .AOB(net_105), .AO(SMT1), .VDDIO(VDDIO));
LS1 I488 ( .A(OEN), .AOB(net_143), .AO(OE1B_1), .VDDIO(VDDIO));
not INPROUT2_A ( NROUT2_1, NROUT1_1);
not INPROUT1_A ( NROUT1_1, NROUT0_1);
not IPROUT2_A ( PROUT2_1, PROUT1_1);
not IPROUT1_A ( PROUT1_1, PROUT0_1);
nor INROUT0_A ( NROUT0_1, DO1, OE1B_1);
NAND2_25OD33 IPROUT0_A ( .A(DO1), .VDDIO(VDDIO), .Y(PROUT0_1),
     .B(net_143));
NAND2_25OD33 I481 ( .A(OE1B_1), .VDDIO(VDDIO), .Y(net200), .B(PU2));
LS3U I490 ( .A(REN), .AOB(PU2), .VDDIO(VDDIO));
DION_11_LPRVT  D8 ( .PLUS(gnd_), .MINUS(REN));
DION_11_LPRVT  D11 ( .PLUS(gnd_), .MINUS(DO));
DION_11_LPRVT  D10 ( .PLUS(gnd_), .MINUS(IE));
DION_11_LPRVT  D19 ( .PLUS(gnd_), .MINUS(OEN));
N_25OD33_LP  N4 ( .D(gnd_), .B(gnd_), .G(SMT1), .S(net_174));
N_25OD33_LP  N44 ( .D(gnd_), .B(gnd_), .G(gnd_), .S(PGATE));
N_25OD33_LP  Ntiegnd ( .D(PAD), .B(gnd_), .G(gnd_), .S(gnd_));
N_25OD33_LP  NM00 ( .D(PAD), .B(gnd_), .G(NROUT2_1), .S(gnd_));
N_25OD33_LP  N5 ( .D(net_174), .B(gnd_), .G(PGATE), .S(DV));
P_25OD33_LP  PUP1 ( .D(VDDIO), .B(VDDIO), .G(net200), .S(PGATE));
P_25OD33_LP  P40 ( .D(VDDIO), .B(VDDIO), .G(VDDIO), .S(PGATE));
P_25OD33_LP  P2 ( .D(VDDIO), .B(VDDIO), .G(SMT1), .S(DV));
P_25OD33_LP  P0 ( .D(VDDIO), .B(VDDIO), .G(PGATE), .S(DV));
P_25OD33_LP  PM4 ( .D(VDDIO), .B(VDDIO), .G(net_181), .S(DV));
P_25OD33_LP  PM0 ( .D(PAD), .B(VDDIO), .G(PROUT2_1), .S(VDDIO));
RNPPO_LP_pcell2460 RRNW0 ( .B(VDDIO), .MINUS(PAD), .PLUS(PGATE));

endmodule
// Library - ice384chip, Cell - IO_top_bank_ice384, View - schematic
// LAST TIME SAVED: Jan  9 18:56:47 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module IO_top_bank_ice384 ( padin_t, pad_t, vpp, vppin, ie, padeb_t,
     pado_t, ren );

inout  vpp, vppin;


output [11:0]  padin_t;

inout [11:0]  pad_t;

input [11:0]  ie;
input [11:0]  ren;
input [11:0]  padeb_t;
input [11:0]  pado_t;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net53;

wire  [3:0]  net62;

wire  [4:0]  net44;



SDDIOBREAK_sbt_a I211 ( .VDDIO(vddp_));
SDDIOBREAK_sbt_a I213 ( .VDDIO(vddio_0));
pvpp vppfast_t ( .vppin(vppin), .vpp(vpp));
SVSS_sbt_a GND_VDDIO_2_1_ ( .VDDIO(vddio_0));
SVSS_sbt_a GND_VDDIO_2_0_ ( .VDDIO(vddio_0));
SVDDIO_sbt_a VDDIO_2_0_ ( .VDDIO(vddio_0));
SVDDIO_sbt_a VDDIO_2_2_ ( .VDDIO(vddio_0));
SVDDIO_sbt_a VDDIO_2_1_ ( .VDDIO(vddio_0));
SVDD_sbt_a VCC_1_ ( );
SVDD_sbt_a VCC_0_ ( );
tielo4x tielo4x ( .tielo(tiegnd_toppad));
SUMB_sbt_HX IO_3_ ( .OEN(padeb_t[3]), .IE(ie[3]), .REN(ren[3]),
     .DO(pado_t[3]), .PAD(pad_t[3]), .DI(padin_t[3]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net62[0]));
SUMB_sbt_HX IO_2_ ( .OEN(padeb_t[2]), .IE(ie[2]), .REN(ren[2]),
     .DO(pado_t[2]), .PAD(pad_t[2]), .DI(padin_t[2]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net62[1]));
SUMB_sbt_HX IO_1_ ( .OEN(padeb_t[1]), .IE(ie[1]), .REN(ren[1]),
     .DO(pado_t[1]), .PAD(pad_t[1]), .DI(padin_t[1]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net62[2]));
SUMB_sbt_HX IO_0_ ( .OEN(padeb_t[0]), .IE(ie[0]), .REN(ren[0]),
     .DO(pado_t[0]), .PAD(pad_t[0]), .DI(padin_t[0]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net62[3]));
SUMB_sbt_HX IO_4_ ( .OEN(padeb_t[4]), .IE(ie[4]), .REN(ren[4]),
     .DO(pado_t[4]), .PAD(pad_t[4]), .DI(padin_t[4]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net35));
SUMB_sbt_HX IO_11_ ( .OEN(padeb_t[11]), .IE(ie[11]), .REN(ren[11]),
     .DO(pado_t[11]), .PAD(pad_t[11]), .DI(padin_t[11]),
     .VDDIO(vddio_0), .nor_in(tiegnd_toppad), .PGATE(net44[0]));
SUMB_sbt_HX IO_10_ ( .OEN(padeb_t[10]), .IE(ie[10]), .REN(ren[10]),
     .DO(pado_t[10]), .PAD(pad_t[10]), .DI(padin_t[10]),
     .VDDIO(vddio_0), .nor_in(tiegnd_toppad), .PGATE(net44[1]));
SUMB_sbt_HX IO_9_ ( .OEN(padeb_t[9]), .IE(ie[9]), .REN(ren[9]),
     .DO(pado_t[9]), .PAD(pad_t[9]), .DI(padin_t[9]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net44[2]));
SUMB_sbt_HX IO_8_ ( .OEN(padeb_t[8]), .IE(ie[8]), .REN(ren[8]),
     .DO(pado_t[8]), .PAD(pad_t[8]), .DI(padin_t[8]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net44[3]));
SUMB_sbt_HX IO_7_ ( .OEN(padeb_t[7]), .IE(ie[7]), .REN(ren[7]),
     .DO(pado_t[7]), .PAD(pad_t[7]), .DI(padin_t[7]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net44[4]));
SUMB_sbt_HX IO_6_ ( .OEN(padeb_t[6]), .IE(ie[6]), .REN(ren[6]),
     .DO(pado_t[6]), .PAD(pad_t[6]), .DI(padin_t[6]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net53[0]));
SUMB_sbt_HX IO_5_ ( .OEN(padeb_t[5]), .IE(ie[5]), .REN(ren[5]),
     .DO(pado_t[5]), .PAD(pad_t[5]), .DI(padin_t[5]), .VDDIO(vddio_0),
     .nor_in(tiegnd_toppad), .PGATE(net53[1]));

endmodule
// Library - umc40nm_io, Cell - SUMB_sbt_8mA_PD, View - schematic
// LAST TIME SAVED: Sep 26 17:00:22 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module SUMB_sbt_8mA_PD ( DI, PGATE, PAD, DO, IE, OEN, REN, VDDIO,
     nor_in );
output  DI, PGATE;

inout  PAD;

input  DO, IE, OEN, REN, VDDIO, nor_in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



RNPPO_LP_pcell2460 RRNW0 ( .B(VDDIO), .MINUS(PAD), .PLUS(PGATE));
P_25OD33_LP  P40 ( .D(VDDIO), .B(VDDIO), .G(VDDIO), .S(PGATE));
P_25OD33_LP  P2 ( .D(VDDIO), .B(VDDIO), .G(SMT1), .S(DV));
P_25OD33_LP  PM1 ( .D(PAD), .B(VDDIO), .G(VDDIO), .S(VDDIO));
P_25OD33_LP  P0 ( .D(VDDIO), .B(VDDIO), .G(PGATE), .S(DV));
P_25OD33_LP  PM4 ( .D(VDDIO), .B(VDDIO), .G(net_132), .S(DV));
P_25OD33_LP  PM0 ( .D(PAD), .B(VDDIO), .G(PROUT2_1), .S(VDDIO));
N_25OD33_LP  NM0 ( .D(gnd_), .B(gnd_), .G(net200), .S(PGATE));
N_25OD33_LP  N4 ( .D(gnd_), .B(gnd_), .G(SMT1), .S(net_153));
N_25OD33_LP  N44 ( .D(gnd_), .B(gnd_), .G(gnd_), .S(PGATE));
N_25OD33_LP  Ntiegnd ( .D(PAD), .B(gnd_), .G(gnd_), .S(gnd_));
N_25OD33_LP  NM00 ( .D(PAD), .B(gnd_), .G(NROUT2_1), .S(gnd_));
N_25OD33_LP  N5 ( .D(net_153), .B(gnd_), .G(PGATE), .S(DV));
DION_11_LPRVT  D19 ( .PLUS(gnd_), .MINUS(OEN));
DION_11_LPRVT  D8 ( .PLUS(gnd_), .MINUS(REN));
DION_11_LPRVT  D11 ( .PLUS(gnd_), .MINUS(DO));
DION_11_LPRVT  D10 ( .PLUS(gnd_), .MINUS(IE));
LS3U I490 ( .A(REN), .AOB(PU2), .VDDIO(VDDIO));
NAND2_25OD33 IPROUT0_A ( .A(DO1), .VDDIO(VDDIO), .Y(PROUT0_1),
     .B(net_176));
NAND2_25OD33 I481 ( .A(OE1B_1), .VDDIO(VDDIO), .Y(net_0180), .B(PU2));
nor INROUT0_A ( NROUT0_1, DO1, OE1B_1);
not INPROUT2_A ( NROUT2_1, NROUT1_1);
not IPROUT1_A ( PROUT1_1, PROUT0_1);
not I78 ( net200, net_0180);
not INPROUT1_A ( NROUT1_1, NROUT0_1);
not IPROUT2_A ( PROUT2_1, PROUT1_1);
LS1 I493 ( .A(IE), .AOB(net_208), .AO(SMT1), .VDDIO(VDDIO));
LS1 I488 ( .A(OEN), .AOB(net_176), .AO(OE1B_1), .VDDIO(VDDIO));
LS41 I580 ( .A(DV), .DV2(net_202), .AOB(DI), .VDDIO(VDDIO),
     .net044(net_132), .nor_in(nor_in));
LS21 I489 ( .A(DO), .AO(DO1), .VDDIO(VDDIO));

endmodule
// Library - umc40nm_io, Cell - SCORNER_sbt_a, View - schematic
// LAST TIME SAVED: Jan 17 18:29:57 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module SCORNER_sbt_a ( VDDIO );
input  VDDIO;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



DIOP_25_LP  D1 ( .PLUS(gnd_), .MINUS(VDDIO));
P_25OD33_LP  PM3 ( .D(net_1260), .B(VDDIO), .G(net_1259), .S(VDDIO));
N_25OD33_LP  NM2 ( .D(VDDIO), .B(gnd_), .G(net_1260), .S(gnd_));
N_25OD33_LP  NM0 ( .D(gnd_), .B(gnd_), .G(net_1259), .S(gnd_));
N_25OD33_LP  NM1 ( .D(net_1260), .B(gnd_), .G(net_1259), .S(gnd_));
RNPPO_LP_pcell2461 R0 ( .B(vdd_), .MINUS(net39), .PLUS(VDDIO));
RNPPO_LP_pcell2462 R2 ( .B(gnd_), .MINUS(net36), .PLUS(net39));
RNPPO_LP_pcell2462 R3 ( .B(VDDIO), .MINUS(net_1259), .PLUS(net36));

endmodule
// Library - leafcell, Cell - tiehi4x, View - schematic
// LAST TIME SAVED: Aug  3 19:21:04 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module tiehi4x ( tiehi );
output  tiehi;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));
N_11_LPHVT  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd2vdd25, View - schematic
// LAST TIME SAVED: Aug  3 19:29:06 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M1 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
P_25_LP  M2 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
P_25_LP  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));
P_25_LP  M0 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
N_25_LP  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
N_25_LP  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_bgen, View - schematic
// LAST TIME SAVED: Aug  3 19:29:11 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_testdec_bgen ( dec_ok, dec_bias, dec_det, testdec_en_b,
     testdec_prec_b );
output  dec_ok;

inout  dec_bias, dec_det;

input  testdec_en_b, testdec_prec_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPRVT  M16 ( .D(net76), .B(vdd_), .G(testdec_en_b), .S(vdd_));
P_11_LPRVT  M18_1_ ( .D(dec_bias_sup), .B(vdd_), .G(testdec_en_b),
     .S(vdd_));
P_11_LPRVT  M18_0_ ( .D(dec_bias_sup), .B(vdd_), .G(testdec_en_b),
     .S(vdd_));
P_11_LPRVT  M9_2_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p),
     .S(dec_bias_sup));
P_11_LPRVT  M9_1_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p),
     .S(dec_bias_sup));
P_11_LPRVT  M9_0_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p),
     .S(dec_bias_sup));
P_11_LPRVT  M19 ( .D(ngate), .B(vdd_), .G(testdec_en_b), .S(net76));
P_11_LPRVT  M8 ( .D(dec_bias_p), .B(vdd_), .G(dec_bias_p),
     .S(dec_bias_sup));
N_11_LPRVT  M13 ( .D(dec_bias), .B(GND_), .G(testdec_en_b), .S(gnd_));
N_11_LPRVT  M6 ( .D(dec_bias), .B(GND_), .G(dec_bias), .S(gnd_));
N_11_LPRVT  M7 ( .D(dec_bias_p), .B(GND_), .G(dec_bias), .S(gnd_));
N_11_LPRVT  M14 ( .D(ngate), .B(GND_), .G(dec_bias), .S(gnd_));
N_11_LPRVT  M15 ( .D(ngate), .B(GND_), .G(testdec_en_b), .S(gnd_));
N_11_LPRVT  M10 ( .D(dec_bias_sup), .B(GND_), .G(ngate), .S(dec_bias));
P_11_LPHVT  M0 ( .D(dec_det), .B(vdd_), .G(testdec_prec_b), .S(vdd_));
N_11_LPHVT  M4 ( .D(dec_det), .B(GND_), .G(testdec_en_b), .S(gnd_));
inv_hvt I134 ( .A(dec_det), .Y(dec_ok));

endmodule
// Library - ice384chip, Cell - IO_rgt_bank_ice384, View - schematic
// LAST TIME SAVED: Jan  9 18:47:44 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module IO_rgt_bank_ice384 ( padin_r, trstb_int, pad_r, TRSTb, ie,
     padeb_r, pado_r, ren );
output  trstb_int;


input  TRSTb;

output [15:0]  padin_r;

inout [15:0]  pad_r;

input [16:0]  ren;
input [15:0]  pado_r;
input [15:0]  padeb_r;
input [15:0]  ie;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net79;

wire  [3:0]  net32;

wire  [6:0]  net31;



SUMB_sbt_8mA_PD I213 ( .OEN(tievdd_rgtpad), .IE(tievdd_rgtpad),
     .REN(ren[16]), .DO(tignd_rgtpad), .PAD(TRSTb), .DI(trstb_int),
     .VDDIO(vddio_1), .PGATE(net33), .nor_in(tignd_rgtpad));
SDDIOBREAK_sbt_a PCT ( .VDDIO(vddio_1));
SCORNER_sbt_a PC_R_TOP ( .VDDIO(vddp_));
SCORNER_sbt_a PC_R_BOT ( .VDDIO(vddio_1));
SVSS_sbt_a GND_VDDIOR_1_ ( .VDDIO(vddio_1));
SVSS_sbt_a GND_VDDIOR_0_ ( .VDDIO(vddio_1));
SVDDIO_sbt_a VDDIO ( .VDDIO(vddp_));
SVDDIO_sbt_a VDDIO_2_1_ ( .VDDIO(vddio_1));
SVDDIO_sbt_a VDDIO_2_0_ ( .VDDIO(vddio_1));
tiehi4x tiehi4x ( .tiehi(tievdd_rgtpad));
tielo4x tielo4x ( .tielo(tignd_rgtpad));
SUMB_sbt_HX IO_3_ ( .OEN(padeb_r[3]), .IE(ie[3]), .REN(ren[3]),
     .DO(pado_r[3]), .PAD(pad_r[3]), .DI(padin_r[3]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net32[0]));
SUMB_sbt_HX IO_2_ ( .OEN(padeb_r[2]), .IE(ie[2]), .REN(ren[2]),
     .DO(pado_r[2]), .PAD(pad_r[2]), .DI(padin_r[2]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net32[1]));
SUMB_sbt_HX IO_1_ ( .OEN(padeb_r[1]), .IE(ie[1]), .REN(ren[1]),
     .DO(pado_r[1]), .PAD(pad_r[1]), .DI(padin_r[1]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net32[2]));
SUMB_sbt_HX IO_0_ ( .OEN(padeb_r[0]), .IE(ie[0]), .REN(ren[0]),
     .DO(pado_r[0]), .PAD(pad_r[0]), .DI(padin_r[0]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net32[3]));
SUMB_sbt_HX IO_4_ ( .OEN(padeb_r[4]), .IE(ie[4]), .REN(ren[4]),
     .DO(pado_r[4]), .PAD(pad_r[4]), .DI(padin_r[4]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net30));
SUMB_sbt_HX IO_15_ ( .OEN(padeb_r[15]), .IE(ie[15]), .REN(ren[15]),
     .DO(pado_r[15]), .PAD(pad_r[15]), .DI(padin_r[15]),
     .VDDIO(vddio_1), .nor_in(tignd_rgtpad), .PGATE(net31[0]));
SUMB_sbt_HX IO_14_ ( .OEN(padeb_r[14]), .IE(ie[14]), .REN(ren[14]),
     .DO(pado_r[14]), .PAD(pad_r[14]), .DI(padin_r[14]),
     .VDDIO(vddio_1), .nor_in(tignd_rgtpad), .PGATE(net31[1]));
SUMB_sbt_HX IO_13_ ( .OEN(padeb_r[13]), .IE(ie[13]), .REN(ren[13]),
     .DO(pado_r[13]), .PAD(pad_r[13]), .DI(padin_r[13]),
     .VDDIO(vddio_1), .nor_in(tignd_rgtpad), .PGATE(net31[2]));
SUMB_sbt_HX IO_12_ ( .OEN(padeb_r[12]), .IE(ie[12]), .REN(ren[12]),
     .DO(pado_r[12]), .PAD(pad_r[12]), .DI(padin_r[12]),
     .VDDIO(vddio_1), .nor_in(tignd_rgtpad), .PGATE(net31[3]));
SUMB_sbt_HX IO_11_ ( .OEN(padeb_r[11]), .IE(ie[11]), .REN(ren[11]),
     .DO(pado_r[11]), .PAD(pad_r[11]), .DI(padin_r[11]),
     .VDDIO(vddio_1), .nor_in(tignd_rgtpad), .PGATE(net31[4]));
SUMB_sbt_HX IO_10_ ( .OEN(padeb_r[10]), .IE(ie[10]), .REN(ren[10]),
     .DO(pado_r[10]), .PAD(pad_r[10]), .DI(padin_r[10]),
     .VDDIO(vddio_1), .nor_in(tignd_rgtpad), .PGATE(net31[5]));
SUMB_sbt_HX IO_9_ ( .OEN(padeb_r[9]), .IE(ie[9]), .REN(ren[9]),
     .DO(pado_r[9]), .PAD(pad_r[9]), .DI(padin_r[9]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net31[6]));
SUMB_sbt_HX IO_8_ ( .OEN(padeb_r[8]), .IE(ie[8]), .REN(ren[8]),
     .DO(pado_r[8]), .PAD(pad_r[8]), .DI(padin_r[8]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net79[0]));
SUMB_sbt_HX IO_7_ ( .OEN(padeb_r[7]), .IE(ie[7]), .REN(ren[7]),
     .DO(pado_r[7]), .PAD(pad_r[7]), .DI(padin_r[7]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net79[1]));
SUMB_sbt_HX IO_6_ ( .OEN(padeb_r[6]), .IE(ie[6]), .REN(ren[6]),
     .DO(pado_r[6]), .PAD(pad_r[6]), .DI(padin_r[6]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net79[2]));
SUMB_sbt_HX IO_5_ ( .OEN(padeb_r[5]), .IE(ie[5]), .REN(ren[5]),
     .DO(pado_r[5]), .PAD(pad_r[5]), .DI(padin_r[5]), .VDDIO(vddio_1),
     .nor_in(tignd_rgtpad), .PGATE(net79[3]));

endmodule
// Library - ice384chip, Cell - io_r2rinbuf_comptbl, View - schematic
// LAST TIME SAVED: Oct  9 20:55:59 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module io_r2rinbuf_comptbl ( out, vddio, cbit[2], cbit[3], cbit[4],
     in_neg_25, in_pos_25, tiegnd );
output  out;

inout  vddio;

input  in_neg_25, in_pos_25, tiegnd;

input [4:2]  cbit;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M36 ( .D(net085), .B(GND_), .G(tiegnd), .S(net152));
N_25_LP  M28 ( .D(net152), .B(GND_), .G(en_25), .S(net137));
N_25_LP  M30 ( .D(net137), .B(GND_), .G(en_25), .S(gnd_));
N_25_LP  X13 ( .D(net0141), .B(GND_), .G(in_pos_25), .S(net152));
N_25_LP  M31 ( .D(net0182), .B(GND_), .G(tiegnd), .S(net0141));
N_25_LP  M34 ( .D(net087), .B(GND_), .G(tiegnd), .S(net152));
N_25_LP  M35 ( .D(net086), .B(GND_), .G(tiegnd), .S(net145));
N_25_LP  M27 ( .D(net145), .B(GND_), .G(in_neg_25), .S(net152));
P_25_LP  M13 ( .D(sa_out), .B(vddio), .G(net145), .S(vddio));
P_25_LP  M17 ( .D(net105), .B(net126), .G(in_neg_25), .S(net126));
P_25_LP  M19 ( .D(net126), .B(vddio), .G(en_b_25), .S(vddio));
P_25_LP  M7 ( .D(net0141), .B(vddio), .G(net0141), .S(vddio));
P_25_LP  M6 ( .D(net105), .B(vddio), .G(net0141), .S(vddio));
P_25_LP  M18 ( .D(sa_out), .B(net126), .G(in_pos_25), .S(net126));
P_25_LP  M5 ( .D(net145), .B(vddio), .G(net145), .S(vddio));
N_11_LPHVT  M22 ( .D(net105), .B(GND_), .G(tiegnd), .S(net0113));
N_11_LPHVT  M20 ( .D(sa_out), .B(GND_), .G(sa_out), .S(sa_out_inv));
N_11_LPHVT  M23 ( .D(sa_out), .B(GND_), .G(tiegnd), .S(net0117));
N_11_LPHVT  M11 ( .D(sa_out), .B(gnd_), .G(net105), .S(gnd_));
N_11_LPHVT  M16 ( .D(net105), .B(gnd_), .G(net105), .S(gnd_));
N_11_LPHVT  M21 ( .D(sa_out_inv), .B(gnd_), .G(sa_out), .S(gnd_));
nor3_hvt I56 ( .B(net081), .Y(net78), .A(cbit[3]), .C(cbit[2]));
ml_ls_vdd2vdd25 I173 ( .in(net78), .sup(vddio), .out_vddio_b(en_b_25),
     .out_vddio(en_25), .in_b(net82));
inv_hvt I298 ( .A(net86), .Y(out));
inv_hvt I295 ( .A(net78), .Y(net82));
inv_hvt I296 ( .A(net82), .Y(sa_out_inv));
inv_hvt I55 ( .A(cbit[4]), .Y(net081));
inv_hvt I66 ( .A(sa_out_inv), .Y(net86));

endmodule
// Library - ice384chip, Cell - PLVDS_pair_HX, View - schematic
// LAST TIME SAVED: Dec  6 14:01:26 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module PLVDS_pair_HX ( c_n, c_p, PAD_n, PAD_p, cbit, i_n, i_p, oen_n,
     oen_p, tiegnd, vddio );
output  c_n, c_p;

inout  PAD_n, PAD_p;

input  i_n, i_p, oen_n, oen_p, tiegnd, vddio;

input [4:0]  cbit;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



io_r2rinbuf_comptbl r2r_buf ( indiff, vddio, cbit[3], cbit[2], cbit[4],
     in_padn_1, in_padp_0, tiegnd);
SUMB_sbt_HX I_ppart_0 ( .OEN(oen_p), .IE(cbit[3]), .REN(cbit[1]),
     .DO(i_p), .PAD(PAD_p), .DI(c_p), .VDDIO(vddio), .nor_in(indiff),
     .PGATE(in_padp_0));
SUMB_sbt_HX I_npart_1 ( .DO(i_n), .DI(c_n), .nor_in(tiegnd),
     .PGATE(in_padn_1), .IE(cbit[2]), .VDDIO(vddio), .REN(cbit[0]),
     .PAD(PAD_n), .OEN(oen_n));

endmodule
// Library - ice384chip, Cell - IO_lft_bank_ice384, View - schematic
// LAST TIME SAVED: Jan 17 11:40:04 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module IO_lft_bank_ice384 ( padin_l, pad_l, ie, lvds_en, padeb_l,
     pado_l, ren );



output [15:0]  padin_l;

inout [15:0]  pad_l;

input [15:0]  ren;
input [15:0]  ie;
input [7:0]  lvds_en;
input [15:0]  pado_l;
input [15:0]  padeb_l;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



SVDD_sbt_a VCC ( );
PLVDS_pair_HX IO_PAIR_1_0 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[0]), .oen_n(padeb_l[1]), .PAD_n(pad_l[1]),
     .c_p(padin_l[0]), .c_n(padin_l[1]), .PAD_p(pad_l[0]),
     .i_n(pado_l[1]), .i_p(pado_l[0]), .cbit({lvds_en[0], ie[0], ie[1],
     ren[0], ren[1]}));
PLVDS_pair_HX IO_PAIR_5_4 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[4]), .oen_n(padeb_l[5]), .PAD_n(pad_l[5]),
     .c_p(padin_l[4]), .c_n(padin_l[5]), .PAD_p(pad_l[4]),
     .i_n(pado_l[5]), .i_p(pado_l[4]), .cbit({lvds_en[2], ie[4], ie[5],
     ren[4], ren[5]}));
PLVDS_pair_HX IO_PAIR_3_2 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[2]), .oen_n(padeb_l[3]), .PAD_n(pad_l[3]),
     .c_p(padin_l[2]), .c_n(padin_l[3]), .PAD_p(pad_l[2]),
     .i_n(pado_l[3]), .i_p(pado_l[2]), .cbit({lvds_en[1], ie[2], ie[3],
     ren[2], ren[3]}));
PLVDS_pair_HX IO_PAIR_9_8 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[8]), .oen_n(padeb_l[9]), .PAD_n(pad_l[9]),
     .c_p(padin_l[8]), .c_n(padin_l[9]), .PAD_p(pad_l[8]),
     .i_n(pado_l[9]), .i_p(pado_l[8]), .cbit({lvds_en[4], ie[8], ie[9],
     ren[8], ren[9]}));
PLVDS_pair_HX IO_PAIR_11_10 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[10]), .oen_n(padeb_l[11]), .PAD_n(pad_l[11]),
     .c_p(padin_l[10]), .c_n(padin_l[11]), .PAD_p(pad_l[10]),
     .i_n(pado_l[11]), .i_p(pado_l[10]), .cbit({lvds_en[5], ie[10],
     ie[11], ren[10], ren[11]}));
PLVDS_pair_HX IO_PAIR_13_12 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[12]), .oen_n(padeb_l[13]), .PAD_n(pad_l[13]),
     .c_p(padin_l[12]), .c_n(padin_l[13]), .PAD_p(pad_l[12]),
     .i_n(pado_l[13]), .i_p(pado_l[12]), .cbit({lvds_en[6], ie[12],
     ie[13], ren[12], ren[13]}));
PLVDS_pair_HX IO_PAIR_15_14 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[14]), .oen_n(padeb_l[15]), .PAD_n(pad_l[15]),
     .c_p(padin_l[14]), .c_n(padin_l[15]), .PAD_p(pad_l[14]),
     .i_n(pado_l[15]), .i_p(pado_l[14]), .cbit({lvds_en[7], ie[14],
     ie[15], ren[14], ren[15]}));
PLVDS_pair_HX IO_PAIR_7_6 ( .tiegnd(tignd_lftpad), .vddio(vddio_3),
     .oen_p(padeb_l[6]), .oen_n(padeb_l[7]), .PAD_n(pad_l[7]),
     .c_p(padin_l[6]), .c_n(padin_l[7]), .PAD_p(pad_l[6]),
     .i_n(pado_l[7]), .i_p(pado_l[6]), .cbit({lvds_en[3], ie[6], ie[7],
     ren[6], ren[7]}));
SCORNER_sbt_a CRNER_BOT_LFT ( .VDDIO(vddio_3));
SCORNER_sbt_a CRNER_TOP_LFT ( .VDDIO(vddio_3));
SVSS_sbt_a GND_2 ( .VDDIO(vddio_3));
SVSS_sbt_a GND ( .VDDIO(vddio_3));
SVDDIO_sbt_a VDDIO_1 ( .VDDIO(vddio_3));
SVDDIO_sbt_a VCCIO_2 ( .VDDIO(vddio_3));
tielo4x tielo4x ( .tielo(tignd_lftpad));

endmodule
// Library - ice384chip, Cell - IO_bot_bank_ice384, View - schematic
// LAST TIME SAVED: Jan 17 11:40:45 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module IO_bot_bank_ice384 ( cdone_int, creset_b_int, padin_b, cdone,
     pad_b, vddio_2, vddio_spi, cdone_out, creset_b, ie, padeb_b,
     pado_b, ren );
output  cdone_int, creset_b_int;

inout  cdone, vddio_2, vddio_spi;

input  cdone_out, creset_b;

output [11:0]  padin_b;

inout [11:0]  pad_b;

input [11:0]  ie;
input [11:0]  pado_b;
input [11:0]  ren;
input [11:0]  padeb_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  net45;

wire  [1:0]  net72;

wire  [1:0]  net36;

wire  [1:0]  net81;



SDDIOBREAK_sbt_a I211 ( .VDDIO(vddio_spi));
SDDIOBREAK_sbt_a I207 ( .VDDIO(vddio_2));
SDDIOBREAK_sbt_a I205 ( .VDDIO(vddio_2));
SVSS_sbt_a GND_VDDIO_2 ( .VDDIO(vddio_2));
SVSS_sbt_a GND_SPI ( .VDDIO(vddio_spi));
SVDDIO_sbt_a VDDIO_2_1_ ( .VDDIO(vddio_2));
SVDDIO_sbt_a VDDIO_2_0_ ( .VDDIO(vddio_2));
SVDDIO_sbt_a VDDIO_SPI ( .VDDIO(vddio_spi));
SVDD_sbt_a VCC_1_ ( );
SVDD_sbt_a VCC_0_ ( );
tiehi4x tiehi4x ( .tiehi(tievdd_botpad));
tielo4x tielo4x ( .tielo(tiegnd_botpad));
SUMB_sbt_HX IO_5_ ( .OEN(padeb_b[5]), .IE(ie[5]), .REN(ren[5]),
     .DO(pado_b[5]), .PAD(pad_b[5]), .DI(padin_b[5]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net45[0]));
SUMB_sbt_HX IO_4_ ( .OEN(padeb_b[4]), .IE(ie[4]), .REN(ren[4]),
     .DO(pado_b[4]), .PAD(pad_b[4]), .DI(padin_b[4]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net45[1]));
SUMB_sbt_HX IO_3_ ( .OEN(padeb_b[3]), .IE(ie[3]), .REN(ren[3]),
     .DO(pado_b[3]), .PAD(pad_b[3]), .DI(padin_b[3]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net45[2]));
SUMB_sbt_HX IO_2_ ( .OEN(padeb_b[2]), .IE(ie[2]), .REN(ren[2]),
     .DO(pado_b[2]), .PAD(pad_b[2]), .DI(padin_b[2]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net45[3]));
SUMB_sbt_HX IO_1_ ( .OEN(padeb_b[1]), .IE(ie[1]), .REN(ren[1]),
     .DO(pado_b[1]), .PAD(pad_b[1]), .DI(padin_b[1]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net45[4]));
SUMB_sbt_HX IO_0_ ( .OEN(padeb_b[0]), .IE(ie[0]), .REN(ren[0]),
     .DO(pado_b[0]), .PAD(pad_b[0]), .DI(padin_b[0]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net45[5]));
SUMB_sbt_HX IO_CONE ( .OEN(cdone_out), .IE(tievdd_botpad),
     .REN(tiegnd_botpad), .DO(tiegnd_botpad), .PAD(cdone),
     .DI(cdone_int), .VDDIO(vddio_2), .nor_in(tiegnd_botpad),
     .PGATE(net052));
SUMB_sbt_HX IO_CRST ( .OEN(tievdd_botpad), .IE(tievdd_botpad),
     .REN(tiegnd_botpad), .DO(tiegnd_botpad), .PAD(creset_b),
     .DI(creset_b_int), .VDDIO(vddio_2), .nor_in(tiegnd_botpad),
     .PGATE(net061));
SUMB_sbt_HX IO_9_ ( .OEN(padeb_b[9]), .IE(ie[9]), .REN(ren[9]),
     .DO(pado_b[9]), .PAD(pad_b[9]), .DI(padin_b[9]),
     .VDDIO(vddio_spi), .nor_in(tiegnd_botpad), .PGATE(net72[0]));
SUMB_sbt_HX IO_8_ ( .OEN(padeb_b[8]), .IE(ie[8]), .REN(ren[8]),
     .DO(pado_b[8]), .PAD(pad_b[8]), .DI(padin_b[8]),
     .VDDIO(vddio_spi), .nor_in(tiegnd_botpad), .PGATE(net72[1]));
SUMB_sbt_HX IO_11_ ( .OEN(padeb_b[11]), .IE(ie[11]), .REN(ren[11]),
     .DO(pado_b[11]), .PAD(pad_b[11]), .DI(padin_b[11]),
     .VDDIO(vddio_spi), .nor_in(tiegnd_botpad), .PGATE(net36[0]));
SUMB_sbt_HX IO_10_ ( .OEN(padeb_b[10]), .IE(ie[10]), .REN(ren[10]),
     .DO(pado_b[10]), .PAD(pad_b[10]), .DI(padin_b[10]),
     .VDDIO(vddio_spi), .nor_in(tiegnd_botpad), .PGATE(net36[1]));
SUMB_sbt_HX IO_7_ ( .OEN(padeb_b[7]), .IE(ie[7]), .REN(ren[7]),
     .DO(pado_b[7]), .PAD(pad_b[7]), .DI(padin_b[7]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net81[0]));
SUMB_sbt_HX IO_6_ ( .OEN(padeb_b[6]), .IE(ie[6]), .REN(ren[6]),
     .DO(pado_b[6]), .PAD(pad_b[6]), .DI(padin_b[6]), .VDDIO(vddio_2),
     .nor_in(tiegnd_botpad), .PGATE(net81[1]));

endmodule
// Library - ice384chip, Cell - padring_ice384, View - schematic
// LAST TIME SAVED: Jan  3 16:45:18 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module padring_ice384 ( cdone_int, creset_b_int, padin_b, padin_l,
     padin_r, padin_t, trstb_int, cdone, pad_b, pad_l, pad_r, pad_t,
     vddio_23, vddio_spi, vpp, vppin, TRSTb, cdone_out, creset_b, ie_b,
     ie_l, ie_r, ie_t, lvds_en, padeb_b, padeb_l, padeb_r, padeb_t,
     pado_b, pado_l, pado_r, pado_t, ren_b, ren_l, ren_r, ren_t );
output  cdone_int, creset_b_int, trstb_int;

inout  cdone, vddio_23, vddio_spi, vpp, vppin;

input  TRSTb, cdone_out, creset_b;

output [15:0]  padin_r;
output [15:0]  padin_l;
output [11:0]  padin_b;
output [11:0]  padin_t;

inout [15:0]  pad_l;
inout [11:0]  pad_t;
inout [15:0]  pad_r;
inout [11:0]  pad_b;

input [15:0]  pado_l;
input [11:0]  ren_t;
input [7:0]  lvds_en;
input [15:0]  pado_r;
input [11:0]  padeb_b;
input [11:0]  ren_b;
input [16:0]  ren_r;
input [15:0]  ie_r;
input [15:0]  ie_l;
input [11:0]  ie_t;
input [11:0]  ie_b;
input [11:0]  pado_t;
input [15:0]  padeb_l;
input [15:0]  ren_l;
input [11:0]  padeb_t;
input [15:0]  padeb_r;
input [11:0]  pado_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



IO_top_bank_ice384 IO_TOP_BANK ( .ren(ren_t[11:0]),
     .pado_t(pado_t[11:0]), .padeb_t(padeb_t[11:0]), .ie(ie_t[11:0]),
     .padin_t(padin_t[11:0]), .vppin(vppin), .vpp(vpp),
     .pad_t(pad_t[11:0]));
IO_rgt_bank_ice384 IO_RGT_BANK ( .ren(ren_r[16:0]),
     .pado_r(pado_r[15:0]), .padeb_r(padeb_r[15:0]), .ie(ie_r[15:0]),
     .TRSTb(TRSTb), .trstb_int(trstb_int), .padin_r(padin_r[15:0]),
     .pad_r(pad_r[15:0]));
IO_lft_bank_ice384 IO_LEFT_BANK ( .lvds_en(lvds_en[7:0]),
     .ren(ren_l[15:0]), .pado_l(pado_l[15:0]), .padeb_l(padeb_l[15:0]),
     .ie(ie_l[15:0]), .padin_l(padin_l[15:0]), .pad_l(pad_l[15:0]));
IO_bot_bank_ice384 IO_BOT_BANK ( .vddio_2(vddio_23),
     .creset_b_int(creset_b_int), .creset_b(creset_b),
     .ren(ren_b[11:0]), .pado_b(pado_b[11:0]), .cdone_out(cdone_out),
     .padeb_b(padeb_b[11:0]), .ie(ie_b[11:0]), .padin_b(padin_b[11:0]),
     .cdone_int(cdone_int), .vddio_spi(vddio_spi), .pad_b(pad_b[11:0]),
     .cdone(cdone));

endmodule
// Library - ice384chip, Cell - ring_route_ice384, View - schematic
// LAST TIME SAVED: Dec 14 15:09:34 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module ring_route_ice384 ( bs_en0, ceb0, end_of_startup, gint_hz, gsr,
     hiz_b0, j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, .cdsNet0(last_rsr[1]),
     .cdsNet0(last_rsr[0]), .cdsNet0(last_rsr[3]),
     .cdsNet0(last_rsr[2]), md_spi_b, mode0, mux_jtag_sel_b, padin_b,
     padin_l, padin_r, padin_t, pgate_l, pgate_r, reset_b_l, reset_b_r,
     sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, trstb_pad, update0, vdd_cntl_l,
     vdd_cntl_r, wl_l, wl_r, bl_bot, bl_top, cdone, pad_b, pad_l,
     pad_r, pad_t, vpp, creset_b, fromsdo, ie_b, ie_l, ie_r, ie_t,
     lvds_en, padeb_b, padeb_l, padeb_r, padeb_t, pado_b, pado_l,
     pado_r, pado_t, ren_b, ren_l, ren_r, ren_t, spi_ss_in_bbank,
     tck_pad, tdi_pad, tms_pad, trstb );
output  bs_en0, ceb0, end_of_startup, gint_hz, gsr, hiz_b0, j_tck,
     j_tdi, jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, mux_jtag_sel_b, sdo_enable, shift0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, totdopad, trstb_pad, update0;

inout  cdone, vpp;

input  creset_b, fromsdo, tck_pad, tdi_pad, tms_pad, trstb;

output [11:0]  padin_t;
output [159:0]  reset_b_l;
output [159:0]  wl_r;
output [11:0]  padin_b;
output [159:0]  vdd_cntl_l;
output [15:0]  padin_r;
output [159:0]  reset_b_r;
output [159:0]  vdd_cntl_r;
output [159:0]  pgate_l;
output [15:0]  padin_l;
output [159:0]  pgate_r;
output [159:0]  wl_l;
output [3:0]  last_rsr;

inout [363:0]  bl_bot;
inout [11:0]  pad_t;
inout [15:0]  pad_l;
inout [363:0]  bl_top;
inout [15:0]  pad_r;
inout [11:0]  pad_b;

input [4:0]  spi_ss_in_bbank;
input [7:0]  lvds_en;
input [11:0]  pado_b;
input [11:0]  pado_t;
input [15:0]  ren_l;
input [11:0]  ie_t;
input [11:0]  ren_t;
input [15:0]  padeb_r;
input [15:0]  pado_l;
input [11:0]  padeb_b;
input [16:0]  ren_r;
input [15:0]  padeb_l;
input [15:0]  pado_r;
input [11:0]  ie_b;
input [15:0]  ie_r;
input [11:0]  ren_b;
input [11:0]  padeb_t;
input [15:0]  ie_l;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ring_route00_ice384 I_ring_route00_ice384 ( .wl_r(wl_r[159:0]),
     .wl_l(wl_l[159:0]), .vdd_cntl_r(vdd_cntl_r[159:0]),
     .vdd_cntl_l(vdd_cntl_l[159:0]), .reset_b_r(reset_b_r[159:0]),
     .reset_b_l(reset_b_l[159:0]), .pgate_r(pgate_r[159:0]),
     .pgate_l(pgate_l[159:0]), .bl_top(bl_top[363:0]),
     .bl_bot(bl_bot[363:0]), .spi_ss_in_bbank(spi_ss_in_bbank[4:0]),
     .trstb_pad(trstb_pad), .tms_pad(tms_pad), .tdi_pad(tdi_pad),
     .tck_pad(tck_pad), .fromsdo(fromsdo), .creset_b_int(creset_b_int),
     .vddio_bottombank(vddio_bottombank), .vddio_spi(vddio_spi),
     .cdone_in(cdone_in), .vppin(vppin), .update0(update0),
     .tdo_pad(totdopad), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .spi_clk_out(spi_clk_out), .shift0(shift0),
     .sdo_enable(sdo_enable), .mode0(mode0), .md_spi_b(md_spi_b),
     .last_rsr(last_rsr[3:0]),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .j_tdi(j_tdi), .j_tck(j_tck), .mux_jtag_sel_b(mux_jtag_sel_b),
     .hiz_b0(hiz_b0), .gsr(gsr), .gint_hz(gint_hz),
     .end_of_startup(end_of_startup), .ceb0(ceb0),
     .cdone_out(cdone_out), .bs_en0(bs_en0));
padring_ice384 I_padring_ice384 ( .lvds_en(lvds_en[7:0]),
     .ren_r(ren_r[16:0]), .ren_t(ren_t[11:0]), .ren_l(ren_l[15:0]),
     .ren_b(ren_b[11:0]), .pado_t(pado_t[11:0]), .pado_r(pado_r[15:0]),
     .pado_l(pado_l[15:0]), .pado_b(pado_b[11:0]),
     .padeb_t(padeb_t[11:0]), .padeb_r(padeb_r[15:0]),
     .padeb_l(padeb_l[15:0]), .padeb_b(padeb_b[11:0]),
     .ie_t(ie_t[11:0]), .ie_r(ie_r[15:0]), .ie_l(ie_l[15:0]),
     .ie_b(ie_b[11:0]), .TRSTb(trstb), .trstb_int(trstb_pad),
     .padin_t(padin_t[11:0]), .padin_r(padin_r[15:0]),
     .padin_l(padin_l[15:0]), .padin_b(padin_b[11:0]),
     .pad_t(pad_t[11:0]), .pad_r(pad_r[15:0]), .pad_l(pad_l[15:0]),
     .pad_b(pad_b[11:0]), .vddio_23(vddio_bottombank), .vppin(vppin),
     .creset_b(creset_b), .cdone_out(cdone_out),
     .creset_b_int(creset_b_int), .vpp(vpp), .cdone(cdone),
     .cdone_int(cdone_in), .vddio_spi(vddio_spi));

endmodule
// Library - ice8chip, Cell - clk_quad_buf_ice8p, View - schematic
// LAST TIME SAVED: Aug 12 09:03:48 2010
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module clk_quad_buf_ice8p ( clko, clki );
output  clko;

input  clki;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_lvt I19 ( .A(clkb), .Y(clko));
inv_lvt I22 ( .A(clki), .Y(clkb));

endmodule
// Library - ice8chip, Cell - clk_quad_buf_x8_ice8p, View - schematic
// LAST TIME SAVED: Jun 24 14:46:09 2010
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module clk_quad_buf_x8_ice8p ( clko, clki );


output [7:0]  clko;

input [7:0]  clki;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



clk_quad_buf_ice8p I_clk_quad_buf_ice8p_7_ ( .clki(clki[7]),
     .clko(clko[7]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_6_ ( .clki(clki[6]),
     .clko(clko[6]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_5_ ( .clki(clki[5]),
     .clko(clko[5]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_4_ ( .clki(clki[4]),
     .clko(clko[4]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_3_ ( .clki(clki[3]),
     .clko(clko[3]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_2_ ( .clki(clki[2]),
     .clko(clko[2]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_1_ ( .clki(clki[1]),
     .clko(clko[1]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_0_ ( .clki(clki[0]),
     .clko(clko[0]));

endmodule
// Library - ice384chip, Cell - quad_clk_drv_l, View - schematic
// LAST TIME SAVED: Jan 13 16:45:09 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module quad_clk_drv_l ( glb_in_0, glb_in_1, glb_in_2, glb_in_3, gclk );


output [7:0]  glb_in_1;
output [7:0]  glb_in_3;
output [7:0]  glb_in_0;
output [7:0]  glb_in_2;

input [7:0]  gclk;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net528;



clk_quad_buf_x8_ice8p I397 ( .clko(glb_in_1[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));
clk_quad_buf_x8_ice8p I398 ( .clko(glb_in_0[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));
clk_quad_buf_x8_ice8p I394 ( .clko(glb_in_3[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));
clk_quad_buf_x8_ice8p I395 ( .clko({net528[0], net528[1], net528[2],
     net528[3], net528[4], net528[5], net528[6], net528[7]}),
     .clki(gclk[7:0]));
clk_quad_buf_x8_ice8p I396 ( .clko(glb_in_2[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_logic_8f_sbb, View -
//schematic
// LAST TIME SAVED: Aug  3 19:28:58 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_8f_sbb ( out_hv_winv, out_hv_woinv, in );
output  out_hv_winv, out_hv_woinv;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_pump_a_clkdly I141 ( .in(net262), .out(net270));
ml_pump_a_clkdly I219 ( .in(net266), .out(net268));
ml_ls_vdd2vdd25 I144 ( .in(net266), .sup(vddp_),
     .out_vddio_b(out_hv_winv), .out_vddio(net279), .in_b(net258));
ml_ls_vdd2vdd25 I148 ( .in(net262), .sup(vddp_),
     .out_vddio_b(out_hv_woinv), .out_vddio(net274), .in_b(net255));
nor2_hvt I140 ( .A(net268), .B(in), .Y(net255));
nor2_hvt I227 ( .A(net264), .B(net270), .Y(net258));
inv_hvt I225 ( .A(net258), .Y(net266));
inv_hvt I134 ( .A(in), .Y(net264));
inv_hvt I226 ( .A(net255), .Y(net262));

endmodule
// Library - ice384chip, Cell - quad_clk_drv, View - schematic
// LAST TIME SAVED: Jan 13 16:36:22 2012
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module quad_clk_drv ( glb_in_0, glb_in_1, glb_in_2, glb_in_3, gclk );


output [7:0]  glb_in_0;
output [7:0]  glb_in_3;
output [7:0]  glb_in_2;
output [7:0]  glb_in_1;

input [7:0]  gclk;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net528;



clk_quad_buf_x8_ice8p I397 ( .clko(glb_in_2[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));
clk_quad_buf_x8_ice8p I398 ( .clko(glb_in_3[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));
clk_quad_buf_x8_ice8p I394 ( .clko(glb_in_0[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));
clk_quad_buf_x8_ice8p I395 ( .clko({net528[0], net528[1], net528[2],
     net528[3], net528[4], net528[5], net528[6], net528[7]}),
     .clki(gclk[7:0]));
clk_quad_buf_x8_ice8p I396 ( .clko(glb_in_1[7:0]), .clki({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7]}));

endmodule
// Library - xpmem, Cell - cram2x2, View - schematic
// LAST TIME SAVED: Jul 30 23:15:00 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module cram2x2 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [3:0]  q;
output [3:0]  q_b;

inout [1:0]  bl;

input [1:0]  r_vdd;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



eh_cram_cell_4 I_1_10 ( .q_b(q_b[1]), .q(q[1]), .wl(wl[0]), .bl(bl[1]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I_2_01 ( .q_b(q_b[2]), .q(q[2]), .wl(wl[1]), .bl(bl[0]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));
eh_cram_cell_4 I_0_00 ( .q_b(q_b[0]), .q(q[0]), .wl(wl[0]), .bl(bl[0]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I_3_11 ( .q_b(q_b[3]), .q(q[3]), .wl(wl[1]), .bl(bl[1]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));

endmodule
// Library - ice8chip, Cell - cram_2x2x2_ice8p, View - schematic
// LAST TIME SAVED: Jul 30 23:15:00 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module cram_2x2x2_ice8p ( q, q_b, bl, pgate_l, pgate_r, r_gnd_l,
     r_gnd_r, reset_l, reset_r, wl_l, wl_r );



output [7:0]  q_b;
output [7:0]  q;

inout [3:0]  bl;

input [1:0]  pgate_l;
input [1:0]  wl_r;
input [1:0]  r_gnd_r;
input [1:0]  pgate_r;
input [1:0]  wl_l;
input [1:0]  r_gnd_l;
input [1:0]  reset_l;
input [1:0]  reset_r;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



cram2x2 I_mem_r ( .bl(bl[3:2]), .q_b(q_b[7:4]), .reset(reset_r[1:0]),
     .q(q[7:4]), .wl(wl_r[1:0]), .r_vdd(r_gnd_r[1:0]),
     .pgate(pgate_r[1:0]));
cram2x2 I_mem_l ( .bl(bl[1:0]), .q_b(q_b[3:0]), .reset(reset_l[1:0]),
     .q(q[3:0]), .wl(wl_l[1:0]), .r_vdd(r_gnd_l[1:0]),
     .pgate(pgate_l[1:0]));

endmodule
// Library - ice384chip, Cell - ice384_cram_row78col4, View - schematic
// LAST TIME SAVED: Nov 21 18:40:10 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module ice384_cram_row78col4 ( bl, pgate_l, pgate_r, reset_l, reset_r,
     vdd_cntl_l, vdd_cntl_r, wl_l, wl_r );


inout [3:0]  bl;

input [77:0]  vdd_cntl_l;
input [77:0]  pgate_l;
input [77:0]  reset_l;
input [77:0]  wl_l;
input [77:0]  wl_r;
input [77:0]  vdd_cntl_r;
input [77:0]  reset_r;
input [77:0]  pgate_r;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [77:0]  r_gnd_r;

wire  [77:0]  r_gnd_l;

wire  [311:0]  net40;

wire  [311:0]  net39;



P_11_LPHVT  M0_77_ ( .D(r_gnd_r[77]), .B(vdd_), .G(vdd_cntl_r[77]),
     .S(vdd_));
P_11_LPHVT  M0_76_ ( .D(r_gnd_r[76]), .B(vdd_), .G(vdd_cntl_r[76]),
     .S(vdd_));
P_11_LPHVT  M0_75_ ( .D(r_gnd_r[75]), .B(vdd_), .G(vdd_cntl_r[75]),
     .S(vdd_));
P_11_LPHVT  M0_74_ ( .D(r_gnd_r[74]), .B(vdd_), .G(vdd_cntl_r[74]),
     .S(vdd_));
P_11_LPHVT  M0_73_ ( .D(r_gnd_r[73]), .B(vdd_), .G(vdd_cntl_r[73]),
     .S(vdd_));
P_11_LPHVT  M0_72_ ( .D(r_gnd_r[72]), .B(vdd_), .G(vdd_cntl_r[72]),
     .S(vdd_));
P_11_LPHVT  M0_71_ ( .D(r_gnd_r[71]), .B(vdd_), .G(vdd_cntl_r[71]),
     .S(vdd_));
P_11_LPHVT  M0_70_ ( .D(r_gnd_r[70]), .B(vdd_), .G(vdd_cntl_r[70]),
     .S(vdd_));
P_11_LPHVT  M0_69_ ( .D(r_gnd_r[69]), .B(vdd_), .G(vdd_cntl_r[69]),
     .S(vdd_));
P_11_LPHVT  M0_68_ ( .D(r_gnd_r[68]), .B(vdd_), .G(vdd_cntl_r[68]),
     .S(vdd_));
P_11_LPHVT  M0_67_ ( .D(r_gnd_r[67]), .B(vdd_), .G(vdd_cntl_r[67]),
     .S(vdd_));
P_11_LPHVT  M0_66_ ( .D(r_gnd_r[66]), .B(vdd_), .G(vdd_cntl_r[66]),
     .S(vdd_));
P_11_LPHVT  M0_65_ ( .D(r_gnd_r[65]), .B(vdd_), .G(vdd_cntl_r[65]),
     .S(vdd_));
P_11_LPHVT  M0_64_ ( .D(r_gnd_r[64]), .B(vdd_), .G(vdd_cntl_r[64]),
     .S(vdd_));
P_11_LPHVT  M0_63_ ( .D(r_gnd_r[63]), .B(vdd_), .G(vdd_cntl_r[63]),
     .S(vdd_));
P_11_LPHVT  M0_62_ ( .D(r_gnd_r[62]), .B(vdd_), .G(vdd_cntl_r[62]),
     .S(vdd_));
P_11_LPHVT  M0_61_ ( .D(r_gnd_r[61]), .B(vdd_), .G(vdd_cntl_r[61]),
     .S(vdd_));
P_11_LPHVT  M0_60_ ( .D(r_gnd_r[60]), .B(vdd_), .G(vdd_cntl_r[60]),
     .S(vdd_));
P_11_LPHVT  M0_59_ ( .D(r_gnd_r[59]), .B(vdd_), .G(vdd_cntl_r[59]),
     .S(vdd_));
P_11_LPHVT  M0_58_ ( .D(r_gnd_r[58]), .B(vdd_), .G(vdd_cntl_r[58]),
     .S(vdd_));
P_11_LPHVT  M0_57_ ( .D(r_gnd_r[57]), .B(vdd_), .G(vdd_cntl_r[57]),
     .S(vdd_));
P_11_LPHVT  M0_56_ ( .D(r_gnd_r[56]), .B(vdd_), .G(vdd_cntl_r[56]),
     .S(vdd_));
P_11_LPHVT  M0_55_ ( .D(r_gnd_r[55]), .B(vdd_), .G(vdd_cntl_r[55]),
     .S(vdd_));
P_11_LPHVT  M0_54_ ( .D(r_gnd_r[54]), .B(vdd_), .G(vdd_cntl_r[54]),
     .S(vdd_));
P_11_LPHVT  M0_53_ ( .D(r_gnd_r[53]), .B(vdd_), .G(vdd_cntl_r[53]),
     .S(vdd_));
P_11_LPHVT  M0_52_ ( .D(r_gnd_r[52]), .B(vdd_), .G(vdd_cntl_r[52]),
     .S(vdd_));
P_11_LPHVT  M0_51_ ( .D(r_gnd_r[51]), .B(vdd_), .G(vdd_cntl_r[51]),
     .S(vdd_));
P_11_LPHVT  M0_50_ ( .D(r_gnd_r[50]), .B(vdd_), .G(vdd_cntl_r[50]),
     .S(vdd_));
P_11_LPHVT  M0_49_ ( .D(r_gnd_r[49]), .B(vdd_), .G(vdd_cntl_r[49]),
     .S(vdd_));
P_11_LPHVT  M0_48_ ( .D(r_gnd_r[48]), .B(vdd_), .G(vdd_cntl_r[48]),
     .S(vdd_));
P_11_LPHVT  M0_47_ ( .D(r_gnd_r[47]), .B(vdd_), .G(vdd_cntl_r[47]),
     .S(vdd_));
P_11_LPHVT  M0_46_ ( .D(r_gnd_r[46]), .B(vdd_), .G(vdd_cntl_r[46]),
     .S(vdd_));
P_11_LPHVT  M0_45_ ( .D(r_gnd_r[45]), .B(vdd_), .G(vdd_cntl_r[45]),
     .S(vdd_));
P_11_LPHVT  M0_44_ ( .D(r_gnd_r[44]), .B(vdd_), .G(vdd_cntl_r[44]),
     .S(vdd_));
P_11_LPHVT  M0_43_ ( .D(r_gnd_r[43]), .B(vdd_), .G(vdd_cntl_r[43]),
     .S(vdd_));
P_11_LPHVT  M0_42_ ( .D(r_gnd_r[42]), .B(vdd_), .G(vdd_cntl_r[42]),
     .S(vdd_));
P_11_LPHVT  M0_41_ ( .D(r_gnd_r[41]), .B(vdd_), .G(vdd_cntl_r[41]),
     .S(vdd_));
P_11_LPHVT  M0_40_ ( .D(r_gnd_r[40]), .B(vdd_), .G(vdd_cntl_r[40]),
     .S(vdd_));
P_11_LPHVT  M0_39_ ( .D(r_gnd_r[39]), .B(vdd_), .G(vdd_cntl_r[39]),
     .S(vdd_));
P_11_LPHVT  M0_38_ ( .D(r_gnd_r[38]), .B(vdd_), .G(vdd_cntl_r[38]),
     .S(vdd_));
P_11_LPHVT  M0_37_ ( .D(r_gnd_r[37]), .B(vdd_), .G(vdd_cntl_r[37]),
     .S(vdd_));
P_11_LPHVT  M0_36_ ( .D(r_gnd_r[36]), .B(vdd_), .G(vdd_cntl_r[36]),
     .S(vdd_));
P_11_LPHVT  M0_35_ ( .D(r_gnd_r[35]), .B(vdd_), .G(vdd_cntl_r[35]),
     .S(vdd_));
P_11_LPHVT  M0_34_ ( .D(r_gnd_r[34]), .B(vdd_), .G(vdd_cntl_r[34]),
     .S(vdd_));
P_11_LPHVT  M0_33_ ( .D(r_gnd_r[33]), .B(vdd_), .G(vdd_cntl_r[33]),
     .S(vdd_));
P_11_LPHVT  M0_32_ ( .D(r_gnd_r[32]), .B(vdd_), .G(vdd_cntl_r[32]),
     .S(vdd_));
P_11_LPHVT  M0_31_ ( .D(r_gnd_r[31]), .B(vdd_), .G(vdd_cntl_r[31]),
     .S(vdd_));
P_11_LPHVT  M0_30_ ( .D(r_gnd_r[30]), .B(vdd_), .G(vdd_cntl_r[30]),
     .S(vdd_));
P_11_LPHVT  M0_29_ ( .D(r_gnd_r[29]), .B(vdd_), .G(vdd_cntl_r[29]),
     .S(vdd_));
P_11_LPHVT  M0_28_ ( .D(r_gnd_r[28]), .B(vdd_), .G(vdd_cntl_r[28]),
     .S(vdd_));
P_11_LPHVT  M0_27_ ( .D(r_gnd_r[27]), .B(vdd_), .G(vdd_cntl_r[27]),
     .S(vdd_));
P_11_LPHVT  M0_26_ ( .D(r_gnd_r[26]), .B(vdd_), .G(vdd_cntl_r[26]),
     .S(vdd_));
P_11_LPHVT  M0_25_ ( .D(r_gnd_r[25]), .B(vdd_), .G(vdd_cntl_r[25]),
     .S(vdd_));
P_11_LPHVT  M0_24_ ( .D(r_gnd_r[24]), .B(vdd_), .G(vdd_cntl_r[24]),
     .S(vdd_));
P_11_LPHVT  M0_23_ ( .D(r_gnd_r[23]), .B(vdd_), .G(vdd_cntl_r[23]),
     .S(vdd_));
P_11_LPHVT  M0_22_ ( .D(r_gnd_r[22]), .B(vdd_), .G(vdd_cntl_r[22]),
     .S(vdd_));
P_11_LPHVT  M0_21_ ( .D(r_gnd_r[21]), .B(vdd_), .G(vdd_cntl_r[21]),
     .S(vdd_));
P_11_LPHVT  M0_20_ ( .D(r_gnd_r[20]), .B(vdd_), .G(vdd_cntl_r[20]),
     .S(vdd_));
P_11_LPHVT  M0_19_ ( .D(r_gnd_r[19]), .B(vdd_), .G(vdd_cntl_r[19]),
     .S(vdd_));
P_11_LPHVT  M0_18_ ( .D(r_gnd_r[18]), .B(vdd_), .G(vdd_cntl_r[18]),
     .S(vdd_));
P_11_LPHVT  M0_17_ ( .D(r_gnd_r[17]), .B(vdd_), .G(vdd_cntl_r[17]),
     .S(vdd_));
P_11_LPHVT  M0_16_ ( .D(r_gnd_r[16]), .B(vdd_), .G(vdd_cntl_r[16]),
     .S(vdd_));
P_11_LPHVT  M0_15_ ( .D(r_gnd_r[15]), .B(vdd_), .G(vdd_cntl_r[15]),
     .S(vdd_));
P_11_LPHVT  M0_14_ ( .D(r_gnd_r[14]), .B(vdd_), .G(vdd_cntl_r[14]),
     .S(vdd_));
P_11_LPHVT  M0_13_ ( .D(r_gnd_r[13]), .B(vdd_), .G(vdd_cntl_r[13]),
     .S(vdd_));
P_11_LPHVT  M0_12_ ( .D(r_gnd_r[12]), .B(vdd_), .G(vdd_cntl_r[12]),
     .S(vdd_));
P_11_LPHVT  M0_11_ ( .D(r_gnd_r[11]), .B(vdd_), .G(vdd_cntl_r[11]),
     .S(vdd_));
P_11_LPHVT  M0_10_ ( .D(r_gnd_r[10]), .B(vdd_), .G(vdd_cntl_r[10]),
     .S(vdd_));
P_11_LPHVT  M0_9_ ( .D(r_gnd_r[9]), .B(vdd_), .G(vdd_cntl_r[9]),
     .S(vdd_));
P_11_LPHVT  M0_8_ ( .D(r_gnd_r[8]), .B(vdd_), .G(vdd_cntl_r[8]),
     .S(vdd_));
P_11_LPHVT  M0_7_ ( .D(r_gnd_r[7]), .B(vdd_), .G(vdd_cntl_r[7]),
     .S(vdd_));
P_11_LPHVT  M0_6_ ( .D(r_gnd_r[6]), .B(vdd_), .G(vdd_cntl_r[6]),
     .S(vdd_));
P_11_LPHVT  M0_5_ ( .D(r_gnd_r[5]), .B(vdd_), .G(vdd_cntl_r[5]),
     .S(vdd_));
P_11_LPHVT  M0_4_ ( .D(r_gnd_r[4]), .B(vdd_), .G(vdd_cntl_r[4]),
     .S(vdd_));
P_11_LPHVT  M0_3_ ( .D(r_gnd_r[3]), .B(vdd_), .G(vdd_cntl_r[3]),
     .S(vdd_));
P_11_LPHVT  M0_2_ ( .D(r_gnd_r[2]), .B(vdd_), .G(vdd_cntl_r[2]),
     .S(vdd_));
P_11_LPHVT  M0_1_ ( .D(r_gnd_r[1]), .B(vdd_), .G(vdd_cntl_r[1]),
     .S(vdd_));
P_11_LPHVT  M0_0_ ( .D(r_gnd_r[0]), .B(vdd_), .G(vdd_cntl_r[0]),
     .S(vdd_));
P_11_LPHVT  M3_77_ ( .D(r_gnd_l[77]), .B(vdd_), .G(vdd_cntl_l[77]),
     .S(vdd_));
P_11_LPHVT  M3_76_ ( .D(r_gnd_l[76]), .B(vdd_), .G(vdd_cntl_l[76]),
     .S(vdd_));
P_11_LPHVT  M3_75_ ( .D(r_gnd_l[75]), .B(vdd_), .G(vdd_cntl_l[75]),
     .S(vdd_));
P_11_LPHVT  M3_74_ ( .D(r_gnd_l[74]), .B(vdd_), .G(vdd_cntl_l[74]),
     .S(vdd_));
P_11_LPHVT  M3_73_ ( .D(r_gnd_l[73]), .B(vdd_), .G(vdd_cntl_l[73]),
     .S(vdd_));
P_11_LPHVT  M3_72_ ( .D(r_gnd_l[72]), .B(vdd_), .G(vdd_cntl_l[72]),
     .S(vdd_));
P_11_LPHVT  M3_71_ ( .D(r_gnd_l[71]), .B(vdd_), .G(vdd_cntl_l[71]),
     .S(vdd_));
P_11_LPHVT  M3_70_ ( .D(r_gnd_l[70]), .B(vdd_), .G(vdd_cntl_l[70]),
     .S(vdd_));
P_11_LPHVT  M3_69_ ( .D(r_gnd_l[69]), .B(vdd_), .G(vdd_cntl_l[69]),
     .S(vdd_));
P_11_LPHVT  M3_68_ ( .D(r_gnd_l[68]), .B(vdd_), .G(vdd_cntl_l[68]),
     .S(vdd_));
P_11_LPHVT  M3_67_ ( .D(r_gnd_l[67]), .B(vdd_), .G(vdd_cntl_l[67]),
     .S(vdd_));
P_11_LPHVT  M3_66_ ( .D(r_gnd_l[66]), .B(vdd_), .G(vdd_cntl_l[66]),
     .S(vdd_));
P_11_LPHVT  M3_65_ ( .D(r_gnd_l[65]), .B(vdd_), .G(vdd_cntl_l[65]),
     .S(vdd_));
P_11_LPHVT  M3_64_ ( .D(r_gnd_l[64]), .B(vdd_), .G(vdd_cntl_l[64]),
     .S(vdd_));
P_11_LPHVT  M3_63_ ( .D(r_gnd_l[63]), .B(vdd_), .G(vdd_cntl_l[63]),
     .S(vdd_));
P_11_LPHVT  M3_62_ ( .D(r_gnd_l[62]), .B(vdd_), .G(vdd_cntl_l[62]),
     .S(vdd_));
P_11_LPHVT  M3_61_ ( .D(r_gnd_l[61]), .B(vdd_), .G(vdd_cntl_l[61]),
     .S(vdd_));
P_11_LPHVT  M3_60_ ( .D(r_gnd_l[60]), .B(vdd_), .G(vdd_cntl_l[60]),
     .S(vdd_));
P_11_LPHVT  M3_59_ ( .D(r_gnd_l[59]), .B(vdd_), .G(vdd_cntl_l[59]),
     .S(vdd_));
P_11_LPHVT  M3_58_ ( .D(r_gnd_l[58]), .B(vdd_), .G(vdd_cntl_l[58]),
     .S(vdd_));
P_11_LPHVT  M3_57_ ( .D(r_gnd_l[57]), .B(vdd_), .G(vdd_cntl_l[57]),
     .S(vdd_));
P_11_LPHVT  M3_56_ ( .D(r_gnd_l[56]), .B(vdd_), .G(vdd_cntl_l[56]),
     .S(vdd_));
P_11_LPHVT  M3_55_ ( .D(r_gnd_l[55]), .B(vdd_), .G(vdd_cntl_l[55]),
     .S(vdd_));
P_11_LPHVT  M3_54_ ( .D(r_gnd_l[54]), .B(vdd_), .G(vdd_cntl_l[54]),
     .S(vdd_));
P_11_LPHVT  M3_53_ ( .D(r_gnd_l[53]), .B(vdd_), .G(vdd_cntl_l[53]),
     .S(vdd_));
P_11_LPHVT  M3_52_ ( .D(r_gnd_l[52]), .B(vdd_), .G(vdd_cntl_l[52]),
     .S(vdd_));
P_11_LPHVT  M3_51_ ( .D(r_gnd_l[51]), .B(vdd_), .G(vdd_cntl_l[51]),
     .S(vdd_));
P_11_LPHVT  M3_50_ ( .D(r_gnd_l[50]), .B(vdd_), .G(vdd_cntl_l[50]),
     .S(vdd_));
P_11_LPHVT  M3_49_ ( .D(r_gnd_l[49]), .B(vdd_), .G(vdd_cntl_l[49]),
     .S(vdd_));
P_11_LPHVT  M3_48_ ( .D(r_gnd_l[48]), .B(vdd_), .G(vdd_cntl_l[48]),
     .S(vdd_));
P_11_LPHVT  M3_47_ ( .D(r_gnd_l[47]), .B(vdd_), .G(vdd_cntl_l[47]),
     .S(vdd_));
P_11_LPHVT  M3_46_ ( .D(r_gnd_l[46]), .B(vdd_), .G(vdd_cntl_l[46]),
     .S(vdd_));
P_11_LPHVT  M3_45_ ( .D(r_gnd_l[45]), .B(vdd_), .G(vdd_cntl_l[45]),
     .S(vdd_));
P_11_LPHVT  M3_44_ ( .D(r_gnd_l[44]), .B(vdd_), .G(vdd_cntl_l[44]),
     .S(vdd_));
P_11_LPHVT  M3_43_ ( .D(r_gnd_l[43]), .B(vdd_), .G(vdd_cntl_l[43]),
     .S(vdd_));
P_11_LPHVT  M3_42_ ( .D(r_gnd_l[42]), .B(vdd_), .G(vdd_cntl_l[42]),
     .S(vdd_));
P_11_LPHVT  M3_41_ ( .D(r_gnd_l[41]), .B(vdd_), .G(vdd_cntl_l[41]),
     .S(vdd_));
P_11_LPHVT  M3_40_ ( .D(r_gnd_l[40]), .B(vdd_), .G(vdd_cntl_l[40]),
     .S(vdd_));
P_11_LPHVT  M3_39_ ( .D(r_gnd_l[39]), .B(vdd_), .G(vdd_cntl_l[39]),
     .S(vdd_));
P_11_LPHVT  M3_38_ ( .D(r_gnd_l[38]), .B(vdd_), .G(vdd_cntl_l[38]),
     .S(vdd_));
P_11_LPHVT  M3_37_ ( .D(r_gnd_l[37]), .B(vdd_), .G(vdd_cntl_l[37]),
     .S(vdd_));
P_11_LPHVT  M3_36_ ( .D(r_gnd_l[36]), .B(vdd_), .G(vdd_cntl_l[36]),
     .S(vdd_));
P_11_LPHVT  M3_35_ ( .D(r_gnd_l[35]), .B(vdd_), .G(vdd_cntl_l[35]),
     .S(vdd_));
P_11_LPHVT  M3_34_ ( .D(r_gnd_l[34]), .B(vdd_), .G(vdd_cntl_l[34]),
     .S(vdd_));
P_11_LPHVT  M3_33_ ( .D(r_gnd_l[33]), .B(vdd_), .G(vdd_cntl_l[33]),
     .S(vdd_));
P_11_LPHVT  M3_32_ ( .D(r_gnd_l[32]), .B(vdd_), .G(vdd_cntl_l[32]),
     .S(vdd_));
P_11_LPHVT  M3_31_ ( .D(r_gnd_l[31]), .B(vdd_), .G(vdd_cntl_l[31]),
     .S(vdd_));
P_11_LPHVT  M3_30_ ( .D(r_gnd_l[30]), .B(vdd_), .G(vdd_cntl_l[30]),
     .S(vdd_));
P_11_LPHVT  M3_29_ ( .D(r_gnd_l[29]), .B(vdd_), .G(vdd_cntl_l[29]),
     .S(vdd_));
P_11_LPHVT  M3_28_ ( .D(r_gnd_l[28]), .B(vdd_), .G(vdd_cntl_l[28]),
     .S(vdd_));
P_11_LPHVT  M3_27_ ( .D(r_gnd_l[27]), .B(vdd_), .G(vdd_cntl_l[27]),
     .S(vdd_));
P_11_LPHVT  M3_26_ ( .D(r_gnd_l[26]), .B(vdd_), .G(vdd_cntl_l[26]),
     .S(vdd_));
P_11_LPHVT  M3_25_ ( .D(r_gnd_l[25]), .B(vdd_), .G(vdd_cntl_l[25]),
     .S(vdd_));
P_11_LPHVT  M3_24_ ( .D(r_gnd_l[24]), .B(vdd_), .G(vdd_cntl_l[24]),
     .S(vdd_));
P_11_LPHVT  M3_23_ ( .D(r_gnd_l[23]), .B(vdd_), .G(vdd_cntl_l[23]),
     .S(vdd_));
P_11_LPHVT  M3_22_ ( .D(r_gnd_l[22]), .B(vdd_), .G(vdd_cntl_l[22]),
     .S(vdd_));
P_11_LPHVT  M3_21_ ( .D(r_gnd_l[21]), .B(vdd_), .G(vdd_cntl_l[21]),
     .S(vdd_));
P_11_LPHVT  M3_20_ ( .D(r_gnd_l[20]), .B(vdd_), .G(vdd_cntl_l[20]),
     .S(vdd_));
P_11_LPHVT  M3_19_ ( .D(r_gnd_l[19]), .B(vdd_), .G(vdd_cntl_l[19]),
     .S(vdd_));
P_11_LPHVT  M3_18_ ( .D(r_gnd_l[18]), .B(vdd_), .G(vdd_cntl_l[18]),
     .S(vdd_));
P_11_LPHVT  M3_17_ ( .D(r_gnd_l[17]), .B(vdd_), .G(vdd_cntl_l[17]),
     .S(vdd_));
P_11_LPHVT  M3_16_ ( .D(r_gnd_l[16]), .B(vdd_), .G(vdd_cntl_l[16]),
     .S(vdd_));
P_11_LPHVT  M3_15_ ( .D(r_gnd_l[15]), .B(vdd_), .G(vdd_cntl_l[15]),
     .S(vdd_));
P_11_LPHVT  M3_14_ ( .D(r_gnd_l[14]), .B(vdd_), .G(vdd_cntl_l[14]),
     .S(vdd_));
P_11_LPHVT  M3_13_ ( .D(r_gnd_l[13]), .B(vdd_), .G(vdd_cntl_l[13]),
     .S(vdd_));
P_11_LPHVT  M3_12_ ( .D(r_gnd_l[12]), .B(vdd_), .G(vdd_cntl_l[12]),
     .S(vdd_));
P_11_LPHVT  M3_11_ ( .D(r_gnd_l[11]), .B(vdd_), .G(vdd_cntl_l[11]),
     .S(vdd_));
P_11_LPHVT  M3_10_ ( .D(r_gnd_l[10]), .B(vdd_), .G(vdd_cntl_l[10]),
     .S(vdd_));
P_11_LPHVT  M3_9_ ( .D(r_gnd_l[9]), .B(vdd_), .G(vdd_cntl_l[9]),
     .S(vdd_));
P_11_LPHVT  M3_8_ ( .D(r_gnd_l[8]), .B(vdd_), .G(vdd_cntl_l[8]),
     .S(vdd_));
P_11_LPHVT  M3_7_ ( .D(r_gnd_l[7]), .B(vdd_), .G(vdd_cntl_l[7]),
     .S(vdd_));
P_11_LPHVT  M3_6_ ( .D(r_gnd_l[6]), .B(vdd_), .G(vdd_cntl_l[6]),
     .S(vdd_));
P_11_LPHVT  M3_5_ ( .D(r_gnd_l[5]), .B(vdd_), .G(vdd_cntl_l[5]),
     .S(vdd_));
P_11_LPHVT  M3_4_ ( .D(r_gnd_l[4]), .B(vdd_), .G(vdd_cntl_l[4]),
     .S(vdd_));
P_11_LPHVT  M3_3_ ( .D(r_gnd_l[3]), .B(vdd_), .G(vdd_cntl_l[3]),
     .S(vdd_));
P_11_LPHVT  M3_2_ ( .D(r_gnd_l[2]), .B(vdd_), .G(vdd_cntl_l[2]),
     .S(vdd_));
P_11_LPHVT  M3_1_ ( .D(r_gnd_l[1]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
P_11_LPHVT  M3_0_ ( .D(r_gnd_l[0]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));
cram_2x2x2_ice8p I_mem2x2x2t_38_ ( .wl_r(wl_r[77:76]),
     .wl_l(wl_l[77:76]), .reset_r(reset_r[77:76]),
     .reset_l(reset_l[77:76]), .pgate_r(pgate_r[77:76]),
     .pgate_l(pgate_l[77:76]), .q_b({net39[0], net39[1], net39[2],
     net39[3], net39[4], net39[5], net39[6], net39[7]}), .q({net40[0],
     net40[1], net40[2], net40[3], net40[4], net40[5], net40[6],
     net40[7]}), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[77:76]),
     .r_gnd_r(r_gnd_r[77:76]));
cram_2x2x2_ice8p I_mem2x2x2t_37_ ( .wl_r(wl_r[75:74]),
     .wl_l(wl_l[75:74]), .reset_r(reset_r[75:74]),
     .reset_l(reset_l[75:74]), .pgate_r(pgate_r[75:74]),
     .pgate_l(pgate_l[75:74]), .q_b({net39[8], net39[9], net39[10],
     net39[11], net39[12], net39[13], net39[14], net39[15]}),
     .q({net40[8], net40[9], net40[10], net40[11], net40[12],
     net40[13], net40[14], net40[15]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[75:74]), .r_gnd_r(r_gnd_r[75:74]));
cram_2x2x2_ice8p I_mem2x2x2t_36_ ( .wl_r(wl_r[73:72]),
     .wl_l(wl_l[73:72]), .reset_r(reset_r[73:72]),
     .reset_l(reset_l[73:72]), .pgate_r(pgate_r[73:72]),
     .pgate_l(pgate_l[73:72]), .q_b({net39[16], net39[17], net39[18],
     net39[19], net39[20], net39[21], net39[22], net39[23]}),
     .q({net40[16], net40[17], net40[18], net40[19], net40[20],
     net40[21], net40[22], net40[23]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[73:72]), .r_gnd_r(r_gnd_r[73:72]));
cram_2x2x2_ice8p I_mem2x2x2t_35_ ( .wl_r(wl_r[71:70]),
     .wl_l(wl_l[71:70]), .reset_r(reset_r[71:70]),
     .reset_l(reset_l[71:70]), .pgate_r(pgate_r[71:70]),
     .pgate_l(pgate_l[71:70]), .q_b({net39[24], net39[25], net39[26],
     net39[27], net39[28], net39[29], net39[30], net39[31]}),
     .q({net40[24], net40[25], net40[26], net40[27], net40[28],
     net40[29], net40[30], net40[31]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[71:70]), .r_gnd_r(r_gnd_r[71:70]));
cram_2x2x2_ice8p I_mem2x2x2t_34_ ( .wl_r(wl_r[69:68]),
     .wl_l(wl_l[69:68]), .reset_r(reset_r[69:68]),
     .reset_l(reset_l[69:68]), .pgate_r(pgate_r[69:68]),
     .pgate_l(pgate_l[69:68]), .q_b({net39[32], net39[33], net39[34],
     net39[35], net39[36], net39[37], net39[38], net39[39]}),
     .q({net40[32], net40[33], net40[34], net40[35], net40[36],
     net40[37], net40[38], net40[39]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[69:68]), .r_gnd_r(r_gnd_r[69:68]));
cram_2x2x2_ice8p I_mem2x2x2t_33_ ( .wl_r(wl_r[67:66]),
     .wl_l(wl_l[67:66]), .reset_r(reset_r[67:66]),
     .reset_l(reset_l[67:66]), .pgate_r(pgate_r[67:66]),
     .pgate_l(pgate_l[67:66]), .q_b({net39[40], net39[41], net39[42],
     net39[43], net39[44], net39[45], net39[46], net39[47]}),
     .q({net40[40], net40[41], net40[42], net40[43], net40[44],
     net40[45], net40[46], net40[47]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[67:66]), .r_gnd_r(r_gnd_r[67:66]));
cram_2x2x2_ice8p I_mem2x2x2t_32_ ( .wl_r(wl_r[65:64]),
     .wl_l(wl_l[65:64]), .reset_r(reset_r[65:64]),
     .reset_l(reset_l[65:64]), .pgate_r(pgate_r[65:64]),
     .pgate_l(pgate_l[65:64]), .q_b({net39[48], net39[49], net39[50],
     net39[51], net39[52], net39[53], net39[54], net39[55]}),
     .q({net40[48], net40[49], net40[50], net40[51], net40[52],
     net40[53], net40[54], net40[55]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[65:64]), .r_gnd_r(r_gnd_r[65:64]));
cram_2x2x2_ice8p I_mem2x2x2t_31_ ( .wl_r(wl_r[63:62]),
     .wl_l(wl_l[63:62]), .reset_r(reset_r[63:62]),
     .reset_l(reset_l[63:62]), .pgate_r(pgate_r[63:62]),
     .pgate_l(pgate_l[63:62]), .q_b({net39[56], net39[57], net39[58],
     net39[59], net39[60], net39[61], net39[62], net39[63]}),
     .q({net40[56], net40[57], net40[58], net40[59], net40[60],
     net40[61], net40[62], net40[63]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[63:62]), .r_gnd_r(r_gnd_r[63:62]));
cram_2x2x2_ice8p I_mem2x2x2t_30_ ( .wl_r(wl_r[61:60]),
     .wl_l(wl_l[61:60]), .reset_r(reset_r[61:60]),
     .reset_l(reset_l[61:60]), .pgate_r(pgate_r[61:60]),
     .pgate_l(pgate_l[61:60]), .q_b({net39[64], net39[65], net39[66],
     net39[67], net39[68], net39[69], net39[70], net39[71]}),
     .q({net40[64], net40[65], net40[66], net40[67], net40[68],
     net40[69], net40[70], net40[71]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[61:60]), .r_gnd_r(r_gnd_r[61:60]));
cram_2x2x2_ice8p I_mem2x2x2t_29_ ( .wl_r(wl_r[59:58]),
     .wl_l(wl_l[59:58]), .reset_r(reset_r[59:58]),
     .reset_l(reset_l[59:58]), .pgate_r(pgate_r[59:58]),
     .pgate_l(pgate_l[59:58]), .q_b({net39[72], net39[73], net39[74],
     net39[75], net39[76], net39[77], net39[78], net39[79]}),
     .q({net40[72], net40[73], net40[74], net40[75], net40[76],
     net40[77], net40[78], net40[79]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[59:58]), .r_gnd_r(r_gnd_r[59:58]));
cram_2x2x2_ice8p I_mem2x2x2t_28_ ( .wl_r(wl_r[57:56]),
     .wl_l(wl_l[57:56]), .reset_r(reset_r[57:56]),
     .reset_l(reset_l[57:56]), .pgate_r(pgate_r[57:56]),
     .pgate_l(pgate_l[57:56]), .q_b({net39[80], net39[81], net39[82],
     net39[83], net39[84], net39[85], net39[86], net39[87]}),
     .q({net40[80], net40[81], net40[82], net40[83], net40[84],
     net40[85], net40[86], net40[87]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[57:56]), .r_gnd_r(r_gnd_r[57:56]));
cram_2x2x2_ice8p I_mem2x2x2t_27_ ( .wl_r(wl_r[55:54]),
     .wl_l(wl_l[55:54]), .reset_r(reset_r[55:54]),
     .reset_l(reset_l[55:54]), .pgate_r(pgate_r[55:54]),
     .pgate_l(pgate_l[55:54]), .q_b({net39[88], net39[89], net39[90],
     net39[91], net39[92], net39[93], net39[94], net39[95]}),
     .q({net40[88], net40[89], net40[90], net40[91], net40[92],
     net40[93], net40[94], net40[95]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[55:54]), .r_gnd_r(r_gnd_r[55:54]));
cram_2x2x2_ice8p I_mem2x2x2t_26_ ( .wl_r(wl_r[53:52]),
     .wl_l(wl_l[53:52]), .reset_r(reset_r[53:52]),
     .reset_l(reset_l[53:52]), .pgate_r(pgate_r[53:52]),
     .pgate_l(pgate_l[53:52]), .q_b({net39[96], net39[97], net39[98],
     net39[99], net39[100], net39[101], net39[102], net39[103]}),
     .q({net40[96], net40[97], net40[98], net40[99], net40[100],
     net40[101], net40[102], net40[103]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[53:52]), .r_gnd_r(r_gnd_r[53:52]));
cram_2x2x2_ice8p I_mem2x2x2t_25_ ( .wl_r(wl_r[51:50]),
     .wl_l(wl_l[51:50]), .reset_r(reset_r[51:50]),
     .reset_l(reset_l[51:50]), .pgate_r(pgate_r[51:50]),
     .pgate_l(pgate_l[51:50]), .q_b({net39[104], net39[105],
     net39[106], net39[107], net39[108], net39[109], net39[110],
     net39[111]}), .q({net40[104], net40[105], net40[106], net40[107],
     net40[108], net40[109], net40[110], net40[111]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[51:50]), .r_gnd_r(r_gnd_r[51:50]));
cram_2x2x2_ice8p I_mem2x2x2t_24_ ( .wl_r(wl_r[49:48]),
     .wl_l(wl_l[49:48]), .reset_r(reset_r[49:48]),
     .reset_l(reset_l[49:48]), .pgate_r(pgate_r[49:48]),
     .pgate_l(pgate_l[49:48]), .q_b({net39[112], net39[113],
     net39[114], net39[115], net39[116], net39[117], net39[118],
     net39[119]}), .q({net40[112], net40[113], net40[114], net40[115],
     net40[116], net40[117], net40[118], net40[119]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[49:48]), .r_gnd_r(r_gnd_r[49:48]));
cram_2x2x2_ice8p I_mem2x2x2t_23_ ( .wl_r(wl_r[47:46]),
     .wl_l(wl_l[47:46]), .reset_r(reset_r[47:46]),
     .reset_l(reset_l[47:46]), .pgate_r(pgate_r[47:46]),
     .pgate_l(pgate_l[47:46]), .q_b({net39[120], net39[121],
     net39[122], net39[123], net39[124], net39[125], net39[126],
     net39[127]}), .q({net40[120], net40[121], net40[122], net40[123],
     net40[124], net40[125], net40[126], net40[127]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[47:46]), .r_gnd_r(r_gnd_r[47:46]));
cram_2x2x2_ice8p I_mem2x2x2t_22_ ( .wl_r(wl_r[45:44]),
     .wl_l(wl_l[45:44]), .reset_r(reset_r[45:44]),
     .reset_l(reset_l[45:44]), .pgate_r(pgate_r[45:44]),
     .pgate_l(pgate_l[45:44]), .q_b({net39[128], net39[129],
     net39[130], net39[131], net39[132], net39[133], net39[134],
     net39[135]}), .q({net40[128], net40[129], net40[130], net40[131],
     net40[132], net40[133], net40[134], net40[135]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[45:44]), .r_gnd_r(r_gnd_r[45:44]));
cram_2x2x2_ice8p I_mem2x2x2t_21_ ( .wl_r(wl_r[43:42]),
     .wl_l(wl_l[43:42]), .reset_r(reset_r[43:42]),
     .reset_l(reset_l[43:42]), .pgate_r(pgate_r[43:42]),
     .pgate_l(pgate_l[43:42]), .q_b({net39[136], net39[137],
     net39[138], net39[139], net39[140], net39[141], net39[142],
     net39[143]}), .q({net40[136], net40[137], net40[138], net40[139],
     net40[140], net40[141], net40[142], net40[143]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[43:42]), .r_gnd_r(r_gnd_r[43:42]));
cram_2x2x2_ice8p I_mem2x2x2t_20_ ( .wl_r(wl_r[41:40]),
     .wl_l(wl_l[41:40]), .reset_r(reset_r[41:40]),
     .reset_l(reset_l[41:40]), .pgate_r(pgate_r[41:40]),
     .pgate_l(pgate_l[41:40]), .q_b({net39[144], net39[145],
     net39[146], net39[147], net39[148], net39[149], net39[150],
     net39[151]}), .q({net40[144], net40[145], net40[146], net40[147],
     net40[148], net40[149], net40[150], net40[151]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[41:40]), .r_gnd_r(r_gnd_r[41:40]));
cram_2x2x2_ice8p I_mem2x2x2t_19_ ( .wl_r(wl_r[39:38]),
     .wl_l(wl_l[39:38]), .reset_r(reset_r[39:38]),
     .reset_l(reset_l[39:38]), .pgate_r(pgate_r[39:38]),
     .pgate_l(pgate_l[39:38]), .q_b({net39[152], net39[153],
     net39[154], net39[155], net39[156], net39[157], net39[158],
     net39[159]}), .q({net40[152], net40[153], net40[154], net40[155],
     net40[156], net40[157], net40[158], net40[159]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[39:38]), .r_gnd_r(r_gnd_r[39:38]));
cram_2x2x2_ice8p I_mem2x2x2t_18_ ( .wl_r(wl_r[37:36]),
     .wl_l(wl_l[37:36]), .reset_r(reset_r[37:36]),
     .reset_l(reset_l[37:36]), .pgate_r(pgate_r[37:36]),
     .pgate_l(pgate_l[37:36]), .q_b({net39[160], net39[161],
     net39[162], net39[163], net39[164], net39[165], net39[166],
     net39[167]}), .q({net40[160], net40[161], net40[162], net40[163],
     net40[164], net40[165], net40[166], net40[167]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[37:36]), .r_gnd_r(r_gnd_r[37:36]));
cram_2x2x2_ice8p I_mem2x2x2t_17_ ( .wl_r(wl_r[35:34]),
     .wl_l(wl_l[35:34]), .reset_r(reset_r[35:34]),
     .reset_l(reset_l[35:34]), .pgate_r(pgate_r[35:34]),
     .pgate_l(pgate_l[35:34]), .q_b({net39[168], net39[169],
     net39[170], net39[171], net39[172], net39[173], net39[174],
     net39[175]}), .q({net40[168], net40[169], net40[170], net40[171],
     net40[172], net40[173], net40[174], net40[175]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[35:34]), .r_gnd_r(r_gnd_r[35:34]));
cram_2x2x2_ice8p I_mem2x2x2t_16_ ( .wl_r(wl_r[33:32]),
     .wl_l(wl_l[33:32]), .reset_r(reset_r[33:32]),
     .reset_l(reset_l[33:32]), .pgate_r(pgate_r[33:32]),
     .pgate_l(pgate_l[33:32]), .q_b({net39[176], net39[177],
     net39[178], net39[179], net39[180], net39[181], net39[182],
     net39[183]}), .q({net40[176], net40[177], net40[178], net40[179],
     net40[180], net40[181], net40[182], net40[183]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[33:32]), .r_gnd_r(r_gnd_r[33:32]));
cram_2x2x2_ice8p I_mem2x2x2t_15_ ( .wl_r(wl_r[31:30]),
     .wl_l(wl_l[31:30]), .reset_r(reset_r[31:30]),
     .reset_l(reset_l[31:30]), .pgate_r(pgate_r[31:30]),
     .pgate_l(pgate_l[31:30]), .q_b({net39[184], net39[185],
     net39[186], net39[187], net39[188], net39[189], net39[190],
     net39[191]}), .q({net40[184], net40[185], net40[186], net40[187],
     net40[188], net40[189], net40[190], net40[191]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[31:30]), .r_gnd_r(r_gnd_r[31:30]));
cram_2x2x2_ice8p I_mem2x2x2t_14_ ( .wl_r(wl_r[29:28]),
     .wl_l(wl_l[29:28]), .reset_r(reset_r[29:28]),
     .reset_l(reset_l[29:28]), .pgate_r(pgate_r[29:28]),
     .pgate_l(pgate_l[29:28]), .q_b({net39[192], net39[193],
     net39[194], net39[195], net39[196], net39[197], net39[198],
     net39[199]}), .q({net40[192], net40[193], net40[194], net40[195],
     net40[196], net40[197], net40[198], net40[199]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[29:28]), .r_gnd_r(r_gnd_r[29:28]));
cram_2x2x2_ice8p I_mem2x2x2t_13_ ( .wl_r(wl_r[27:26]),
     .wl_l(wl_l[27:26]), .reset_r(reset_r[27:26]),
     .reset_l(reset_l[27:26]), .pgate_r(pgate_r[27:26]),
     .pgate_l(pgate_l[27:26]), .q_b({net39[200], net39[201],
     net39[202], net39[203], net39[204], net39[205], net39[206],
     net39[207]}), .q({net40[200], net40[201], net40[202], net40[203],
     net40[204], net40[205], net40[206], net40[207]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[27:26]), .r_gnd_r(r_gnd_r[27:26]));
cram_2x2x2_ice8p I_mem2x2x2t_12_ ( .wl_r(wl_r[25:24]),
     .wl_l(wl_l[25:24]), .reset_r(reset_r[25:24]),
     .reset_l(reset_l[25:24]), .pgate_r(pgate_r[25:24]),
     .pgate_l(pgate_l[25:24]), .q_b({net39[208], net39[209],
     net39[210], net39[211], net39[212], net39[213], net39[214],
     net39[215]}), .q({net40[208], net40[209], net40[210], net40[211],
     net40[212], net40[213], net40[214], net40[215]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[25:24]), .r_gnd_r(r_gnd_r[25:24]));
cram_2x2x2_ice8p I_mem2x2x2t_11_ ( .wl_r(wl_r[23:22]),
     .wl_l(wl_l[23:22]), .reset_r(reset_r[23:22]),
     .reset_l(reset_l[23:22]), .pgate_r(pgate_r[23:22]),
     .pgate_l(pgate_l[23:22]), .q_b({net39[216], net39[217],
     net39[218], net39[219], net39[220], net39[221], net39[222],
     net39[223]}), .q({net40[216], net40[217], net40[218], net40[219],
     net40[220], net40[221], net40[222], net40[223]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[23:22]), .r_gnd_r(r_gnd_r[23:22]));
cram_2x2x2_ice8p I_mem2x2x2t_10_ ( .wl_r(wl_r[21:20]),
     .wl_l(wl_l[21:20]), .reset_r(reset_r[21:20]),
     .reset_l(reset_l[21:20]), .pgate_r(pgate_r[21:20]),
     .pgate_l(pgate_l[21:20]), .q_b({net39[224], net39[225],
     net39[226], net39[227], net39[228], net39[229], net39[230],
     net39[231]}), .q({net40[224], net40[225], net40[226], net40[227],
     net40[228], net40[229], net40[230], net40[231]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[21:20]), .r_gnd_r(r_gnd_r[21:20]));
cram_2x2x2_ice8p I_mem2x2x2t_9_ ( .wl_r(wl_r[19:18]),
     .wl_l(wl_l[19:18]), .reset_r(reset_r[19:18]),
     .reset_l(reset_l[19:18]), .pgate_r(pgate_r[19:18]),
     .pgate_l(pgate_l[19:18]), .q_b({net39[232], net39[233],
     net39[234], net39[235], net39[236], net39[237], net39[238],
     net39[239]}), .q({net40[232], net40[233], net40[234], net40[235],
     net40[236], net40[237], net40[238], net40[239]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[19:18]), .r_gnd_r(r_gnd_r[19:18]));
cram_2x2x2_ice8p I_mem2x2x2t_8_ ( .wl_r(wl_r[17:16]),
     .wl_l(wl_l[17:16]), .reset_r(reset_r[17:16]),
     .reset_l(reset_l[17:16]), .pgate_r(pgate_r[17:16]),
     .pgate_l(pgate_l[17:16]), .q_b({net39[240], net39[241],
     net39[242], net39[243], net39[244], net39[245], net39[246],
     net39[247]}), .q({net40[240], net40[241], net40[242], net40[243],
     net40[244], net40[245], net40[246], net40[247]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[17:16]), .r_gnd_r(r_gnd_r[17:16]));
cram_2x2x2_ice8p I_mem2x2x2t_7_ ( .wl_r(wl_r[15:14]),
     .wl_l(wl_l[15:14]), .reset_r(reset_r[15:14]),
     .reset_l(reset_l[15:14]), .pgate_r(pgate_r[15:14]),
     .pgate_l(pgate_l[15:14]), .q_b({net39[248], net39[249],
     net39[250], net39[251], net39[252], net39[253], net39[254],
     net39[255]}), .q({net40[248], net40[249], net40[250], net40[251],
     net40[252], net40[253], net40[254], net40[255]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[15:14]), .r_gnd_r(r_gnd_r[15:14]));
cram_2x2x2_ice8p I_mem2x2x2t_6_ ( .wl_r(wl_r[13:12]),
     .wl_l(wl_l[13:12]), .reset_r(reset_r[13:12]),
     .reset_l(reset_l[13:12]), .pgate_r(pgate_r[13:12]),
     .pgate_l(pgate_l[13:12]), .q_b({net39[256], net39[257],
     net39[258], net39[259], net39[260], net39[261], net39[262],
     net39[263]}), .q({net40[256], net40[257], net40[258], net40[259],
     net40[260], net40[261], net40[262], net40[263]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[13:12]), .r_gnd_r(r_gnd_r[13:12]));
cram_2x2x2_ice8p I_mem2x2x2t_5_ ( .wl_r(wl_r[11:10]),
     .wl_l(wl_l[11:10]), .reset_r(reset_r[11:10]),
     .reset_l(reset_l[11:10]), .pgate_r(pgate_r[11:10]),
     .pgate_l(pgate_l[11:10]), .q_b({net39[264], net39[265],
     net39[266], net39[267], net39[268], net39[269], net39[270],
     net39[271]}), .q({net40[264], net40[265], net40[266], net40[267],
     net40[268], net40[269], net40[270], net40[271]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[11:10]), .r_gnd_r(r_gnd_r[11:10]));
cram_2x2x2_ice8p I_mem2x2x2t_4_ ( .wl_r(wl_r[9:8]), .wl_l(wl_l[9:8]),
     .reset_r(reset_r[9:8]), .reset_l(reset_l[9:8]),
     .pgate_r(pgate_r[9:8]), .pgate_l(pgate_l[9:8]), .q_b({net39[272],
     net39[273], net39[274], net39[275], net39[276], net39[277],
     net39[278], net39[279]}), .q({net40[272], net40[273], net40[274],
     net40[275], net40[276], net40[277], net40[278], net40[279]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[9:8]), .r_gnd_r(r_gnd_r[9:8]));
cram_2x2x2_ice8p I_mem2x2x2t_3_ ( .wl_r(wl_r[7:6]), .wl_l(wl_l[7:6]),
     .reset_r(reset_r[7:6]), .reset_l(reset_l[7:6]),
     .pgate_r(pgate_r[7:6]), .pgate_l(pgate_l[7:6]), .q_b({net39[280],
     net39[281], net39[282], net39[283], net39[284], net39[285],
     net39[286], net39[287]}), .q({net40[280], net40[281], net40[282],
     net40[283], net40[284], net40[285], net40[286], net40[287]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[7:6]), .r_gnd_r(r_gnd_r[7:6]));
cram_2x2x2_ice8p I_mem2x2x2t_2_ ( .wl_r(wl_r[5:4]), .wl_l(wl_l[5:4]),
     .reset_r(reset_r[5:4]), .reset_l(reset_l[5:4]),
     .pgate_r(pgate_r[5:4]), .pgate_l(pgate_l[5:4]), .q_b({net39[288],
     net39[289], net39[290], net39[291], net39[292], net39[293],
     net39[294], net39[295]}), .q({net40[288], net40[289], net40[290],
     net40[291], net40[292], net40[293], net40[294], net40[295]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[5:4]), .r_gnd_r(r_gnd_r[5:4]));
cram_2x2x2_ice8p I_mem2x2x2t_1_ ( .wl_r(wl_r[3:2]), .wl_l(wl_l[3:2]),
     .reset_r(reset_r[3:2]), .reset_l(reset_l[3:2]),
     .pgate_r(pgate_r[3:2]), .pgate_l(pgate_l[3:2]), .q_b({net39[296],
     net39[297], net39[298], net39[299], net39[300], net39[301],
     net39[302], net39[303]}), .q({net40[296], net40[297], net40[298],
     net40[299], net40[300], net40[301], net40[302], net40[303]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[3:2]), .r_gnd_r(r_gnd_r[3:2]));
cram_2x2x2_ice8p I_mem2x2x2t_0_ ( .wl_r(wl_r[1:0]), .wl_l(wl_l[1:0]),
     .reset_r(reset_r[1:0]), .reset_l(reset_l[1:0]),
     .pgate_r(pgate_r[1:0]), .pgate_l(pgate_l[1:0]), .q_b({net39[304],
     net39[305], net39[306], net39[307], net39[308], net39[309],
     net39[310], net39[311]}), .q({net40[304], net40[305], net40[306],
     net40[307], net40[308], net40[309], net40[310], net40[311]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[1:0]), .r_gnd_r(r_gnd_r[1:0]));

endmodule
// Library - xpmem, Cell - cram2x2x5, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module cram2x2x5 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [19:0]  q;
output [19:0]  q_b;

inout [9:0]  bl;

input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  r_gnd;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - sbox11to9_p2_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:57 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox11to9_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  b;

input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_l10 ( .prog(prog), .in6(t[4]), .in5(t[10]), .in4(r[2]),
     .in3(r[10]), .in2(r[7]), .in1(b[10]), .in0(b[5]), .out(l[10]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t10 ( .prog(prog), .in6(r[4]), .in5(r[10]), .in4(b[2]),
     .in3(b[10]), .in2(b[7]), .in1(l[10]), .in0(l[5]), .out(t[10]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t11 ( .prog(prog), .in6(r[5]), .in5(r[11]), .in4(b[3]),
     .in3(b[11]), .in2(b[8]), .in1(l[11]), .in0(l[6]), .out(t[11]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t9 ( .prog(prog), .in6(r[3]), .in5(r[9]), .in4(b[1]),
     .in3(b[9]), .in2(b[6]), .in1(l[9]), .in0(l[4]), .out(t[9]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l11 ( .prog(prog), .in6(t[5]), .in5(t[11]), .in4(r[3]),
     .in3(r[11]), .in2(r[8]), .in1(b[11]), .in0(b[6]), .out(l[11]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l9 ( .prog(prog), .in6(t[3]), .in5(t[9]), .in4(r[1]),
     .in3(r[9]), .in2(r[6]), .in1(b[9]), .in0(b[4]), .out(l[9]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox11to9_p1_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:57 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox11to9_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  b;
inout [11:0]  t;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_r10 ( .prog(prog), .in6(b[4]), .in5(b[10]), .in4(l[2]),
     .in3(l[10]), .in2(l[7]), .in1(t[10]), .in0(t[5]), .out(r[10]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b10 ( .prog(prog), .in6(l[4]), .in5(l[10]), .in4(t[2]),
     .in3(t[10]), .in2(t[7]), .in1(r[10]), .in0(r[5]), .out(b[10]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b11 ( .prog(prog), .in6(l[5]), .in5(l[11]), .in4(t[3]),
     .in3(t[11]), .in2(t[8]), .in1(r[11]), .in0(r[6]), .out(b[11]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b9 ( .prog(prog), .in6(l[3]), .in5(l[9]), .in4(t[1]),
     .in3(t[9]), .in2(t[6]), .in1(r[9]), .in0(r[4]), .out(b[9]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r11 ( .prog(prog), .in6(b[5]), .in5(b[11]), .in4(l[3]),
     .in3(l[11]), .in2(l[8]), .in1(t[11]), .in0(t[6]), .out(r[11]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r9 ( .prog(prog), .in6(b[3]), .in5(b[9]), .in4(l[1]),
     .in3(l[9]), .in2(l[6]), .in1(t[9]), .in0(t[4]), .out(r[9]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox8to6_p2_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:58 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox8to6_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  t;

input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I554 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_l7 ( .prog(prog), .in6(t[1]), .in5(t[7]), .in4(r[11]),
     .in3(r[7]), .in2(r[4]), .in1(b[7]), .in0(b[2]), .out(l[7]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t7 ( .prog(prog), .in6(r[1]), .in5(r[7]), .in4(b[11]),
     .in3(b[7]), .in2(b[4]), .in1(l[7]), .in0(l[2]), .out(t[7]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t8 ( .prog(prog), .in6(r[2]), .in5(r[8]), .in4(b[0]),
     .in3(b[8]), .in2(b[5]), .in1(l[8]), .in0(l[3]), .out(t[8]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t6 ( .prog(prog), .in6(r[0]), .in5(r[6]), .in4(b[10]),
     .in3(b[6]), .in2(b[3]), .in1(l[6]), .in0(l[1]), .out(t[6]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l8 ( .prog(prog), .in6(t[2]), .in5(t[8]), .in4(r[0]),
     .in3(r[8]), .in2(r[5]), .in1(b[8]), .in0(b[3]), .out(l[8]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l6 ( .prog(prog), .in6(t[0]), .in5(t[6]), .in4(r[10]),
     .in3(r[6]), .in2(r[3]), .in1(b[6]), .in0(b[1]), .out(l[6]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox8to6_p1_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:58 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox8to6_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  t;
inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_r7 ( .prog(prog), .in6(b[1]), .in5(b[7]), .in4(l[11]),
     .in3(l[7]), .in2(l[4]), .in1(t[7]), .in0(t[2]), .out(r[7]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b7 ( .prog(prog), .in6(l[1]), .in5(l[7]), .in4(t[11]),
     .in3(t[7]), .in2(t[4]), .in1(r[7]), .in0(r[2]), .out(b[7]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b8 ( .prog(prog), .in6(l[2]), .in5(l[8]), .in4(t[0]),
     .in3(t[8]), .in2(t[5]), .in1(r[8]), .in0(r[3]), .out(b[8]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b6 ( .prog(prog), .in6(l[0]), .in5(l[6]), .in4(t[10]),
     .in3(t[6]), .in2(t[3]), .in1(r[6]), .in0(r[1]), .out(b[6]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r8 ( .prog(prog), .in6(b[2]), .in5(b[8]), .in4(l[0]),
     .in3(l[8]), .in2(l[5]), .in1(t[8]), .in0(t[3]), .out(r[8]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r6 ( .prog(prog), .in6(b[0]), .in5(b[6]), .in4(l[10]),
     .in3(l[6]), .in2(l[3]), .in1(t[6]), .in0(t[1]), .out(r[6]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox5to3_p2_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:57 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox5to3_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;
inout [9:0]  bl;
inout [11:0]  t;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  reset_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_l4 ( .prog(prog), .in6(t[10]), .in5(t[4]), .in4(r[8]),
     .in3(r[4]), .in2(r[1]), .in1(b[4]), .in0(b[11]), .out(l[4]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t4 ( .prog(prog), .in6(r[10]), .in5(r[4]), .in4(b[8]),
     .in3(b[4]), .in2(b[1]), .in1(l[4]), .in0(l[11]), .out(t[4]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t5 ( .prog(prog), .in6(r[11]), .in5(r[5]), .in4(b[9]),
     .in3(b[5]), .in2(b[2]), .in1(l[5]), .in0(l[0]), .out(t[5]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t3 ( .prog(prog), .in6(r[9]), .in5(r[3]), .in4(b[7]),
     .in3(b[3]), .in2(b[0]), .in1(l[3]), .in0(l[10]), .out(t[3]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l5 ( .prog(prog), .in6(t[11]), .in5(t[5]), .in4(r[9]),
     .in3(r[5]), .in2(r[2]), .in1(b[5]), .in0(b[0]), .out(l[5]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l3 ( .prog(prog), .in6(t[9]), .in5(t[3]), .in4(r[7]),
     .in3(r[3]), .in2(r[0]), .in1(b[3]), .in0(b[10]), .out(l[3]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - sbtlibn65lp, Cell - oai2211x2_hvt, View - schematic
// LAST TIME SAVED: Aug  3 19:21:56 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module oai2211x2_hvt ( Y, A0, A1, B0, B1, C0, D0 );
output  Y;

input  A0, A1, B0, B1, C0, D0;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M2 ( .D(Y), .B(VDD_), .G(C0), .S(vdd_));
P_11_LPHVT  M18 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
P_11_LPHVT  M8 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
P_11_LPHVT  M19 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
P_11_LPHVT  M7 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));
P_11_LPHVT  M12 ( .D(Y), .B(VDD_), .G(D0), .S(vdd_));
N_11_LPHVT  M10 ( .D(net040), .B(GND_), .G(A1), .S(net024));
N_11_LPHVT  M13 ( .D(net040), .B(GND_), .G(A0), .S(net024));
N_11_LPHVT  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
N_11_LPHVT  M11 ( .D(Y), .B(GND_), .G(C0), .S(net044));
N_11_LPHVT  M0 ( .D(net044), .B(GND_), .G(D0), .S(net040));
N_11_LPHVT  M1 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));

endmodule
// Library - leafcell, Cell - sbox5to3_p1_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:57 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox5to3_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  b;
inout [11:0]  l;

input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_r4 ( .prog(prog), .in6(b[10]), .in5(b[4]), .in4(l[8]),
     .in3(l[4]), .in2(l[1]), .in1(t[4]), .in0(t[11]), .out(r[4]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b4 ( .prog(prog), .in6(l[10]), .in5(l[4]), .in4(t[8]),
     .in3(t[4]), .in2(t[1]), .in1(r[4]), .in0(r[11]), .out(b[4]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b5 ( .prog(prog), .in6(l[11]), .in5(l[5]), .in4(t[9]),
     .in3(t[5]), .in2(t[2]), .in1(r[5]), .in0(r[0]), .out(b[5]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b3 ( .prog(prog), .in6(l[9]), .in5(l[3]), .in4(t[7]),
     .in3(t[3]), .in2(t[0]), .in1(r[3]), .in0(r[10]), .out(b[3]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r5 ( .prog(prog), .in6(b[11]), .in5(b[5]), .in4(l[9]),
     .in3(l[5]), .in2(l[2]), .in1(t[5]), .in0(t[0]), .out(r[5]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r3 ( .prog(prog), .in6(b[9]), .in5(b[3]), .in4(l[7]),
     .in3(l[3]), .in2(l[0]), .in1(t[3]), .in0(t[10]), .out(r[3]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox2to0_p2_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:57 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox2to0_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  b;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_l1 ( .prog(prog), .in6(t[7]), .in5(t[1]), .in4(r[5]),
     .in3(r[1]), .in2(r[10]), .in1(b[1]), .in0(b[8]), .out(l[1]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_l0 ( .prog(prog), .in6(t[6]), .in5(t[0]), .in4(r[4]),
     .in3(r[0]), .in2(r[9]), .in1(b[0]), .in0(b[7]), .out(l[0]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));
sbox7to1_220 I_t1 ( .prog(prog), .in6(r[7]), .in5(r[1]), .in4(b[5]),
     .in3(b[1]), .in2(b[10]), .in1(l[1]), .in0(l[8]), .out(t[1]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_l2 ( .prog(prog), .in6(t[8]), .in5(t[2]), .in4(r[6]),
     .in3(r[2]), .in2(r[11]), .in1(b[2]), .in0(b[9]), .out(l[2]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_t2 ( .prog(prog), .in6(r[8]), .in5(r[2]), .in4(b[6]),
     .in3(b[2]), .in2(b[11]), .in1(l[2]), .in0(l[9]), .out(t[2]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t0 ( .prog(prog), .in6(r[6]), .in5(r[0]), .in4(b[4]),
     .in3(b[0]), .in2(b[9]), .in1(l[0]), .in0(l[7]), .out(t[0]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));

endmodule
// Library - leafcell, Cell - sbox2to0_p1_v2, View - schematic
// LAST TIME SAVED: Jul 30 21:54:57 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox2to0_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  l;
inout [11:0]  t;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_r1 ( .prog(prog), .in6(b[7]), .in5(b[1]), .in4(l[5]),
     .in3(l[1]), .in2(l[10]), .in1(t[1]), .in0(t[8]), .out(r[1]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_r0 ( .prog(prog), .in6(b[6]), .in5(b[0]), .in4(l[4]),
     .in3(l[0]), .in2(l[9]), .in1(t[0]), .in0(t[7]), .out(r[0]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));
sbox7to1_220 I_b1 ( .prog(prog), .in6(l[7]), .in5(l[1]), .in4(t[5]),
     .in3(t[1]), .in2(t[10]), .in1(r[1]), .in0(r[8]), .out(b[1]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_r2 ( .prog(prog), .in6(b[8]), .in5(b[2]), .in4(l[6]),
     .in3(l[2]), .in2(l[11]), .in1(t[2]), .in0(t[9]), .out(r[2]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_b2 ( .prog(prog), .in6(l[8]), .in5(l[2]), .in4(t[6]),
     .in3(t[2]), .in2(t[11]), .in1(r[2]), .in0(r[9]), .out(b[2]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b0 ( .prog(prog), .in6(l[6]), .in5(l[0]), .in4(t[4]),
     .in3(t[0]), .in2(t[9]), .in1(r[0]), .in0(r[7]), .out(b[0]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));

endmodule
// Library - leafcell, Cell - span4_switchandmem_v3, View - schematic
// LAST TIME SAVED: Jul 30 21:54:58 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module span4_switchandmem_v3 ( c, cc, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [15:8]  cc;
output [7:0]  c;

inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  t;
inout [9:0]  bl;
inout [11:0]  l;

input [15:0]  pgate;
input [15:0]  reset_b;
input [15:0]  wl;
input [15:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  n5;

wire  [19:0]  n4;

wire  [19:0]  n0;

wire  [19:0]  n6;

wire  [19:0]  n1;

wire  [19:0]  n7;

wire  [19:0]  n2;

wire  [19:0]  n3;

wire  [19:0]  net0250;

wire  [19:0]  net0248;

wire  [19:0]  net0245;

wire  [19:0]  net0241;

wire  [19:0]  net0236;

wire  [19:0]  net0189;

wire  [19:0]  net0177;

wire  [19:0]  net0201;



sbox11to9_p2_v2 I_sbox11to9_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0241[0], net0241[1], net0241[2], net0241[3],
     net0241[4], net0241[5], net0241[6], net0241[7], net0241[8],
     net0241[9], net0241[10], net0241[11], net0241[12], net0241[13],
     net0241[14], net0241[15], net0241[16], net0241[17], net0241[18],
     net0241[19]}), .cbit({n7[19:8], cc[15], n7[6], cc[14], n7[4:0]}),
     .wl(wl[15:14]), .vdd_cntl(vdd_cntl[15:14]),
     .reset_b(reset_b[15:14]), .pgate(pgate[15:14]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox11to9_p1_v2 I_sbox11to9_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0236[0], net0236[1], net0236[2], net0236[3],
     net0236[4], net0236[5], net0236[6], net0236[7], net0236[8],
     net0236[9], net0236[10], net0236[11], net0236[12], net0236[13],
     net0236[14], net0236[15], net0236[16], net0236[17], net0236[18],
     net0236[19]}), .cbit({n6[19:8], cc[13], n6[6], cc[12], n6[4:0]}),
     .wl(wl[13:12]), .vdd_cntl(vdd_cntl[13:12]),
     .reset_b(reset_b[13:12]), .pgate(pgate[13:12]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox8to6_p2_v2 I_sbox8to6_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0248[0], net0248[1], net0248[2], net0248[3],
     net0248[4], net0248[5], net0248[6], net0248[7], net0248[8],
     net0248[9], net0248[10], net0248[11], net0248[12], net0248[13],
     net0248[14], net0248[15], net0248[16], net0248[17], net0248[18],
     net0248[19]}), .cbit({n5[19:8], cc[11], n5[6], cc[10], n5[4:0]}),
     .wl(wl[11:10]), .vdd_cntl(vdd_cntl[11:10]),
     .reset_b(reset_b[11:10]), .pgate(pgate[11:10]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox8to6_p1_v2 I_sbox8to6_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0177[0], net0177[1], net0177[2], net0177[3],
     net0177[4], net0177[5], net0177[6], net0177[7], net0177[8],
     net0177[9], net0177[10], net0177[11], net0177[12], net0177[13],
     net0177[14], net0177[15], net0177[16], net0177[17], net0177[18],
     net0177[19]}), .cbit({n4[19:8], cc[9], n4[6], cc[8], n4[4:0]}),
     .wl(wl[9:8]), .vdd_cntl(vdd_cntl[9:8]), .reset_b(reset_b[9:8]),
     .pgate(pgate[9:8]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox5to3_p2_v2 I_sbox5to3_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0189[0], net0189[1], net0189[2], net0189[3],
     net0189[4], net0189[5], net0189[6], net0189[7], net0189[8],
     net0189[9], net0189[10], net0189[11], net0189[12], net0189[13],
     net0189[14], net0189[15], net0189[16], net0189[17], net0189[18],
     net0189[19]}), .cbit({n3[19:8], c[7], n3[6], c[6], n3[4:0]}),
     .wl(wl[7:6]), .vdd_cntl(vdd_cntl[7:6]), .reset_b(reset_b[7:6]),
     .pgate(pgate[7:6]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox5to3_p1_v2 I_sbox5to3_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0201[0], net0201[1], net0201[2], net0201[3],
     net0201[4], net0201[5], net0201[6], net0201[7], net0201[8],
     net0201[9], net0201[10], net0201[11], net0201[12], net0201[13],
     net0201[14], net0201[15], net0201[16], net0201[17], net0201[18],
     net0201[19]}), .cbit({n2[19:8], c[5], n2[6], c[4], n2[4:0]}),
     .wl(wl[5:4]), .vdd_cntl(vdd_cntl[5:4]), .reset_b(reset_b[5:4]),
     .pgate(pgate[5:4]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox2to0_p2_v2 I_sbox2to0_p2_v2 ( .b(b[11:0]), .cbitb({net0245[0],
     net0245[1], net0245[2], net0245[3], net0245[4], net0245[5],
     net0245[6], net0245[7], net0245[8], net0245[9], net0245[10],
     net0245[11], net0245[12], net0245[13], net0245[14], net0245[15],
     net0245[16], net0245[17], net0245[18], net0245[19]}),
     .cbit({n1[19:8], c[3], n1[6], c[2], n1[4:0]}), .wl(wl[3:2]),
     .vdd_cntl(vdd_cntl[3:2]), .reset_b(reset_b[3:2]), .prog(prog),
     .pgate(pgate[3:2]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox2to0_p1_v2 I_sbox2to0_p1_v2 ( .cbitb({net0250[0], net0250[1],
     net0250[2], net0250[3], net0250[4], net0250[5], net0250[6],
     net0250[7], net0250[8], net0250[9], net0250[10], net0250[11],
     net0250[12], net0250[13], net0250[14], net0250[15], net0250[16],
     net0250[17], net0250[18], net0250[19]}), .cbit({n0[19:8], c[1],
     n0[6], c[0], n0[4:0]}), .wl(wl[1:0]), .vdd_cntl(vdd_cntl[1:0]),
     .reset_b(reset_b[1:0]), .prog(prog), .pgate(pgate[1:0]),
     .t(t[11:0]), .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]), .b(b[11:0]));

endmodule
// Library - leafcell, Cell - span4_ice8p, View - schematic
// LAST TIME SAVED: Jul 30 21:54:58 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module span4_ice8p ( bram_cbit, ccntrl_cbit, bl, sp4_h_l, sp4_h_r,
     sp4_v_b, sp4_v_t, pgate, prog, reset_b, vdd_cntl, wl );


input  prog;

output [7:0]  bram_cbit;
output [7:0]  ccntrl_cbit;

inout [9:0]  bl;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_t;
inout [47:0]  sp4_h_r;

input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  reset_b;
input [15:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  sp4_h_r_mid;

wire  [11:0]  sp4_v_b_mid;



RM6  R1_27_ ( .MINUS(sp4_h_r[47]), .PLUS(sp4_h_l[34]));
RM6  R1_26_ ( .MINUS(sp4_h_r[46]), .PLUS(sp4_h_l[35]));
RM6  R1_25_ ( .MINUS(sp4_h_r[45]), .PLUS(sp4_h_l[32]));
RM6  R1_24_ ( .MINUS(sp4_h_r[44]), .PLUS(sp4_h_l[33]));
RM6  R1_23_ ( .MINUS(sp4_h_r[43]), .PLUS(sp4_h_l[30]));
RM6  R1_22_ ( .MINUS(sp4_h_r[42]), .PLUS(sp4_h_l[31]));
RM6  R1_21_ ( .MINUS(sp4_h_r[41]), .PLUS(sp4_h_l[28]));
RM6  R1_20_ ( .MINUS(sp4_h_r[40]), .PLUS(sp4_h_l[29]));
RM6  R1_19_ ( .MINUS(sp4_h_r[39]), .PLUS(sp4_h_l[26]));
RM6  R1_18_ ( .MINUS(sp4_h_r[38]), .PLUS(sp4_h_l[27]));
RM6  R1_17_ ( .MINUS(sp4_h_r[37]), .PLUS(sp4_h_l[24]));
RM6  R1_16_ ( .MINUS(sp4_h_r[36]), .PLUS(sp4_h_l[25]));
RM6  R1_15_ ( .MINUS(sp4_h_r[35]), .PLUS(sp4_h_l[22]));
RM6  R1_14_ ( .MINUS(sp4_h_r[34]), .PLUS(sp4_h_l[23]));
RM6  R1_13_ ( .MINUS(sp4_h_r[23]), .PLUS(sp4_h_l[10]));
RM6  R1_12_ ( .MINUS(sp4_h_r[22]), .PLUS(sp4_h_l[11]));
RM6  R1_11_ ( .MINUS(sp4_h_r_mid[11]), .PLUS(sp4_h_l[46]));
RM6  R1_10_ ( .MINUS(sp4_h_r_mid[10]), .PLUS(sp4_h_l[47]));
RM6  R1_9_ ( .MINUS(sp4_h_r_mid[9]), .PLUS(sp4_h_l[44]));
RM6  R1_8_ ( .MINUS(sp4_h_r_mid[8]), .PLUS(sp4_h_l[45]));
RM6  R1_7_ ( .MINUS(sp4_h_r_mid[7]), .PLUS(sp4_h_l[42]));
RM6  R1_6_ ( .MINUS(sp4_h_r_mid[6]), .PLUS(sp4_h_l[43]));
RM6  R1_5_ ( .MINUS(sp4_h_r_mid[5]), .PLUS(sp4_h_l[40]));
RM6  R1_4_ ( .MINUS(sp4_h_r_mid[4]), .PLUS(sp4_h_l[41]));
RM6  R1_3_ ( .MINUS(sp4_h_r_mid[3]), .PLUS(sp4_h_l[38]));
RM6  R1_2_ ( .MINUS(sp4_h_r_mid[2]), .PLUS(sp4_h_l[39]));
RM6  R1_1_ ( .MINUS(sp4_h_r_mid[1]), .PLUS(sp4_h_l[36]));
RM6  R1_0_ ( .MINUS(sp4_h_r_mid[0]), .PLUS(sp4_h_l[37]));
RM6  R2_19_ ( .MINUS(sp4_h_r[33]), .PLUS(sp4_h_l[20]));
RM6  R2_18_ ( .MINUS(sp4_h_r[32]), .PLUS(sp4_h_l[21]));
RM6  R2_17_ ( .MINUS(sp4_h_r[31]), .PLUS(sp4_h_l[18]));
RM6  R2_16_ ( .MINUS(sp4_h_r[30]), .PLUS(sp4_h_l[19]));
RM6  R2_15_ ( .MINUS(sp4_h_r[29]), .PLUS(sp4_h_l[16]));
RM6  R2_14_ ( .MINUS(sp4_h_r[28]), .PLUS(sp4_h_l[17]));
RM6  R2_13_ ( .MINUS(sp4_h_r[27]), .PLUS(sp4_h_l[14]));
RM6  R2_12_ ( .MINUS(sp4_h_r[26]), .PLUS(sp4_h_l[15]));
RM6  R2_11_ ( .MINUS(sp4_h_r[25]), .PLUS(sp4_h_l[12]));
RM6  R2_10_ ( .MINUS(sp4_h_r[24]), .PLUS(sp4_h_l[13]));
RM6  R2_9_ ( .MINUS(sp4_h_r[21]), .PLUS(sp4_h_l[8]));
RM6  R2_8_ ( .MINUS(sp4_h_r[20]), .PLUS(sp4_h_l[9]));
RM6  R2_7_ ( .MINUS(sp4_h_r[19]), .PLUS(sp4_h_l[6]));
RM6  R2_6_ ( .MINUS(sp4_h_r[18]), .PLUS(sp4_h_l[7]));
RM6  R2_5_ ( .MINUS(sp4_h_r[17]), .PLUS(sp4_h_l[4]));
RM6  R2_4_ ( .MINUS(sp4_h_r[16]), .PLUS(sp4_h_l[5]));
RM6  R2_3_ ( .MINUS(sp4_h_r[15]), .PLUS(sp4_h_l[2]));
RM6  R2_2_ ( .MINUS(sp4_h_r[14]), .PLUS(sp4_h_l[3]));
RM6  R2_1_ ( .MINUS(sp4_h_r[13]), .PLUS(sp4_h_l[0]));
RM6  R2_0_ ( .MINUS(sp4_h_r[12]), .PLUS(sp4_h_l[1]));
RM7  R0_47_ ( .MINUS(sp4_v_b[47]), .PLUS(sp4_v_t[34]));
RM7  R0_46_ ( .MINUS(sp4_v_b[46]), .PLUS(sp4_v_t[35]));
RM7  R0_45_ ( .MINUS(sp4_v_b[45]), .PLUS(sp4_v_t[32]));
RM7  R0_44_ ( .MINUS(sp4_v_b[44]), .PLUS(sp4_v_t[33]));
RM7  R0_43_ ( .MINUS(sp4_v_b[43]), .PLUS(sp4_v_t[30]));
RM7  R0_42_ ( .MINUS(sp4_v_b[42]), .PLUS(sp4_v_t[31]));
RM7  R0_41_ ( .MINUS(sp4_v_b[41]), .PLUS(sp4_v_t[28]));
RM7  R0_40_ ( .MINUS(sp4_v_b[40]), .PLUS(sp4_v_t[29]));
RM7  R0_39_ ( .MINUS(sp4_v_b[39]), .PLUS(sp4_v_t[26]));
RM7  R0_38_ ( .MINUS(sp4_v_b[38]), .PLUS(sp4_v_t[27]));
RM7  R0_37_ ( .MINUS(sp4_v_b[37]), .PLUS(sp4_v_t[24]));
RM7  R0_36_ ( .MINUS(sp4_v_b[36]), .PLUS(sp4_v_t[25]));
RM7  R0_35_ ( .MINUS(sp4_v_b[35]), .PLUS(sp4_v_t[22]));
RM7  R0_34_ ( .MINUS(sp4_v_b[34]), .PLUS(sp4_v_t[23]));
RM7  R0_33_ ( .MINUS(sp4_v_b[33]), .PLUS(sp4_v_t[20]));
RM7  R0_32_ ( .MINUS(sp4_v_b[32]), .PLUS(sp4_v_t[21]));
RM7  R0_31_ ( .MINUS(sp4_v_b[31]), .PLUS(sp4_v_t[18]));
RM7  R0_30_ ( .MINUS(sp4_v_b[30]), .PLUS(sp4_v_t[19]));
RM7  R0_29_ ( .MINUS(sp4_v_b[29]), .PLUS(sp4_v_t[16]));
RM7  R0_28_ ( .MINUS(sp4_v_b[28]), .PLUS(sp4_v_t[17]));
RM7  R0_27_ ( .MINUS(sp4_v_b[27]), .PLUS(sp4_v_t[14]));
RM7  R0_26_ ( .MINUS(sp4_v_b[26]), .PLUS(sp4_v_t[15]));
RM7  R0_25_ ( .MINUS(sp4_v_b[25]), .PLUS(sp4_v_t[12]));
RM7  R0_24_ ( .MINUS(sp4_v_b[24]), .PLUS(sp4_v_t[13]));
RM7  R0_23_ ( .MINUS(sp4_v_b[23]), .PLUS(sp4_v_t[10]));
RM7  R0_22_ ( .MINUS(sp4_v_b[22]), .PLUS(sp4_v_t[11]));
RM7  R0_21_ ( .MINUS(sp4_v_b[21]), .PLUS(sp4_v_t[8]));
RM7  R0_20_ ( .MINUS(sp4_v_b[20]), .PLUS(sp4_v_t[9]));
RM7  R0_19_ ( .MINUS(sp4_v_b[19]), .PLUS(sp4_v_t[6]));
RM7  R0_18_ ( .MINUS(sp4_v_b[18]), .PLUS(sp4_v_t[7]));
RM7  R0_17_ ( .MINUS(sp4_v_b[17]), .PLUS(sp4_v_t[4]));
RM7  R0_16_ ( .MINUS(sp4_v_b[16]), .PLUS(sp4_v_t[5]));
RM7  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[2]));
RM7  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[3]));
RM7  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[0]));
RM7  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[1]));
RM7  R0_11_ ( .MINUS(sp4_v_b_mid[11]), .PLUS(sp4_v_t[46]));
RM7  R0_10_ ( .MINUS(sp4_v_b_mid[10]), .PLUS(sp4_v_t[47]));
RM7  R0_9_ ( .MINUS(sp4_v_b_mid[9]), .PLUS(sp4_v_t[44]));
RM7  R0_8_ ( .MINUS(sp4_v_b_mid[8]), .PLUS(sp4_v_t[45]));
RM7  R0_7_ ( .MINUS(sp4_v_b_mid[7]), .PLUS(sp4_v_t[42]));
RM7  R0_6_ ( .MINUS(sp4_v_b_mid[6]), .PLUS(sp4_v_t[43]));
RM7  R0_5_ ( .MINUS(sp4_v_b_mid[5]), .PLUS(sp4_v_t[40]));
RM7  R0_4_ ( .MINUS(sp4_v_b_mid[4]), .PLUS(sp4_v_t[41]));
RM7  R0_3_ ( .MINUS(sp4_v_b_mid[3]), .PLUS(sp4_v_t[38]));
RM7  R0_2_ ( .MINUS(sp4_v_b_mid[2]), .PLUS(sp4_v_t[39]));
RM7  R0_1_ ( .MINUS(sp4_v_b_mid[1]), .PLUS(sp4_v_t[36]));
RM7  R0_0_ ( .MINUS(sp4_v_b_mid[0]), .PLUS(sp4_v_t[37]));
span4_switchandmem_v3 I_span4_switchandmem_rev ( .cc(ccntrl_cbit[7:0]),
     .c(bram_cbit[7:0]), .wl(wl[15:0]), .vdd_cntl(vdd_cntl[15:0]),
     .reset_b(reset_b[15:0]), .prog(prog), .pgate(pgate[15:0]),
     .t(sp4_v_b_mid[11:0]), .r(sp4_h_r[11:0]), .l(sp4_h_r_mid[11:0]),
     .bl(bl[9:0]), .b(sp4_v_b[11:0]));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev0, View - schematic
// LAST TIME SAVED: Jul 30 23:15:00 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module clkmandcmuxrev0 ( clk, clkb, glb2local, s_r, cbit, cbitb,
     glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, min0, min1,
     min2, min3, prog );
output  clk, clkb, s_r;

input  prog;

output [3:0]  glb2local;

input [7:0]  min1;
input [7:0]  min3;
input [7:0]  min0;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g0;
input [7:0]  min2;
input [5:0]  lc_trk_g3;
input [31:0]  cbit;
input [31:0]  cbitb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



clk_mux12to1_icc I_clkmux12to1 ( .prog(prog), .min({lc_trk_g3[1],
     lc_trk_g2[0], lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}),
     .clk(clk), .clkb(clkb), .cbitb({cbitb[31], cbitb[4], cbitb[3],
     cbitb[2], cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3],
     cbit[2], cbit[1], cbit[0]}), .cenb(ceb));
clk_mux8to1 I_clkmux8to1_0 ( .prog(prog), .inmuxo(glb2local[0]),
     .min(min3[7:0]), .cbit(cbit[16:13]), .cbitb(cbitb[16:13]));
clk_mux8to1 I_clkmux8to1_1 ( .prog(prog), .inmuxo(glb2local[1]),
     .min(min2[7:0]), .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I_clkmux8to1_3 ( .prog(prog), .inmuxo(glb2local[3]),
     .min(min0[7:0]), .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));
clk_mux8to1 I_clkmux8to1_2 ( .prog(prog), .inmuxo(glb2local[2]),
     .min(min1[7:0]), .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
ce_clkm8to1 I_cemux8to1 ( .cbitb(cbitb[8:5]), .min({lc_trk_g3[3],
     lc_trk_g2[2], lc_trk_g1[3], lc_trk_g0[2], glb_netwk[7],
     glb_netwk[5], glb_netwk[3], glb_netwk[1]}), .cbit(cbit[8:5]),
     .moutb(ceb), .prog(prog));
sr_clkm8to1 I_srmux8to1 ( .cbitb(cbitb[12:9]), .min({lc_trk_g3[5],
     lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4], glb_netwk[6],
     glb_netwk[4], glb_netwk[2], glb_netwk[0]}), .cbit(cbit[12:9]),
     .mout(s_r), .prog(prog));

endmodule
// Library - leafcell, Cell - sbox1, View - schematic
// LAST TIME SAVED: Jul 30 21:54:57 2011
// NETLIST TIME: Jan 18 18:48:19 2012
`timescale 1ns / 1ns 

module sbox1 ( b, l, r, t, c, cb, prog );
inout  b, l, r, t;

input  prog;

input [7:0]  c;
input [7:0]  cb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



sbox1m3to1_icc I232 ( .in2(r), .cb(cb[7:6]), .op(t), .in0(l), .in1(b),
     .c(c[7:6]), .prog(prog));
sbox1m3to1_icc I230 ( .in2(r), .cb(cb[3:2]), .op(l), .in0(b), .in1(t),
     .c(c[3:2]), .prog(prog));
sbox1m3to1_icc I226 ( .in2(r), .cb(cb[1:0]), .op(b), .in0(l), .in1(t),
     .c(c[1:0]), .prog(prog));
sbox1m3to1_icc I231 ( .in2(b), .cb(cb[5:4]), .op(r), .in0(l), .in1(t),
     .c(c[5:4]), .prog(prog));

endmodule
// Library - xpmem, Cell - cram16x4, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module cram16x4 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [63:0]  q_b;
output [63:0]  q;

inout [3:0]  bl;

input [15:0]  wl;
input [15:0]  r_gnd;
input [15:0]  pgate;
input [15:0]  reset_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



cram2x2 I16_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[1:0]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[15:14]));
cram2x2 I16_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[1:0]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[13:12]));
cram2x2 I16_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[1:0]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[11:10]));
cram2x2 I16_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[1:0]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[9:8]));
cram2x2 I16_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[1:0]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[7:6]));
cram2x2 I16_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[1:0]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[5:4]));
cram2x2 I16_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[1:0]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[3:2]));
cram2x2 I16_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[3:2]), .q_b(q_b[63:60]),
     .q(q[63:60]), .wl(wl[15:14]));
cram2x2 Imstake_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[3:2]), .q_b(q_b[59:56]),
     .q(q[59:56]), .wl(wl[13:12]));
cram2x2 Imstake_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[3:2]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[11:10]));
cram2x2 Imstake_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[3:2]), .q_b(q_b[51:48]), .q(q[51:48]),
     .wl(wl[9:8]));
cram2x2 Imstake_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[3:2]), .q_b(q_b[47:44]), .q(q[47:44]),
     .wl(wl[7:6]));
cram2x2 Imstake_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[3:2]), .q_b(q_b[43:40]), .q(q[43:40]),
     .wl(wl[5:4]));
cram2x2 Imstake_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[3:2]), .q_b(q_b[39:36]), .q(q[39:36]),
     .wl(wl[3:2]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[35:32]), .q(q[35:32]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - misc_module4_v3, View - schematic
// LAST TIME SAVED: Jul 30 21:54:55 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module misc_module4_v3 ( S_R, cbit, cbitb, clk, clkb, glb2local, sp4,
     bl, b, glb_netwk, l, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3,
     m, min0, min1, min2, min3, pgate, prog, r, reset_b, sp12,
     vdd_cntl, wl );
output  S_R, clk, clkb;


input  prog;

output [7:0]  sp4;
output [3:0]  glb2local;
output [63:0]  cbit;
output [63:0]  cbitb;

inout [3:0]  bl;

input [15:0]  vdd_cntl;
input [15:0]  wl;
input [1:0]  m;
input [1:0]  b;
input [5:0]  lc_trk_g2;
input [7:0]  min0;
input [1:0]  r;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g0;
input [7:0]  min2;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g3;
input [7:0]  min1;
input [7:0]  min3;
input [7:0]  sp12;
input [15:0]  pgate;
input [1:0]  l;
input [15:0]  reset_b;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  r_vdd;



P_11_LPHVT  M0_15_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[15]),
     .D(r_vdd[15]));
P_11_LPHVT  M0_14_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[14]),
     .D(r_vdd[14]));
P_11_LPHVT  M0_13_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[13]),
     .D(r_vdd[13]));
P_11_LPHVT  M0_12_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[12]),
     .D(r_vdd[12]));
P_11_LPHVT  M0_11_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[11]),
     .D(r_vdd[11]));
P_11_LPHVT  M0_10_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[10]),
     .D(r_vdd[10]));
P_11_LPHVT  M0_9_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[9]), .D(r_vdd[9]));
P_11_LPHVT  M0_8_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[8]), .D(r_vdd[8]));
P_11_LPHVT  M0_7_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[7]), .D(r_vdd[7]));
P_11_LPHVT  M0_6_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[6]), .D(r_vdd[6]));
P_11_LPHVT  M0_5_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[5]), .D(r_vdd[5]));
P_11_LPHVT  M0_4_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[4]), .D(r_vdd[4]));
P_11_LPHVT  M0_3_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[3]), .D(r_vdd[3]));
P_11_LPHVT  M0_2_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[2]), .D(r_vdd[2]));
P_11_LPHVT  M0_1_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[1]), .D(r_vdd[1]));
P_11_LPHVT  M0_0_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl[0]), .D(r_vdd[0]));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
clkmandcmuxrev0 I_clkmandcmuxrev0 ( .prog(progd),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]), .clk(clk),
     .clkb(clkb), .glb_netwk(glb_netwk[7:0]), .s_r(S_R),
     .glb2local(glb2local[3:0]), .cbit({cbit[2], cbit[1], cbit[0],
     cbit[27], cbit[25], cbit[26], cbit[24], cbit[23], cbit[21],
     cbit[22], cbit[20], cbit[19], cbit[17], cbit[18], cbit[16],
     cbit[15], cbit[13], cbit[14], cbit[12], cbit[31], cbit[29],
     cbit[30], cbit[28], cbit[11], cbit[9], cbit[10], cbit[8],
     cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}), .min2(min2[7:0]),
     .min1(min1[7:0]), .min0(min0[7:0]), .min3(min3[7:0]),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}));
sp12to4 I_sp12to4_7_ ( .prog(progd), .triout(sp4[7]),
     .cbitb(cbitb[62]), .drv(sp12[7]));
sp12to4 I_sp12to4_6_ ( .prog(progd), .triout(sp4[6]),
     .cbitb(cbitb[58]), .drv(sp12[6]));
sp12to4 I_sp12to4_5_ ( .prog(progd), .triout(sp4[5]),
     .cbitb(cbitb[54]), .drv(sp12[5]));
sp12to4 I_sp12to4_4_ ( .prog(progd), .triout(sp4[4]),
     .cbitb(cbitb[50]), .drv(sp12[4]));
sp12to4 I_sp12to4_3_ ( .prog(progd), .triout(sp4[3]),
     .cbitb(cbitb[46]), .drv(sp12[3]));
sp12to4 I_sp12to4_2_ ( .prog(progd), .triout(sp4[2]),
     .cbitb(cbitb[42]), .drv(sp12[2]));
sp12to4 I_sp12to4_1_ ( .prog(progd), .triout(sp4[1]), .cbitb(cbitb[5]),
     .drv(sp12[1]));
sp12to4 I_sp12to4_0_ ( .prog(progd), .triout(sp4[0]),
     .cbitb(cbitb[34]), .drv(sp12[0]));
sbox1 I_sbox1_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(progd));
sbox1 I_sbox1_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(progd));
cram16x4 I_cram16x4 ( .q(cbit[63:0]), .r_gnd(r_vdd[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));

endmodule
// Library - xpmem, Cell - cram2x2x6, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module cram2x2x6 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [23:0]  q;
output [23:0]  q_b;

inout [11:0]  bl;

input [1:0]  r_gnd;
input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_5_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - sbtlibn65lp, Cell - anor31_hvt, View - schematic
// LAST TIME SAVED: Aug  3 19:21:54 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module anor31_hvt ( Y, A, B, C, D );
output  Y;

input  A, B, C, D;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M4 ( .D(net35), .B(vdd_), .G(A), .S(vdd_));
P_11_LPHVT  M0 ( .D(net35), .B(vdd_), .G(B), .S(vdd_));
P_11_LPHVT  M2 ( .D(net35), .B(vdd_), .G(C), .S(vdd_));
P_11_LPHVT  M3 ( .D(Y), .B(vdd_), .G(D), .S(net35));
N_11_LPHVT  M1 ( .D(Y), .B(gnd_), .G(A), .S(net23));
N_11_LPHVT  M6 ( .D(net030), .B(gnd_), .G(C), .S(gnd_));
N_11_LPHVT  M5 ( .D(net23), .B(gnd_), .G(B), .S(net030));
N_11_LPHVT  M7 ( .D(Y), .B(gnd_), .G(D), .S(gnd_));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_base, View - schematic
// LAST TIME SAVED: Jul 30 21:54:52 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_base ( lc_trk_out, sp4_out, bl, min0, min1, min2,
     min3, pgate, prog, reset_b, sp12_in, vdd_cntl, wl );


input  prog;

output [1:0]  sp4_out;
output [3:0]  lc_trk_out;

inout [11:0]  bl;

input [15:0]  min1;
input [1:0]  vdd_cntl;
input [1:0]  sp12_in;
input [15:0]  min2;
input [15:0]  min0;
input [1:0]  pgate;
input [1:0]  reset_b;
input [15:0]  min3;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  cbitb;

wire  [23:0]  cbit;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net60));
g_mux I_mux2 ( .min(min2[15:0]), .prog(net60), .inmuxo(lc_trk_out[2]),
     .cbit({cbit[16], cbit[17], cbit[20], cbit[23], cbit[21]}),
     .cbitb({cbitb[16], cbitb[17], cbitb[20], cbitb[23], cbitb[21]}));
g_mux I_mux3 ( .min(min3[15:0]), .prog(net60), .inmuxo(lc_trk_out[3]),
     .cbit({cbit[18], cbit[19], cbit[22], cbit[15], cbit[13]}),
     .cbitb({cbitb[18], cbitb[19], cbitb[22], cbitb[15], cbitb[13]}));
g_mux I_mux1 ( .min(min1[15:0]), .prog(net60), .inmuxo(lc_trk_out[1]),
     .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}));
g_mux I_mux0 ( .min(min0[15:0]), .prog(net60), .inmuxo(lc_trk_out[0]),
     .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}));
cram2x2x6 I_mem2x2x6 ( .pgate(pgate[1:0]), .q(cbit[23:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[11:0]), .q_b(cbitb[23:0]));
sp12to4 I_sp12to4_1_ ( .triout(sp4_out[1]), .cbitb(cbitb[11]),
     .drv(sp12_in[1]), .prog(net60));
sp12to4 I_sp12to4_0_ ( .triout(sp4_out[0]), .cbitb(cbitb[9]),
     .drv(sp12_in[0]), .prog(net60));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0a, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g0a ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g0;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [1:0]  wl;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  bot_op;
input [7:0]  top_op;
input [1:0]  pgate;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  rgt_op;
input [7:0]  lft_op;
input [1:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[34], sp4_r_v_b[25]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[33], sp4_r_v_b[26]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[35], sp4_r_v_b[24]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[32], sp4_r_v_b[27]}),
     .sp4_out(sp4_v_b[13:12]), .sp12_in({sp12_v_b[3], sp12_v_b[1]}),
     .lc_trk_out(lc_trk_g0[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0b, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g0b ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, glb2local, lft_op,
     pgate, prog, reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op,
     vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g0;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;

input [7:0]  tnr_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [7:0]  tnl_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [1:0]  wl;
input [7:0]  rgt_op;
input [3:0]  glb2local;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], glb2local[1]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], glb2local[2]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], glb2local[0]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], glb2local[3]}),
     .sp4_out(sp4_v_b[15:14]), .sp12_in({sp12_v_b[7], sp12_v_b[5]}),
     .lc_trk_out(lc_trk_g0[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1a, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g1a ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g1;

inout [11:0]  bl;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_b;

input [7:0]  tnr_op;
input [1:0]  wl;
input [7:0]  tnl_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
input [7:0]  top_op;
input [7:0]  rgt_op;
input [7:0]  lft_op;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[25], sp4_r_v_b[1]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[26], sp4_r_v_b[2]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[24], sp4_r_v_b[0]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[27], sp4_r_v_b[3]}),
     .sp4_out(sp4_v_b[17:16]), .sp12_in({sp12_v_b[11], sp12_v_b[9]}),
     .lc_trk_out(lc_trk_g1[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1b, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g1b ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;

input [1:0]  pgate;
input [7:0]  tnr_op;
input [1:0]  reset_b;
input [7:0]  tnl_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
input [7:0]  top_op;
input [1:0]  wl;
input [7:0]  bnl_op;
input [1:0]  vdd_cntl;
input [7:0]  slf_op;
input [7:0]  rgt_op;
input [7:0]  lft_op;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], sp4_r_v_b[5]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], sp4_r_v_b[6]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], sp4_r_v_b[4]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], sp4_r_v_b[7]}),
     .sp4_out(sp4_v_b[19:18]), .sp12_in({sp12_v_b[15], sp12_v_b[13]}),
     .lc_trk_out(lc_trk_g1[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2a, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g2a ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g2;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_b;

input [1:0]  pgate;
input [7:0]  bot_op;
input [1:0]  reset_b;
input [7:0]  top_op;
input [7:0]  bnr_op;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [1:0]  wl;
input [7:0]  slf_op;
input [1:0]  vdd_cntl;
input [7:0]  rgt_op;
input [7:0]  lft_op;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[33], sp4_r_v_b[9]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[34], sp4_r_v_b[10]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[32], sp4_r_v_b[8]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[35], sp4_r_v_b[11]}),
     .sp4_out(sp4_v_b[21:20]), .sp12_in({sp12_v_b[19], sp12_v_b[17]}),
     .lc_trk_out(lc_trk_g2[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2b, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g2b ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g2;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;

input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  bot_op;
input [7:0]  top_op;
input [7:0]  bnr_op;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  rgt_op;
input [7:0]  lft_op;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[37], sp4_r_v_b[13]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[38], sp4_r_v_b[14]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[36], sp4_r_v_b[12]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[39], sp4_r_v_b[15]}),
     .sp4_out(sp4_v_b[23:22]), .sp12_in({sp12_v_b[23], sp12_v_b[21]}),
     .lc_trk_out(lc_trk_g2[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3a, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g3a ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g3;

inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  bot_op;
input [7:0]  bnr_op;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [1:0]  wl;
input [7:0]  slf_op;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [7:0]  top_op;
input [1:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[41], sp4_r_v_b[17]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[42], sp4_r_v_b[18]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[40], sp4_r_v_b[16]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[43], sp4_r_v_b[19]}),
     .sp4_out(sp4_h_r[13:12]), .sp12_in({sp12_h_r[2], sp12_h_r[0]}),
     .lc_trk_out(lc_trk_g3[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3b, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4_g3b ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g3;

inout [23:0]  sp12_h_r;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_r_v_b;

input [7:0]  top_op;
input [7:0]  bnr_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [7:0]  lft_op;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  bot_op;
input [7:0]  bnl_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base I_gmux_12to4_g3b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[45], sp4_r_v_b[21]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[46], sp4_r_v_b[22]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[44], sp4_r_v_b[20]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[47], sp4_r_v_b[23]}),
     .sp4_out(sp4_h_r[15:14]), .sp12_in({sp12_h_r[6], sp12_h_r[4]}),
     .lc_trk_out(lc_trk_g3[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4, View - schematic
// LAST TIME SAVED: Jul 30 21:54:52 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module gmux_sp12to4 ( lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, bl,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bnl_op, bnr_op,
     bot_op, glb2local, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g3;

inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_h_r;

input [7:0]  lft_op;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  top_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnr_op;
input [3:0]  glb2local;
input [7:0]  bnl_op;
input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  bot_op;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_g0a I_g0_30 ( .vdd_cntl(vdd_cntl[1:0]),
     .pgate(pgate[1:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp12_v_b(sp12_v_b[23:0]), .lc_trk_g0(lc_trk_g0[3:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g0b I_g0_74 ( .vdd_cntl(vdd_cntl[3:2]),
     .pgate(pgate[3:2]), .glb2local(glb2local[3:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .lc_trk_g0(lc_trk_g0[7:4]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[3:2]), .reset_b(reset_b[3:2]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g1a I_g1_30 ( .vdd_cntl(vdd_cntl[5:4]),
     .pgate(pgate[5:4]), .bl(bl[11:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]),
     .lft_op(lft_op[7:0]), .prog(prog), .rgt_op(rgt_op[7:0]),
     .reset_b(reset_b[5:4]), .slf_op(slf_op[7:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .wl(wl[5:4]), .lc_trk_g1(lc_trk_g1[3:0]));
gmux_sp12to4_g1b I_g1_74 ( .vdd_cntl(vdd_cntl[7:6]),
     .pgate(pgate[7:6]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g1(lc_trk_g1[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g2a I_g2_30 ( .vdd_cntl(vdd_cntl[9:8]), .wl(wl[9:8]),
     .reset_b(reset_b[9:8]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[3:0]), .pgate(pgate[9:8]));
gmux_sp12to4_g2b I_g2_74 ( .vdd_cntl(vdd_cntl[11:10]),
     .pgate(pgate[11:10]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[11:10]),
     .reset_b(reset_b[11:10]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g3a I_g3_30 ( .vdd_cntl(vdd_cntl[13:12]), .wl(wl[13:12]),
     .reset_b(reset_b[13:12]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .pgate(pgate[13:12]), .lc_trk_g3(lc_trk_g3[3:0]));
gmux_sp12to4_g3b I_g3_74 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g3(lc_trk_g3[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .prog(prog),
     .bl(bl[11:0]), .reset_b(reset_b[15:14]), .wl(wl[15:14]));

endmodule
// Library - sbtlibn65lp, Cell - oai22x2_hvt, View - schematic
// LAST TIME SAVED: Aug  3 19:21:57 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module oai22x2_hvt ( Y, A0, A1, B0, B1 );
output  Y;

input  A0, A1, B0, B1;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
P_11_LPHVT  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
P_11_LPHVT  M0 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
P_11_LPHVT  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));
N_11_LPHVT  M2 ( .D(Y), .B(GND_), .G(A0), .S(net024));
N_11_LPHVT  M4 ( .D(Y), .B(GND_), .G(A1), .S(net024));
N_11_LPHVT  M1 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
N_11_LPHVT  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));

endmodule
// Library - xpmem, Cell - cram_2x28, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module cram_2x28 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [55:0]  q_b;
output [55:0]  q;

inout [27:0]  bl;

input [1:0]  wl;
input [1:0]  reset;
input [1:0]  r_vdd;
input [1:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



cram2x2 I_mstake_13_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[27:26]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[1:0]));
cram2x2 I_mstake_12_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[25:24]), .q_b(q_b[51:48]),
     .q(q[51:48]), .wl(wl[1:0]));
cram2x2 I_mstake_11_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[23:22]), .q_b(q_b[47:44]),
     .q(q[47:44]), .wl(wl[1:0]));
cram2x2 I_mstake_10_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[21:20]), .q_b(q_b[43:40]),
     .q(q[43:40]), .wl(wl[1:0]));
cram2x2 I_mstake_9_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[19:18]), .q_b(q_b[39:36]),
     .q(q[39:36]), .wl(wl[1:0]));
cram2x2 I_mstake_8_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[17:16]), .q_b(q_b[35:32]),
     .q(q[35:32]), .wl(wl[1:0]));
cram2x2 I_mstake_7_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[15:14]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[1:0]));
cram2x2 I_mstake_6_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[13:12]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[1:0]));
cram2x2 I_mstake_5_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 I_mstake_4_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 I_mstake_3_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 I_mstake_2_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 I_mstake_1_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 I_mstake_0_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - odrv12_30, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module odrv12_30 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_h_r;

input  prog, slfop;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_h_r;

input [11:0]  cbitb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



odrv12 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b[1]));
odrv12 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp12(sp12_v_b[0]));
odrv12 I70 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r));
odrv4 I69_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I71_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[2]));
odrv4 I71_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[1]));
odrv4 I71_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp4(sp4_v_b[0]));
odrv4 I73_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I73_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I73_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - logic_cell_rev, View - schematic
// LAST TIME SAVED: Jul 30 21:54:54 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module logic_cell_rev ( carry_out, out, out_vic, carry_in, cbit, clk,
     clkb, in0, in1, in2, in3, prog, purst, s_r );
output  carry_out, out, out_vic;

input  carry_in, clk, clkb, in0, in1, in2, in3, prog, purst, s_r;

input [20:0]  cbit;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



clut4vic I_clut4 ( .lut4vic(out_vic), .in3b(in3b), .in3(in3),
     .in2b(in2b), .in2(in2), .in1b(in1b), .in1(in1), .in0b(in0b),
     .in0(in0), .cbit(cbit[15:0]), .lut4(LUT4_outd));
o_mux I_o_mux ( .prog(prog), .in1(rego), .in0(LUT4_outd),
     .cbit(cbit[19]), .out(out));
inv_lvt I196 ( .A(in3), .Y(in3b));
inv_lvt I189 ( .A(in0), .Y(in0b));
inv_lvt I194 ( .A(in1), .Y(in1b));
inv_lvt I195 ( .A(in2), .Y(in2b));
carry_logic_nand I_carry_logic ( .vg_en(cbit[20]), .carry_in(carry_in),
     .b_bar(in1b), .b(in1), .a_bar(in2b), .a(in2), .cout(carry_out));
coredffr I_coredffr ( .purst(purst), .d(LUT4_outd), .clkb(clkb),
     .clk(clk), .cbit(cbit[17:16]), .S_R(s_r), .q(rego));

endmodule
// Library - leafcell, Cell - lcmuxod3_0_0, View - schematic
// LAST TIME SAVED: Jul 30 21:54:54 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module lcmuxod3_0_0 ( carry_out, cbit, cbitb, op, op_vic, sp4_h_r,
     sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb,
     min0, min1, min2, min3, op_bot, pgate, prog, purst, reset_b, s_r,
     vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_h_r;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [1:0]  sp12_v_b;
output [2:0]  sp4_h_r;
output [55:0]  cbit;
output [55:0]  cbitb;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;

input [1:0]  pgate;
input [27:0]  bl;
input [1:0]  reset_b;
input [15:0]  min1;
input [1:0]  vdd_cntl;
input [15:0]  min2;
input [15:0]  min3;
input [1:0]  wl;
input [15:0]  min0;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
in_mux_nand_icc I_in2mux_nand ( .cbitb({cbitb[50], cbitb[12],
     cbitb[13], cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50],
     cbit[12], cbit[13], cbit[16], cbit[19], cbit[17]}),
     .op_bot(op_bot), .prog(prog), .inmuxo(in2), .min(min2[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_30 I_odrv30 ( .slfop(op), .prog(prog),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53], cbitb[55],
     cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44], cbitb[46],
     cbitb[43], cbitb[41], cbitb[42], cbitb[40]}), .sp12_h_r(sp12_h_r),
     .sp12_v_b(sp12_v_b[1:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));

endmodule
// Library - leafcell, Cell - lcmuxod3_0, View - schematic
// LAST TIME SAVED: Jul 30 21:54:54 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module lcmuxod3_0 ( carry_out, op, op_vic, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, op_bot, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_h_r;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min2;
input [27:0]  bl;
input [15:0]  min0;
input [15:0]  min1;
input [1:0]  reset_b;
input [15:0]  min3;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
in_mux_nand_icc I_in2mux_nand ( .cbitb({cbitb[50], cbitb[12],
     cbitb[13], cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50],
     cbit[12], cbit[13], cbit[16], cbit[19], cbit[17]}),
     .op_bot(op_bot), .prog(prog), .inmuxo(in2), .min(min2[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_30 I_odrv30 ( .slfop(op), .prog(prog),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53], cbitb[55],
     cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44], cbitb[46],
     cbitb[43], cbitb[41], cbitb[42], cbitb[40]}), .sp12_h_r(sp12_h_r),
     .sp12_v_b(sp12_v_b[1:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));

endmodule
// Library - leafcell, Cell - odrv12_74, View - schematic
// LAST TIME SAVED: Jul 30 23:15:01 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module odrv12_74 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_v_b;

input  prog, slfop;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [1:0]  sp12_h_r;
output [2:0]  sp4_h_r;

input [11:0]  cbitb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



odrv12 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp12(sp12_h_r[1]));
odrv12 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r[0]));
odrv12 I71 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b));
odrv4 I68_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I68_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I68_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I70_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp4(sp4_v_b[2]));
odrv4 I70_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[1]));
odrv4 I70_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[0]));
odrv4 I72_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - lcmuxod7_4, View - schematic
// LAST TIME SAVED: Jul 30 21:54:54 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module lcmuxod7_4 ( carry_out, op, op_vic, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, op_bot, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_v_b;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [1:0]  sp12_h_r;
output [2:0]  sp4_v_b;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;

input [15:0]  min3;
input [15:0]  min0;
input [27:0]  bl;
input [15:0]  min1;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [15:0]  min2;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [55:0]  cbitb;

wire  [55:0]  cbit;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
in_mux_nand_icc I_in2mux ( .cbitb({cbitb[50], cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50], cbit[12],
     cbit[13], cbit[16], cbit[19], cbit[17]}), .op_bot(op_bot),
     .prog(prog), .inmuxo(in2), .min(min2[15:0]));
in_mux_icc I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux_icc I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14],
     cbit[15], cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14],
     cbitb[15], cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux_icc I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5],
     cbit[4], cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4],
     cbitb[1], cbitb[2], cbitb[0]}), .min(min0[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_74 I_odrv74 ( .slfop(op), .prog(prog), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));

endmodule
// Library - leafcell, Cell - lccol_rev0, View - schematic
// LAST TIME SAVED: Jul 30 21:54:53 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module lccol_rev0 ( carry_out, op_vic, slf_op, bl, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, cin2local, clk, clkb, lc_trk_g0,
     lc_trk_g1, lc_trk_g2, lc_trk_g3, op_bot, pgate, prog, purst,
     reset_b, s_r, vdd_cntl, wl );
output  carry_out, op_vic;


input  cin2local, clk, clkb, op_bot, prog, purst, s_r;

output [7:0]  slf_op;

inout [27:0]  bl;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;

input [15:0]  reset_b;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g2;
input [7:0]  lc_trk_g3;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbitb;

wire  [55:0]  cbit;



lcmuxod3_0_0 I_LC_00 ( .cbitb(cbitb[55:0]), .cbit(cbit[55:0]),
     .op_bot(op_bot), .op_vic(net0118), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .carry_out(c_01),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], cin}),
     .reset_b(reset_b[1:0]), .vdd_cntl(vdd_cntl[1:0]), .wl(wl[1:0]),
     .op(slf_op[0]), .s_r(s_r), .sp4_h_r({sp4_h_r[32], sp4_h_r[16],
     sp4_h_r[0]}), .sp12_v_b({sp12_v_b[16], sp12_v_b[0]}),
     .sp4_r_v_b({sp4_r_v_b[33], sp4_r_v_b[17], sp4_r_v_b[1]}),
     .sp4_v_b({sp4_v_b[32], sp4_v_b[16], sp4_v_b[0]}), .carry_in(cin),
     .sp12_h_r(sp12_h_r[8]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[1:0]), .prog(prog));
lcmuxod3_0 I_LC_02 ( .op_bot(net0166), .op_vic(net094),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .carry_out(c_23), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_12}),
     .reset_b(reset_b[5:4]), .vdd_cntl(vdd_cntl[5:4]), .wl(wl[5:4]),
     .op(slf_op[2]), .s_r(s_r), .sp4_h_r({sp4_h_r[36], sp4_h_r[20],
     sp4_h_r[4]}), .sp12_v_b({sp12_v_b[20], sp12_v_b[4]}),
     .sp4_r_v_b({sp4_r_v_b[37], sp4_r_v_b[21], sp4_r_v_b[5]}),
     .sp4_v_b({sp4_v_b[36], sp4_v_b[20], sp4_v_b[4]}), .carry_in(c_12),
     .sp12_h_r(sp12_h_r[12]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[5:4]), .prog(prog));
lcmuxod3_0 I_LC_03 ( .op_bot(net094), .op_vic(net0142),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .carry_out(c_34), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_23}),
     .reset_b(reset_b[7:6]), .vdd_cntl(vdd_cntl[7:6]), .wl(wl[7:6]),
     .op(slf_op[3]), .s_r(s_r), .sp4_h_r({sp4_h_r[38], sp4_h_r[22],
     sp4_h_r[6]}), .sp12_v_b({sp12_v_b[22], sp12_v_b[6]}),
     .sp4_r_v_b({sp4_r_v_b[39], sp4_r_v_b[23], sp4_r_v_b[7]}),
     .sp4_v_b({sp4_v_b[38], sp4_v_b[22], sp4_v_b[6]}), .carry_in(c_23),
     .sp12_h_r(sp12_h_r[14]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[7:6]), .prog(prog));
lcmuxod3_0 I_LC_01 ( .op_bot(net0118), .op_vic(net0166),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .carry_out(c_12), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_01}),
     .reset_b(reset_b[3:2]), .vdd_cntl(vdd_cntl[3:2]), .wl(wl[3:2]),
     .op(slf_op[1]), .s_r(s_r), .sp4_h_r({sp4_h_r[34], sp4_h_r[18],
     sp4_h_r[2]}), .sp12_v_b({sp12_v_b[18], sp12_v_b[2]}),
     .sp4_r_v_b({sp4_r_v_b[35], sp4_r_v_b[19], sp4_r_v_b[3]}),
     .sp4_v_b({sp4_v_b[34], sp4_v_b[18], sp4_v_b[2]}), .carry_in(c_01),
     .sp12_h_r(sp12_h_r[10]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[3:2]), .prog(prog));
lcmuxod7_4 I_LC_07 ( .op_vic(op_vic), .op_bot(net0261), .bl(bl[27:0]),
     .reset_b(reset_b[15:14]), .purst(purst), .wl(wl[15:14]),
     .vdd_cntl(vdd_cntl[15:14]), .sp4_r_v_b({sp4_r_v_b[47],
     sp4_r_v_b[31], sp4_r_v_b[15]}), .sp4_h_r({sp4_h_r[46],
     sp4_h_r[30], sp4_h_r[14]}), .sp4_v_b({sp4_v_b[46], sp4_v_b[30],
     sp4_v_b[14]}), .pgate(pgate[15:14]), .sp12_h_r({sp12_h_r[22],
     sp12_h_r[6]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_67}),
     .carry_out(carry_out), .op(slf_op[7]), .s_r(s_r),
     .sp12_v_b(sp12_v_b[14]), .clk(clk), .carry_in(c_67),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clkb(clkb), .prog(prog));
lcmuxod7_4 I_LC_04 ( .op_vic(net0213), .op_bot(net0142), .prog(prog),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_34}), .clkb(clkb),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .purst(purst),
     .sp4_h_r({sp4_h_r[40], sp4_h_r[24], sp4_h_r[8]}),
     .sp4_r_v_b({sp4_r_v_b[41], sp4_r_v_b[25], sp4_r_v_b[9]}),
     .sp12_v_b(sp12_v_b[8]), .reset_b(reset_b[9:8]),
     .vdd_cntl(vdd_cntl[9:8]), .bl(bl[27:0]), .pgate(pgate[9:8]),
     .wl(wl[9:8]), .sp4_v_b({sp4_v_b[40], sp4_v_b[24], sp4_v_b[8]}),
     .sp12_h_r({sp12_h_r[16], sp12_h_r[0]}), .carry_out(c_45),
     .carry_in(c_34), .op(slf_op[4]));
lcmuxod7_4 I_LC_05 ( .op_vic(net0237), .op_bot(net0213), .prog(prog),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_45}), .clkb(clkb),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .purst(purst),
     .sp4_h_r({sp4_h_r[42], sp4_h_r[26], sp4_h_r[10]}),
     .sp4_r_v_b({sp4_r_v_b[43], sp4_r_v_b[27], sp4_r_v_b[11]}),
     .sp12_v_b(sp12_v_b[10]), .reset_b(reset_b[11:10]),
     .vdd_cntl(vdd_cntl[11:10]), .bl(bl[27:0]), .pgate(pgate[11:10]),
     .wl(wl[11:10]), .sp4_v_b({sp4_v_b[42], sp4_v_b[26], sp4_v_b[10]}),
     .sp12_h_r({sp12_h_r[18], sp12_h_r[2]}), .carry_out(c_56),
     .carry_in(c_45), .op(slf_op[5]));
lcmuxod7_4 I_LC_06 ( .op_vic(net0261), .op_bot(net0237), .prog(prog),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_56}), .clkb(clkb),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .purst(purst),
     .sp4_h_r({sp4_h_r[44], sp4_h_r[28], sp4_h_r[12]}),
     .sp4_r_v_b({sp4_r_v_b[45], sp4_r_v_b[29], sp4_r_v_b[13]}),
     .sp12_v_b(sp12_v_b[12]), .reset_b(reset_b[13:12]),
     .vdd_cntl(vdd_cntl[13:12]), .bl(bl[27:0]), .pgate(pgate[13:12]),
     .wl(wl[13:12]), .sp4_v_b({sp4_v_b[44], sp4_v_b[28], sp4_v_b[12]}),
     .sp12_h_r({sp12_h_r[20], sp12_h_r[4]}), .carry_out(c_67),
     .carry_in(c_56), .op(slf_op[6]));
mux_4carry I_carry_cnt ( .cin(cin2local), .lcl_cin(cin),
     .cbitb({cbitb[45], cbitb[48]}), .prog(prog), .cbit({cbit[45],
     cbit[48]}));

endmodule
// Library - ice1chip, Cell - ltile4_ice1f, View - schematic
// LAST TIME SAVED: Jul 30 21:53:45 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ltile4_ice1f ( carry_out, cntl_cbit, op_vic, slf_op, bl,
     sp4_h_l, sp4_h_r, sp4_r_v_b, sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r,
     sp12_v_b, sp12_v_t, bnl_op, bnr_op, bot_op, carry_in, glb_netwk,
     lft_op, op_bot, pgate, prog, purst, reset_b, rgt_op, tnl_op,
     tnr_op, top_op, vdd_cntl, wl );
output  carry_out, op_vic;


input  carry_in, op_bot, prog, purst;

output [7:0]  slf_op;
output [7:0]  cntl_cbit;

inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_t;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_t;
inout [23:0]  sp12_h_l;
inout [53:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  top_op;
input [15:0]  pgate;
input [7:0]  lft_op;
input [7:0]  bot_op;
input [7:0]  glb_netwk;
input [7:0]  tnr_op;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [7:0]  bnl_op;
input [15:0]  reset_b;
input [7:0]  bnr_op;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net187;

wire  [63:0]  cbitb_c;

wire  [63:0]  cbit_c;

wire  [3:0]  net_glb2local;

wire  [1:0]  sp12_h_r_mid;

wire  [7:0]  lc_trk_g3;

wire  [7:0]  lc_trk_g2;

wire  [1:0]  sp12_v_b_mid;

wire  [7:0]  net188;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



RM7  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
RM7  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
RM7  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
RM7  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
RM7  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
RM7  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
RM7  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
RM7  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
RM7  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
RM7  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
RM7  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
RM7  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
RM7  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
RM7  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
RM7  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
RM7  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
RM7  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
RM7  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
RM7  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
RM7  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
RM7  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
RM7  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
RM7  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
RM7  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
RM8  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
RM8  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
RM8  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
RM8  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
RM8  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
RM8  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
RM8  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
RM8  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
RM8  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
RM8  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
RM8  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
RM8  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
RM8  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
RM8  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
RM8  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
RM8  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
RM8  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
RM8  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
RM8  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
RM8  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
RM8  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
RM8  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
RM8  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
RM8  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
inv_hvt I97 ( .A(purst), .Y(purstb));
inv_hvt I98 ( .A(purstb), .Y(purstd));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(progd));
span4_ice8p I_sp4_sw ( .bram_cbit({net188[0], net188[1], net188[2],
     net188[3], net188[4], net188[5], net188[6], net188[7]}),
     .ccntrl_cbit({net187[0], net187[1], net187[2], net187[3],
     net187[4], net187[5], net187[6], net187[7]}),
     .sp4_h_l(sp4_h_l[47:0]), .bl(bl[13:4]), .wl({wl[14], wl[15],
     wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4],
     wl[5], wl[2], wl[3], wl[0], wl[1]}), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_t(sp4_v_t[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .prog(progd));
misc_module4_v3 I_misc ( .cbitb(cbitb_c[63:0]), .cbit({cbit_c[63:61],
     cntl_cbit[7], cbit_c[59:57], cntl_cbit[6], cbit_c[55:53],
     cntl_cbit[5], cbit_c[51:49], cntl_cbit[4], cbit_c[47:45],
     cntl_cbit[3], cbit_c[43:41], cntl_cbit[2], cbit_c[39:33],
     cntl_cbit[1], cbit_c[31:4], cntl_cbit[0], cbit_c[2:0]}),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .lc_trk_g1(lc_trk_g1[5:0]), .glb2local(net_glb2local[3:0]),
     .clkb(clkb), .bl(bl[3:0]), .min2(glb_netwk[7:0]),
     .min3(glb_netwk[7:0]), .min1(glb_netwk[7:0]),
     .min0(glb_netwk[7:0]), .glb_netwk(glb_netwk[7:0]),
     .lc_trk_g0(lc_trk_g0[5:0]), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .sp4(sp4_h_r[23:16]), .l(sp12_h_r_mid[1:0]),
     .S_R(s_r), .clk(clk), .b(sp12_v_b[1:0]), .r(sp12_h_r[1:0]),
     .m(sp12_v_b_mid[1:0]), .prog(progd), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18],
     sp12_h_r[16], sp12_h_r[14], sp12_h_r[12], sp12_h_r[10],
     sp12_h_r[8]}), .reset_b({reset_b[14], reset_b[15], reset_b[12],
     reset_b[13], reset_b[10], reset_b[11], reset_b[8], reset_b[9],
     reset_b[6], reset_b[7], reset_b[4], reset_b[5], reset_b[2],
     reset_b[3], reset_b[0], reset_b[1]}), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}));
gmux_sp12to4 I_gmux_sp12to4 ( .reset_b({reset_b[14], reset_b[15],
     reset_b[12], reset_b[13], reset_b[10], reset_b[11], reset_b[8],
     reset_b[9], reset_b[6], reset_b[7], reset_b[4], reset_b[5],
     reset_b[2], reset_b[3], reset_b[0], reset_b[1]}),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .lft_op(lft_op[7:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .glb2local(net_glb2local[3:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .bnr_op(bnr_op[7:0]), .lc_trk_g2(lc_trk_g2[7:0]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .bl(bl[25:14]), .lc_trk_g3(lc_trk_g3[7:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .prog(progd));
lccol_rev0 I_lccol_rev0 ( .op_bot(op_bot), .op_vic(op_vic),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .wl({wl[14], wl[15], wl[12], wl[13],
     wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2],
     wl[3], wl[0], wl[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .s_r(s_r), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .prog(progd), .purst(purstd), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .clkb(clkb), .clk(clk),
     .cin2local(carry_in), .slf_op(slf_op[7:0]), .carry_out(carry_out),
     .sp12_v_b(sp12_v_b[23:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .bl(bl[53:26]));

endmodule
// Library - ice384chip, Cell - lt_1x4_bot_ice384, View - schematic
// LAST TIME SAVED: Nov 10 17:52:15 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module lt_1x4_bot_ice384 ( carry_out, op_vic, slf_op_01, slf_op_02,
     slf_op_03, slf_op_04, bl, glb_netwk, pgate, reset_b, sp4_h_l_01,
     sp4_h_l_02, sp4_h_l_03, sp4_h_l_04, sp4_h_r_01, sp4_h_r_02,
     sp4_h_r_03, sp4_h_r_04, sp4_r_v_b_01, sp4_r_v_b_02, sp4_r_v_b_03,
     sp4_r_v_b_04, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03, sp4_v_b_04,
     sp4_v_t_04, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04,
     sp12_h_r_01, sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_v_b_01,
     sp12_v_t_04, vdd_cntl, wl, bnl_op_01, bnr_op_01, bot_op_01,
     carry_in, lc_bot, lft_op_01, lft_op_02, lft_op_03, lft_op_04,
     prog, purst, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04,
     tnl_op_04, tnr_op_04, top_op_04 );
output  carry_out, op_vic;


input  carry_in, lc_bot, prog, purst;

output [7:0]  slf_op_01;
output [7:0]  slf_op_04;
output [7:0]  slf_op_02;
output [7:0]  slf_op_03;

inout [47:0]  sp4_h_l_04;
inout [23:0]  sp12_v_b_01;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_h_r_01;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_v_b_02;
inout [23:0]  sp12_v_t_04;
inout [53:0]  bl;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_v_t_04;
inout [47:0]  sp4_r_v_b_01;
inout [23:0]  sp12_h_r_01;
inout [23:0]  sp12_h_l_02;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_r_v_b_02;
inout [63:0]  reset_b;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_h_l_03;
inout [63:0]  wl;
inout [63:0]  vdd_cntl;
inout [63:0]  pgate;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_03;
inout [7:0]  glb_netwk;

input [7:0]  lft_op_01;
input [7:0]  tnr_op_04;
input [7:0]  tnl_op_04;
input [7:0]  bnr_op_01;
input [7:0]  lft_op_02;
input [7:0]  rgt_op_04;
input [7:0]  lft_op_03;
input [7:0]  top_op_04;
input [7:0]  bot_op_01;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_04;
input [7:0]  bnl_op_01;
input [7:0]  rgt_op_02;
input [7:0]  rgt_op_01;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net1087;

wire  [7:0]  net0437;

wire  [23:0]  net1130;

wire  [23:0]  net1068;

wire  [7:0]  net1056;

wire  [23:0]  net1099;

wire  [7:0]  net1118;



ltile4_ice1f I_LT03 ( .cntl_cbit({net1056[0], net1056[1], net1056[2],
     net1056[3], net1056[4], net1056[5], net1056[6], net1056[7]}),
     .op_bot(net1089), .op_vic(net1058), .prog(prog),
     .carry_out(net1060), .lft_op(lft_op_03[7:0]),
     .sp12_h_l(sp12_h_l_03[23:0]), .sp4_h_l(sp4_h_l_03[47:0]),
     .sp4_v_b(sp4_v_b_03[47:0]), .sp12_v_b({net1099[0], net1099[1],
     net1099[2], net1099[3], net1099[4], net1099[5], net1099[6],
     net1099[7], net1099[8], net1099[9], net1099[10], net1099[11],
     net1099[12], net1099[13], net1099[14], net1099[15], net1099[16],
     net1099[17], net1099[18], net1099[19], net1099[20], net1099[21],
     net1099[22], net1099[23]}), .sp12_h_r(sp12_h_r_03[23:0]),
     .sp4_h_r(sp4_h_r_03[47:0]), .sp12_v_t({net1068[0], net1068[1],
     net1068[2], net1068[3], net1068[4], net1068[5], net1068[6],
     net1068[7], net1068[8], net1068[9], net1068[10], net1068[11],
     net1068[12], net1068[13], net1068[14], net1068[15], net1068[16],
     net1068[17], net1068[18], net1068[19], net1068[20], net1068[21],
     net1068[22], net1068[23]}), .sp4_v_t(sp4_v_b_04[47:0]),
     .sp4_r_v_b(sp4_r_v_b_03[47:0]), .wl(wl[47:32]),
     .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net1091), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4_ice1f I_LT04 ( .cntl_cbit({net0437[0], net0437[1], net0437[2],
     net0437[3], net0437[4], net0437[5], net0437[6], net0437[7]}),
     .op_bot(net1058), .op_vic(op_vic), .prog(prog),
     .carry_out(carry_out), .lft_op(lft_op_04[7:0]),
     .sp12_h_l(sp12_h_l_04[23:0]), .sp4_h_l(sp4_h_l_04[47:0]),
     .sp4_v_b(sp4_v_b_04[47:0]), .sp12_v_b({net1068[0], net1068[1],
     net1068[2], net1068[3], net1068[4], net1068[5], net1068[6],
     net1068[7], net1068[8], net1068[9], net1068[10], net1068[11],
     net1068[12], net1068[13], net1068[14], net1068[15], net1068[16],
     net1068[17], net1068[18], net1068[19], net1068[20], net1068[21],
     net1068[22], net1068[23]}), .sp12_h_r(sp12_h_r_04[23:0]),
     .sp4_h_r(sp4_h_r_04[47:0]), .sp12_v_t(sp12_v_t_04[23:0]),
     .sp4_v_t(sp4_v_t_04[47:0]), .sp4_r_v_b(sp4_r_v_b_04[47:0]),
     .wl(wl[63:48]), .top_op(top_op_04[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net1060), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(tnr_op_04[7:0]),
     .tnl_op(tnl_op_04[7:0]));
ltile4_ice1f I_LT01 ( .cntl_cbit({net1118[0], net1118[1], net1118[2],
     net1118[3], net1118[4], net1118[5], net1118[6], net1118[7]}),
     .op_bot(lc_bot), .op_vic(net1120), .prog(prog),
     .carry_out(net1122), .lft_op(lft_op_01[7:0]),
     .sp12_h_l(sp12_h_l_01[23:0]), .sp4_h_l(sp4_h_l_01[47:0]),
     .sp4_v_b(sp4_v_b_01[47:0]), .sp12_v_b(sp12_v_b_01[23:0]),
     .sp12_h_r(sp12_h_r_01[23:0]), .sp4_h_r(sp4_h_r_01[47:0]),
     .sp12_v_t({net1130[0], net1130[1], net1130[2], net1130[3],
     net1130[4], net1130[5], net1130[6], net1130[7], net1130[8],
     net1130[9], net1130[10], net1130[11], net1130[12], net1130[13],
     net1130[14], net1130[15], net1130[16], net1130[17], net1130[18],
     net1130[19], net1130[20], net1130[21], net1130[22], net1130[23]}),
     .sp4_v_t(sp4_v_b_02[47:0]), .sp4_r_v_b(sp4_r_v_b_01[47:0]),
     .wl(wl[15:0]), .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4_ice1f I_LT02 ( .cntl_cbit({net1087[0], net1087[1], net1087[2],
     net1087[3], net1087[4], net1087[5], net1087[6], net1087[7]}),
     .op_bot(net1120), .op_vic(net1089), .prog(prog),
     .carry_out(net1091), .lft_op(lft_op_02[7:0]),
     .sp12_h_l(sp12_h_l_02[23:0]), .sp4_h_l(sp4_h_l_02[47:0]),
     .sp4_v_b(sp4_v_b_02[47:0]), .sp12_v_b({net1130[0], net1130[1],
     net1130[2], net1130[3], net1130[4], net1130[5], net1130[6],
     net1130[7], net1130[8], net1130[9], net1130[10], net1130[11],
     net1130[12], net1130[13], net1130[14], net1130[15], net1130[16],
     net1130[17], net1130[18], net1130[19], net1130[20], net1130[21],
     net1130[22], net1130[23]}), .sp12_h_r(sp12_h_r_02[23:0]),
     .sp4_h_r(sp4_h_r_02[47:0]), .sp12_v_t({net1099[0], net1099[1],
     net1099[2], net1099[3], net1099[4], net1099[5], net1099[6],
     net1099[7], net1099[8], net1099[9], net1099[10], net1099[11],
     net1099[12], net1099[13], net1099[14], net1099[15], net1099[16],
     net1099[17], net1099[18], net1099[19], net1099[20], net1099[21],
     net1099[22], net1099[23]}), .sp4_v_t(sp4_v_b_03[47:0]),
     .sp4_r_v_b(sp4_r_v_b_02[47:0]), .wl(wl[31:16]),
     .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net1122), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_logic_1f, View - schematic
// LAST TIME SAVED: Aug  3 19:28:57 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_1f ( dec_trim, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, s_rd, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25, yp1_sel,
     yp2_sel, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, yp21_b_low_b, yp_test, vdd_tieh,
     fsm_blkadd, fsm_coladd, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     tm_allbank_sel, tm_tcol, ysup_25 );
output  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp21_b_low_b;

inout  vdd_tieh;

input  fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h,
     fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec,
     fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis, tm_allbank_sel,
     tm_tcol, ysup_25;

output [3:0]  s_rd;
output [7:5]  dec_trim;
output [3:0]  sbhv_high_25;
output [7:0]  yp3_sel;
output [1:0]  yp_test;
output [3:0]  sb25_high_25;
output [3:0]  sb25_gnd_25;
output [5:0]  yp1_sel;
output [3:0]  sbhv_gnd_25;
output [7:0]  yp2_sel;

input [2:0]  fsm_trim_rrefpgm;
input [2:0]  fsm_trim_rrefrd;
input [9:0]  fsm_coladd;
input [1:0]  fsm_rowadd;
input [3:0]  fsm_blkadd;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net561;

wire  [5:0]  yp1_sel_b;

wire  [3:0]  sb25low_b;

wire  [7:0]  yp2_sel_b;

wire  [7:0]  yp3_sel_b;

wire  [3:0]  sbhvlow_b;

wire  [9:0]  yadd_b;

wire  [7:5]  dec_trim_b;

wire  [3:0]  s_rd_b;

wire  [1:0]  yp_test_b;

wire  [2:0]  tdec_b;

wire  [2:0]  tdec;

wire  [1:0]  xadd_b;

wire  [1:0]  xadd;

wire  [9:0]  yadd;



inv_25 I104 ( .IN(net302), .OUT(en_blinhi_pgm_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I285 ( .IN(net311), .OUT(yp3_b_low_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I284 ( .IN(net306), .OUT(yp3_b_high_odd_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I283 ( .IN(net316), .OUT(yp3_b_high_even_b_ysup_25),
     .P(ysup_25), .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
ml_core_ctrl_logic_8f_sbb Isb25_3_ ( .in(sb25low_b[3]),
     .out_hv_woinv(sb25_gnd_25[3]), .out_hv_winv(sb25_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isb25_2_ ( .in(sb25low_b[2]),
     .out_hv_woinv(sb25_gnd_25[2]), .out_hv_winv(sb25_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isb25_1_ ( .in(sb25low_b[1]),
     .out_hv_woinv(sb25_gnd_25[1]), .out_hv_winv(sb25_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isb25_0_ ( .in(sb25low_b[0]),
     .out_hv_woinv(sb25_gnd_25[0]), .out_hv_winv(sb25_high_25[0]));
ml_core_ctrl_logic_8f_sbb Isbhv_3_ ( .in(sbhvlow_b[3]),
     .out_hv_woinv(sbhv_gnd_25[3]), .out_hv_winv(sbhv_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isbhv_2_ ( .in(sbhvlow_b[2]),
     .out_hv_woinv(sbhv_gnd_25[2]), .out_hv_winv(sbhv_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isbhv_1_ ( .in(sbhvlow_b[1]),
     .out_hv_woinv(sbhv_gnd_25[1]), .out_hv_winv(sbhv_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isbhv_0_ ( .in(sbhvlow_b[0]),
     .out_hv_woinv(sbhv_gnd_25[0]), .out_hv_winv(sbhv_high_25[0]));
ml_ls_vdd25_nor2 I106 ( .in(net343), .sup(ysup_25),
     .out_vddio_b(net301), .out_vddio(net302), .in_b(en_blinhi_pgm_b));
ml_ls_vdd25_nor2 I68 ( .in(net576), .sup(ysup_25),
     .out_vddio_b(net306), .out_vddio(net307), .in_b(net308));
ml_ls_vdd25_nor2 I192 ( .in(net396), .sup(ysup_25),
     .out_vddio_b(net311), .out_vddio(net312), .in_b(net544));
ml_ls_vdd25_nor2 I65 ( .in(net571), .sup(ysup_25),
     .out_vddio_b(net316), .out_vddio(net317), .in_b(net318));
exor2_hvt I151_3_ ( .A(net561[0]), .Y(sb25low_b[3]), .B(pgm_hvact_b));
exor2_hvt I151_2_ ( .A(net561[1]), .Y(sb25low_b[2]), .B(pgm_hvact_b));
exor2_hvt I151_1_ ( .A(net561[2]), .Y(sb25low_b[1]), .B(pgm_hvact_b));
exor2_hvt I151_0_ ( .A(net561[3]), .Y(sb25low_b[0]), .B(pgm_hvact_b));
mux2_hvt I152 ( .in1(net504), .in0(net514), .out(ensb25_dec),
     .sel(pgm_hvact));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(tdec[2]), .sel(ref_pgm));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(tdec[1]), .sel(ref_pgm));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(tdec[0]), .sel(ref_pgm));
oai21x2_hvt I55 ( .A1(sa_bl_to_blsa), .Y(net331), .A0(blk_dec),
     .B0(ymux_dis_b));
nor3_hvt I324 ( .B(fsm_tm_testdec), .Y(net335), .A(fsm_tm_allbl_l),
     .C(fsm_tm_allbl_h));
nor3_hvt I321 ( .B(fsm_tm_allbl_h), .Y(net339), .A(nvcmen_buf_b),
     .C(yp3_b_high_b));
nor4_hvt I326 ( .B(fsm_tm_allbl_l), .Y(net343), .D(nvcmen_buf_b),
     .A(net384), .C(fsm_tm_allbl_l));
nor4_hvt I327 ( .B(fsm_tm_allbl_h), .Y(ymux_dis_b), .D(net405),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_h));
nand3_hvt I227 ( .Y(net352), .B(pgm_hvact), .C(fsm_tm_allwl_h),
     .A(fsm_lshven));
nand3_hvt I236_3_ ( .Y(s_rd_b[3]), .B(xadd[0]), .C(en_rdp),
     .A(xadd[1]));
nand3_hvt I236_2_ ( .Y(s_rd_b[2]), .B(xadd_b[0]), .C(en_rdp),
     .A(xadd[1]));
nand3_hvt I236_1_ ( .Y(s_rd_b[1]), .B(xadd[0]), .C(en_rdp),
     .A(xadd_b[1]));
nand3_hvt I236_0_ ( .Y(s_rd_b[0]), .B(xadd_b[0]), .C(en_rdp),
     .A(xadd_b[1]));
nand3_hvt I230 ( .Y(pgm_hvact_b), .B(fsm_pgm), .C(net502),
     .A(fsm_lshven));
nand3_hvt I232 ( .Y(net364), .B(sa_bl_to_blsa), .C(tm_allwl_l_b),
     .A(fsm_vpxaset));
nand3_hvt I233 ( .Y(net368), .B(net492), .C(nvcmen_buf), .A(net387));
nand3_hvt I234_7_ ( .Y(dec_trim_b[7]), .B(tdec[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I234_6_ ( .Y(dec_trim_b[6]), .B(tdec[1]), .C(tdec_b[0]),
     .A(tdec[2]));
nand3_hvt I234_5_ ( .Y(dec_trim_b[5]), .B(tdec_b[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I231_7_ ( .Y(yp2_sel_b[7]), .B(yadd[4]), .C(yadd[3]),
     .A(yadd[5]));
nand3_hvt I231_6_ ( .Y(yp2_sel_b[6]), .B(yadd[4]), .C(yadd_b[3]),
     .A(yadd[5]));
nand3_hvt I231_5_ ( .Y(yp2_sel_b[5]), .B(yadd_b[4]), .C(yadd[3]),
     .A(yadd[5]));
nand3_hvt I231_4_ ( .Y(yp2_sel_b[4]), .B(yadd_b[4]), .C(yadd_b[3]),
     .A(yadd[5]));
nand3_hvt I231_3_ ( .Y(yp2_sel_b[3]), .B(yadd[4]), .C(yadd[3]),
     .A(yadd_b[5]));
nand3_hvt I231_2_ ( .Y(yp2_sel_b[2]), .B(yadd[4]), .C(yadd_b[3]),
     .A(yadd_b[5]));
nand3_hvt I231_1_ ( .Y(yp2_sel_b[1]), .B(yadd_b[4]), .C(yadd[3]),
     .A(yadd_b[5]));
nand3_hvt I231_0_ ( .Y(yp2_sel_b[0]), .B(yadd_b[4]), .C(yadd_b[3]),
     .A(yadd_b[5]));
nand2_hvt I299 ( .A(fsm_tm_rd_mode), .Y(one_blk_sel_b), .B(blk_dec));
nand2_hvt I301 ( .A(pgm_hvact), .Y(net384), .B(pgm_hvact));
nand2_hvt I293 ( .A(fsm_lshven), .Y(net387), .B(pgm_hvact));
nand2_hvt I297 ( .A(blk_dec_b), .Y(blk_dec), .B(tm_pgm_rd_allblk_n));
nand2_hvt I296 ( .A(blk_dec), .Y(net393), .B(fsm_pgmien));
nand2_hvt I294 ( .A(net387), .Y(net396), .B(net335));
nand2_hvt I298 ( .A(all_blk_sel_b), .Y(sa_bl_to_blsa),
     .B(one_blk_sel_b));
nand2_hvt I300 ( .A(tm_allwl_l_b), .Y(net503), .B(blk_dec));
nand2_hvt I295 ( .A(fsm_nvcmen), .Y(net405), .B(fsm_lshven));
nand2_hvt I291_1_ ( .A(yadd[0]), .Y(yp_test_b[1]), .B(ymux_test_en));
nand2_hvt I291_0_ ( .A(yadd_b[0]), .Y(yp_test_b[0]), .B(ymux_test_en));
nand2_hvt I245 ( .A(rd_and_vfy), .Y(all_blk_sel_b), .B(net536));
nand4_hvt I306 ( .D(fsm_blkadd[0]), .A(fsm_blkadd[3]),
     .C(fsm_blkadd[1]), .Y(blk_dec_b), .B(fsm_blkadd[2]));
nand4_hvt I307_5_ ( .D(yadd[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[5]), .B(yadd[8]));
nand4_hvt I307_4_ ( .D(yadd_b[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[4]), .B(yadd[8]));
nand4_hvt I304_7_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[7]), .B(yadd[2]));
nand4_hvt I304_6_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[6]), .B(yadd[2]));
nand4_hvt I304_5_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[5]), .B(yadd[2]));
nand4_hvt I304_4_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[4]), .B(yadd[2]));
nand4_hvt I304_3_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[3]), .B(yadd_b[2]));
nand4_hvt I304_2_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[2]), .B(yadd_b[2]));
nand4_hvt I304_1_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[1]), .B(yadd_b[2]));
nand4_hvt I304_0_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[0]), .B(yadd_b[2]));
nand4_hvt I239 ( .D(fsm_tm_rprd), .Y(net429), .B(fsm_lshven),
     .C(nvcmen_buf), .A(rd_and_vfy));
nand4_hvt I308 ( .D(fsm_lshven), .A(tm_allwl_l_b), .C(pgm_hvact),
     .Y(net436), .B(blk_dec));
nor2_hvt I316_5_ ( .A(yp1_sel_b[5]), .B(tm_tcol), .Y(yp1_sel[5]));
nor2_hvt I316_4_ ( .A(yp1_sel_b[4]), .B(tm_tcol), .Y(yp1_sel[4]));
nor2_hvt I310 ( .A(fsm_pgmvfy), .B(fsm_pgm), .Y(net443));
nor2_hvt I315 ( .A(net331), .B(net530), .Y(ymux_test_en));
nor2_hvt I312 ( .A(net579), .B(net532), .Y(net449));
nor2_hvt I319 ( .A(fsm_rd), .B(fsm_pgmvfy), .Y(net452));
nor2_hvt I328 ( .A(net331), .B(tm_tcol), .Y(ymux_en_core));
nor2_hvt I317_3_ ( .A(yp1_sel_b[3]), .B(tm_tcol), .Y(yp1_sel[3]));
nor2_hvt I317_2_ ( .A(yp1_sel_b[2]), .B(tm_tcol), .Y(yp1_sel[2]));
nor2_hvt I317_1_ ( .A(yp1_sel_b[1]), .B(tm_tcol), .Y(yp1_sel[1]));
nor2_hvt I317_0_ ( .A(yp1_sel_b[0]), .B(tm_tcol), .Y(yp1_sel[0]));
nor2_hvt I313 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I318 ( .A(fsm_tm_rd_mode), .B(fsm_pgmvfy), .Y(net464));
anor21_hvt I119_1_ ( .A(fsm_rowadd[1]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I119_0_ ( .A(fsm_rowadd[0]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
anor21_hvt I109 ( .A(pgm_hvact), .B(fsm_tm_allwl_h), .Y(net505),
     .C(nvcmen_buf_b));
inv_hvt I271_9_ ( .A(yadd[9]), .Y(yadd_b[9]));
inv_hvt I272_9_ ( .A(vdd_tieh), .Y(yadd[9]));
inv_hvt I247 ( .A(net452), .Y(rd_and_vfy));
inv_hvt I265 ( .A(net464), .Y(net484));
inv_hvt I323 ( .A(fsm_tm_allbl_l), .Y(yp3_b_high_b));
inv_hvt I237_3_ ( .A(s_rd_b[3]), .Y(s_rd[3]));
inv_hvt I237_2_ ( .A(s_rd_b[2]), .Y(s_rd[2]));
inv_hvt I237_1_ ( .A(s_rd_b[1]), .Y(s_rd[1]));
inv_hvt I237_0_ ( .A(s_rd_b[0]), .Y(s_rd[0]));
inv_hvt I252_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I252_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I200 ( .A(fsm_tm_testdec), .Y(net492));
inv_hvt I261 ( .A(net393), .Y(sa_bl_to_pgm_glb));
inv_hvt I271_8_ ( .A(yadd_b[8]), .Y(yadd[8]));
inv_hvt I271_7_ ( .A(yadd_b[7]), .Y(yadd[7]));
inv_hvt I271_6_ ( .A(yadd_b[6]), .Y(yadd[6]));
inv_hvt I271_5_ ( .A(yadd_b[5]), .Y(yadd[5]));
inv_hvt I271_4_ ( .A(yadd_b[4]), .Y(yadd[4]));
inv_hvt I271_3_ ( .A(yadd_b[3]), .Y(yadd[3]));
inv_hvt I271_2_ ( .A(yadd_b[2]), .Y(yadd[2]));
inv_hvt I271_1_ ( .A(yadd_b[1]), .Y(yadd[1]));
inv_hvt I271_0_ ( .A(yadd_b[0]), .Y(yadd[0]));
inv_hvt I268 ( .A(net579), .Y(vddp_rd_overw));
inv_hvt I260 ( .A(nvcmen_buf_b), .Y(nvcmen_buf));
inv_hvt I254 ( .A(net576), .Y(net308));
inv_hvt I278 ( .A(fsm_pgmvfy), .Y(net502));
inv_hvt I281 ( .A(net503), .Y(net504));
inv_hvt I279 ( .A(net505), .Y(net506));
inv_hvt I251 ( .A(net352), .Y(net508));
inv_hvt I258 ( .A(net368), .Y(yp21_b_low_b));
inv_hvt I263 ( .A(fsm_nvcmen), .Y(nvcmen_buf_b));
inv_hvt I280 ( .A(net364), .Y(net514));
inv_hvt I264 ( .A(tm_allbank_sel), .Y(tm_pgm_rd_allblk_n));
inv_hvt I250 ( .A(net436), .Y(net518));
inv_hvt I241 ( .A(net429), .Y(en_rdp));
inv_hvt I255 ( .A(net343), .Y(en_blinhi_pgm_b));
inv_hvt I249 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I277 ( .A(pgm_hvact_b), .Y(pgm_hvact));
inv_hvt I266 ( .A(net443), .Y(ref_pgm));
inv_hvt I259 ( .A(tm_tcol), .Y(net530));
inv_hvt I267 ( .A(fsm_multibl_read), .Y(net532));
inv_hvt I262 ( .A(all_blk_sel_b), .Y(net534));
inv_hvt I272_8_ ( .A(fsm_coladd[8]), .Y(yadd_b[8]));
inv_hvt I272_7_ ( .A(fsm_coladd[7]), .Y(yadd_b[7]));
inv_hvt I272_6_ ( .A(fsm_coladd[6]), .Y(yadd_b[6]));
inv_hvt I272_5_ ( .A(fsm_coladd[5]), .Y(yadd_b[5]));
inv_hvt I272_4_ ( .A(fsm_coladd[4]), .Y(yadd_b[4]));
inv_hvt I272_3_ ( .A(fsm_coladd[3]), .Y(yadd_b[3]));
inv_hvt I272_2_ ( .A(fsm_coladd[2]), .Y(yadd_b[2]));
inv_hvt I272_1_ ( .A(fsm_coladd[1]), .Y(yadd_b[1]));
inv_hvt I272_0_ ( .A(fsm_coladd[0]), .Y(yadd_b[0]));
inv_hvt I201 ( .A(fsm_tm_rd_mode), .Y(net536));
inv_hvt I270_2_ ( .A(tdec[2]), .Y(tdec_b[2]));
inv_hvt I270_1_ ( .A(tdec[1]), .Y(tdec_b[1]));
inv_hvt I270_0_ ( .A(tdec[0]), .Y(tdec_b[0]));
inv_hvt I273_7_ ( .A(yp2_sel_b[7]), .Y(yp2_sel[7]));
inv_hvt I273_6_ ( .A(yp2_sel_b[6]), .Y(yp2_sel[6]));
inv_hvt I273_5_ ( .A(yp2_sel_b[5]), .Y(yp2_sel[5]));
inv_hvt I273_4_ ( .A(yp2_sel_b[4]), .Y(yp2_sel[4]));
inv_hvt I273_3_ ( .A(yp2_sel_b[3]), .Y(yp2_sel[3]));
inv_hvt I273_2_ ( .A(yp2_sel_b[2]), .Y(yp2_sel[2]));
inv_hvt I273_1_ ( .A(yp2_sel_b[1]), .Y(yp2_sel[1]));
inv_hvt I273_0_ ( .A(yp2_sel_b[0]), .Y(yp2_sel[0]));
inv_hvt I256_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I256_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I256_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I257 ( .A(net396), .Y(net544));
inv_hvt I274_7_ ( .A(yp3_sel_b[7]), .Y(yp3_sel[7]));
inv_hvt I274_6_ ( .A(yp3_sel_b[6]), .Y(yp3_sel[6]));
inv_hvt I274_5_ ( .A(yp3_sel_b[5]), .Y(yp3_sel[5]));
inv_hvt I274_4_ ( .A(yp3_sel_b[4]), .Y(yp3_sel[4]));
inv_hvt I274_3_ ( .A(yp3_sel_b[3]), .Y(yp3_sel[3]));
inv_hvt I274_2_ ( .A(yp3_sel_b[2]), .Y(yp3_sel[2]));
inv_hvt I274_1_ ( .A(yp3_sel_b[1]), .Y(yp3_sel[1]));
inv_hvt I274_0_ ( .A(yp3_sel_b[0]), .Y(yp3_sel[0]));
inv_hvt I253 ( .A(net571), .Y(net318));
inv_hvt I275_1_ ( .A(yp_test_b[1]), .Y(yp_test[1]));
inv_hvt I275_0_ ( .A(yp_test_b[0]), .Y(yp_test[0]));
oai2211x2_hvt I86_3_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[3]), .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai2211x2_hvt I86_2_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[2]), .A0(yadd[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
oai2211x2_hvt I86_1_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[1]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd[6]));
oai2211x2_hvt I86_0_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[0]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
anor31_hvt I155_3_ ( .A(ensb25_dec), .D(net506), .B(xadd[1]),
     .Y(net561[0]), .C(xadd[0]));
anor31_hvt I155_2_ ( .A(ensb25_dec), .D(net506), .B(xadd[1]),
     .Y(net561[1]), .C(xadd_b[0]));
anor31_hvt I155_1_ ( .A(ensb25_dec), .D(net506), .B(xadd_b[1]),
     .Y(net561[2]), .C(xadd[0]));
anor31_hvt I155_0_ ( .A(ensb25_dec), .D(net506), .B(xadd_b[1]),
     .Y(net561[3]), .C(xadd_b[0]));
anor31_hvt I121_3_ ( .A(net518), .D(net508), .B(xadd[1]),
     .Y(sbhvlow_b[3]), .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net518), .D(net508), .B(xadd[1]),
     .Y(sbhvlow_b[2]), .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net518), .D(net508), .B(xadd_b[1]),
     .Y(sbhvlow_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net518), .D(net508), .B(xadd_b[1]),
     .Y(sbhvlow_b[0]), .C(xadd_b[0]));
anor31_hvt I107 ( .A(fsm_tm_testdec), .D(net339), .B(nvcmen_buf),
     .Y(net571), .C(yadd[0]));
anor31_hvt I108 ( .A(fsm_tm_testdec), .D(net339), .B(nvcmen_buf),
     .Y(net576), .C(yadd_b[0]));
oai22x2_hvt I93 ( .A1(net534), .Y(net579), .A0(net484),
     .B0(fsm_nv_rri_trim), .B1(fsm_nv_sisi_ui));

endmodule
// Library - ice8chip, Cell - tckbufx32_ice8p, View - schematic
// LAST TIME SAVED: Aug 13 15:04:42 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module tckbufx32_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_lvt I_inv_lvt_1 ( .A(in), .Y(net4));
inv_lvt Iinv_lvt_2 ( .A(net4), .Y(out));

endmodule
// Library - ice8chip, Cell - fabric_buf_ice8p, View - schematic
// LAST TIME SAVED: Aug 13 15:11:11 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module fabric_buf_ice8p ( f_out, f_in );
output  f_out;

input  f_in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_lvt I_inv_lvt_2 ( .A(net6), .Y(f_out));
inv_lvt I_inv_lvt_1 ( .A(f_in), .Y(net6));

endmodule
// Library - io, Cell - ioin_mux_v3, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioin_mux_v3 ( inmuxo, cbit,
     cbitb, min[7:0], prog );
output  inmuxo;

input  prog;

input [3:0]  cbitb;
input [3:0]  cbit;
input [7:0]  min;
supply1 vdd_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

nor2_lvt I282 ( .A(prog), .Y(en), .B(cbitb[3]));
inv_lvt I281 ( .A(inmuxob), .Y(inmuxo));
nand2_lvt I_nand2 ( .A(st2), .Y(inmuxob), .B(en));
txgate_lvt I285 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I289 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I286 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I283 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_lvt I292 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I293 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I291 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I294 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I287 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I290 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I288 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I295 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I284 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc_v0, View - schematic
// LAST TIME SAVED: Aug  3 19:20:28 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc_v0 ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  spi;
output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  padin;
input [7:0]  min1;
input [1:0]  wl;
input [1:0]  pgate;
input [7:0]  min0;
input [1:0]  reset;
input [7:0]  min2;
input [1:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ioin_mux_v3 I_ioin_mux_bankcntl ( bankcntl, {cbit[11], cbit[8], cbit[9],
     cbit[10]}, {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0],
     prog);
ioin_mux_v3 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v3 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
inv_lvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_lvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
nor2_lvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_lvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nand2inv_v0, View - schematic
// LAST TIME SAVED: Aug  3 19:20:28 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioinmx2nand2inv_v0 ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [7:0]  min0;
input [1:0]  wl;
input [1:0]  pgate;
input [7:0]  min1;
input [1:0]  reset;
input [7:0]  ce;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ioin_mux_v3 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v3 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
nand2_lvt I180 ( .A(update_b), .Y(updt), .B(bs_en));
inv_lvt I181 ( .A(update), .Y(update_b));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioin_mux_v2, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioin_mux_v2 ( inmuxo, cbit,
     cbitb, min[7:0], prog );
output  inmuxo;

input  prog;

input [3:0]  cbit;
input [7:0]  min;
input [3:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

nor2_lvt I_nor2_lvt ( .A(prog), .Y(en), .B(cbitb[3]));
inv_lvt I281 ( .A(inmuxob), .Y(inmuxo));
nand2_lvt I_nand2 ( .A(st2), .Y(inmuxob), .B(en));
txgate_lvt I285 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I289 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I286 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I283 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_lvt I292 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I293 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I291 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I294 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I287 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I290 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I288 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I295 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I284 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));

endmodule
// Library - io, Cell - ioinmx1mux2_v1, View - schematic
// LAST TIME SAVED: Aug  3 19:20:28 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioinmx1mux2_v1 ( clk, ti, bl, ce, ceb, min, pgate, prog, reset,
     vdd_cntl, wl );
output  clk, ti;


input  ceb, prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [11:0]  ce;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
input [7:0]  min;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clk_mux12to1_icc I_clk_mux12to1 ( .prog(prog), .min(ce[11:0]),
     .clk(clk), .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7],
     cbitb[10], cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7],
     cbit[10], cbit[6], cbit[4]}), .cenb(ceb));
ioin_mux_v2 I_ioin_mux ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1mem, View - schematic
// LAST TIME SAVED: Aug  3 19:20:31 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module sbox1mem ( b, bl, l, r, t, pgate, prog, reset, vdd_cntl, wl );
inout  b, l, r, t;

input  prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  reset;
input [1:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbitb;

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox1m3to1_icc I232 ( .in2(r), .cb({cbitb[3], cbitb[6]}), .op(t),
     .in0(l), .in1(b), .c({cbit[3], cbit[6]}), .prog(prog));
sbox1m3to1_icc I230 ( .in2(r), .cb({cbitb[1], cbitb[4]}), .op(l),
     .in0(b), .in1(t), .c({cbit[1], cbit[4]}), .prog(prog));
sbox1m3to1_icc I226 ( .in2(r), .cb({cbitb[8], cbitb[5]}), .op(b),
     .in0(l), .in1(t), .c({cbit[8], cbit[5]}), .prog(prog));
sbox1m3to1_icc I231 ( .in2(b), .cb({cbitb[10], cbitb[7]}), .op(r),
     .in0(l), .in1(t), .c({cbit[10], cbit[7]}), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc_v4, View - schematic
// LAST TIME SAVED: Dec  7 10:50:25 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module sbox1_colbdlc_v4 ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [5:0]  ti;

inout [5:0]  bl;
inout [3:0]  r;
inout [3:0]  l;
inout [3:0]  sp4_v_b;
inout [3:0]  t_mid;

input [1:0]  oeb;
input [7:0]  min1;
input [1:0]  padin;
input [7:0]  min3;
input [7:0]  min4;
input [7:0]  min6;
input [11:0]  clk_in;
input [1:0]  out;
input [7:0]  min0;
input [11:0]  inclk_in;
input [1:0]  spioeb;
input [1:0]  spiout;
input [7:0]  ceb_in;
input [15:0]  reset;
input [7:0]  min2;
input [15:0]  vdd_cntl;
input [7:0]  min5;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spioob;

wire  [1:0]  spioo;

wire  [1:0]  oeboo;

wire  [1:0]  oeboob;



ioinmx2nor2invx2bdlc_v0 I5 ( .vdd_cntl(vdd_cntl[5:4]),
     .min2(min6[7:0]), .bankcntl(fabric_out), .bl(bl[5:0]),
     .prog(prog), .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx2nand2inv_v0 I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
ioinmx1mux2_v1 I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .ti(ti[2]), .min(min2[7:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]));
ioinmx1mux2_v1 I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .ti(ti[5]), .min(min5[7:0]), .wl(wl[15:14]), .reset(reset[15:14]),
     .pgate(pgate[15:14]));
inv_lvt I_inv_2_1_ ( .A(spioob[1]), .Y(pado[1]));
inv_lvt I_inv_2_0_ ( .A(spioob[0]), .Y(pado[0]));
inv_lvt I9_1_ ( .A(oeboo[1]), .Y(oeboob[1]));
inv_lvt I9_0_ ( .A(oeboo[0]), .Y(oeboob[0]));
inv_lvt I8_1_ ( .A(oeboob[1]), .Y(padeb[1]));
inv_lvt I8_0_ ( .A(oeboob[0]), .Y(padeb[0]));
inv_lvt inv_1_1_ ( .A(spioo[1]), .Y(spioob[1]));
inv_lvt inv_1_0_ ( .A(spioo[0]), .Y(spioob[0]));
mux2x1_hvt I10_1_ ( .in1(oeb[1]), .in0(spioeb[1]), .out(oeboo[1]),
     .sel(cdone_in));
mux2x1_hvt I10_0_ ( .in1(oeb[0]), .in0(spioeb[0]), .out(oeboo[0]),
     .sel(cdone_in));
mux2x1_hvt I_emux_1_ ( .in1(out[1]), .in0(spiout[1]), .out(spioo[1]),
     .sel(cdone_in));
mux2x1_hvt I_emux_0_ ( .in1(out[0]), .in0(spiout[0]), .out(spioo[0]),
     .sel(cdone_in));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - io, Cell - io_gmux_x2v3, View - schematic
// LAST TIME SAVED: Aug  3 19:20:26 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_gmux_x2v3 ( .cbit_colcntl({cbit[11], cbit[9]}), gout, bl,
     min0, min1, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [1:0]  gout;
output [11:0]  cbit;

inout [5:0]  bl;

input [15:0]  min0;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [15:0]  min1;
input [1:0]  wl;
input [1:0]  reset;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux I_g_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux I_g_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - umc40lp, Cell - RNPPO_LP, View - schematic
// LAST TIME SAVED: Jan 18 18:48:10 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module RNPPO_LP_pcell2460 ( MINUS, PLUS, B );
inout  MINUS, PLUS;

input  B;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



primRes3  R0 ( .MINUS(MINUS), .PLUS(PLUS), .B(B));

endmodule
// Library - io, Cell - io_gmux_x16bare_v4, View - schematic
// LAST TIME SAVED: Aug 25 13:36:24 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_gmux_x16bare_v4 ( cbit_colcntl, lc_trk_g0, lc_trk_g1, bl,
     min0, min1, min2, min3, min4, min5, min6, min7, min8, min9, min10,
     min11, min12, min13, min14, min15, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [7:0]  cbit_colcntl;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g1;

inout [5:0]  bl;

input [15:0]  min9;
input [15:0]  min12;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min0;
input [15:0]  min7;
input [15:0]  min5;
input [15:0]  min3;
input [15:0]  min4;
input [15:0]  min10;
input [15:0]  min6;
input [15:0]  min8;
input [15:0]  min15;
input [15:0]  min14;
input [15:0]  min11;
input [15:0]  reset;
input [15:0]  min2;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net187;

wire  [1:0]  net114;

wire  [1:0]  net124;

wire  [1:0]  net188;



io_gmux_x2v3 I_io_gmux_x2_7 ( .cbit_colcntl({net114[0], net114[1]}),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[15:14]));
io_gmux_x2v3 I_io_gmux_x2_6 ( .cbit_colcntl({net124[0], net124[1]}),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[13:12]));
io_gmux_x2v3 I_io_gmux_x2_2 ( .cbit_colcntl(cbit_colcntl[5:4]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[5:4]));
io_gmux_x2v3 I_io_gmux_x2_0 ( .cbit_colcntl(cbit_colcntl[1:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[1:0]));
io_gmux_x2v3 _io_gmux_x2_1 ( .cbit_colcntl(cbit_colcntl[3:2]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[3:2]));
io_gmux_x2v3 I_io_gmux_x2_4 ( .cbit_colcntl({net187[0], net187[1]}),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[9:8]));
io_gmux_x2v3 I_io_gmux_x2_5 ( .cbit_colcntl({net188[0], net188[1]}),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[11:10]));
io_gmux_x2v3 I_io_gmux_x2_3 ( .cbit_colcntl(cbit_colcntl[7:6]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[7:6]));

endmodule
// Library - io, Cell - io_odrv4x5, View - schematic
// LAST TIME SAVED: Aug  3 19:20:26 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_odrv4x5 ( cbit, sp4_out, bl, pgate, prog,
     reset, slfop, vdd_cntl, wl );


input  prog, slfop;

output [4:0]  sp4_out;
output [7:5]  cbit;

inout [3:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  cbitb;

wire  [1:0]  r_vdd;

wire [7:0] cbit_int;
assign cbit[7:5] = cbit_int[7:5];

pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv4 I_odrv_4_ ( .cbitb(cbitb[4]), .sp4(sp4_out[4]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_3_ ( .cbitb(cbitb[3]), .sp4(sp4_out[3]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_2_ ( .cbitb(cbitb[2]), .sp4(sp4_out[2]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_1_ ( .cbitb(cbitb[1]), .sp4(sp4_out[1]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_0_ ( .cbitb(cbitb[0]), .sp4(sp4_out[0]), .slfop(slfop),
     .prog(prog));
cram2x2 Icram2x2_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset[1:0]), .q(cbit_int[7:4]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));
cram2x2 Icram2x2_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset[1:0]), .q(cbit_int[3:0]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - io_col_odrv4_x40bare_v3, View - schematic
// LAST TIME SAVED: Jun  2 10:03:19 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_col_odrv4_x40bare_v3 ( cf, bl, sp4_h_l,
     sp4_v_b, dout0, dout1,
     pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [23:0]  cf;

inout [3:0]  bl;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_b;

input [0:1]  dout1;
input [0:1]  dout0;
input [15:0]  wl;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

io_odrv4x5 I_io_odrv4x5_6 ( cf[20:18], {sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6]}, bl[3:0], pgate[13:12],
     prog, reset[13:12], dout1[1], vdd_cntl[13:12], wl[13:12]);
io_odrv4x5 I_io_odrv4x5_4 ( cf[14:12], {sp4_h_l[36], sp4_h_l[28],
     sp4_h_l[20], sp4_h_l[12], sp4_h_l[4]}, bl[3:0], pgate[9:8], prog,
     reset[9:8], dout0[1], vdd_cntl[9:8], wl[9:8]);
io_odrv4x5 I_io_odrv4x5_7 ( cf[23:21], {sp4_v_b[15], sp4_v_b[11],
     sp4_v_b[7], sp4_v_b[3], sp4_h_l[46]}, bl[3:0], pgate[15:14], prog,
     reset[15:14], dout1[1], vdd_cntl[15:14], wl[15:14]);
io_odrv4x5 I_io_odrv4x5_3 ( cf[11:9], {sp4_v_b[13], sp4_v_b[9],
     sp4_v_b[5], sp4_v_b[1], sp4_h_l[42]}, bl[3:0], pgate[7:6], prog,
     reset[7:6], dout1[0], vdd_cntl[7:6], wl[7:6]);
io_odrv4x5 I_io_odrv4x5_2 ( cf[8:6], {sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2]}, bl[3:0], pgate[5:4], prog,
     reset[5:4], dout1[0], vdd_cntl[5:4], wl[5:4]);
io_odrv4x5 I_io_odrv4x5_0 ( cf[2:0], {sp4_h_l[32], sp4_h_l[24],
     sp4_h_l[16], sp4_h_l[8], sp4_h_l[0]}, bl[3:0], pgate[1:0], prog,
     reset[1:0], dout0[0], vdd_cntl[1:0], wl[1:0]);
io_odrv4x5 I_io_odrv4x5_1 ( cf[5:3], {sp4_v_b[12], sp4_v_b[8],
     sp4_v_b[4], sp4_v_b[0], sp4_h_l[40]}, bl[3:0], pgate[3:2], prog,
     reset[3:2], dout0[0], vdd_cntl[3:2], wl[3:2]);
io_odrv4x5 I_io_odrv4x5_5 ( cf[17:15], {sp4_v_b[14], sp4_v_b[10],
     sp4_v_b[6], sp4_v_b[2], sp4_h_l[44]}, bl[3:0], pgate[11:10], prog,
     reset[11:10], dout0[1], vdd_cntl[11:10], wl[11:10]);

endmodule
// Library - io, Cell - insel1_lvt_imp, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module insel1_lvt_imp ( out, in0, in1, in2, in3, sb, sel );
output  out;

input  in0, in1, in2, in3;

input [1:0]  sel;
input [1:0]  sb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I39 ( .in(in3), .out(outd23), .pp(sb[0]), .nn(sel[0]));
txgate_lvt I40 ( .in(in2), .out(outd23), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I33 ( .in(outd01), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_lvt I_txgate1 ( .in(in1), .out(outd01), .pp(sb[0]),
     .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(outd01), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(outd23), .out(out), .pp(sb[1]), .nn(sel[1]));

endmodule
// Library - io, Cell - cebdffrqn, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module cebdffrqn ( q, qn, ceb, clk, d, r );
output  q, qn;

input  ceb, clk, d, r;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_lvt I43 ( .A(so), .Y(low_s));
inv_lvt I50 ( .A(clkb), .Y(clkd));
inv_lvt Iinv_ckfb ( .A(clatb), .Y(net50));
inv_lvt I40 ( .A(r), .Y(rstb));
inv_lvt I_q_inv ( .A(qn), .Y(q));
inv_lvt I39 ( .A(net77), .Y(qn));
txgate_lvt I52 ( .in(so), .out(mi), .pp(clkb), .nn(clkd));
txgate_lvt I44 ( .in(d), .out(si), .pp(clkd), .nn(clkb));
txgate_lvt I51 ( .in(si), .out(low_s), .pp(clkb), .nn(clkd));
txgate_lvt I53 ( .in(mi), .out(qn), .pp(clkd), .nn(clkb));
nand2_lvt I290 ( .A(clk), .Y(clkb), .B(clatb));
nand2_lvt I42 ( .A(si), .Y(so), .B(rstb));
nor2_lvt INAND2_m ( .A(r), .B(mi), .Y(net77));
anor21_lvt I54 ( .A(net50), .B(clk), .Y(clatb), .C(ceb));

endmodule
// Library - io, Cell - dffrckb, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module dffrckb ( q, qn, clk, d, e, r );
output  q, qn;

input  clk, d, e, r;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



oai21x2_lvt I57 ( .A1(clk), .Y(clat), .A0(clatb), .B0(e));
nor2_lvt I48 ( .B(clat), .A(clk), .Y(clkb));
nand2_lvt I54 ( .A(rstb), .Y(qn), .B(q));
nand2_lvt I42 ( .A(si), .B(rstb), .Y(so));
txgate_lvt I59 ( .in(d), .out(si), .pp(clkb), .nn(clkd));
txgate_lvt I64 ( .in(low_s), .out(si), .pp(clkd), .nn(clkb));
txgate_lvt I62 ( .in(qn), .out(mi), .pp(clkb), .nn(clkd));
txgate_lvt I60 ( .in(so), .out(mi), .pp(clkd), .nn(clkb));
inv_lvt I55 ( .A(mi), .Y(q));
inv_lvt I50 ( .A(clkb), .Y(clkd));
inv_lvt I56 ( .A(clat), .Y(clatb));
inv_lvt I43 ( .A(so), .Y(low_s));
inv_lvt I40 ( .A(r), .Y(rstb));

endmodule
// Library - io, Cell - in_logic_v1_imp, View - schematic
// LAST TIME SAVED: Jun 24 11:06:20 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module in_logic_v1_imp ( dout0, dout1, sdo, bs_en, cbit, cbitb, ceb,
     clk, cntl, din, mode, rstio, sdi, shift, tclk, ud );
output  dout0, dout1, sdo;

input  bs_en, ceb, clk, cntl, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbitb;
input [1:0]  cbit;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



insel1_lvt_imp I_insel1 ( .in1(dinb), .in0(regb), .out(reg_),
     .sb({cbit1b, cbitb[0]}), .sel({cbit1, cbit[0]}), .in2(net037),
     .in3(net037));
mux2x1_hvt I_mux_mode ( .sel(mode), .in1(udd), .in0(reg_),
     .out(doutb));
mux2x1_hvt I_mux_clk ( .in1(tclk), .in0(clk), .out(ck2r0),
     .sel(bs_en));
mux2x1_hvt I_mux_data ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
mux2x1_hvt I_mux2_btw ( .in1(sdo), .in0(din), .out(net056),
     .sel(bs_en));
nand2_lvt I188 ( .A(cntl), .Y(cbit1b), .B(cbit[1]));
inv_lvt I_inv_dout0 ( .A(doutb), .Y(dout0));
inv_lvt I_inv_dout1 ( .A(udd), .Y(dout1));
inv_lvt I185 ( .A(cbit1b), .Y(cbit1));
inv_lvt I186 ( .A(dout0), .Y(net037));
inv_lvt I172 ( .A(din), .Y(dinb));
cebdffrqn I_dff0 ( .ceb(ceb), .clk(ck2r0), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff1 ( .e(ud), .clk(ck2r0), .qn(udd), .r(rstio), .q(net060),
     .d(net056));

endmodule
// Library - io, Cell - in_logic_v3_imp, View - schematic
// LAST TIME SAVED: Aug  3 19:20:23 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module in_logic_v3_imp ( dout0, dout1, sdo, sp12, bl, bs_en, ceb, clk,
     cntl, din, mode, pgate, prog, reset, rstio, sdi, shift, slfop,
     tclk, ud, vdd_cntl, wl );
output  dout0, dout1, sdo, sp12;


input  bs_en, ceb, clk, cntl, din, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



P_11_LPHVT  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
P_11_LPHVT  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
in_logic_v1_imp I_in_logic ( .ceb(ceb), .rstio(rstio), .din(din),
     .cntl(cntl), .dout1(dout1), .dout0(dout0), .shift(shift), .ud(ud),
     .clk(clk), .sdo(sdo), .sdi(sdi), .cbit({cbit[0], cbit[1]}),
     .cbitb({cbitb[0], cbitb[1]}), .tclk(tclk), .bs_en(bs_en),
     .mode(mode));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[3]), .sp12(sp12),
     .prog(prog));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - outsel1_lvt, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module outsel1_lvt ( out, clk, in0, in1, in2, sb, sel );
output  out;

input  clk, in0, in1, in2;

input [1:0]  sel;
input [1:0]  sb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_lvt I41 ( .A(in1), .Y(net036));
inv_lvt I40 ( .A(clk), .Y(clkb));
txgate_lvt I33 ( .in(whatever), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_lvt I_txgate1 ( .in(net036), .out(whatever), .pp(sb[0]),
     .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(whatever), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(ddr), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_lvt I38 ( .in(in2), .out(ddr), .pp(clkb), .nn(clk));
txgate_lvt I39 ( .in(in1), .out(ddr), .pp(clk), .nn(clkb));

endmodule
// Library - io, Cell - out_logic_v1, View - schematic
// LAST TIME SAVED: Aug 13 11:02:21 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module out_logic_v1 ( dout, sdo, bs_en, cbit, cbitb, ceb, clk, ddr0,
     ddr1, mode, rstio, sdi, shift, tclk, ud );
output  dout, sdo;

input  bs_en, ceb, clk, ddr0, ddr1, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



outsel1_lvt I169 ( .clk(ddrclk), .in2(udb), .sb(cbitb[1:0]),
     .sel(cbit[1:0]), .in1(net094), .in0(dinb), .out(muxob));
mux2x1_hvt I170 ( .sel(mode), .in1(udb), .in0(muxob), .out(doutb));
mux2x1_hvt I177 ( .in1(tclk), .in0(clk), .out(mux4clk), .sel(bs_en));
mux2x1_hvt I173 ( .in1(sdi), .in0(ddr0), .out(dd), .sel(shift));
mux2x1_hvt I176 ( .in1(sdo), .in0(ddr1), .out(mux4d), .sel(bs_en));
nor2_lvt I179 ( .A(mux4clk), .B(cbit[0]), .Y(ddrclk));
inv_lvt I171 ( .A(doutb), .Y(dout));
inv_lvt I172 ( .A(ddr0), .Y(dinb));
cebdffrqn I_reg0 ( .ceb(ceb), .clk(mux4clk), .qn(net094), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_reg1 ( .e(ud), .clk(mux4clk), .qn(udb), .r(rstio), .q(net44),
     .d(mux4d));

endmodule
// Library - NVCM_40nm, Cell - ml_dff_nvcm, View - schematic
// LAST TIME SAVED: Aug  3 19:29:00 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_dff_nvcm ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I132 ( .A(clk_b), .Y(clk_buf));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I146 ( .A(net57), .Y(Q));
inv_hvt I147 ( .A(net60), .Y(QN));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net64), .Y(net57));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net64), .Y(net53));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net60), .Y(net57));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net53));
nor2_hvt I129 ( .A(net57), .B(R), .Y(net60));
nor2_hvt I125 ( .A(net53), .B(R), .Y(net64));

endmodule
// Library - io, Cell - out_logic_v3, View - schematic
// LAST TIME SAVED: Aug  3 19:20:30 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module out_logic_v3 ( dout, sdo, sp12, bl, bs_en, ceb, clk, ddr0, ddr1,
     mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk, ud,
     vdd_cntl, wl );
output  dout, sdo, sp12;


input  bs_en, ceb, clk, ddr0, ddr1, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;

wire  [3:0]  cbit;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
out_logic_v1 I_outlogic_v1 ( .shift(shift), .ud(ud), .clk(clk),
     .sdo(sdo), .sdi(sdi), .ceb(ceb), .cbit({cbit[2], cbit[3]}),
     .cbitb({cbitb[2], cbitb[3]}), .dout(dout), .ddr0(ddr0),
     .tclk(tclk), .bs_en(bs_en), .rstio(rstio), .ddr1(ddr1),
     .mode(mode));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
odrv12 I_odrv12 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp12(sp12));

endmodule
// Library - io, Cell - ioesel_lvt, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioesel_lvt ( out, in0, in1, sb, sel );
output  out;

input  in0, in1;

input [1:0]  sb;
input [1:0]  sel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_lvt I38 ( .A(sel[0]), .Y(net017));
txgate_lvt I33 ( .in(mid), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_lvt I_txgate1 ( .in(in1), .out(mid), .pp(sb[0]), .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(mid), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(net017), .out(out), .pp(sel[1]), .nn(sb[1]));

endmodule
// Library - io, Cell - ioe_logic_v1, View - schematic
// LAST TIME SAVED: Aug 13 14:52:51 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioe_logic_v1 ( outb, sdo, bs_en, cbit, cbitb, ceb, clk, din,
     mode, rstio, sdi, shift, tclk, ud );
output  outb, sdo;

input  bs_en, ceb, clk, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ioesel_lvt I_ioe_mux2 ( .sb(cbitb[1:0]), .sel(cbit[1:0]), .in1(regb),
     .in0(dinb), .out(regmuxb));
mux2x1_hvt I175 ( .in1(tclk), .in0(clk), .out(net039), .sel(bs_en));
mux2x1_hvt I170 ( .sel(mode), .in1(udd), .in0(regmuxb), .out(outb));
mux2x1_hvt I173 ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
inv_lvt I172 ( .A(din), .Y(dinb));
cebdffrqn I_dff_1 ( .ceb(ceb), .clk(net039), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff_2 ( .e(ud), .clk(net039), .qn(udd), .r(rstio), .q(net44),
     .d(sdo));

endmodule
// Library - io, Cell - ioe_logic_v3, View - schematic
// LAST TIME SAVED: Aug  3 19:20:27 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioe_logic_v3 ( padeb, sdo, sp12, bl, bs_en, ceb, clk, din,
     hiz_b, mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk,
     ud, vdd_cntl, wl );
output  padeb, sdo, sp12;


input  bs_en, ceb, clk, din, hiz_b, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbit;

wire  [3:0]  cbitb;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
inv_lvt I_inv ( .A(oeb), .Y(oed));
nand2_lvt I_nand2 ( .A(oed), .Y(padeb), .B(hiz_b));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
ioe_logic_v1 I_ioe_logic ( .shift(shift), .ud(ud), .clk(clk),
     .sdo(sdo), .sdi(sdi), .cbit(cbit[3:2]), .din(din),
     .cbitb(cbitb[3:2]), .ceb(ceb), .rstio(rstio), .bs_en(bs_en),
     .tclk(tclk), .outb(oeb), .mode(mode));
odrv12 I_odrv12x2 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp12(sp12));

endmodule
// Library - io, Cell - odrv12x3, View - schematic
// LAST TIME SAVED: Aug  3 19:20:30 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module odrv12x3 ( sp12, bl, pgate, prog, reset, slfop, vdd_cntl, wl );


input  prog;

output [2:0]  sp12;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [2:0]  slfop;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12_2_ ( .slfop(slfop[2]), .cbitb(cbitb[2]),
     .sp12(sp12[2]), .prog(prog));
odrv12 I_odrv12_1_ ( .slfop(slfop[1]), .cbitb(cbitb[1]),
     .sp12(sp12[1]), .prog(prog));
odrv12 I_odrv12_0_ ( .slfop(slfop[0]), .cbitb(cbitb[0]),
     .sp12(sp12[0]), .prog(prog));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioe_col2_v3, View - schematic
// LAST TIME SAVED: May 12 17:42:20 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioe_col2_v3 ( dout, padeb, pado, sdo, sp12_h_l, bl, bs_en, ceb,
     hiz_b, hold, inclk, mode, outclk, padin, pgate, prog, reset,
     rstio, sdi, shift, tclk, ti, update, vdd_cntl, wl );
output  sdo;


input  bs_en, ceb, hiz_b, hold, inclk, mode, outclk, prog, rstio, sdi,
     shift, tclk, update;

output [1:0]  pado;
output [23:0]  sp12_h_l;
output [3:0]  dout;
output [1:0]  padeb;

inout [1:0]  bl;

input [1:0]  padin;
input [5:0]  ti;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



in_logic_v3_imp I_in1 ( .slfop(dout[3]), .shift(shift),
     .dout1(dout[3]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[2]), .sp12(sp12_h_l[14]), .wl(wl[13:12]),
     .ceb(ceb), .reset(reset[13:12]), .sdo(s4), .sdi(s3),
     .vdd_cntl(vdd_cntl[13:12]), .pgate(pgate[13:12]), .din(padin[1]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode),
     .rstio(rstio));
in_logic_v3_imp I_in0 ( .slfop(dout[0]), .shift(shift),
     .dout1(dout[1]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[0]), .sp12(sp12_h_l[8]), .wl(wl[3:2]),
     .ceb(ceb), .reset(reset[3:2]), .sdo(s1), .sdi(s0),
     .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]), .din(padin[0]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode),
     .rstio(rstio));
out_logic_v3 I_out1 ( .shift(shift), .slfop(dout[3]), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .sp12(sp12_h_l[6]),
     .wl(wl[11:10]), .ceb(ceb), .reset(reset[11:10]), .sdo(s3),
     .sdi(s2), .vdd_cntl(vdd_cntl[11:10]), .pgate(pgate[11:10]),
     .dout(pado[1]), .tclk(tclk), .bs_en(bs_en), .rstio(rstio),
     .ddr1(ti[5]), .mode(mode), .ddr0(ti[4]));
out_logic_v3 I_out0 ( .shift(shift), .slfop(dout[0]), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .sp12(sp12_h_l[0]),
     .wl(wl[1:0]), .ceb(ceb), .reset(reset[1:0]), .sdo(s0), .sdi(sdi),
     .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]), .dout(pado[0]),
     .tclk(tclk), .bs_en(bs_en), .rstio(rstio), .ddr1(ti[2]),
     .mode(mode), .ddr0(ti[1]));
ioe_logic_v3 I_ioe0 ( .shift(shift), .hiz_b(hiz_b), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .padeb(padeb[0]),
     .slfop(dout[0]), .sp12(sp12_h_l[16]), .wl(wl[5:4]), .ceb(ceb),
     .reset(reset[5:4]), .sdo(s2), .sdi(s1), .pgate(pgate[5:4]),
     .din(ti[0]), .tclk(tclk), .vdd_cntl(vdd_cntl[5:4]), .bs_en(bs_en),
     .mode(mode), .rstio(rstio));
ioe_logic_v3 I_ioe1 ( .shift(shift), .hiz_b(hiz_b), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .padeb(padeb[1]),
     .slfop(dout[3]), .sp12(sp12_h_l[22]), .wl(wl[15:14]), .ceb(ceb),
     .reset(reset[15:14]), .sdo(sdo), .sdi(s4), .pgate(pgate[15:14]),
     .din(ti[3]), .tclk(tclk), .vdd_cntl(vdd_cntl[15:14]),
     .bs_en(bs_en), .mode(mode), .rstio(rstio));
odrv12x3 I_odrv12x3_1 ( .bl(bl[1:0]), .wl(wl[7:6]), .reset(reset[7:6]),
     .pgate(pgate[7:6]), .slfop({dout[1], dout[1], dout[1]}),
     .sp12({sp12_h_l[18], sp12_h_l[10], sp12_h_l[2]}),
     .vdd_cntl(vdd_cntl[7:6]), .prog(prog));
odrv12x3 I_odrv12x3_2 ( .bl(bl[1:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]), .slfop({dout[2], dout[2], dout[2]}),
     .sp12({sp12_h_l[20], sp12_h_l[12], sp12_h_l[4]}),
     .vdd_cntl(vdd_cntl[9:8]), .prog(prog));

endmodule
// Library - ice8chip, Cell - io_col4_lft_ice8p_v2, View - schematic
// LAST TIME SAVED: Aug  3 19:20:04 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_col4_lft_ice8p_v2 ( cbit_colcntl, cf, fabric_out, padeb,
     pado, sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t,
     sp12_h_l, bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold,
     lft_op, mode, padin, pgate, prog, r, reset, sdi, shift, spioeb,
     spiout, tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [7:0]  cbit_colcntl;
output [1:0]  pado;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;
output [1:0]  padeb;
output [23:0]  cf;

inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;

input [1:0]  spioeb;
input [15:0]  wl;
input [15:0]  reset;
input [15:0]  pgate;
input [7:0]  bnl_op;
input [7:0]  tnl_op;
input [15:0]  vdd_cntl;
input [7:0]  glb_netwk;
input [1:0]  spiout;
input [1:0]  padin;
input [7:0]  lft_op;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [1:0]  om;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [3:0]  t_mid;



RM7  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
RM7  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
RM7  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
RM7  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
RM7  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
RM7  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
RM7  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
RM7  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
RM7  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
RM7  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
RM7  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
RM7  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
RM7  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
RM7  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
RM7  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
RM7  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
sbox1_colbdlc_v4 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_gmux_x16bare_v4 I_io_gmux_x16bare_v4 (
     .cbit_colcntl(cbit_colcntl[7:0]), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));

endmodule
// Library - ice384chip, Cell - io_lft_bot_1x4_ice384, View - schematic
// LAST TIME SAVED: Nov 11 14:59:11 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_lft_bot_1x4_ice384 ( cf_l, fabric_out_03, fabric_out_04,
     padeb, pado, sdo, slf_op_01, slf_op_02, slf_op_03, slf_op_04,
     tclk_o, SP4_h_l_01, SP4_h_l_02, SP4_h_l_03, SP4_h_l_04,
     SP12_h_l_01, SP12_h_l_02, SP12_h_l_03, SP12_h_l_04, bl, glb_netwk,
     pgate, reset_b, sp4_v_b_00_01, sp4_v_t_04, vdd_cntl, wl,
     bnr_op_00_01, bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu0_b,
     last_rsr, mode, padin, prog, r, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, sdi, shift, tclk, tnr_op_04, update );
output  fabric_out_03, fabric_out_04, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu0_b, mode, prog,
     r, sdi, shift, tclk, update;

output [3:0]  slf_op_04;
output [3:0]  slf_op_03;
output [3:0]  slf_op_01;
output [3:0]  slf_op_02;
output [7:0]  padeb;
output [7:0]  pado;
output [95:0]  cf_l;

inout [47:0]  SP4_h_l_02;
inout [23:0]  SP12_h_l_02;
inout [47:0]  SP4_h_l_04;
inout [15:0]  sp4_v_t_04;
inout [47:0]  SP4_h_l_03;
inout [47:0]  SP4_h_l_01;
inout [23:0]  SP12_h_l_04;
inout [23:0]  SP12_h_l_01;
inout [17:0]  bl;
inout [63:0]  vdd_cntl;
inout [63:0]  reset_b;
inout [63:0]  wl;
inout [7:0]  glb_netwk;
inout [23:0]  SP12_h_l_03;
inout [63:0]  pgate;
inout [15:0]  sp4_v_b_00_01;

input [7:0]  rgt_op_04;
input [7:0]  bnr_op_00_01;
input [7:0]  rgt_op_01;
input [7:0]  tnr_op_04;
input [7:0]  rgt_op_03;
input [7:0]  padin;
input [7:0]  rgt_op_02;
input [0:0]  last_rsr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net0626;

wire  [15:0]  net937;

wire  [7:0]  net1008;

wire  [1:0]  net1005;

wire  [15:0]  net901;

wire  [1:0]  net1009;

wire  [7:0]  net884;

wire  [7:0]  net1007;

wire  [15:0]  net865;

wire  [1:0]  net1014;

wire  [1:0]  net1002;



tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
fabric_buf_ice8p I172 ( .f_in(net955), .f_out(fabric_out_03));
fabric_buf_ice8p I171 ( .f_in(net0473), .f_out(fabric_out_04));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
io_col4_lft_ice8p_v2 I_io_00_02 ( .cbit_colcntl({net1007[0],
     net1007[1], net1007[2], net1007[3], net1007[4], net1007[5],
     net1007[6], net1007[7]}), .ceb(ceb), .sdo(net887), .sdi(net851),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin(padin[3:2]),
     .pado(pado[3:2]), .padeb(padeb[3:2]), .sp4_v_t({net865[0],
     net865[1], net865[2], net865[3], net865[4], net865[5], net865[6],
     net865[7], net865[8], net865[9], net865[10], net865[11],
     net865[12], net865[13], net865[14], net865[15]}),
     .sp4_h_l(SP4_h_l_02[47:0]), .sp12_h_l(SP12_h_l_02[23:0]),
     .prog(prog), .spi_ss_in_b({net1014[0], net1014[1]}),
     .tnl_op(rgt_op_03[7:0]), .lft_op(rgt_op_02[7:0]),
     .bnl_op(rgt_op_01[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15]}), .wl(wl[31:16]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(net883));
io_col4_lft_ice8p_v2 I_io_00_01 ( .cbit_colcntl({net884[0], net884[1],
     net884[2], net884[3], net884[4], net884[5], net884[6],
     net884[7]}), .ceb(ceb), .sdo(sdo), .sdi(net887), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin(padin[1:0]),
     .pado(pado[1:0]), .padeb(padeb[1:0]), .sp4_v_t({net901[0],
     net901[1], net901[2], net901[3], net901[4], net901[5], net901[6],
     net901[7], net901[8], net901[9], net901[10], net901[11],
     net901[12], net901[13], net901[14], net901[15]}),
     .sp4_h_l(SP4_h_l_01[47:0]), .sp12_h_l(SP12_h_l_01[23:0]),
     .prog(prog), .spi_ss_in_b({net1005[0], net1005[1]}),
     .tnl_op(rgt_op_02[7:0]), .lft_op(rgt_op_01[7:0]),
     .bnl_op(bnr_op_00_01[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_00_01[15:0]),
     .wl(wl[15:0]), .cf(cf_l[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk[7:0]), .hold(hold), .fabric_out(net0546));
io_col4_lft_ice8p_v2 I_io_00_03 ( .cbit_colcntl({net1008[0],
     net1008[1], net1008[2], net1008[3], net1008[4], net1008[5],
     net1008[6], net1008[7]}), .ceb(ceb), .sdo(net851), .sdi(net923),
     .spiout({tiegnd, last_rsr[0]}),
     .cdone_in(jtag_rowtest_mode_rowu0_b), .spioeb({tievdd, tiegnd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin(padin[5:4]),
     .pado(pado[5:4]), .padeb(padeb[5:4]), .sp4_v_t({net937[0],
     net937[1], net937[2], net937[3], net937[4], net937[5], net937[6],
     net937[7], net937[8], net937[9], net937[10], net937[11],
     net937[12], net937[13], net937[14], net937[15]}),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b({net1009[0], net1009[1]}),
     .tnl_op(rgt_op_04[7:0]), .lft_op(rgt_op_03[7:0]),
     .bnl_op(rgt_op_02[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b({net865[0], net865[1], net865[2],
     net865[3], net865[4], net865[5], net865[6], net865[7], net865[8],
     net865[9], net865[10], net865[11], net865[12], net865[13],
     net865[14], net865[15]}), .wl(wl[47:32]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(net955));
io_col4_lft_ice8p_v2 I_io_00_04 ( .cbit_colcntl({net0626[0],
     net0626[1], net0626[2], net0626[3], net0626[4], net0626[5],
     net0626[6], net0626[7]}), .ceb(ceb), .sdo(net923), .sdi(sdi),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin(padin[7:6]),
     .pado(pado[7:6]), .padeb(padeb[7:6]), .sp4_v_t(sp4_v_t_04[15:0]),
     .sp4_h_l(SP4_h_l_04[47:0]), .sp12_h_l(SP12_h_l_04[23:0]),
     .prog(prog), .spi_ss_in_b({net1002[0], net1002[1]}),
     .tnl_op(tnr_op_04[7:0]), .lft_op(rgt_op_04[7:0]),
     .bnl_op(rgt_op_03[7:0]), .pgate(pgate[63:48]),
     .reset(reset_b[63:48]), .sp4_v_b({net937[0], net937[1], net937[2],
     net937[3], net937[4], net937[5], net937[6], net937[7], net937[8],
     net937[9], net937[10], net937[11], net937[12], net937[13],
     net937[14], net937[15]}), .wl(wl[63:48]), .cf(cf_l[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(net0473));

endmodule
// Library - leafcell, Cell - bram_bufferx4x6, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module bram_bufferx4x6 ( out, in );
output  out;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I4 ( .in(d1), .out(d2));
bram_bufferx4 I5 ( .in(d2), .out(d3));
bram_bufferx4 I6 ( .in(d3), .out(d4));
bram_bufferx4 I7 ( .in(d4), .out(out));
bram_bufferx4 I3 ( .in(d0), .out(d1));
bram_bufferx4 I0 ( .in(in), .out(d0));

endmodule
// Library - leafcell, Cell - lowla_modified, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module lowla_modified ( lao, clk, min );
output  lao;

input  clk, min;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I249 ( .in(lao), .out(st2), .pp(cbitb), .nn(clkd));
txgate_hvt I248 ( .in(min), .out(st2), .pp(clkd), .nn(cbitb));
inv_hvt I289 ( .A(net29), .Y(lao));
inv_hvt I290 ( .A(st2), .Y(net29));
inv_hvt I_inv ( .A(clk), .Y(cbitb));
inv_hvt I_inv3 ( .A(cbitb), .Y(clkd));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_resref_40nm, View - schematic
// LAST TIME SAVED: Sep 24 16:17:12 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_sa_resref_40nm ( bl_in, bl_out, ref );
inout  bl_in, bl_out;

inout [3:0]  ref;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



RNPPO_LP_pcell2460 R9 ( .B(gnd_), .MINUS(ref[3]), .PLUS(ref[2]));
RNPPO_LP_pcell2460 R11 ( .B(gnd_), .MINUS(ref[1]), .PLUS(ref[0]));
RNPPO_LP_pcell2460 R18 ( .B(gnd_), .MINUS(net41), .PLUS(bl_in));
RNPPO_LP_pcell2460 R10 ( .B(gnd_), .MINUS(ref[2]), .PLUS(ref[1]));
RNPPO_LP_pcell2460 R7 ( .B(gnd_), .MINUS(ref[0]), .PLUS(net41));
RNPPO_LP_pcell2460 R24 ( .B(gnd_), .MINUS(bl_out), .PLUS(ref[3]));

endmodule
// Library - ice8chip, Cell - scan_buf_ice8p, View - schematic
// LAST TIME SAVED: Jun 28 09:23:39 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module scan_buf_ice8p ( bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo,
     shift_o, tclk_o, update_o, bs_en_i, ceb_i, hiz_b_i, mode_i, r_i,
     sdi, shift_i, tclk_i, update_i );
output  bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo, shift_o, tclk_o,
     update_o;

input  bs_en_i, ceb_i, hiz_b_i, mode_i, r_i, sdi, shift_i, tclk_i,
     update_i;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



tckbufx32_ice8p I_tclkbuf ( .in(tclk_i), .out(tclk_o));
bram_bufferx4 I_bs_enbuf ( .in(bs_en_i), .out(bs_en_o));
bram_bufferx4 I_cebbuf ( .in(ceb_i), .out(ceb_o));
bram_bufferx4 I_modebuf ( .in(mode_i), .out(mode_o));
bram_bufferx4 I_hiz_bbuf ( .in(hiz_b_i), .out(hiz_b_o));
bram_bufferx4 I_updatebuf ( .in(update_i), .out(update_o));
bram_bufferx4 I_shiftbuf ( .in(shift_i), .out(shift_o));
bram_bufferx4 I_rbuf ( .in(r_i), .out(r_o));
bram_bufferx4x6 I_sdibuf ( .in(sdi), .out(sdi_2));
lowla_modified I_lowla ( .clk(tclk_i), .min(sdi_2), .lao(sdo));

endmodule
// Library - io, Cell - io_gmux_x2v2, View - schematic
// LAST TIME SAVED: Aug  3 19:20:26 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_gmux_x2v2 ( .cbitb_colcntl({cbitb[11], cbitb[9]}), gout, bl,
     min0, min1, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [1:0]  gout;
output [11:0]  cbitb;

inout [5:0]  bl;

input [15:0]  min0;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [15:0]  min1;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux I_g_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux I_g_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare_v3, View - schematic
// LAST TIME SAVED: Jun  2 10:52:40 2010
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module io_gmux_x16bare_v3 ( cbitb_colcntl, lc_trk_g0, lc_trk_g1, bl,
     min0, min1, min2, min3, min4, min5, min6, min7, min8, min9, min10,
     min11, min12, min13, min14, min15, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  cbitb_colcntl;

inout [5:0]  bl;

input [15:0]  min7;
input [15:0]  min0;
input [15:0]  min9;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min15;
input [15:0]  min3;
input [15:0]  min14;
input [15:0]  min12;
input [15:0]  min6;
input [15:0]  min8;
input [15:0]  min5;
input [15:0]  min4;
input [15:0]  min11;
input [15:0]  min10;
input [15:0]  vdd_cntl;
input [15:0]  min2;
input [15:0]  reset;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net114;

wire  [1:0]  net187;

wire  [1:0]  net188;

wire  [1:0]  net124;



io_gmux_x2v2 I_io_gmux_x2_7 ( .cbitb_colcntl({net114[0], net114[1]}),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[15:14]));
io_gmux_x2v2 I_io_gmux_x2_6 ( .cbitb_colcntl({net124[0], net124[1]}),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[13:12]));
io_gmux_x2v2 I_io_gmux_x2_2 ( .cbitb_colcntl(cbitb_colcntl[5:4]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[5:4]));
io_gmux_x2v2 I_io_gmux_x2_0 ( .cbitb_colcntl(cbitb_colcntl[1:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[1:0]));
io_gmux_x2v2 _io_gmux_x2_1 ( .cbitb_colcntl(cbitb_colcntl[3:2]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[3:2]));
io_gmux_x2v2 I_io_gmux_x2_4 ( .cbitb_colcntl({net187[0], net187[1]}),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[9:8]));
io_gmux_x2v2 I_io_gmux_x2_5 ( .cbitb_colcntl({net188[0], net188[1]}),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[11:10]));
io_gmux_x2v2 I_io_gmux_x2_3 ( .cbitb_colcntl(cbitb_colcntl[7:6]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[7:6]));

endmodule
// Library - io, Cell - ioinmx1mux2_imp, View - schematic
// LAST TIME SAVED: Aug  3 19:20:28 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioinmx1mux2_imp ( clk, mo, ti, bl, cdone_in, ce, ceb, in, min,
     pgate, prog, reset, spi, vdd_cntl, wl );
output  clk, ti;


input  cdone_in, ceb, prog;

output [1:0]  mo;

inout [5:0]  bl;

input [1:0]  spi;
input [11:0]  ce;
input [7:0]  min;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  in;
input [1:0]  vdd_cntl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  moo;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  mob;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
mux2x1_hvt I_emux_1_ ( .in1(in[1]), .in0(spi[1]), .out(moo[1]),
     .sel(cdone_in));
mux2x1_hvt I_emux_0_ ( .in1(in[0]), .in0(spi[0]), .out(moo[0]),
     .sel(cdone_in));
inv_lvt inv_1_1_ ( .A(moo[1]), .Y(mob[1]));
inv_lvt inv_1_0_ ( .A(moo[0]), .Y(mob[0]));
inv_lvt I_inv_2_1_ ( .A(mob[1]), .Y(mo[1]));
inv_lvt I_inv_2_0_ ( .A(mob[0]), .Y(mo[0]));
ioin_mux_v2 I_ioin_mux ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);
clk_mux12to1 I_clk_mux12to1 ( .prog(prog), .min(ce[11:0]), .clk(clk),
     .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7], cbitb[10],
     cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7], cbit[10],
     cbit[6], cbit[4]}), .cenb(ceb));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc, View - schematic
// LAST TIME SAVED: Aug  3 19:20:28 2011
// NETLIST TIME: Jan 18 18:48:20 2012
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  spi;
output [1:0]  ti;

inout [5:0]  bl;

input [7:0]  min2;
input [7:0]  min1;
input [1:0]  vdd_cntl;
input [7:0]  min0;
input [1:0]  padin;
input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
inv_lvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_lvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
nor2_lvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_lvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
ioin_mux_v2 I_ioin_mux_bankcntl ( bankcntl, {cbit[11], cbit[8], cbit[9],
     cbit[10]}, {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0],
     prog);
ioin_mux_v2 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v2 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nand2inv, View - schematic
// LAST TIME SAVED: Aug  3 19:20:28 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module ioinmx2nand2inv ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [7:0]  min0;
input [1:0]  pgate;
input [7:0]  ce;
input [7:0]  min1;
input [1:0]  reset;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



P_11_LPHVT  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
P_11_LPHVT  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
nand2_lvt I180 ( .A(update_b), .Y(updt), .B(bs_en));
inv_lvt I181 ( .A(update), .Y(update_b));
ioin_mux_v2 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v2 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc_v3, View - schematic
// LAST TIME SAVED: May 12 17:30:59 2010
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module sbox1_colbdlc_v3 ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  spi_ss_in_b;
output [1:0]  padeb;
output [5:0]  ti;
output [1:0]  pado;

inout [5:0]  bl;
inout [3:0]  t_mid;
inout [3:0]  sp4_v_b;
inout [3:0]  l;
inout [3:0]  r;

input [1:0]  out;
input [1:0]  padin;
input [11:0]  clk_in;
input [7:0]  min5;
input [1:0]  spiout;
input [7:0]  ceb_in;
input [7:0]  min4;
input [11:0]  inclk_in;
input [7:0]  min2;
input [1:0]  oeb;
input [7:0]  min1;
input [1:0]  spioeb;
input [7:0]  min3;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  min0;
input [7:0]  min6;
input [15:0]  wl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ioinmx1mux2_imp I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .in(out[1:0]), .ti(ti[2]), .min(min2[7:0]), .spi(spiout[1:0]),
     .wl(wl[9:8]), .reset(reset[9:8]), .pgate(pgate[9:8]),
     .cdone_in(cdone_in), .mo(pado[1:0]));
ioinmx1mux2_imp I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .in(oeb[1:0]), .ti(ti[5]), .min(min5[7:0]), .spi(spioeb[1:0]),
     .wl(wl[15:14]), .reset(reset[15:14]), .pgate(pgate[15:14]),
     .cdone_in(cdone_in), .mo(padeb[1:0]));
ioinmx2nor2invx2bdlc I5 ( .vdd_cntl(vdd_cntl[5:4]), .min2(min6[7:0]),
     .bankcntl(fabric_out), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx2nand2inv I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - ice8chip, Cell - io_col4_bot_ice8p, View - schematic
// LAST TIME SAVED: Aug  3 19:20:03 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_col4_bot_ice8p ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [23:0]  cf;
output [3:0]  slf_op;
output [1:0]  pado;

inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_b;
inout [15:0]  sp4_v_t;

input [1:0]  padin;
input [1:0]  spioeb;
input [1:0]  spiout;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  wl;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  glb_netwk;
input [15:0]  reset;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [7:0]  net225;



RM6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
RM6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
RM6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
RM6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
RM6  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
RM6  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
RM6  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
RM6  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
RM6  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
RM6  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
RM6  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
RM6  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
RM6  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
RM6  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
RM6  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
RM6  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
inv_lvt I_inv1 ( .A(prog), .Y(progb));
inv_lvt I_inv2 ( .A(progb), .Y(progd));
io_gmux_x16bare_v3 I_io_gmux_x16bare_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .cbitb_colcntl({net225[0], net225[1], net225[2], net225[3],
     net225[4], net225[5], net225[6], net225[7]}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
sbox1_colbdlc_v3 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));

endmodule
// Library - ice384chip, Cell - io_bot_lft_1x3_ice384, View - schematic
// LAST TIME SAVED: Nov 16 16:05:55 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_bot_lft_1x3_ice384 ( bs_en_o, ceb_o, cf_bot_l,
     fabric_out_02_00, fabric_out_03_00, hiz_b_o, mode_o, padeb_b_l,
     pado_b_l, r_o, sdo, shift_o, slf_op_01_00, slf_op_02_00,
     slf_op_03_00, tclk_o, update_o, bl_01, bl_02, bl_03,
     sp4_h_l_01_00, sp4_h_r_03_00, sp4_v_b_01_00, sp4_v_b_02_00,
     sp4_v_b_03_00, sp12_v_b_01_00, sp12_v_b_02_00, sp12_v_b_03_00,
     bnl_op_01_00, bs_en_i, ceb_i, glb_net_01, glb_net_02, glb_net_03,
     hiz_b_i, hold_b_l, lft_op_01_00, lft_op_02_00, lft_op_03_00,
     mode_i, padin_b_l, pgate_l, prog, r_i, reset_l, sdi, shift_i,
     tclk_i, tnr_op_03_00, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_02_00, fabric_out_03_00, hiz_b_o,
     mode_o, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_03_00;
output [3:0]  slf_op_02_00;
output [5:0]  pado_b_l;
output [5:0]  padeb_b_l;
output [71:0]  cf_bot_l;
output [3:0]  slf_op_01_00;

inout [47:0]  sp4_v_b_01_00;
inout [23:0]  sp12_v_b_01_00;
inout [15:0]  sp4_h_r_03_00;
inout [47:0]  sp4_v_b_03_00;
inout [47:0]  sp4_v_b_02_00;
inout [53:0]  bl_02;
inout [53:0]  bl_03;
inout [53:0]  bl_01;
inout [23:0]  sp12_v_b_03_00;
inout [15:0]  sp4_h_l_01_00;
inout [23:0]  sp12_v_b_02_00;

input [7:0]  glb_net_01;
input [7:0]  glb_net_03;
input [15:0]  reset_l;
input [7:0]  bnl_op_01_00;
input [15:0]  wl_l;
input [15:0]  pgate_l;
input [7:0]  lft_op_01_00;
input [7:0]  lft_op_03_00;
input [5:0]  padin_b_l;
input [7:0]  tnr_op_03_00;
input [15:0]  vdd_cntl_l;
input [7:0]  lft_op_02_00;
input [7:0]  glb_net_02;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net519;

wire  [1:0]  net312;

wire  [15:0]  net378;

wire  [1:0]  net382;

wire  [15:0]  net343;



fabric_buf_ice8p I362 ( .f_in(net0179), .f_out(fabric_out_03_00));
fabric_buf_ice8p I785 ( .f_in(net0181), .f_out(fabric_out_02_00));
scan_buf_ice8p I_scanbuf_bl ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net284), .shift_o(shift_o),
     .sdo(net286), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_bot_ice8p I_IO_02_00 ( .sdo(net327), .sdi(net362),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net378[0], net378[1], net378[2], net378[3],
     net378[4], net378[5], net378[6], net378[7], net378[8], net378[9],
     net378[10], net378[11], net378[12], net378[13], net378[14],
     net378[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_b_l[3:2]), .pado(pado_b_l[3:2]),
     .padeb(padeb_b_l[3:2]), .sp4_v_b({net343[0], net343[1], net343[2],
     net343[3], net343[4], net343[5], net343[6], net343[7], net343[8],
     net343[9], net343[10], net343[11], net343[12], net343[13],
     net343[14], net343[15]}), .sp4_h_l(sp4_v_b_02_00[47:0]),
     .sp12_h_l(sp12_v_b_02_00[23:0]), .prog(prog),
     .spi_ss_in_b({net312[0], net312[1]}), .tnl_op(lft_op_01_00[7:0]),
     .lft_op(lft_op_02_00[7:0]), .bnl_op(lft_op_03_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_02[5],
     bl_02[4], bl_02[37], bl_02[36], bl_02[35], bl_02[34], bl_02[33],
     bl_02[32], bl_02[14], bl_02[20], bl_02[19], bl_02[18], bl_02[17],
     bl_02[16], bl_02[27], bl_02[26], bl_02[25], bl_02[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[47:24]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_02_00[3:0]),
     .glb_netwk(glb_net_02[7:0]), .hold(hold_b_l),
     .fabric_out(net0181));
io_col4_bot_ice8p I_IO_01_00 ( .sdo(net362), .sdi(net286),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_01_00[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b_l[1:0]),
     .pado(pado_b_l[1:0]), .padeb(padeb_b_l[1:0]), .sp4_v_b({net378[0],
     net378[1], net378[2], net378[3], net378[4], net378[5], net378[6],
     net378[7], net378[8], net378[9], net378[10], net378[11],
     net378[12], net378[13], net378[14], net378[15]}),
     .sp4_h_l(sp4_v_b_01_00[47:0]), .sp12_h_l(sp12_v_b_01_00[23:0]),
     .prog(prog), .spi_ss_in_b({net382[0], net382[1]}),
     .tnl_op(bnl_op_01_00[7:0]), .lft_op(lft_op_01_00[7:0]),
     .bnl_op(lft_op_02_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[23:0]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_00[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_b_l), .fabric_out(net0310));
io_col4_bot_ice8p I_IO_03_00 ( .sdo(sdo), .sdi(net327),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net343[0], net343[1], net343[2], net343[3],
     net343[4], net343[5], net343[6], net343[7], net343[8], net343[9],
     net343[10], net343[11], net343[12], net343[13], net343[14],
     net343[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_b_l[5:4]), .pado(pado_b_l[5:4]),
     .padeb(padeb_b_l[5:4]), .sp4_v_b(sp4_h_r_03_00[15:0]),
     .sp4_h_l(sp4_v_b_03_00[47:0]), .sp12_h_l(sp12_v_b_03_00[23:0]),
     .prog(prog), .spi_ss_in_b({net519[0], net519[1]}),
     .tnl_op(lft_op_02_00[7:0]), .lft_op(lft_op_03_00[7:0]),
     .bnl_op(tnr_op_03_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[71:48]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_00[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_b_l), .fabric_out(net0179));
tckbufx32_ice8p I354 ( .in(net284), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));

endmodule
// Library - leafcell, Cell - pinlatbuf12p, View - schematic
// LAST TIME SAVED: Jul 30 23:15:00 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module pinlatbuf12p ( cout, cbit, icegate, pad_in, prog );
output  cout;

input  cbit, icegate, pad_in, prog;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I_txgate_lvt_2 ( .in(cout), .out(net13), .pp(net046),
     .nn(net17));
txgate_lvt I_txgate_lvt_1 ( .in(pad_in), .out(net13), .pp(net17),
     .nn(net046));
nand2_lvt I_nand2_lvt ( .A(net19), .Y(net044), .B(net13));
nand2_lvt I5 ( .A(icegate), .Y(net046), .B(cbit));
inv_lvt I6 ( .A(net046), .Y(net17));
inv_lvt I24 ( .A(prog), .Y(net19));
inv_lvt I_inv_lvt ( .A(net044), .Y(cout));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_restop_40nm, View - schematic
// LAST TIME SAVED: Sep 24 16:17:49 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_sa_restop_40nm ( bl_bot, bl_top );
inout  bl_bot, bl_top;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



RNPPO_LP_pcell2460 R24 ( .B(gnd_), .MINUS(bl_top), .PLUS(net66));
RNPPO_LP_pcell2460 R23 ( .B(gnd_), .MINUS(net66), .PLUS(bl_bot));

endmodule
// Library - leafcell, Cell - pinlatbuf12p_1, View - schematic
// LAST TIME SAVED: Jul 30 23:15:02 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module pinlatbuf12p_1 ( cout, cbit, icegate, pad_in, prog );
output  cout;

input  cbit, icegate, pad_in, prog;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I_txgate_lvt_2 ( .in(cout), .out(net13), .pp(net046),
     .nn(net17));
txgate_lvt I_txgate_lvt_1 ( .in(pad_in), .out(net13), .pp(net17),
     .nn(net046));
inv_lvt I6 ( .A(net046), .Y(net17));
inv_lvt I24 ( .A(prog), .Y(net19));
inv_lvt I_inv_lvt ( .A(net044), .Y(cout));
nand2_lvt I_nand2_lvt ( .A(net19), .Y(net044), .B(net13));
nand2_lvt I5 ( .A(icegate), .Y(net046), .B(cbit));

endmodule
// Library - ice384chip, Cell - quad_bl_ice384, View - schematic
// LAST TIME SAVED: Dec  5 14:02:36 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module quad_bl_ice384 ( bs_en_o, carry_out_01_04, carry_out_02_04,
     carry_out_03_04, ceb_o, cf_b_l, cf_l, fabric_out_00_03,
     fabric_out_00_04, fabric_out_02_00, fabric_out_03_00, hiz_b_o,
     mode_o, op_vic_01_04, op_vic_02_04, op_vic_03_04, padeb_b_l,
     padeb_l_b, padin_00_04b, padin_03_00b, pado_b_l, pado_l_b, r_o,
     sdo, shift_o, slf_op_00_04, slf_op_01_04, slf_op_02_04,
     slf_op_03_00, slf_op_03_01, slf_op_03_02, slf_op_03_03,
     slf_op_03_04, tclk_o, update_o, bl, pgate_l, reset_b_l,
     sp4_h_r_03_00, sp4_h_r_03_01, sp4_h_r_03_02, sp4_h_r_03_03,
     sp4_h_r_03_04, sp4_r_v_b_03_01, sp4_r_v_b_03_02, sp4_r_v_b_03_03,
     sp4_r_v_b_03_04, sp4_v_t_00_04, sp4_v_t_01_04, sp4_v_t_02_04,
     sp4_v_t_03_04, sp12_h_r_03_01, sp12_h_r_03_02, sp12_h_r_03_03,
     sp12_h_r_03_04, sp12_v_t_01_04, sp12_v_t_02_04, sp12_v_t_03_04,
     vdd_cntl_l, wl_l, bnr_op_03_01, bs_en_i, ceb_i, glb_in_0,
     glb_in_1, glb_in_2, glb_in_3, hiz_b_i, hold_b_l, hold_l_b,
     jtag_rowtest_mode_rowu0_b, last_rsr, mode_i, padin_b_l, padin_l_b,
     prog, purst, r_i, rgt_op_03_01, rgt_op_03_02, rgt_op_03_03,
     rgt_op_03_04, sdi, shift_i, tclk_i, tnl_op_01_04, tnl_op_02_04,
     tnl_op_03_04, tnr_op_00_04, tnr_op_01_04, tnr_op_02_04,
     tnr_op_03_04, top_op_01_04, top_op_02_04, top_op_03_04, update_i
     );
output  bs_en_o, carry_out_01_04, carry_out_02_04, carry_out_03_04,
     ceb_o, fabric_out_00_03, fabric_out_00_04, fabric_out_02_00,
     fabric_out_03_00, hiz_b_o, mode_o, op_vic_01_04, op_vic_02_04,
     op_vic_03_04, padin_00_04b, padin_03_00b, r_o, sdo, shift_o,
     tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_l, hold_l_b,
     jtag_rowtest_mode_rowu0_b, mode_i, prog, purst, r_i, sdi, shift_i,
     tclk_i, update_i;

output [7:0]  slf_op_03_04;
output [5:0]  pado_b_l;
output [7:0]  slf_op_02_04;
output [5:0]  padeb_b_l;
output [7:0]  slf_op_03_03;
output [7:0]  slf_op_01_04;
output [95:0]  cf_l;
output [71:0]  cf_b_l;
output [3:0]  slf_op_03_00;
output [7:0]  slf_op_03_02;
output [3:0]  slf_op_00_04;
output [7:0]  pado_l_b;
output [7:0]  padeb_l_b;
output [7:0]  slf_op_03_01;

inout [47:0]  sp4_h_r_03_03;
inout [47:0]  sp4_r_v_b_03_03;
inout [47:0]  sp4_v_t_03_04;
inout [47:0]  sp4_r_v_b_03_02;
inout [47:0]  sp4_r_v_b_03_01;
inout [23:0]  sp12_v_t_01_04;
inout [47:0]  sp4_h_r_03_04;
inout [23:0]  sp12_v_t_03_04;
inout [15:0]  sp4_v_t_00_04;
inout [15:0]  sp4_h_r_03_00;
inout [47:0]  sp4_h_r_03_02;
inout [47:0]  sp4_v_t_01_04;
inout [23:0]  sp12_h_r_03_01;
inout [47:0]  sp4_h_r_03_01;
inout [47:0]  sp4_r_v_b_03_04;
inout [23:0]  sp12_v_t_02_04;
inout [23:0]  sp12_h_r_03_03;
inout [79:0]  reset_b_l;
inout [47:0]  sp4_v_t_02_04;
inout [79:0]  wl_l;
inout [179:0]  bl;
inout [23:0]  sp12_h_r_03_04;
inout [79:0]  vdd_cntl_l;
inout [79:0]  pgate_l;
inout [23:0]  sp12_h_r_03_02;

input [7:0]  top_op_01_04;
input [7:0]  top_op_03_04;
input [7:0]  glb_in_2;
input [7:0]  glb_in_3;
input [7:0]  top_op_02_04;
input [7:0]  rgt_op_03_03;
input [7:0]  tnl_op_01_04;
input [7:0]  tnl_op_02_04;
input [7:0]  rgt_op_03_04;
input [7:0]  tnr_op_01_04;
input [7:0]  rgt_op_03_01;
input [7:0]  rgt_op_03_02;
input [7:0]  glb_in_1;
input [7:0]  tnl_op_03_04;
input [7:0]  glb_in_0;
input [7:0]  padin_l_b;
input [5:0]  padin_b_l;
input [3:0]  bnr_op_03_01;
input [0:0]  last_rsr;
input [7:0]  tnr_op_00_04;
input [7:0]  tnr_op_02_04;
input [7:0]  tnr_op_03_04;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  slf_op_02_00;

wire  [3:0]  slf_op_01_00;

wire  [3:0]  slf_op_00_01;

wire  [7:7]  padinlat_l_b;

wire  [3:0]  slf_op_00_02;

wire  [3:0]  slf_op_00_03;

wire  [5:5]  padinlat_b_l;

wire  [15:0]  net515;

wire  [47:0]  net355;

wire  [7:0]  net589;

wire  [47:0]  net587;

wire  [23:0]  net538;

wire  [47:0]  net608;

wire  [7:0]  net590;

wire  [23:0]  net539;

wire  [47:0]  net487;

wire  [47:0]  net524;

wire  [47:0]  net473;

wire  [47:0]  net521;

wire  [23:0]  net353;

wire  [47:0]  net361;

wire  [23:0]  net537;

wire  [47:0]  net582;

wire  [23:0]  net541;

wire  [47:0]  net470;

wire  [47:0]  net362;

wire  [7:0]  net518;

wire  [23:0]  net352;

wire  [47:0]  net471;

wire  [47:0]  net522;

wire  [23:0]  net465;

wire  [47:0]  net588;

wire  [47:0]  net357;

wire  [23:0]  net350;

wire  [47:0]  net474;

wire  [23:0]  net464;

wire  [47:0]  net475;

wire  [47:0]  net359;

wire  [23:0]  net466;

wire  [23:0]  net583;

wire  [23:0]  net351;

wire  [47:0]  net486;

wire  [47:0]  net476;

wire  [7:0]  net447;

wire  [47:0]  net356;

wire  [47:0]  net360;

wire  [7:0]  net526;

wire  [23:0]  net575;

wire  [7:0]  net445;

wire  [47:0]  net523;

wire  [47:0]  net469;

wire  [23:0]  net467;

wire  [23:0]  net561;



lt_1x4_bot_ice384 I805 ( .rgt_op_03(slf_op_03_03[7:0]),
     .slf_op_02({net447[0], net447[1], net447[2], net447[3], net447[4],
     net447[5], net447[6], net447[7]}), .rgt_op_02(slf_op_03_02[7:0]),
     .rgt_op_01(slf_op_03_01[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(slf_op_01_04[7:0]), .lft_op_03({net526[0], net526[1],
     net526[2], net526[3], net526[4], net526[5], net526[6],
     net526[7]}), .lft_op_02({net518[0], net518[1], net518[2],
     net518[3], net518[4], net518[5], net518[6], net518[7]}),
     .lft_op_01({net589[0], net589[1], net589[2], net589[3], net589[4],
     net589[5], net589[6], net589[7]}), .rgt_op_04(slf_op_03_04[7:0]),
     .carry_in(tiegnd_bl), .bnl_op_01({slf_op_01_00[3],
     slf_op_01_00[2], slf_op_01_00[1], slf_op_01_00[0],
     slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0]}), .slf_op_04(slf_op_02_04[7:0]),
     .slf_op_03({net445[0], net445[1], net445[2], net445[3], net445[4],
     net445[5], net445[6], net445[7]}), .slf_op_01({net590[0],
     net590[1], net590[2], net590[3], net590[4], net590[5], net590[6],
     net590[7]}), .sp4_h_l_04({net473[0], net473[1], net473[2],
     net473[3], net473[4], net473[5], net473[6], net473[7], net473[8],
     net473[9], net473[10], net473[11], net473[12], net473[13],
     net473[14], net473[15], net473[16], net473[17], net473[18],
     net473[19], net473[20], net473[21], net473[22], net473[23],
     net473[24], net473[25], net473[26], net473[27], net473[28],
     net473[29], net473[30], net473[31], net473[32], net473[33],
     net473[34], net473[35], net473[36], net473[37], net473[38],
     net473[39], net473[40], net473[41], net473[42], net473[43],
     net473[44], net473[45], net473[46], net473[47]}),
     .carry_out(carry_out_02_04), .vdd_cntl(vdd_cntl_l[79:16]),
     .sp12_h_r_04({net350[0], net350[1], net350[2], net350[3],
     net350[4], net350[5], net350[6], net350[7], net350[8], net350[9],
     net350[10], net350[11], net350[12], net350[13], net350[14],
     net350[15], net350[16], net350[17], net350[18], net350[19],
     net350[20], net350[21], net350[22], net350[23]}),
     .sp12_h_r_03({net351[0], net351[1], net351[2], net351[3],
     net351[4], net351[5], net351[6], net351[7], net351[8], net351[9],
     net351[10], net351[11], net351[12], net351[13], net351[14],
     net351[15], net351[16], net351[17], net351[18], net351[19],
     net351[20], net351[21], net351[22], net351[23]}),
     .sp12_h_r_02({net352[0], net352[1], net352[2], net352[3],
     net352[4], net352[5], net352[6], net352[7], net352[8], net352[9],
     net352[10], net352[11], net352[12], net352[13], net352[14],
     net352[15], net352[16], net352[17], net352[18], net352[19],
     net352[20], net352[21], net352[22], net352[23]}),
     .sp12_h_r_01({net353[0], net353[1], net353[2], net353[3],
     net353[4], net353[5], net353[6], net353[7], net353[8], net353[9],
     net353[10], net353[11], net353[12], net353[13], net353[14],
     net353[15], net353[16], net353[17], net353[18], net353[19],
     net353[20], net353[21], net353[22], net353[23]}),
     .sp4_v_b_01({net587[0], net587[1], net587[2], net587[3],
     net587[4], net587[5], net587[6], net587[7], net587[8], net587[9],
     net587[10], net587[11], net587[12], net587[13], net587[14],
     net587[15], net587[16], net587[17], net587[18], net587[19],
     net587[20], net587[21], net587[22], net587[23], net587[24],
     net587[25], net587[26], net587[27], net587[28], net587[29],
     net587[30], net587[31], net587[32], net587[33], net587[34],
     net587[35], net587[36], net587[37], net587[38], net587[39],
     net587[40], net587[41], net587[42], net587[43], net587[44],
     net587[45], net587[46], net587[47]}), .sp4_r_v_b_04({net355[0],
     net355[1], net355[2], net355[3], net355[4], net355[5], net355[6],
     net355[7], net355[8], net355[9], net355[10], net355[11],
     net355[12], net355[13], net355[14], net355[15], net355[16],
     net355[17], net355[18], net355[19], net355[20], net355[21],
     net355[22], net355[23], net355[24], net355[25], net355[26],
     net355[27], net355[28], net355[29], net355[30], net355[31],
     net355[32], net355[33], net355[34], net355[35], net355[36],
     net355[37], net355[38], net355[39], net355[40], net355[41],
     net355[42], net355[43], net355[44], net355[45], net355[46],
     net355[47]}), .sp4_r_v_b_03({net356[0], net356[1], net356[2],
     net356[3], net356[4], net356[5], net356[6], net356[7], net356[8],
     net356[9], net356[10], net356[11], net356[12], net356[13],
     net356[14], net356[15], net356[16], net356[17], net356[18],
     net356[19], net356[20], net356[21], net356[22], net356[23],
     net356[24], net356[25], net356[26], net356[27], net356[28],
     net356[29], net356[30], net356[31], net356[32], net356[33],
     net356[34], net356[35], net356[36], net356[37], net356[38],
     net356[39], net356[40], net356[41], net356[42], net356[43],
     net356[44], net356[45], net356[46], net356[47]}),
     .sp4_r_v_b_02({net357[0], net357[1], net357[2], net357[3],
     net357[4], net357[5], net357[6], net357[7], net357[8], net357[9],
     net357[10], net357[11], net357[12], net357[13], net357[14],
     net357[15], net357[16], net357[17], net357[18], net357[19],
     net357[20], net357[21], net357[22], net357[23], net357[24],
     net357[25], net357[26], net357[27], net357[28], net357[29],
     net357[30], net357[31], net357[32], net357[33], net357[34],
     net357[35], net357[36], net357[37], net357[38], net357[39],
     net357[40], net357[41], net357[42], net357[43], net357[44],
     net357[45], net357[46], net357[47]}), .sp4_r_v_b_01({net588[0],
     net588[1], net588[2], net588[3], net588[4], net588[5], net588[6],
     net588[7], net588[8], net588[9], net588[10], net588[11],
     net588[12], net588[13], net588[14], net588[15], net588[16],
     net588[17], net588[18], net588[19], net588[20], net588[21],
     net588[22], net588[23], net588[24], net588[25], net588[26],
     net588[27], net588[28], net588[29], net588[30], net588[31],
     net588[32], net588[33], net588[34], net588[35], net588[36],
     net588[37], net588[38], net588[39], net588[40], net588[41],
     net588[42], net588[43], net588[44], net588[45], net588[46],
     net588[47]}), .sp4_h_r_04({net359[0], net359[1], net359[2],
     net359[3], net359[4], net359[5], net359[6], net359[7], net359[8],
     net359[9], net359[10], net359[11], net359[12], net359[13],
     net359[14], net359[15], net359[16], net359[17], net359[18],
     net359[19], net359[20], net359[21], net359[22], net359[23],
     net359[24], net359[25], net359[26], net359[27], net359[28],
     net359[29], net359[30], net359[31], net359[32], net359[33],
     net359[34], net359[35], net359[36], net359[37], net359[38],
     net359[39], net359[40], net359[41], net359[42], net359[43],
     net359[44], net359[45], net359[46], net359[47]}),
     .sp4_h_r_03({net360[0], net360[1], net360[2], net360[3],
     net360[4], net360[5], net360[6], net360[7], net360[8], net360[9],
     net360[10], net360[11], net360[12], net360[13], net360[14],
     net360[15], net360[16], net360[17], net360[18], net360[19],
     net360[20], net360[21], net360[22], net360[23], net360[24],
     net360[25], net360[26], net360[27], net360[28], net360[29],
     net360[30], net360[31], net360[32], net360[33], net360[34],
     net360[35], net360[36], net360[37], net360[38], net360[39],
     net360[40], net360[41], net360[42], net360[43], net360[44],
     net360[45], net360[46], net360[47]}), .sp4_h_r_02({net361[0],
     net361[1], net361[2], net361[3], net361[4], net361[5], net361[6],
     net361[7], net361[8], net361[9], net361[10], net361[11],
     net361[12], net361[13], net361[14], net361[15], net361[16],
     net361[17], net361[18], net361[19], net361[20], net361[21],
     net361[22], net361[23], net361[24], net361[25], net361[26],
     net361[27], net361[28], net361[29], net361[30], net361[31],
     net361[32], net361[33], net361[34], net361[35], net361[36],
     net361[37], net361[38], net361[39], net361[40], net361[41],
     net361[42], net361[43], net361[44], net361[45], net361[46],
     net361[47]}), .sp4_h_r_01({net362[0], net362[1], net362[2],
     net362[3], net362[4], net362[5], net362[6], net362[7], net362[8],
     net362[9], net362[10], net362[11], net362[12], net362[13],
     net362[14], net362[15], net362[16], net362[17], net362[18],
     net362[19], net362[20], net362[21], net362[22], net362[23],
     net362[24], net362[25], net362[26], net362[27], net362[28],
     net362[29], net362[30], net362[31], net362[32], net362[33],
     net362[34], net362[35], net362[36], net362[37], net362[38],
     net362[39], net362[40], net362[41], net362[42], net362[43],
     net362[44], net362[45], net362[46], net362[47]}),
     .sp4_h_l_03({net474[0], net474[1], net474[2], net474[3],
     net474[4], net474[5], net474[6], net474[7], net474[8], net474[9],
     net474[10], net474[11], net474[12], net474[13], net474[14],
     net474[15], net474[16], net474[17], net474[18], net474[19],
     net474[20], net474[21], net474[22], net474[23], net474[24],
     net474[25], net474[26], net474[27], net474[28], net474[29],
     net474[30], net474[31], net474[32], net474[33], net474[34],
     net474[35], net474[36], net474[37], net474[38], net474[39],
     net474[40], net474[41], net474[42], net474[43], net474[44],
     net474[45], net474[46], net474[47]}), .sp4_h_l_02({net475[0],
     net475[1], net475[2], net475[3], net475[4], net475[5], net475[6],
     net475[7], net475[8], net475[9], net475[10], net475[11],
     net475[12], net475[13], net475[14], net475[15], net475[16],
     net475[17], net475[18], net475[19], net475[20], net475[21],
     net475[22], net475[23], net475[24], net475[25], net475[26],
     net475[27], net475[28], net475[29], net475[30], net475[31],
     net475[32], net475[33], net475[34], net475[35], net475[36],
     net475[37], net475[38], net475[39], net475[40], net475[41],
     net475[42], net475[43], net475[44], net475[45], net475[46],
     net475[47]}), .sp4_h_l_01({net476[0], net476[1], net476[2],
     net476[3], net476[4], net476[5], net476[6], net476[7], net476[8],
     net476[9], net476[10], net476[11], net476[12], net476[13],
     net476[14], net476[15], net476[16], net476[17], net476[18],
     net476[19], net476[20], net476[21], net476[22], net476[23],
     net476[24], net476[25], net476[26], net476[27], net476[28],
     net476[29], net476[30], net476[31], net476[32], net476[33],
     net476[34], net476[35], net476[36], net476[37], net476[38],
     net476[39], net476[40], net476[41], net476[42], net476[43],
     net476[44], net476[45], net476[46], net476[47]}), .bl(bl[125:72]),
     .bot_op_01({slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0], slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0]}), .sp12_h_l_01({net467[0],
     net467[1], net467[2], net467[3], net467[4], net467[5], net467[6],
     net467[7], net467[8], net467[9], net467[10], net467[11],
     net467[12], net467[13], net467[14], net467[15], net467[16],
     net467[17], net467[18], net467[19], net467[20], net467[21],
     net467[22], net467[23]}), .sp12_h_l_02({net466[0], net466[1],
     net466[2], net466[3], net466[4], net466[5], net466[6], net466[7],
     net466[8], net466[9], net466[10], net466[11], net466[12],
     net466[13], net466[14], net466[15], net466[16], net466[17],
     net466[18], net466[19], net466[20], net466[21], net466[22],
     net466[23]}), .sp12_h_l_03({net465[0], net465[1], net465[2],
     net465[3], net465[4], net465[5], net465[6], net465[7], net465[8],
     net465[9], net465[10], net465[11], net465[12], net465[13],
     net465[14], net465[15], net465[16], net465[17], net465[18],
     net465[19], net465[20], net465[21], net465[22], net465[23]}),
     .sp12_h_l_04({net464[0], net464[1], net464[2], net464[3],
     net464[4], net464[5], net464[6], net464[7], net464[8], net464[9],
     net464[10], net464[11], net464[12], net464[13], net464[14],
     net464[15], net464[16], net464[17], net464[18], net464[19],
     net464[20], net464[21], net464[22], net464[23]}),
     .sp4_v_b_04({net469[0], net469[1], net469[2], net469[3],
     net469[4], net469[5], net469[6], net469[7], net469[8], net469[9],
     net469[10], net469[11], net469[12], net469[13], net469[14],
     net469[15], net469[16], net469[17], net469[18], net469[19],
     net469[20], net469[21], net469[22], net469[23], net469[24],
     net469[25], net469[26], net469[27], net469[28], net469[29],
     net469[30], net469[31], net469[32], net469[33], net469[34],
     net469[35], net469[36], net469[37], net469[38], net469[39],
     net469[40], net469[41], net469[42], net469[43], net469[44],
     net469[45], net469[46], net469[47]}), .sp4_v_b_03({net470[0],
     net470[1], net470[2], net470[3], net470[4], net470[5], net470[6],
     net470[7], net470[8], net470[9], net470[10], net470[11],
     net470[12], net470[13], net470[14], net470[15], net470[16],
     net470[17], net470[18], net470[19], net470[20], net470[21],
     net470[22], net470[23], net470[24], net470[25], net470[26],
     net470[27], net470[28], net470[29], net470[30], net470[31],
     net470[32], net470[33], net470[34], net470[35], net470[36],
     net470[37], net470[38], net470[39], net470[40], net470[41],
     net470[42], net470[43], net470[44], net470[45], net470[46],
     net470[47]}), .sp4_v_b_02({net471[0], net471[1], net471[2],
     net471[3], net471[4], net471[5], net471[6], net471[7], net471[8],
     net471[9], net471[10], net471[11], net471[12], net471[13],
     net471[14], net471[15], net471[16], net471[17], net471[18],
     net471[19], net471[20], net471[21], net471[22], net471[23],
     net471[24], net471[25], net471[26], net471[27], net471[28],
     net471[29], net471[30], net471[31], net471[32], net471[33],
     net471[34], net471[35], net471[36], net471[37], net471[38],
     net471[39], net471[40], net471[41], net471[42], net471[43],
     net471[44], net471[45], net471[46], net471[47]}),
     .bnr_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .top_op_04(top_op_02_04[7:0]),
     .sp12_v_t_04(sp12_v_t_02_04[23:0]), .tnl_op_04(tnl_op_02_04[7:0]),
     .pgate(pgate_l[79:16]), .reset_b(reset_b_l[79:16]),
     .wl(wl_l[79:16]), .tnr_op_04(tnr_op_02_04[7:0]),
     .sp4_v_t_04(sp4_v_t_02_04[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_02_04), .sp12_v_b_01({net575[0], net575[1],
     net575[2], net575[3], net575[4], net575[5], net575[6], net575[7],
     net575[8], net575[9], net575[10], net575[11], net575[12],
     net575[13], net575[14], net575[15], net575[16], net575[17],
     net575[18], net575[19], net575[20], net575[21], net575[22],
     net575[23]}), .glb_netwk(glb_in_2[7:0]));
lt_1x4_bot_ice384 I806 ( .rgt_op_03(rgt_op_03_03[7:0]),
     .slf_op_02(slf_op_03_02[7:0]), .rgt_op_02(rgt_op_03_02[7:0]),
     .rgt_op_01(rgt_op_03_01[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(slf_op_02_04[7:0]), .lft_op_03({net445[0], net445[1],
     net445[2], net445[3], net445[4], net445[5], net445[6],
     net445[7]}), .lft_op_02({net447[0], net447[1], net447[2],
     net447[3], net447[4], net447[5], net447[6], net447[7]}),
     .lft_op_01({net590[0], net590[1], net590[2], net590[3], net590[4],
     net590[5], net590[6], net590[7]}), .rgt_op_04(rgt_op_03_04[7:0]),
     .carry_in(tiegnd_bl), .bnl_op_01({slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0],
     slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0]}), .slf_op_04(slf_op_03_04[7:0]),
     .slf_op_03(slf_op_03_03[7:0]), .slf_op_01(slf_op_03_01[7:0]),
     .sp4_h_l_04({net359[0], net359[1], net359[2], net359[3],
     net359[4], net359[5], net359[6], net359[7], net359[8], net359[9],
     net359[10], net359[11], net359[12], net359[13], net359[14],
     net359[15], net359[16], net359[17], net359[18], net359[19],
     net359[20], net359[21], net359[22], net359[23], net359[24],
     net359[25], net359[26], net359[27], net359[28], net359[29],
     net359[30], net359[31], net359[32], net359[33], net359[34],
     net359[35], net359[36], net359[37], net359[38], net359[39],
     net359[40], net359[41], net359[42], net359[43], net359[44],
     net359[45], net359[46], net359[47]}), .carry_out(carry_out_03_04),
     .vdd_cntl(vdd_cntl_l[79:16]), .sp12_h_r_04(sp12_h_r_03_04[23:0]),
     .sp12_h_r_03(sp12_h_r_03_03[23:0]),
     .sp12_h_r_02(sp12_h_r_03_02[23:0]),
     .sp12_h_r_01(sp12_h_r_03_01[23:0]), .sp4_v_b_01({net588[0],
     net588[1], net588[2], net588[3], net588[4], net588[5], net588[6],
     net588[7], net588[8], net588[9], net588[10], net588[11],
     net588[12], net588[13], net588[14], net588[15], net588[16],
     net588[17], net588[18], net588[19], net588[20], net588[21],
     net588[22], net588[23], net588[24], net588[25], net588[26],
     net588[27], net588[28], net588[29], net588[30], net588[31],
     net588[32], net588[33], net588[34], net588[35], net588[36],
     net588[37], net588[38], net588[39], net588[40], net588[41],
     net588[42], net588[43], net588[44], net588[45], net588[46],
     net588[47]}), .sp4_r_v_b_04(sp4_r_v_b_03_04[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_03_03[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_03_02[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_03_01[47:0]),
     .sp4_h_r_04(sp4_h_r_03_04[47:0]),
     .sp4_h_r_03(sp4_h_r_03_03[47:0]),
     .sp4_h_r_02(sp4_h_r_03_02[47:0]),
     .sp4_h_r_01(sp4_h_r_03_01[47:0]), .sp4_h_l_03({net360[0],
     net360[1], net360[2], net360[3], net360[4], net360[5], net360[6],
     net360[7], net360[8], net360[9], net360[10], net360[11],
     net360[12], net360[13], net360[14], net360[15], net360[16],
     net360[17], net360[18], net360[19], net360[20], net360[21],
     net360[22], net360[23], net360[24], net360[25], net360[26],
     net360[27], net360[28], net360[29], net360[30], net360[31],
     net360[32], net360[33], net360[34], net360[35], net360[36],
     net360[37], net360[38], net360[39], net360[40], net360[41],
     net360[42], net360[43], net360[44], net360[45], net360[46],
     net360[47]}), .sp4_h_l_02({net361[0], net361[1], net361[2],
     net361[3], net361[4], net361[5], net361[6], net361[7], net361[8],
     net361[9], net361[10], net361[11], net361[12], net361[13],
     net361[14], net361[15], net361[16], net361[17], net361[18],
     net361[19], net361[20], net361[21], net361[22], net361[23],
     net361[24], net361[25], net361[26], net361[27], net361[28],
     net361[29], net361[30], net361[31], net361[32], net361[33],
     net361[34], net361[35], net361[36], net361[37], net361[38],
     net361[39], net361[40], net361[41], net361[42], net361[43],
     net361[44], net361[45], net361[46], net361[47]}),
     .sp4_h_l_01({net362[0], net362[1], net362[2], net362[3],
     net362[4], net362[5], net362[6], net362[7], net362[8], net362[9],
     net362[10], net362[11], net362[12], net362[13], net362[14],
     net362[15], net362[16], net362[17], net362[18], net362[19],
     net362[20], net362[21], net362[22], net362[23], net362[24],
     net362[25], net362[26], net362[27], net362[28], net362[29],
     net362[30], net362[31], net362[32], net362[33], net362[34],
     net362[35], net362[36], net362[37], net362[38], net362[39],
     net362[40], net362[41], net362[42], net362[43], net362[44],
     net362[45], net362[46], net362[47]}), .bl(bl[179:126]),
     .bot_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .sp12_h_l_01({net353[0],
     net353[1], net353[2], net353[3], net353[4], net353[5], net353[6],
     net353[7], net353[8], net353[9], net353[10], net353[11],
     net353[12], net353[13], net353[14], net353[15], net353[16],
     net353[17], net353[18], net353[19], net353[20], net353[21],
     net353[22], net353[23]}), .sp12_h_l_02({net352[0], net352[1],
     net352[2], net352[3], net352[4], net352[5], net352[6], net352[7],
     net352[8], net352[9], net352[10], net352[11], net352[12],
     net352[13], net352[14], net352[15], net352[16], net352[17],
     net352[18], net352[19], net352[20], net352[21], net352[22],
     net352[23]}), .sp12_h_l_03({net351[0], net351[1], net351[2],
     net351[3], net351[4], net351[5], net351[6], net351[7], net351[8],
     net351[9], net351[10], net351[11], net351[12], net351[13],
     net351[14], net351[15], net351[16], net351[17], net351[18],
     net351[19], net351[20], net351[21], net351[22], net351[23]}),
     .sp12_h_l_04({net350[0], net350[1], net350[2], net350[3],
     net350[4], net350[5], net350[6], net350[7], net350[8], net350[9],
     net350[10], net350[11], net350[12], net350[13], net350[14],
     net350[15], net350[16], net350[17], net350[18], net350[19],
     net350[20], net350[21], net350[22], net350[23]}),
     .sp4_v_b_04({net355[0], net355[1], net355[2], net355[3],
     net355[4], net355[5], net355[6], net355[7], net355[8], net355[9],
     net355[10], net355[11], net355[12], net355[13], net355[14],
     net355[15], net355[16], net355[17], net355[18], net355[19],
     net355[20], net355[21], net355[22], net355[23], net355[24],
     net355[25], net355[26], net355[27], net355[28], net355[29],
     net355[30], net355[31], net355[32], net355[33], net355[34],
     net355[35], net355[36], net355[37], net355[38], net355[39],
     net355[40], net355[41], net355[42], net355[43], net355[44],
     net355[45], net355[46], net355[47]}), .sp4_v_b_03({net356[0],
     net356[1], net356[2], net356[3], net356[4], net356[5], net356[6],
     net356[7], net356[8], net356[9], net356[10], net356[11],
     net356[12], net356[13], net356[14], net356[15], net356[16],
     net356[17], net356[18], net356[19], net356[20], net356[21],
     net356[22], net356[23], net356[24], net356[25], net356[26],
     net356[27], net356[28], net356[29], net356[30], net356[31],
     net356[32], net356[33], net356[34], net356[35], net356[36],
     net356[37], net356[38], net356[39], net356[40], net356[41],
     net356[42], net356[43], net356[44], net356[45], net356[46],
     net356[47]}), .sp4_v_b_02({net357[0], net357[1], net357[2],
     net357[3], net357[4], net357[5], net357[6], net357[7], net357[8],
     net357[9], net357[10], net357[11], net357[12], net357[13],
     net357[14], net357[15], net357[16], net357[17], net357[18],
     net357[19], net357[20], net357[21], net357[22], net357[23],
     net357[24], net357[25], net357[26], net357[27], net357[28],
     net357[29], net357[30], net357[31], net357[32], net357[33],
     net357[34], net357[35], net357[36], net357[37], net357[38],
     net357[39], net357[40], net357[41], net357[42], net357[43],
     net357[44], net357[45], net357[46], net357[47]}),
     .bnr_op_01({bnr_op_03_01[3], bnr_op_03_01[2], bnr_op_03_01[1],
     bnr_op_03_01[0], bnr_op_03_01[3], bnr_op_03_01[2],
     bnr_op_03_01[1], bnr_op_03_01[0]}), .top_op_04(top_op_03_04[7:0]),
     .sp12_v_t_04(sp12_v_t_03_04[23:0]), .tnl_op_04(tnl_op_03_04[7:0]),
     .pgate(pgate_l[79:16]), .reset_b(reset_b_l[79:16]),
     .wl(wl_l[79:16]), .tnr_op_04(tnr_op_03_04[7:0]),
     .sp4_v_t_04(sp4_v_t_03_04[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_03_04), .sp12_v_b_01({net583[0], net583[1],
     net583[2], net583[3], net583[4], net583[5], net583[6], net583[7],
     net583[8], net583[9], net583[10], net583[11], net583[12],
     net583[13], net583[14], net583[15], net583[16], net583[17],
     net583[18], net583[19], net583[20], net583[21], net583[22],
     net583[23]}), .glb_netwk(glb_in_3[7:0]));
lt_1x4_bot_ice384 I804 ( .rgt_op_03({net445[0], net445[1], net445[2],
     net445[3], net445[4], net445[5], net445[6], net445[7]}),
     .slf_op_02({net518[0], net518[1], net518[2], net518[3], net518[4],
     net518[5], net518[6], net518[7]}), .rgt_op_02({net447[0],
     net447[1], net447[2], net447[3], net447[4], net447[5], net447[6],
     net447[7]}), .rgt_op_01({net590[0], net590[1], net590[2],
     net590[3], net590[4], net590[5], net590[6], net590[7]}),
     .purst(purst), .prog(prog), .lft_op_04({slf_op_00_04[3],
     slf_op_00_04[2], slf_op_00_04[1], slf_op_00_04[0],
     slf_op_00_04[3], slf_op_00_04[2], slf_op_00_04[1],
     slf_op_00_04[0]}), .lft_op_03({slf_op_00_03[3], slf_op_00_03[2],
     slf_op_00_03[1], slf_op_00_03[0], slf_op_00_03[3],
     slf_op_00_03[2], slf_op_00_03[1], slf_op_00_03[0]}),
     .lft_op_02({slf_op_00_02[3], slf_op_00_02[2], slf_op_00_02[1],
     slf_op_00_02[0], slf_op_00_02[3], slf_op_00_02[2],
     slf_op_00_02[1], slf_op_00_02[0]}), .lft_op_01({slf_op_00_01[3],
     slf_op_00_01[2], slf_op_00_01[1], slf_op_00_01[0],
     slf_op_00_01[3], slf_op_00_01[2], slf_op_00_01[1],
     slf_op_00_01[0]}), .rgt_op_04(slf_op_02_04[7:0]),
     .carry_in(tiegnd_bl), .bnl_op_01({tiegnd_bl, tiegnd_bl, tiegnd_bl,
     tiegnd_bl, tiegnd_bl, tiegnd_bl, tiegnd_bl, tiegnd_bl}),
     .slf_op_04(slf_op_01_04[7:0]), .slf_op_03({net526[0], net526[1],
     net526[2], net526[3], net526[4], net526[5], net526[6],
     net526[7]}), .slf_op_01({net589[0], net589[1], net589[2],
     net589[3], net589[4], net589[5], net589[6], net589[7]}),
     .sp4_h_l_04({net522[0], net522[1], net522[2], net522[3],
     net522[4], net522[5], net522[6], net522[7], net522[8], net522[9],
     net522[10], net522[11], net522[12], net522[13], net522[14],
     net522[15], net522[16], net522[17], net522[18], net522[19],
     net522[20], net522[21], net522[22], net522[23], net522[24],
     net522[25], net522[26], net522[27], net522[28], net522[29],
     net522[30], net522[31], net522[32], net522[33], net522[34],
     net522[35], net522[36], net522[37], net522[38], net522[39],
     net522[40], net522[41], net522[42], net522[43], net522[44],
     net522[45], net522[46], net522[47]}), .carry_out(carry_out_01_04),
     .vdd_cntl(vdd_cntl_l[79:16]), .sp12_h_r_04({net464[0], net464[1],
     net464[2], net464[3], net464[4], net464[5], net464[6], net464[7],
     net464[8], net464[9], net464[10], net464[11], net464[12],
     net464[13], net464[14], net464[15], net464[16], net464[17],
     net464[18], net464[19], net464[20], net464[21], net464[22],
     net464[23]}), .sp12_h_r_03({net465[0], net465[1], net465[2],
     net465[3], net465[4], net465[5], net465[6], net465[7], net465[8],
     net465[9], net465[10], net465[11], net465[12], net465[13],
     net465[14], net465[15], net465[16], net465[17], net465[18],
     net465[19], net465[20], net465[21], net465[22], net465[23]}),
     .sp12_h_r_02({net466[0], net466[1], net466[2], net466[3],
     net466[4], net466[5], net466[6], net466[7], net466[8], net466[9],
     net466[10], net466[11], net466[12], net466[13], net466[14],
     net466[15], net466[16], net466[17], net466[18], net466[19],
     net466[20], net466[21], net466[22], net466[23]}),
     .sp12_h_r_01({net467[0], net467[1], net467[2], net467[3],
     net467[4], net467[5], net467[6], net467[7], net467[8], net467[9],
     net467[10], net467[11], net467[12], net467[13], net467[14],
     net467[15], net467[16], net467[17], net467[18], net467[19],
     net467[20], net467[21], net467[22], net467[23]}),
     .sp4_v_b_01({net582[0], net582[1], net582[2], net582[3],
     net582[4], net582[5], net582[6], net582[7], net582[8], net582[9],
     net582[10], net582[11], net582[12], net582[13], net582[14],
     net582[15], net582[16], net582[17], net582[18], net582[19],
     net582[20], net582[21], net582[22], net582[23], net582[24],
     net582[25], net582[26], net582[27], net582[28], net582[29],
     net582[30], net582[31], net582[32], net582[33], net582[34],
     net582[35], net582[36], net582[37], net582[38], net582[39],
     net582[40], net582[41], net582[42], net582[43], net582[44],
     net582[45], net582[46], net582[47]}), .sp4_r_v_b_04({net469[0],
     net469[1], net469[2], net469[3], net469[4], net469[5], net469[6],
     net469[7], net469[8], net469[9], net469[10], net469[11],
     net469[12], net469[13], net469[14], net469[15], net469[16],
     net469[17], net469[18], net469[19], net469[20], net469[21],
     net469[22], net469[23], net469[24], net469[25], net469[26],
     net469[27], net469[28], net469[29], net469[30], net469[31],
     net469[32], net469[33], net469[34], net469[35], net469[36],
     net469[37], net469[38], net469[39], net469[40], net469[41],
     net469[42], net469[43], net469[44], net469[45], net469[46],
     net469[47]}), .sp4_r_v_b_03({net470[0], net470[1], net470[2],
     net470[3], net470[4], net470[5], net470[6], net470[7], net470[8],
     net470[9], net470[10], net470[11], net470[12], net470[13],
     net470[14], net470[15], net470[16], net470[17], net470[18],
     net470[19], net470[20], net470[21], net470[22], net470[23],
     net470[24], net470[25], net470[26], net470[27], net470[28],
     net470[29], net470[30], net470[31], net470[32], net470[33],
     net470[34], net470[35], net470[36], net470[37], net470[38],
     net470[39], net470[40], net470[41], net470[42], net470[43],
     net470[44], net470[45], net470[46], net470[47]}),
     .sp4_r_v_b_02({net471[0], net471[1], net471[2], net471[3],
     net471[4], net471[5], net471[6], net471[7], net471[8], net471[9],
     net471[10], net471[11], net471[12], net471[13], net471[14],
     net471[15], net471[16], net471[17], net471[18], net471[19],
     net471[20], net471[21], net471[22], net471[23], net471[24],
     net471[25], net471[26], net471[27], net471[28], net471[29],
     net471[30], net471[31], net471[32], net471[33], net471[34],
     net471[35], net471[36], net471[37], net471[38], net471[39],
     net471[40], net471[41], net471[42], net471[43], net471[44],
     net471[45], net471[46], net471[47]}), .sp4_r_v_b_01({net587[0],
     net587[1], net587[2], net587[3], net587[4], net587[5], net587[6],
     net587[7], net587[8], net587[9], net587[10], net587[11],
     net587[12], net587[13], net587[14], net587[15], net587[16],
     net587[17], net587[18], net587[19], net587[20], net587[21],
     net587[22], net587[23], net587[24], net587[25], net587[26],
     net587[27], net587[28], net587[29], net587[30], net587[31],
     net587[32], net587[33], net587[34], net587[35], net587[36],
     net587[37], net587[38], net587[39], net587[40], net587[41],
     net587[42], net587[43], net587[44], net587[45], net587[46],
     net587[47]}), .sp4_h_r_04({net473[0], net473[1], net473[2],
     net473[3], net473[4], net473[5], net473[6], net473[7], net473[8],
     net473[9], net473[10], net473[11], net473[12], net473[13],
     net473[14], net473[15], net473[16], net473[17], net473[18],
     net473[19], net473[20], net473[21], net473[22], net473[23],
     net473[24], net473[25], net473[26], net473[27], net473[28],
     net473[29], net473[30], net473[31], net473[32], net473[33],
     net473[34], net473[35], net473[36], net473[37], net473[38],
     net473[39], net473[40], net473[41], net473[42], net473[43],
     net473[44], net473[45], net473[46], net473[47]}),
     .sp4_h_r_03({net474[0], net474[1], net474[2], net474[3],
     net474[4], net474[5], net474[6], net474[7], net474[8], net474[9],
     net474[10], net474[11], net474[12], net474[13], net474[14],
     net474[15], net474[16], net474[17], net474[18], net474[19],
     net474[20], net474[21], net474[22], net474[23], net474[24],
     net474[25], net474[26], net474[27], net474[28], net474[29],
     net474[30], net474[31], net474[32], net474[33], net474[34],
     net474[35], net474[36], net474[37], net474[38], net474[39],
     net474[40], net474[41], net474[42], net474[43], net474[44],
     net474[45], net474[46], net474[47]}), .sp4_h_r_02({net475[0],
     net475[1], net475[2], net475[3], net475[4], net475[5], net475[6],
     net475[7], net475[8], net475[9], net475[10], net475[11],
     net475[12], net475[13], net475[14], net475[15], net475[16],
     net475[17], net475[18], net475[19], net475[20], net475[21],
     net475[22], net475[23], net475[24], net475[25], net475[26],
     net475[27], net475[28], net475[29], net475[30], net475[31],
     net475[32], net475[33], net475[34], net475[35], net475[36],
     net475[37], net475[38], net475[39], net475[40], net475[41],
     net475[42], net475[43], net475[44], net475[45], net475[46],
     net475[47]}), .sp4_h_r_01({net476[0], net476[1], net476[2],
     net476[3], net476[4], net476[5], net476[6], net476[7], net476[8],
     net476[9], net476[10], net476[11], net476[12], net476[13],
     net476[14], net476[15], net476[16], net476[17], net476[18],
     net476[19], net476[20], net476[21], net476[22], net476[23],
     net476[24], net476[25], net476[26], net476[27], net476[28],
     net476[29], net476[30], net476[31], net476[32], net476[33],
     net476[34], net476[35], net476[36], net476[37], net476[38],
     net476[39], net476[40], net476[41], net476[42], net476[43],
     net476[44], net476[45], net476[46], net476[47]}),
     .sp4_h_l_03({net521[0], net521[1], net521[2], net521[3],
     net521[4], net521[5], net521[6], net521[7], net521[8], net521[9],
     net521[10], net521[11], net521[12], net521[13], net521[14],
     net521[15], net521[16], net521[17], net521[18], net521[19],
     net521[20], net521[21], net521[22], net521[23], net521[24],
     net521[25], net521[26], net521[27], net521[28], net521[29],
     net521[30], net521[31], net521[32], net521[33], net521[34],
     net521[35], net521[36], net521[37], net521[38], net521[39],
     net521[40], net521[41], net521[42], net521[43], net521[44],
     net521[45], net521[46], net521[47]}), .sp4_h_l_02({net523[0],
     net523[1], net523[2], net523[3], net523[4], net523[5], net523[6],
     net523[7], net523[8], net523[9], net523[10], net523[11],
     net523[12], net523[13], net523[14], net523[15], net523[16],
     net523[17], net523[18], net523[19], net523[20], net523[21],
     net523[22], net523[23], net523[24], net523[25], net523[26],
     net523[27], net523[28], net523[29], net523[30], net523[31],
     net523[32], net523[33], net523[34], net523[35], net523[36],
     net523[37], net523[38], net523[39], net523[40], net523[41],
     net523[42], net523[43], net523[44], net523[45], net523[46],
     net523[47]}), .sp4_h_l_01({net524[0], net524[1], net524[2],
     net524[3], net524[4], net524[5], net524[6], net524[7], net524[8],
     net524[9], net524[10], net524[11], net524[12], net524[13],
     net524[14], net524[15], net524[16], net524[17], net524[18],
     net524[19], net524[20], net524[21], net524[22], net524[23],
     net524[24], net524[25], net524[26], net524[27], net524[28],
     net524[29], net524[30], net524[31], net524[32], net524[33],
     net524[34], net524[35], net524[36], net524[37], net524[38],
     net524[39], net524[40], net524[41], net524[42], net524[43],
     net524[44], net524[45], net524[46], net524[47]}), .bl(bl[71:18]),
     .bot_op_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}), .sp12_h_l_01({net539[0],
     net539[1], net539[2], net539[3], net539[4], net539[5], net539[6],
     net539[7], net539[8], net539[9], net539[10], net539[11],
     net539[12], net539[13], net539[14], net539[15], net539[16],
     net539[17], net539[18], net539[19], net539[20], net539[21],
     net539[22], net539[23]}), .sp12_h_l_02({net537[0], net537[1],
     net537[2], net537[3], net537[4], net537[5], net537[6], net537[7],
     net537[8], net537[9], net537[10], net537[11], net537[12],
     net537[13], net537[14], net537[15], net537[16], net537[17],
     net537[18], net537[19], net537[20], net537[21], net537[22],
     net537[23]}), .sp12_h_l_03({net541[0], net541[1], net541[2],
     net541[3], net541[4], net541[5], net541[6], net541[7], net541[8],
     net541[9], net541[10], net541[11], net541[12], net541[13],
     net541[14], net541[15], net541[16], net541[17], net541[18],
     net541[19], net541[20], net541[21], net541[22], net541[23]}),
     .sp12_h_l_04({net538[0], net538[1], net538[2], net538[3],
     net538[4], net538[5], net538[6], net538[7], net538[8], net538[9],
     net538[10], net538[11], net538[12], net538[13], net538[14],
     net538[15], net538[16], net538[17], net538[18], net538[19],
     net538[20], net538[21], net538[22], net538[23]}),
     .sp4_v_b_04({net486[0], net486[1], net486[2], net486[3],
     net486[4], net486[5], net486[6], net486[7], net486[8], net486[9],
     net486[10], net486[11], net486[12], net486[13], net486[14],
     net486[15], net486[16], net486[17], net486[18], net486[19],
     net486[20], net486[21], net486[22], net486[23], net486[24],
     net486[25], net486[26], net486[27], net486[28], net486[29],
     net486[30], net486[31], net486[32], net486[33], net486[34],
     net486[35], net486[36], net486[37], net486[38], net486[39],
     net486[40], net486[41], net486[42], net486[43], net486[44],
     net486[45], net486[46], net486[47]}), .sp4_v_b_03({net487[0],
     net487[1], net487[2], net487[3], net487[4], net487[5], net487[6],
     net487[7], net487[8], net487[9], net487[10], net487[11],
     net487[12], net487[13], net487[14], net487[15], net487[16],
     net487[17], net487[18], net487[19], net487[20], net487[21],
     net487[22], net487[23], net487[24], net487[25], net487[26],
     net487[27], net487[28], net487[29], net487[30], net487[31],
     net487[32], net487[33], net487[34], net487[35], net487[36],
     net487[37], net487[38], net487[39], net487[40], net487[41],
     net487[42], net487[43], net487[44], net487[45], net487[46],
     net487[47]}), .sp4_v_b_02({net608[0], net608[1], net608[2],
     net608[3], net608[4], net608[5], net608[6], net608[7], net608[8],
     net608[9], net608[10], net608[11], net608[12], net608[13],
     net608[14], net608[15], net608[16], net608[17], net608[18],
     net608[19], net608[20], net608[21], net608[22], net608[23],
     net608[24], net608[25], net608[26], net608[27], net608[28],
     net608[29], net608[30], net608[31], net608[32], net608[33],
     net608[34], net608[35], net608[36], net608[37], net608[38],
     net608[39], net608[40], net608[41], net608[42], net608[43],
     net608[44], net608[45], net608[46], net608[47]}),
     .bnr_op_01({slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0], slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0]}), .top_op_04(top_op_01_04[7:0]),
     .sp12_v_t_04(sp12_v_t_01_04[23:0]), .tnl_op_04(tnl_op_01_04[7:0]),
     .pgate(pgate_l[79:16]), .reset_b(reset_b_l[79:16]),
     .wl(wl_l[79:16]), .tnr_op_04(tnr_op_01_04[7:0]),
     .sp4_v_t_04(sp4_v_t_01_04[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_01_04), .sp12_v_b_01({net561[0], net561[1],
     net561[2], net561[3], net561[4], net561[5], net561[6], net561[7],
     net561[8], net561[9], net561[10], net561[11], net561[12],
     net561[13], net561[14], net561[15], net561[16], net561[17],
     net561[18], net561[19], net561[20], net561[21], net561[22],
     net561[23]}), .glb_netwk(glb_in_1[7:0]));
io_lft_bot_1x4_ice384 I803 ( .shift(net502), .bs_en(net503),
     .mode(net504), .sdi(net505), .hiz_b(net506), .prog(prog),
     .hold(hold_l_b), .update(net509), .r(net510),
     .slf_op_01(slf_op_00_01[3:0]), .slf_op_02(slf_op_00_02[3:0]),
     .sdo(net513), .bl({bl[0], bl[1], bl[2], bl[3], bl[4], bl[5],
     bl[6], bl[7], bl[8], bl[9], bl[10], bl[11], bl[12], bl[13],
     bl[14], bl[15], bl[16], bl[17]}), .sp4_v_b_00_01({net515[0],
     net515[1], net515[2], net515[3], net515[4], net515[5], net515[6],
     net515[7], net515[8], net515[9], net515[10], net515[11],
     net515[12], net515[13], net515[14], net515[15]}), .tclk(net516),
     .reset_b(reset_b_l[79:16]), .rgt_op_02({net518[0], net518[1],
     net518[2], net518[3], net518[4], net518[5], net518[6],
     net518[7]}), .slf_op_04(slf_op_00_04[3:0]),
     .slf_op_03(slf_op_00_03[3:0]), .SP4_h_l_03({net521[0], net521[1],
     net521[2], net521[3], net521[4], net521[5], net521[6], net521[7],
     net521[8], net521[9], net521[10], net521[11], net521[12],
     net521[13], net521[14], net521[15], net521[16], net521[17],
     net521[18], net521[19], net521[20], net521[21], net521[22],
     net521[23], net521[24], net521[25], net521[26], net521[27],
     net521[28], net521[29], net521[30], net521[31], net521[32],
     net521[33], net521[34], net521[35], net521[36], net521[37],
     net521[38], net521[39], net521[40], net521[41], net521[42],
     net521[43], net521[44], net521[45], net521[46], net521[47]}),
     .SP4_h_l_04({net522[0], net522[1], net522[2], net522[3],
     net522[4], net522[5], net522[6], net522[7], net522[8], net522[9],
     net522[10], net522[11], net522[12], net522[13], net522[14],
     net522[15], net522[16], net522[17], net522[18], net522[19],
     net522[20], net522[21], net522[22], net522[23], net522[24],
     net522[25], net522[26], net522[27], net522[28], net522[29],
     net522[30], net522[31], net522[32], net522[33], net522[34],
     net522[35], net522[36], net522[37], net522[38], net522[39],
     net522[40], net522[41], net522[42], net522[43], net522[44],
     net522[45], net522[46], net522[47]}), .SP4_h_l_02({net523[0],
     net523[1], net523[2], net523[3], net523[4], net523[5], net523[6],
     net523[7], net523[8], net523[9], net523[10], net523[11],
     net523[12], net523[13], net523[14], net523[15], net523[16],
     net523[17], net523[18], net523[19], net523[20], net523[21],
     net523[22], net523[23], net523[24], net523[25], net523[26],
     net523[27], net523[28], net523[29], net523[30], net523[31],
     net523[32], net523[33], net523[34], net523[35], net523[36],
     net523[37], net523[38], net523[39], net523[40], net523[41],
     net523[42], net523[43], net523[44], net523[45], net523[46],
     net523[47]}), .SP4_h_l_01({net524[0], net524[1], net524[2],
     net524[3], net524[4], net524[5], net524[6], net524[7], net524[8],
     net524[9], net524[10], net524[11], net524[12], net524[13],
     net524[14], net524[15], net524[16], net524[17], net524[18],
     net524[19], net524[20], net524[21], net524[22], net524[23],
     net524[24], net524[25], net524[26], net524[27], net524[28],
     net524[29], net524[30], net524[31], net524[32], net524[33],
     net524[34], net524[35], net524[36], net524[37], net524[38],
     net524[39], net524[40], net524[41], net524[42], net524[43],
     net524[44], net524[45], net524[46], net524[47]}),
     .padin(padin_l_b[7:0]), .rgt_op_03({net526[0], net526[1],
     net526[2], net526[3], net526[4], net526[5], net526[6],
     net526[7]}), .rgt_op_01({net589[0], net589[1], net589[2],
     net589[3], net589[4], net589[5], net589[6], net589[7]}),
     .pado(pado_l_b[7:0]), .padeb(padeb_l_b[7:0]), .cf_l(cf_l[95:0]),
     .vdd_cntl(vdd_cntl_l[79:16]), .pgate(pgate_l[79:16]),
     .wl(wl_l[79:16]),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .tclk_o(net535), .ceb(net536), .SP12_h_l_02({net537[0], net537[1],
     net537[2], net537[3], net537[4], net537[5], net537[6], net537[7],
     net537[8], net537[9], net537[10], net537[11], net537[12],
     net537[13], net537[14], net537[15], net537[16], net537[17],
     net537[18], net537[19], net537[20], net537[21], net537[22],
     net537[23]}), .SP12_h_l_04({net538[0], net538[1], net538[2],
     net538[3], net538[4], net538[5], net538[6], net538[7], net538[8],
     net538[9], net538[10], net538[11], net538[12], net538[13],
     net538[14], net538[15], net538[16], net538[17], net538[18],
     net538[19], net538[20], net538[21], net538[22], net538[23]}),
     .SP12_h_l_01({net539[0], net539[1], net539[2], net539[3],
     net539[4], net539[5], net539[6], net539[7], net539[8], net539[9],
     net539[10], net539[11], net539[12], net539[13], net539[14],
     net539[15], net539[16], net539[17], net539[18], net539[19],
     net539[20], net539[21], net539[22], net539[23]}),
     .fabric_out_03(fabric_out_00_03), .SP12_h_l_03({net541[0],
     net541[1], net541[2], net541[3], net541[4], net541[5], net541[6],
     net541[7], net541[8], net541[9], net541[10], net541[11],
     net541[12], net541[13], net541[14], net541[15], net541[16],
     net541[17], net541[18], net541[19], net541[20], net541[21],
     net541[22], net541[23]}), .tnr_op_04(tnr_op_00_04[7:0]),
     .fabric_out_04(fabric_out_00_04), .glb_netwk(glb_in_0[7:0]),
     .last_rsr(last_rsr[0]), .rgt_op_04(slf_op_01_04[7:0]),
     .bnr_op_00_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}),
     .sp4_v_t_04(sp4_v_t_00_04[15:0]));
io_bot_lft_1x3_ice384 I802 ( .wl_l({wl_l[1], wl_l[0], wl_l[2], wl_l[3],
     wl_l[5], wl_l[4], wl_l[6], wl_l[7], wl_l[9], wl_l[8], wl_l[10],
     wl_l[11], wl_l[13], wl_l[12], wl_l[14], wl_l[15]}),
     .slf_op_01_00(slf_op_01_00[3:0]), .vdd_cntl_l({vdd_cntl_l[1],
     vdd_cntl_l[0], vdd_cntl_l[2], vdd_cntl_l[3], vdd_cntl_l[5],
     vdd_cntl_l[4], vdd_cntl_l[6], vdd_cntl_l[7], vdd_cntl_l[9],
     vdd_cntl_l[8], vdd_cntl_l[10], vdd_cntl_l[11], vdd_cntl_l[13],
     vdd_cntl_l[12], vdd_cntl_l[14], vdd_cntl_l[15]}),
     .update_i(net509), .tclk_i(net535), .shift_i(net502),
     .sdi(net513), .reset_l({reset_b_l[1], reset_b_l[0], reset_b_l[2],
     reset_b_l[3], reset_b_l[5], reset_b_l[4], reset_b_l[6],
     reset_b_l[7], reset_b_l[9], reset_b_l[8], reset_b_l[10],
     reset_b_l[11], reset_b_l[13], reset_b_l[12], reset_b_l[14],
     reset_b_l[15]}), .r_i(net510), .prog(prog), .pgate_l({pgate_l[1],
     pgate_l[0], pgate_l[2], pgate_l[3], pgate_l[5], pgate_l[4],
     pgate_l[6], pgate_l[7], pgate_l[9], pgate_l[8], pgate_l[10],
     pgate_l[11], pgate_l[13], pgate_l[12], pgate_l[14], pgate_l[15]}),
     .mode_i(net504), .sp12_v_b_01_00({net561[0], net561[1], net561[2],
     net561[3], net561[4], net561[5], net561[6], net561[7], net561[8],
     net561[9], net561[10], net561[11], net561[12], net561[13],
     net561[14], net561[15], net561[16], net561[17], net561[18],
     net561[19], net561[20], net561[21], net561[22], net561[23]}),
     .hiz_b_i(net506), .bs_en_i(net503), .update_o(update_o),
     .tclk_o(tclk_o), .shift_o(shift_o), .sdo(sdo), .r_o(r_o),
     .mode_o(mode_o), .hiz_b_o(hiz_b_o), .glb_net_03(glb_in_3[7:0]),
     .glb_net_02(glb_in_2[7:0]), .glb_net_01(glb_in_1[7:0]),
     .bs_en_o(bs_en_o), .sp12_v_b_02_00({net575[0], net575[1],
     net575[2], net575[3], net575[4], net575[5], net575[6], net575[7],
     net575[8], net575[9], net575[10], net575[11], net575[12],
     net575[13], net575[14], net575[15], net575[16], net575[17],
     net575[18], net575[19], net575[20], net575[21], net575[22],
     net575[23]}), .bl_02(bl[125:72]), .bl_01(bl[71:18]),
     .hold_b_l(hold_b_l), .bnl_op_01_00({slf_op_00_01[3],
     slf_op_00_01[2], slf_op_00_01[1], slf_op_00_01[0],
     slf_op_00_01[3], slf_op_00_01[2], slf_op_00_01[1],
     slf_op_00_01[0]}), .cf_bot_l(cf_b_l[71:0]),
     .slf_op_03_00(slf_op_03_00[3:0]), .sp4_v_b_01_00({net582[0],
     net582[1], net582[2], net582[3], net582[4], net582[5], net582[6],
     net582[7], net582[8], net582[9], net582[10], net582[11],
     net582[12], net582[13], net582[14], net582[15], net582[16],
     net582[17], net582[18], net582[19], net582[20], net582[21],
     net582[22], net582[23], net582[24], net582[25], net582[26],
     net582[27], net582[28], net582[29], net582[30], net582[31],
     net582[32], net582[33], net582[34], net582[35], net582[36],
     net582[37], net582[38], net582[39], net582[40], net582[41],
     net582[42], net582[43], net582[44], net582[45], net582[46],
     net582[47]}), .sp12_v_b_03_00({net583[0], net583[1], net583[2],
     net583[3], net583[4], net583[5], net583[6], net583[7], net583[8],
     net583[9], net583[10], net583[11], net583[12], net583[13],
     net583[14], net583[15], net583[16], net583[17], net583[18],
     net583[19], net583[20], net583[21], net583[22], net583[23]}),
     .slf_op_02_00(slf_op_02_00[3:0]),
     .tnr_op_03_00(rgt_op_03_01[7:0]),
     .lft_op_03_00(slf_op_03_01[7:0]), .sp4_v_b_02_00({net587[0],
     net587[1], net587[2], net587[3], net587[4], net587[5], net587[6],
     net587[7], net587[8], net587[9], net587[10], net587[11],
     net587[12], net587[13], net587[14], net587[15], net587[16],
     net587[17], net587[18], net587[19], net587[20], net587[21],
     net587[22], net587[23], net587[24], net587[25], net587[26],
     net587[27], net587[28], net587[29], net587[30], net587[31],
     net587[32], net587[33], net587[34], net587[35], net587[36],
     net587[37], net587[38], net587[39], net587[40], net587[41],
     net587[42], net587[43], net587[44], net587[45], net587[46],
     net587[47]}), .sp4_v_b_03_00({net588[0], net588[1], net588[2],
     net588[3], net588[4], net588[5], net588[6], net588[7], net588[8],
     net588[9], net588[10], net588[11], net588[12], net588[13],
     net588[14], net588[15], net588[16], net588[17], net588[18],
     net588[19], net588[20], net588[21], net588[22], net588[23],
     net588[24], net588[25], net588[26], net588[27], net588[28],
     net588[29], net588[30], net588[31], net588[32], net588[33],
     net588[34], net588[35], net588[36], net588[37], net588[38],
     net588[39], net588[40], net588[41], net588[42], net588[43],
     net588[44], net588[45], net588[46], net588[47]}),
     .lft_op_01_00({net589[0], net589[1], net589[2], net589[3],
     net589[4], net589[5], net589[6], net589[7]}),
     .lft_op_02_00({net590[0], net590[1], net590[2], net590[3],
     net590[4], net590[5], net590[6], net590[7]}),
     .sp4_h_r_03_00(sp4_h_r_03_00[15:0]), .bl_03(bl[179:126]),
     .padin_b_l(padin_b_l[5:0]), .padeb_b_l(padeb_b_l[5:0]),
     .pado_b_l(pado_b_l[5:0]), .fabric_out_02_00(fabric_out_02_00),
     .fabric_out_03_00(fabric_out_03_00), .ceb_o(ceb_o),
     .sp4_h_l_01_00({net515[0], net515[1], net515[2], net515[3],
     net515[4], net515[5], net515[6], net515[7], net515[8], net515[9],
     net515[10], net515[11], net515[12], net515[13], net515[14],
     net515[15]}), .ceb_i(net536));
tielo I450 ( .tielo(tiegnd_bl));
pinlatbuf12p I_pinlatbuf12p_b ( .pad_in(padin_b_l[5]),
     .icegate(hold_l_b), .cbit(cf_b_l[63]), .cout(padinlat_b_l[5]),
     .prog(prog));
scan_buf_ice8p I_scanbuf_8p_ml ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net509), .tclk_o(net516), .shift_o(net502),
     .sdo(net505), .r_o(net510), .mode_o(net504), .hiz_b_o(net506),
     .ceb_o(net536), .bs_en_o(net503));
fabric_buf_ice8p I_fabric_buf8p_25 ( .f_in(padinlat_l_b[7]),
     .f_out(padin_00_04b));
fabric_buf_ice8p I784 ( .f_in(padinlat_b_l[5]), .f_out(padin_03_00b));
pinlatbuf12p_1 I_pinlatbuf12p ( .pad_in(padin_l_b[7]),
     .icegate(hold_l_b), .cbit(cf_l[87]), .cout(padinlat_l_b[7]),
     .prog(prog));

endmodule
// Library - ice8chip, Cell - io_col4_rgt_ice8p_v2, View - schematic
// LAST TIME SAVED: Aug  3 19:20:04 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_col4_rgt_ice8p_v2 ( cbit_colcntl, cf, fabric_out, padeb,
     pado, sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t,
     sp12_h_l, bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold,
     lft_op, mode, padin, pgate, prog, r, reset, sdi, shift, spioeb,
     spiout, tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [7:0]  cbit_colcntl;
output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [1:0]  padeb;
output [3:0]  slf_op;
output [23:0]  cf;

inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;

input [1:0]  padin;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [15:0]  wl;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  tnl_op;
input [1:0]  spioeb;
input [7:0]  glb_netwk;
input [1:0]  spiout;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



RM7  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
RM7  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
RM7  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
RM7  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
RM7  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
RM7  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
RM7  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
RM7  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
RM7  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
RM7  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
RM7  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
RM7  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
RM7  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
RM7  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
RM7  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
RM7  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
sbox1_colbdlc_v4 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_gmux_x16bare_v4 I_io_gmux_x16bare_v4 (
     .cbit_colcntl(cbit_colcntl[7:0]), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});

endmodule
// Library - ice384chip, Cell - io_rgt_bot_1x4_ice384, View - schematic
// LAST TIME SAVED: Jan 12 11:47:06 2012
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_rgt_bot_1x4_ice384 ( cf_r, fabric_out_07_04, padeb, pado,
     sdo, slf_op_07_01, slf_op_07_02, slf_op_07_03, slf_op_07_04,
     tck_pad, tclk_o, tdi_pad, tms_pad, SP4_h_l_07_01, SP4_h_l_07_02,
     SP4_h_l_07_03, SP4_h_l_07_04, SP12_h_l_07_01, SP12_h_l_07_02,
     SP12_h_l_07_03, SP12_h_l_07_04, bl, pgate, reset_b, sp4_v_b_07_01,
     sp4_v_t_07_04, vdd_cntl, wl, bnl_op_07_01, bs_en, ceb, glb_netwk,
     hiz_b, hold, jtag_rowtest_mode_rowu2_b, last_rsr, lft_op_07_01,
     lft_op_07_02, lft_op_07_03, lft_op_07_04, mode, mux_jtag_sel_b,
     padin, prog, r, sdi, sdo_enable, shift, tclk, tnl_op_07_04,
     totdopad, trstb_pad, update );
output  fabric_out_07_04, sdo, tck_pad, tclk_o, tdi_pad, tms_pad;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu2_b, mode,
     mux_jtag_sel_b, prog, r, sdi, sdo_enable, shift, tclk, totdopad,
     trstb_pad, update;

output [3:0]  slf_op_07_04;
output [3:0]  slf_op_07_01;
output [3:0]  slf_op_07_02;
output [3:0]  slf_op_07_03;
output [7:0]  pado;
output [7:0]  padeb;
output [95:0]  cf_r;

inout [47:0]  SP4_h_l_07_02;
inout [23:0]  SP12_h_l_07_03;
inout [47:0]  SP4_h_l_07_01;
inout [15:0]  sp4_v_t_07_04;
inout [15:0]  sp4_v_b_07_01;
inout [23:0]  SP12_h_l_07_01;
inout [23:0]  SP12_h_l_07_04;
inout [23:0]  SP12_h_l_07_02;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_07_03;
inout [47:0]  SP4_h_l_07_04;
inout [63:0]  vdd_cntl;
inout [63:0]  pgate;
inout [63:0]  reset_b;
inout [63:0]  wl;

input [7:0]  lft_op_07_01;
input [7:0]  lft_op_07_02;
input [7:0]  tnl_op_07_04;
input [7:0]  glb_netwk;
input [7:0]  bnl_op_07_01;
input [2:2]  last_rsr;
input [7:0]  lft_op_07_04;
input [7:0]  lft_op_07_03;
input [7:0]  padin;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  net256;

wire  [15:0]  net292;

wire  [1:0]  net217;

wire  [7:0]  net260;

wire  [7:0]  net368;

wire  [7:0]  net296;

wire  [2:0]  net208;

wire  [1:0]  net344;

wire  [35:11]  cf_rp;

wire  [7:0]  net216;

wire  [15:0]  net328;



fabric_buf_ice8p I180 ( .f_in(net370), .f_out(fabric_out_07_04));
mux2_hvt I_mux_jtagcf_2_ ( .in1(cf_rp[35]), .in0(tievdd),
     .out(net208[0]), .sel(mux_jtag_sel_b));
mux2_hvt I_mux_jtagcf_1_ ( .in1(cf_rp[12]), .in0(tievdd),
     .out(net208[1]), .sel(mux_jtag_sel_b));
mux2_hvt I_mux_jtagcf_0_ ( .in1(cf_rp[11]), .in0(tievdd),
     .out(net208[2]), .sel(mux_jtag_sel_b));
bram_bufferx4 I_muxedjtagbuf_2_ ( .in(net208[0]), .out(cf_r[35]));
bram_bufferx4 I_muxedjtagbuf_1_ ( .in(net208[1]), .out(cf_r[12]));
bram_bufferx4 I_muxedjtagbuf_0_ ( .in(net208[2]), .out(cf_r[11]));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tiegnd));
tckbufx32_ice8p I_tmsbuf ( .in(tms), .out(tms_pad));
tckbufx32_ice8p I_tckbuf ( .in(tck), .out(tck_pad));
tckbufx32_ice8p I_tdibuf ( .in(tdi), .out(tdi_pad));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
io_col4_rgt_ice8p_v2 I_io_07_02 ( .slf_op(slf_op_07_02[3:0]),
     .cdone_in(mux_jtag_sel_b), .spioeb({sdo_enable, tievdd}),
     .tnl_op(lft_op_07_03[7:0]), .spi_ss_in_b({nc_ss, tck}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_07_02[23:0]), .spiout({totdopad, tiegnd}),
     .sp4_v_b({net292[0], net292[1], net292[2], net292[3], net292[4],
     net292[5], net292[6], net292[7], net292[8], net292[9], net292[10],
     net292[11], net292[12], net292[13], net292[14], net292[15]}),
     .prog(prog), .cf({cf_r[47:36], cf_rp[35], cf_r[34:24]}),
     .vdd_cntl(vdd_cntl[31:16]), .lft_op(lft_op_07_02[7:0]),
     .padin(padin[3:2]), .mode(mode), .wl(wl[31:16]), .pado(pado[3:2]),
     .sp4_v_t({net256[0], net256[1], net256[2], net256[3], net256[4],
     net256[5], net256[6], net256[7], net256[8], net256[9], net256[10],
     net256[11], net256[12], net256[13], net256[14], net256[15]}),
     .padeb(padeb[3:2]), .reset(reset_b[31:16]), .bl(bl[17:0]),
     .cbit_colcntl({net260[0], net260[1], net260[2], net260[3],
     net260[4], net260[5], net260[6], net260[7]}), .sdo(net261),
     .fabric_out(net219), .glb_netwk(glb_netwk[7:0]),
     .pgate(pgate[31:16]), .sdi(net297), .sp4_h_l(SP4_h_l_07_02[47:0]),
     .bnl_op(lft_op_07_01[7:0]));
io_col4_rgt_ice8p_v2 I_io_07_01 ( .slf_op(slf_op_07_01[3:0]),
     .cdone_in(mux_jtag_sel_b), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_07_02[7:0]), .spi_ss_in_b({tms, tdi}), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_07_01[23:0]),
     .spiout({tiegnd, tiegnd}), .sp4_v_b(sp4_v_b_07_01[15:0]),
     .prog(prog), .cf({cf_r[23:13], cf_rp[12], cf_rp[11], cf_r[10:0]}),
     .vdd_cntl(vdd_cntl[15:0]), .lft_op(lft_op_07_01[7:0]),
     .padin(padin[1:0]), .mode(mode), .wl(wl[15:0]), .pado(pado[1:0]),
     .sp4_v_t({net292[0], net292[1], net292[2], net292[3], net292[4],
     net292[5], net292[6], net292[7], net292[8], net292[9], net292[10],
     net292[11], net292[12], net292[13], net292[14], net292[15]}),
     .padeb(padeb[1:0]), .reset(reset_b[15:0]), .bl(bl[17:0]),
     .cbit_colcntl({net296[0], net296[1], net296[2], net296[3],
     net296[4], net296[5], net296[6], net296[7]}), .sdo(net297),
     .fabric_out(net0296), .glb_netwk(glb_netwk[7:0]),
     .pgate(pgate[15:0]), .sdi(sdi), .sp4_h_l(SP4_h_l_07_01[47:0]),
     .bnl_op(bnl_op_07_01[7:0]));
io_col4_rgt_ice8p_v2 I_io_07_03 ( .slf_op(slf_op_07_03[3:0]),
     .cdone_in(jtag_rowtest_mode_rowu2_b), .spioeb({tievdd, tiegnd}),
     .tnl_op(lft_op_07_04[7:0]), .spi_ss_in_b({net217[0], net217[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_07_03[23:0]), .spiout({tiegnd, last_rsr[2]}),
     .sp4_v_b({net256[0], net256[1], net256[2], net256[3], net256[4],
     net256[5], net256[6], net256[7], net256[8], net256[9], net256[10],
     net256[11], net256[12], net256[13], net256[14], net256[15]}),
     .prog(prog), .cf(cf_r[71:48]), .vdd_cntl(vdd_cntl[47:32]),
     .lft_op(lft_op_07_03[7:0]), .padin(padin[5:4]), .mode(mode),
     .wl(wl[47:32]), .pado(pado[5:4]), .sp4_v_t({net328[0], net328[1],
     net328[2], net328[3], net328[4], net328[5], net328[6], net328[7],
     net328[8], net328[9], net328[10], net328[11], net328[12],
     net328[13], net328[14], net328[15]}), .padeb(padeb[5:4]),
     .reset(reset_b[47:32]), .bl(bl[17:0]), .cbit_colcntl({net216[0],
     net216[1], net216[2], net216[3], net216[4], net216[5], net216[6],
     net216[7]}), .sdo(net333), .fabric_out(net334),
     .glb_netwk(glb_netwk[7:0]), .pgate(pgate[47:32]), .sdi(net261),
     .sp4_h_l(SP4_h_l_07_03[47:0]), .bnl_op(lft_op_07_02[7:0]));
io_col4_rgt_ice8p_v2 I_io_07_04 ( .slf_op(slf_op_07_04[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(tnl_op_07_04[7:0]), .spi_ss_in_b({net344[0], net344[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_07_04[23:0]), .spiout({tiegnd, tiegnd}),
     .sp4_v_b({net328[0], net328[1], net328[2], net328[3], net328[4],
     net328[5], net328[6], net328[7], net328[8], net328[9], net328[10],
     net328[11], net328[12], net328[13], net328[14], net328[15]}),
     .prog(prog), .cf(cf_r[95:72]), .vdd_cntl(vdd_cntl[63:48]),
     .lft_op(lft_op_07_04[7:0]), .padin(padin[7:6]), .mode(mode),
     .wl(wl[63:48]), .pado(pado[7:6]), .sp4_v_t(sp4_v_t_07_04[15:0]),
     .padeb(padeb[7:6]), .reset(reset_b[63:48]), .bl(bl[17:0]),
     .cbit_colcntl({net368[0], net368[1], net368[2], net368[3],
     net368[4], net368[5], net368[6], net368[7]}), .sdo(sdo),
     .fabric_out(net370), .glb_netwk(glb_netwk[7:0]),
     .pgate(pgate[63:48]), .sdi(net333), .sp4_h_l(SP4_h_l_07_04[47:0]),
     .bnl_op(lft_op_07_03[7:0]));

endmodule
// Library - ice384chip, Cell - io_bot_rgt_1x3_ice384, View - schematic
// LAST TIME SAVED: Jan 18 13:09:36 2012
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_bot_rgt_1x3_ice384 ( cf_b_r, fabric_out_04_00, padeb_b_r,
     pado_b_r, sdo_pad, slf_op_04_00, slf_op_05_00, slf_op_06_00,
     spi_ss_in_bbank, bl_04, bl_05, bl_06, sp4_h_l_04_00,
     sp4_h_r_06_00, sp4_v_b_04_00, sp4_v_b_05_00, sp4_v_b_06_00,
     sp12_v_b_04_00, sp12_v_b_05_00, sp12_v_b_06_00, bnl_op_04_00,
     bs_en_i, ceb_i, end_of_startup, glb_net_04, glb_net_05,
     glb_net_06, hiz_b_i, hold_b_r, lft_op_04_00, lft_op_05_00,
     lft_op_06_00, md_spi_b, mode_i, padin_b_r, pgate_r, prog, r_i,
     reset_r, sdi, shift_i, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk_i, tnr_op_06_00, update_i, vdd_cntl_r, wl_r );
output  fabric_out_04_00, sdo_pad;


input  bs_en_i, ceb_i, end_of_startup, hiz_b_i, hold_b_r, md_spi_b,
     mode_i, prog, r_i, sdi, shift_i, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk_i, update_i;

output [3:0]  slf_op_05_00;
output [3:0]  slf_op_04_00;
output [3:0]  slf_op_06_00;
output [4:0]  spi_ss_in_bbank;
output [11:6]  padeb_b_r;
output [11:6]  pado_b_r;
output [71:0]  cf_b_r;

inout [15:0]  sp4_h_l_04_00;
inout [23:0]  sp12_v_b_06_00;
inout [47:0]  sp4_v_b_05_00;
inout [47:0]  sp4_v_b_04_00;
inout [23:0]  sp12_v_b_04_00;
inout [53:0]  bl_06;
inout [47:0]  sp4_v_b_06_00;
inout [15:0]  sp4_h_r_06_00;
inout [23:0]  sp12_v_b_05_00;
inout [53:0]  bl_05;
inout [53:0]  bl_04;

input [7:0]  lft_op_06_00;
input [7:0]  bnl_op_04_00;
input [15:0]  reset_r;
input [15:0]  vdd_cntl_r;
input [7:0]  glb_net_04;
input [15:0]  wl_r;
input [7:0]  tnr_op_06_00;
input [7:0]  glb_net_06;
input [15:0]  pgate_r;
input [11:6]  padin_b_r;
input [7:0]  lft_op_05_00;
input [7:0]  lft_op_04_00;
input [7:0]  glb_net_05;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net0206;

wire  [15:0]  net442;

wire  [15:0]  net407;

wire  [60:11]  cf_b_r_p;

wire  [1:0]  net0197;



lowla_modified I_lowla_modified ( .clk(endtck), .min(net0185),
     .lao(sdo_pad));
bram_bufferx4x6 I_bram_bufferx4x6 ( .in(net0298), .out(net0185));
mux2_hvt I_cfmux_spiss_ck_1_ ( .in1(cf_b_r_p[60]), .in0(tievdd),
     .out(net0197[0]), .sel(end_of_startup));
mux2_hvt I_cfmux_spiss_ck_0_ ( .in1(cf_b_r_p[59]), .in0(tievdd),
     .out(net0197[1]), .sel(end_of_startup));
mux2_hvt I_cfmux_spisdi ( .in1(cf_b_r_p[36]), .in0(tievdd),
     .out(mid_br36), .sel(end_of_startup));
mux2_hvt I_cfmux_coldboot_1_ ( .in1(cf_b_r_p[12]), .in0(tievdd),
     .out(net0206[0]), .sel(end_of_startup));
mux2_hvt I_cfmux_coldboot_0_ ( .in1(cf_b_r_p[11]), .in0(tievdd),
     .out(net0206[1]), .sel(end_of_startup));
bram_bufferx4 I_cfbuf_spiss_ck_1_ ( .in(net0197[0]), .out(cf_b_r[60]));
bram_bufferx4 I_cfbuf_spiss_ck_0_ ( .in(net0197[1]), .out(cf_b_r[59]));
bram_bufferx4 I_buf_spisdi ( .in(mid_br36), .out(cf_b_r[36]));
bram_bufferx4 I_buf_coldboot_1_ ( .in(net0206[0]), .out(cf_b_r[12]));
bram_bufferx4 I_buf_coldboot_0_ ( .in(net0206[1]), .out(cf_b_r[11]));
fabric_buf_ice8p I785 ( .f_in(net460), .f_out(fabric_out_04_00));
scan_buf_ice8p I_scanbuf_bl ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net0219), .tclk_o(net383), .shift_o(net0221),
     .sdo(net385), .r_o(net0223), .mode_o(net0224), .hiz_b_o(net0225),
     .ceb_o(net0226), .bs_en_o(net0227));
io_col4_bot_ice8p I_IO_05_00 ( .sdo(net391), .sdi(net426),
     .spiout({tielow, spi_sdo}), .cdone_in(end_of_startup),
     .spioeb({tievdd, spi_sdo_oe_b}), .sp4_v_t({net442[0], net442[1],
     net442[2], net442[3], net442[4], net442[5], net442[6], net442[7],
     net442[8], net442[9], net442[10], net442[11], net442[12],
     net442[13], net442[14], net442[15]}), .mode(net0224),
     .shift(net0221), .hiz_b(net0225), .r(net0223), .bs_en(net0227),
     .tclk(endtck), .update(net0219), .padin(padin_b_r[9:8]),
     .pado(pado_b_r[9:8]), .padeb(padeb_b_r[9:8]), .sp4_v_b({net407[0],
     net407[1], net407[2], net407[3], net407[4], net407[5], net407[6],
     net407[7], net407[8], net407[9], net407[10], net407[11],
     net407[12], net407[13], net407[14], net407[15]}),
     .sp4_h_l(sp4_v_b_05_00[47:0]), .sp12_h_l(sp12_v_b_05_00[23:0]),
     .prog(prog), .spi_ss_in_b({spi_ss_in_bbank[2], spi_ss_nc}),
     .tnl_op(lft_op_04_00[7:0]), .lft_op(lft_op_05_00[7:0]),
     .bnl_op(lft_op_06_00[7:0]), .pgate(pgate_r[15:0]),
     .reset(reset_r[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_r[15:0]),
     .cf({cf_b_r[47:37], cf_b_r_p[36], cf_b_r[35:24]}), .ceb(net0226),
     .vdd_cntl(vdd_cntl_r[15:0]), .slf_op(slf_op_05_00[3:0]),
     .glb_netwk(glb_net_05[7:0]), .hold(hold_b_r),
     .fabric_out(net371));
io_col4_bot_ice8p I_IO_04_00 ( .sdo(net426), .sdi(net385),
     .spiout({tielow, tielow}), .cdone_in(end_of_startup),
     .spioeb({tievdd, tievdd}), .sp4_v_t(sp4_h_l_04_00[15:0]),
     .mode(net0224), .shift(net0221), .hiz_b(net0225), .r(net0223),
     .bs_en(net0227), .tclk(endtck), .update(net0219),
     .padin(padin_b_r[7:6]), .pado(pado_b_r[7:6]),
     .padeb(padeb_b_r[7:6]), .sp4_v_b({net442[0], net442[1], net442[2],
     net442[3], net442[4], net442[5], net442[6], net442[7], net442[8],
     net442[9], net442[10], net442[11], net442[12], net442[13],
     net442[14], net442[15]}), .sp4_h_l(sp4_v_b_04_00[47:0]),
     .sp12_h_l(sp12_v_b_04_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_bbank[1:0]), .tnl_op(bnl_op_04_00[7:0]),
     .lft_op(lft_op_04_00[7:0]), .bnl_op(lft_op_05_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .bl({bl_04[5],
     bl_04[4], bl_04[37], bl_04[36], bl_04[35], bl_04[34], bl_04[33],
     bl_04[32], bl_04[14], bl_04[20], bl_04[19], bl_04[18], bl_04[17],
     bl_04[16], bl_04[27], bl_04[26], bl_04[25], bl_04[23]}),
     .wl(wl_r[15:0]), .cf({cf_b_r[23:13], cf_b_r_p[12:11],
     cf_b_r[10:0]}), .ceb(net0226), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_04_00[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_b_r), .fabric_out(net460));
io_col4_bot_ice8p I_IO_06_00 ( .sdo(net0298), .sdi(net391),
     .spiout({spi_ss_out, spi_clk_out}), .cdone_in(end_of_startup),
     .spioeb({md_spi_b, md_spi_b}), .sp4_v_t({net407[0], net407[1],
     net407[2], net407[3], net407[4], net407[5], net407[6], net407[7],
     net407[8], net407[9], net407[10], net407[11], net407[12],
     net407[13], net407[14], net407[15]}), .mode(net0224),
     .shift(net0221), .hiz_b(net0225), .r(net0223), .bs_en(net0227),
     .tclk(endtck), .update(net0219), .padin(padin_b_r[11:10]),
     .pado(pado_b_r[11:10]), .padeb(padeb_b_r[11:10]),
     .sp4_v_b(sp4_h_r_06_00[15:0]), .sp4_h_l(sp4_v_b_06_00[47:0]),
     .sp12_h_l(sp12_v_b_06_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_bbank[4:3]), .tnl_op(lft_op_05_00[7:0]),
     .lft_op(lft_op_06_00[7:0]), .bnl_op(tnr_op_06_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_r[15:0]), .cf({cf_b_r[71:61], cf_b_r_p[60:59],
     cf_b_r[58:48]}), .ceb(net0226), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_06_00[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_b_r), .fabric_out(net369));
tckbufx32_ice8p I354 ( .in(net383), .out(endtck));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));

endmodule
// Library - ice384chip, Cell - quad_br_ice384, View - schematic
// LAST TIME SAVED: Dec  6 15:05:48 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module quad_br_ice384 ( bs_en_o, carry_out_04_04, carry_out_05_04,
     carry_out_06_04, ceb_o, cf_b_r, cf_r, fabric_out_04_00,
     fabric_out_07_04, hiz_b_o, mode_o, op_vic_04_04, op_vic_05_04,
     op_vic_06_04, padeb_b_r, padeb_r, padin_04_00a, padin_07_04b,
     pado_b_r, pado_r, r_o, sdo, sdo_pad, shift_o, slf_op_04_00,
     slf_op_04_01, slf_op_04_02, slf_op_04_03, slf_op_04_04,
     slf_op_05_04, slf_op_06_04, slf_op_07_04, spi_ss_in_bbank,
     tck_pad, tclk_o, tdi_pad, tms_pad, update_o, bl, pgate_r,
     reset_b_r, sp4_h_l_04_00, sp4_h_l_04_01, sp4_h_l_04_02,
     sp4_h_l_04_03, sp4_h_l_04_04, sp4_v_b_04_01, sp4_v_b_04_02,
     sp4_v_b_04_03, sp4_v_b_04_04, sp4_v_t_04_04, sp4_v_t_05_04,
     sp4_v_t_06_04, sp4_v_t_07_04, sp12_h_l_04_01, sp12_h_l_04_02,
     sp12_h_l_04_03, sp12_h_l_04_04, sp12_v_t_04_04, sp12_v_t_05_04,
     sp12_v_t_06_04, vdd_cntl_r, wl_r, bnl_op_04_01, bs_en_i, bs_en_mi,
     ceb_i, ceb_mi, end_of_startup, glb_in_4, glb_in_5, glb_in_6,
     glb_in_7, hiz_b_i, hiz_b_mi, hold_b_r, hold_r_b,
     jtag_rowtest_mode_rowu2_b, last_rsr, lft_op_04_01, lft_op_04_02,
     lft_op_04_03, lft_op_04_04, md_spi_b, mode_i, mode_mi,
     mux_jtag_sel_b, padin_b_r, padin_r, prog, purst, r_i, r_mi, sdi,
     sdi_pad, sdo_enable, shift_i, shift_mi, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk_i, tclk_mi, tnl_op_04_04,
     tnl_op_05_04, tnl_op_06_04, tnl_op_07_04, tnr_op_04_04,
     tnr_op_05_04, tnr_op_06_04, top_op_04_04, top_op_05_04,
     top_op_06_04, totdopad, trstb_pad, update_i, update_mi );
output  bs_en_o, carry_out_04_04, carry_out_05_04, carry_out_06_04,
     ceb_o, fabric_out_04_00, fabric_out_07_04, hiz_b_o, mode_o,
     op_vic_04_04, op_vic_05_04, op_vic_06_04, padin_04_00a,
     padin_07_04b, r_o, sdo, sdo_pad, shift_o, tck_pad, tclk_o,
     tdi_pad, tms_pad, update_o;


input  bs_en_i, bs_en_mi, ceb_i, ceb_mi, end_of_startup, hiz_b_i,
     hiz_b_mi, hold_b_r, hold_r_b, jtag_rowtest_mode_rowu2_b, md_spi_b,
     mode_i, mode_mi, mux_jtag_sel_b, prog, purst, r_i, r_mi, sdi,
     sdi_pad, sdo_enable, shift_i, shift_mi, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk_i, tclk_mi, totdopad, trstb_pad,
     update_i, update_mi;

output [7:0]  padeb_r;
output [7:0]  slf_op_04_02;
output [7:0]  slf_op_04_04;
output [11:6]  pado_b_r;
output [7:0]  slf_op_04_03;
output [3:0]  slf_op_04_00;
output [95:0]  cf_r;
output [3:0]  slf_op_07_04;
output [7:0]  slf_op_06_04;
output [11:6]  padeb_b_r;
output [71:0]  cf_b_r;
output [4:0]  spi_ss_in_bbank;
output [7:0]  slf_op_04_01;
output [7:0]  slf_op_05_04;
output [7:0]  pado_r;

inout [15:0]  sp4_v_t_07_04;
inout [47:0]  sp4_h_l_04_01;
inout [23:0]  sp12_h_l_04_03;
inout [23:0]  sp12_v_t_05_04;
inout [23:0]  sp12_v_t_06_04;
inout [47:0]  sp4_v_t_04_04;
inout [47:0]  sp4_v_t_05_04;
inout [47:0]  sp4_h_l_04_03;
inout [179:0]  bl;
inout [47:0]  sp4_v_b_04_02;
inout [79:0]  pgate_r;
inout [79:0]  reset_b_r;
inout [79:0]  vdd_cntl_r;
inout [15:0]  sp4_h_l_04_00;
inout [47:0]  sp4_v_t_06_04;
inout [79:0]  wl_r;
inout [47:0]  sp4_v_b_04_04;
inout [47:0]  sp4_v_b_04_03;
inout [23:0]  sp12_v_t_04_04;
inout [23:0]  sp12_h_l_04_01;
inout [23:0]  sp12_h_l_04_02;
inout [47:0]  sp4_h_l_04_04;
inout [47:0]  sp4_h_l_04_02;
inout [47:0]  sp4_v_b_04_01;
inout [23:0]  sp12_h_l_04_04;

input [7:0]  tnl_op_06_04;
input [7:0]  lft_op_04_04;
input [7:0]  glb_in_7;
input [7:0]  tnr_op_05_04;
input [7:0]  lft_op_04_01;
input [7:0]  tnr_op_04_04;
input [7:0]  top_op_04_04;
input [3:0]  bnl_op_04_01;
input [7:0]  tnl_op_04_04;
input [7:0]  glb_in_5;
input [7:0]  lft_op_04_02;
input [7:0]  glb_in_6;
input [11:6]  padin_b_r;
input [2:2]  last_rsr;
input [7:0]  lft_op_04_03;
input [7:0]  glb_in_4;
input [7:0]  tnl_op_05_04;
input [7:0]  top_op_06_04;
input [7:0]  tnl_op_07_04;
input [7:0]  top_op_05_04;
input [7:0]  padin_r;
input [7:0]  tnr_op_06_04;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [47:0]  net643;

wire  [47:0]  net638;

wire  [3:0]  slf_op_05_00;

wire  [3:0]  slf_op_06_00;

wire  [3:0]  slf_op_07_02;

wire  [3:0]  slf_op_07_03;

wire  [3:0]  slf_op_07_01;

wire  [23:0]  net574;

wire  [47:0]  net583;

wire  [47:0]  net585;

wire  [7:0]  net498;

wire  [7:0]  net500;

wire  [47:0]  net443;

wire  [47:0]  net642;

wire  [23:0]  net610;

wire  [23:0]  net634;

wire  [23:0]  net517;

wire  [47:0]  net524;

wire  [23:0]  net577;

wire  [47:0]  net672;

wire  [7:0]  net614;

wire  [47:0]  net641;

wire  [23:0]  net631;

wire  [47:0]  net526;

wire  [7:0]  net445;

wire  [23:0]  net518;

wire  [47:0]  net527;

wire  [23:0]  net478;

wire  [23:0]  net519;

wire  [47:0]  net529;

wire  [23:0]  net463;

wire  [47:0]  net586;

wire  [7:0]  net451;

wire  [15:0]  net449;

wire  [23:0]  net520;

wire  [23:0]  net575;

wire  [47:0]  net637;

wire  [47:0]  net460;

wire  [23:0]  net633;

wire  [47:0]  net584;

wire  [23:0]  net576;

wire  [47:0]  net522;

wire  [47:0]  net640;

wire  [47:0]  net673;

wire  [47:0]  net523;

wire  [47:0]  net528;

wire  [7:0]  net612;

wire  [47:0]  net670;

wire  [47:0]  net671;

wire  [23:0]  net632;

wire  [47:0]  net636;



scan_buf_ice8p I_scanbuf_8p_br ( .update_i(update_mi),
     .tclk_i(tclk_mi), .shift_i(shift_mi), .sdi(sdi_pad), .r_i(r_mi),
     .mode_i(mode_mi), .hiz_b_i(hiz_b_mi), .ceb_i(ceb_mi),
     .bs_en_i(bs_en_mi), .update_o(update_o), .tclk_o(net379),
     .shift_o(shift_o), .sdo(net381), .r_o(r_o), .mode_o(mode_o),
     .hiz_b_o(hiz_b_o), .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_rgt_bot_1x4_ice384 I809 ( .shift(shift_o), .bs_en(bs_en_o),
     .mode(mode_o), .sdi(net381), .hiz_b(hiz_b_o), .prog(prog),
     .hold(hold_r_b), .update(update_o), .r(r_o), .sdo(sdo),
     .bl(bl[179:162]), .tclk(net379), .trstb_pad(trstb_pad),
     .mux_jtag_sel_b(mux_jtag_sel_b), .sdo_enable(sdo_enable),
     .tclk_o(tclk_o), .ceb(ceb_o), .totdopad(totdopad),
     .tck_pad(tck_pad), .tdi_pad(tdi_pad), .tms_pad(tms_pad),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .last_rsr(last_rsr[2]), .tnl_op_07_04(tnl_op_07_04[7:0]),
     .sp4_v_t_07_04(sp4_v_t_07_04[15:0]), .SP4_h_l_07_01({net586[0],
     net586[1], net586[2], net586[3], net586[4], net586[5], net586[6],
     net586[7], net586[8], net586[9], net586[10], net586[11],
     net586[12], net586[13], net586[14], net586[15], net586[16],
     net586[17], net586[18], net586[19], net586[20], net586[21],
     net586[22], net586[23], net586[24], net586[25], net586[26],
     net586[27], net586[28], net586[29], net586[30], net586[31],
     net586[32], net586[33], net586[34], net586[35], net586[36],
     net586[37], net586[38], net586[39], net586[40], net586[41],
     net586[42], net586[43], net586[44], net586[45], net586[46],
     net586[47]}), .SP4_h_l_07_02({net585[0], net585[1], net585[2],
     net585[3], net585[4], net585[5], net585[6], net585[7], net585[8],
     net585[9], net585[10], net585[11], net585[12], net585[13],
     net585[14], net585[15], net585[16], net585[17], net585[18],
     net585[19], net585[20], net585[21], net585[22], net585[23],
     net585[24], net585[25], net585[26], net585[27], net585[28],
     net585[29], net585[30], net585[31], net585[32], net585[33],
     net585[34], net585[35], net585[36], net585[37], net585[38],
     net585[39], net585[40], net585[41], net585[42], net585[43],
     net585[44], net585[45], net585[46], net585[47]}),
     .SP4_h_l_07_03({net584[0], net584[1], net584[2], net584[3],
     net584[4], net584[5], net584[6], net584[7], net584[8], net584[9],
     net584[10], net584[11], net584[12], net584[13], net584[14],
     net584[15], net584[16], net584[17], net584[18], net584[19],
     net584[20], net584[21], net584[22], net584[23], net584[24],
     net584[25], net584[26], net584[27], net584[28], net584[29],
     net584[30], net584[31], net584[32], net584[33], net584[34],
     net584[35], net584[36], net584[37], net584[38], net584[39],
     net584[40], net584[41], net584[42], net584[43], net584[44],
     net584[45], net584[46], net584[47]}), .SP4_h_l_07_04({net583[0],
     net583[1], net583[2], net583[3], net583[4], net583[5], net583[6],
     net583[7], net583[8], net583[9], net583[10], net583[11],
     net583[12], net583[13], net583[14], net583[15], net583[16],
     net583[17], net583[18], net583[19], net583[20], net583[21],
     net583[22], net583[23], net583[24], net583[25], net583[26],
     net583[27], net583[28], net583[29], net583[30], net583[31],
     net583[32], net583[33], net583[34], net583[35], net583[36],
     net583[37], net583[38], net583[39], net583[40], net583[41],
     net583[42], net583[43], net583[44], net583[45], net583[46],
     net583[47]}), .pgate(pgate_r[79:16]), .wl(wl_r[79:16]),
     .vdd_cntl(vdd_cntl_r[79:16]), .reset_b(reset_b_r[79:16]),
     .slf_op_07_03(slf_op_07_03[3:0]),
     .slf_op_07_01(slf_op_07_01[3:0]),
     .slf_op_07_02(slf_op_07_02[3:0]),
     .slf_op_07_04(slf_op_07_04[3:0]), .glb_netwk(glb_in_7[7:0]),
     .lft_op_07_03({net498[0], net498[1], net498[2], net498[3],
     net498[4], net498[5], net498[6], net498[7]}),
     .lft_op_07_01({net451[0], net451[1], net451[2], net451[3],
     net451[4], net451[5], net451[6], net451[7]}),
     .lft_op_07_02({net500[0], net500[1], net500[2], net500[3],
     net500[4], net500[5], net500[6], net500[7]}),
     .lft_op_07_04(slf_op_06_04[7:0]), .SP12_h_l_07_02({net576[0],
     net576[1], net576[2], net576[3], net576[4], net576[5], net576[6],
     net576[7], net576[8], net576[9], net576[10], net576[11],
     net576[12], net576[13], net576[14], net576[15], net576[16],
     net576[17], net576[18], net576[19], net576[20], net576[21],
     net576[22], net576[23]}), .SP12_h_l_07_03({net575[0], net575[1],
     net575[2], net575[3], net575[4], net575[5], net575[6], net575[7],
     net575[8], net575[9], net575[10], net575[11], net575[12],
     net575[13], net575[14], net575[15], net575[16], net575[17],
     net575[18], net575[19], net575[20], net575[21], net575[22],
     net575[23]}), .SP12_h_l_07_01({net577[0], net577[1], net577[2],
     net577[3], net577[4], net577[5], net577[6], net577[7], net577[8],
     net577[9], net577[10], net577[11], net577[12], net577[13],
     net577[14], net577[15], net577[16], net577[17], net577[18],
     net577[19], net577[20], net577[21], net577[22], net577[23]}),
     .SP12_h_l_07_04({net574[0], net574[1], net574[2], net574[3],
     net574[4], net574[5], net574[6], net574[7], net574[8], net574[9],
     net574[10], net574[11], net574[12], net574[13], net574[14],
     net574[15], net574[16], net574[17], net574[18], net574[19],
     net574[20], net574[21], net574[22], net574[23]}),
     .bnl_op_07_01({slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0], slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0]}), .sp4_v_b_07_01({net449[0],
     net449[1], net449[2], net449[3], net449[4], net449[5], net449[6],
     net449[7], net449[8], net449[9], net449[10], net449[11],
     net449[12], net449[13], net449[14], net449[15]}),
     .fabric_out_07_04(fabric_out_07_04), .padeb(padeb_r[7:0]),
     .pado(pado_r[7:0]), .padin(padin_r[7:0]), .cf_r(cf_r[95:0]));
io_bot_rgt_1x3_ice384 I802 ( .padeb_b_r(padeb_b_r[11:6]),
     .pado_b_r(pado_b_r[11:6]), .padin_b_r(padin_b_r[11:6]),
     .sdo_pad(sdo_pad), .sp4_h_l_04_00(sp4_h_l_04_00[15:0]),
     .bnl_op_04_00(lft_op_04_01[7:0]), .vdd_cntl_r({vdd_cntl_r[1],
     vdd_cntl_r[0], vdd_cntl_r[2], vdd_cntl_r[3], vdd_cntl_r[5],
     vdd_cntl_r[4], vdd_cntl_r[6], vdd_cntl_r[7], vdd_cntl_r[9],
     vdd_cntl_r[8], vdd_cntl_r[10], vdd_cntl_r[11], vdd_cntl_r[13],
     vdd_cntl_r[12], vdd_cntl_r[14], vdd_cntl_r[15]}),
     .sp4_v_b_05_00({net443[0], net443[1], net443[2], net443[3],
     net443[4], net443[5], net443[6], net443[7], net443[8], net443[9],
     net443[10], net443[11], net443[12], net443[13], net443[14],
     net443[15], net443[16], net443[17], net443[18], net443[19],
     net443[20], net443[21], net443[22], net443[23], net443[24],
     net443[25], net443[26], net443[27], net443[28], net443[29],
     net443[30], net443[31], net443[32], net443[33], net443[34],
     net443[35], net443[36], net443[37], net443[38], net443[39],
     net443[40], net443[41], net443[42], net443[43], net443[44],
     net443[45], net443[46], net443[47]}), .cf_b_r(cf_b_r[71:0]),
     .lft_op_05_00({net445[0], net445[1], net445[2], net445[3],
     net445[4], net445[5], net445[6], net445[7]}), .bl_05(bl[107:54]),
     .sp12_v_b_06_00({net610[0], net610[1], net610[2], net610[3],
     net610[4], net610[5], net610[6], net610[7], net610[8], net610[9],
     net610[10], net610[11], net610[12], net610[13], net610[14],
     net610[15], net610[16], net610[17], net610[18], net610[19],
     net610[20], net610[21], net610[22], net610[23]}),
     .sp4_h_r_06_00({net449[0], net449[1], net449[2], net449[3],
     net449[4], net449[5], net449[6], net449[7], net449[8], net449[9],
     net449[10], net449[11], net449[12], net449[13], net449[14],
     net449[15]}), .glb_net_06(glb_in_6[7:0]),
     .lft_op_06_00({net451[0], net451[1], net451[2], net451[3],
     net451[4], net451[5], net451[6], net451[7]}), .bl_06(bl[161:108]),
     .tnr_op_06_00({slf_op_07_01[3], slf_op_07_01[2], slf_op_07_01[1],
     slf_op_07_01[0], slf_op_07_01[3], slf_op_07_01[2],
     slf_op_07_01[1], slf_op_07_01[0]}), .wl_r({wl_r[1], wl_r[0],
     wl_r[2], wl_r[3], wl_r[5], wl_r[4], wl_r[6], wl_r[7], wl_r[9],
     wl_r[8], wl_r[10], wl_r[11], wl_r[13], wl_r[12], wl_r[14],
     wl_r[15]}), .spi_clk_out(spi_clk_out), .spi_ss_out(spi_ss_out),
     .spi_sdo_oe_b(spi_sdo_oe_b), .md_spi_b(md_spi_b),
     .slf_op_06_00(slf_op_06_00[3:0]), .sp4_v_b_06_00({net460[0],
     net460[1], net460[2], net460[3], net460[4], net460[5], net460[6],
     net460[7], net460[8], net460[9], net460[10], net460[11],
     net460[12], net460[13], net460[14], net460[15], net460[16],
     net460[17], net460[18], net460[19], net460[20], net460[21],
     net460[22], net460[23], net460[24], net460[25], net460[26],
     net460[27], net460[28], net460[29], net460[30], net460[31],
     net460[32], net460[33], net460[34], net460[35], net460[36],
     net460[37], net460[38], net460[39], net460[40], net460[41],
     net460[42], net460[43], net460[44], net460[45], net460[46],
     net460[47]}), .glb_net_04(glb_in_4[7:0]),
     .lft_op_04_00(slf_op_04_01[7:0]), .sp12_v_b_04_00({net463[0],
     net463[1], net463[2], net463[3], net463[4], net463[5], net463[6],
     net463[7], net463[8], net463[9], net463[10], net463[11],
     net463[12], net463[13], net463[14], net463[15], net463[16],
     net463[17], net463[18], net463[19], net463[20], net463[21],
     net463[22], net463[23]}), .sp4_v_b_04_00(sp4_v_b_04_01[47:0]),
     .slf_op_04_00(slf_op_04_00[3:0]), .bl_04(bl[53:0]),
     .spi_ss_in_bbank(spi_ss_in_bbank[4:0]), .spi_sdo(spi_sdo),
     .hold_b_r(hold_b_r), .end_of_startup(end_of_startup),
     .reset_r({reset_b_r[1], reset_b_r[0], reset_b_r[2], reset_b_r[3],
     reset_b_r[5], reset_b_r[4], reset_b_r[6], reset_b_r[7],
     reset_b_r[9], reset_b_r[8], reset_b_r[10], reset_b_r[11],
     reset_b_r[13], reset_b_r[12], reset_b_r[14], reset_b_r[15]}),
     .fabric_out_04_00(fabric_out_04_00), .glb_net_05(glb_in_5[7:0]),
     .slf_op_05_00(slf_op_05_00[3:0]), .pgate_r({pgate_r[1],
     pgate_r[0], pgate_r[2], pgate_r[3], pgate_r[5], pgate_r[4],
     pgate_r[6], pgate_r[7], pgate_r[9], pgate_r[8], pgate_r[10],
     pgate_r[11], pgate_r[13], pgate_r[12], pgate_r[14], pgate_r[15]}),
     .sp12_v_b_05_00({net478[0], net478[1], net478[2], net478[3],
     net478[4], net478[5], net478[6], net478[7], net478[8], net478[9],
     net478[10], net478[11], net478[12], net478[13], net478[14],
     net478[15], net478[16], net478[17], net478[18], net478[19],
     net478[20], net478[21], net478[22], net478[23]}),
     .update_i(update_i), .tclk_i(tclk_i), .shift_i(shift_i),
     .sdi(sdi), .r_i(r_i), .prog(prog), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .bs_en_i(bs_en_i), .ceb_i(ceb_i));
lt_1x4_bot_ice384 I805 ( .rgt_op_03({net498[0], net498[1], net498[2],
     net498[3], net498[4], net498[5], net498[6], net498[7]}),
     .slf_op_02({net614[0], net614[1], net614[2], net614[3], net614[4],
     net614[5], net614[6], net614[7]}), .rgt_op_02({net500[0],
     net500[1], net500[2], net500[3], net500[4], net500[5], net500[6],
     net500[7]}), .rgt_op_01({net451[0], net451[1], net451[2],
     net451[3], net451[4], net451[5], net451[6], net451[7]}),
     .purst(purst), .prog(prog), .lft_op_04(slf_op_04_04[7:0]),
     .lft_op_03(slf_op_04_03[7:0]), .lft_op_02(slf_op_04_02[7:0]),
     .lft_op_01(slf_op_04_01[7:0]), .rgt_op_04(slf_op_06_04[7:0]),
     .carry_in(tiegnd_bl), .bnl_op_01({slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0],
     slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0]}), .slf_op_04(slf_op_05_04[7:0]),
     .slf_op_03({net612[0], net612[1], net612[2], net612[3], net612[4],
     net612[5], net612[6], net612[7]}), .slf_op_01({net445[0],
     net445[1], net445[2], net445[3], net445[4], net445[5], net445[6],
     net445[7]}), .sp4_h_l_04({net640[0], net640[1], net640[2],
     net640[3], net640[4], net640[5], net640[6], net640[7], net640[8],
     net640[9], net640[10], net640[11], net640[12], net640[13],
     net640[14], net640[15], net640[16], net640[17], net640[18],
     net640[19], net640[20], net640[21], net640[22], net640[23],
     net640[24], net640[25], net640[26], net640[27], net640[28],
     net640[29], net640[30], net640[31], net640[32], net640[33],
     net640[34], net640[35], net640[36], net640[37], net640[38],
     net640[39], net640[40], net640[41], net640[42], net640[43],
     net640[44], net640[45], net640[46], net640[47]}),
     .carry_out(carry_out_05_04), .vdd_cntl(vdd_cntl_r[79:16]),
     .sp12_h_r_04({net517[0], net517[1], net517[2], net517[3],
     net517[4], net517[5], net517[6], net517[7], net517[8], net517[9],
     net517[10], net517[11], net517[12], net517[13], net517[14],
     net517[15], net517[16], net517[17], net517[18], net517[19],
     net517[20], net517[21], net517[22], net517[23]}),
     .sp12_h_r_03({net518[0], net518[1], net518[2], net518[3],
     net518[4], net518[5], net518[6], net518[7], net518[8], net518[9],
     net518[10], net518[11], net518[12], net518[13], net518[14],
     net518[15], net518[16], net518[17], net518[18], net518[19],
     net518[20], net518[21], net518[22], net518[23]}),
     .sp12_h_r_02({net519[0], net519[1], net519[2], net519[3],
     net519[4], net519[5], net519[6], net519[7], net519[8], net519[9],
     net519[10], net519[11], net519[12], net519[13], net519[14],
     net519[15], net519[16], net519[17], net519[18], net519[19],
     net519[20], net519[21], net519[22], net519[23]}),
     .sp12_h_r_01({net520[0], net520[1], net520[2], net520[3],
     net520[4], net520[5], net520[6], net520[7], net520[8], net520[9],
     net520[10], net520[11], net520[12], net520[13], net520[14],
     net520[15], net520[16], net520[17], net520[18], net520[19],
     net520[20], net520[21], net520[22], net520[23]}),
     .sp4_v_b_01({net443[0], net443[1], net443[2], net443[3],
     net443[4], net443[5], net443[6], net443[7], net443[8], net443[9],
     net443[10], net443[11], net443[12], net443[13], net443[14],
     net443[15], net443[16], net443[17], net443[18], net443[19],
     net443[20], net443[21], net443[22], net443[23], net443[24],
     net443[25], net443[26], net443[27], net443[28], net443[29],
     net443[30], net443[31], net443[32], net443[33], net443[34],
     net443[35], net443[36], net443[37], net443[38], net443[39],
     net443[40], net443[41], net443[42], net443[43], net443[44],
     net443[45], net443[46], net443[47]}), .sp4_r_v_b_04({net522[0],
     net522[1], net522[2], net522[3], net522[4], net522[5], net522[6],
     net522[7], net522[8], net522[9], net522[10], net522[11],
     net522[12], net522[13], net522[14], net522[15], net522[16],
     net522[17], net522[18], net522[19], net522[20], net522[21],
     net522[22], net522[23], net522[24], net522[25], net522[26],
     net522[27], net522[28], net522[29], net522[30], net522[31],
     net522[32], net522[33], net522[34], net522[35], net522[36],
     net522[37], net522[38], net522[39], net522[40], net522[41],
     net522[42], net522[43], net522[44], net522[45], net522[46],
     net522[47]}), .sp4_r_v_b_03({net523[0], net523[1], net523[2],
     net523[3], net523[4], net523[5], net523[6], net523[7], net523[8],
     net523[9], net523[10], net523[11], net523[12], net523[13],
     net523[14], net523[15], net523[16], net523[17], net523[18],
     net523[19], net523[20], net523[21], net523[22], net523[23],
     net523[24], net523[25], net523[26], net523[27], net523[28],
     net523[29], net523[30], net523[31], net523[32], net523[33],
     net523[34], net523[35], net523[36], net523[37], net523[38],
     net523[39], net523[40], net523[41], net523[42], net523[43],
     net523[44], net523[45], net523[46], net523[47]}),
     .sp4_r_v_b_02({net524[0], net524[1], net524[2], net524[3],
     net524[4], net524[5], net524[6], net524[7], net524[8], net524[9],
     net524[10], net524[11], net524[12], net524[13], net524[14],
     net524[15], net524[16], net524[17], net524[18], net524[19],
     net524[20], net524[21], net524[22], net524[23], net524[24],
     net524[25], net524[26], net524[27], net524[28], net524[29],
     net524[30], net524[31], net524[32], net524[33], net524[34],
     net524[35], net524[36], net524[37], net524[38], net524[39],
     net524[40], net524[41], net524[42], net524[43], net524[44],
     net524[45], net524[46], net524[47]}), .sp4_r_v_b_01({net460[0],
     net460[1], net460[2], net460[3], net460[4], net460[5], net460[6],
     net460[7], net460[8], net460[9], net460[10], net460[11],
     net460[12], net460[13], net460[14], net460[15], net460[16],
     net460[17], net460[18], net460[19], net460[20], net460[21],
     net460[22], net460[23], net460[24], net460[25], net460[26],
     net460[27], net460[28], net460[29], net460[30], net460[31],
     net460[32], net460[33], net460[34], net460[35], net460[36],
     net460[37], net460[38], net460[39], net460[40], net460[41],
     net460[42], net460[43], net460[44], net460[45], net460[46],
     net460[47]}), .sp4_h_r_04({net526[0], net526[1], net526[2],
     net526[3], net526[4], net526[5], net526[6], net526[7], net526[8],
     net526[9], net526[10], net526[11], net526[12], net526[13],
     net526[14], net526[15], net526[16], net526[17], net526[18],
     net526[19], net526[20], net526[21], net526[22], net526[23],
     net526[24], net526[25], net526[26], net526[27], net526[28],
     net526[29], net526[30], net526[31], net526[32], net526[33],
     net526[34], net526[35], net526[36], net526[37], net526[38],
     net526[39], net526[40], net526[41], net526[42], net526[43],
     net526[44], net526[45], net526[46], net526[47]}),
     .sp4_h_r_03({net527[0], net527[1], net527[2], net527[3],
     net527[4], net527[5], net527[6], net527[7], net527[8], net527[9],
     net527[10], net527[11], net527[12], net527[13], net527[14],
     net527[15], net527[16], net527[17], net527[18], net527[19],
     net527[20], net527[21], net527[22], net527[23], net527[24],
     net527[25], net527[26], net527[27], net527[28], net527[29],
     net527[30], net527[31], net527[32], net527[33], net527[34],
     net527[35], net527[36], net527[37], net527[38], net527[39],
     net527[40], net527[41], net527[42], net527[43], net527[44],
     net527[45], net527[46], net527[47]}), .sp4_h_r_02({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7], net528[8], net528[9], net528[10], net528[11],
     net528[12], net528[13], net528[14], net528[15], net528[16],
     net528[17], net528[18], net528[19], net528[20], net528[21],
     net528[22], net528[23], net528[24], net528[25], net528[26],
     net528[27], net528[28], net528[29], net528[30], net528[31],
     net528[32], net528[33], net528[34], net528[35], net528[36],
     net528[37], net528[38], net528[39], net528[40], net528[41],
     net528[42], net528[43], net528[44], net528[45], net528[46],
     net528[47]}), .sp4_h_r_01({net529[0], net529[1], net529[2],
     net529[3], net529[4], net529[5], net529[6], net529[7], net529[8],
     net529[9], net529[10], net529[11], net529[12], net529[13],
     net529[14], net529[15], net529[16], net529[17], net529[18],
     net529[19], net529[20], net529[21], net529[22], net529[23],
     net529[24], net529[25], net529[26], net529[27], net529[28],
     net529[29], net529[30], net529[31], net529[32], net529[33],
     net529[34], net529[35], net529[36], net529[37], net529[38],
     net529[39], net529[40], net529[41], net529[42], net529[43],
     net529[44], net529[45], net529[46], net529[47]}),
     .sp4_h_l_03({net641[0], net641[1], net641[2], net641[3],
     net641[4], net641[5], net641[6], net641[7], net641[8], net641[9],
     net641[10], net641[11], net641[12], net641[13], net641[14],
     net641[15], net641[16], net641[17], net641[18], net641[19],
     net641[20], net641[21], net641[22], net641[23], net641[24],
     net641[25], net641[26], net641[27], net641[28], net641[29],
     net641[30], net641[31], net641[32], net641[33], net641[34],
     net641[35], net641[36], net641[37], net641[38], net641[39],
     net641[40], net641[41], net641[42], net641[43], net641[44],
     net641[45], net641[46], net641[47]}), .sp4_h_l_02({net642[0],
     net642[1], net642[2], net642[3], net642[4], net642[5], net642[6],
     net642[7], net642[8], net642[9], net642[10], net642[11],
     net642[12], net642[13], net642[14], net642[15], net642[16],
     net642[17], net642[18], net642[19], net642[20], net642[21],
     net642[22], net642[23], net642[24], net642[25], net642[26],
     net642[27], net642[28], net642[29], net642[30], net642[31],
     net642[32], net642[33], net642[34], net642[35], net642[36],
     net642[37], net642[38], net642[39], net642[40], net642[41],
     net642[42], net642[43], net642[44], net642[45], net642[46],
     net642[47]}), .sp4_h_l_01({net643[0], net643[1], net643[2],
     net643[3], net643[4], net643[5], net643[6], net643[7], net643[8],
     net643[9], net643[10], net643[11], net643[12], net643[13],
     net643[14], net643[15], net643[16], net643[17], net643[18],
     net643[19], net643[20], net643[21], net643[22], net643[23],
     net643[24], net643[25], net643[26], net643[27], net643[28],
     net643[29], net643[30], net643[31], net643[32], net643[33],
     net643[34], net643[35], net643[36], net643[37], net643[38],
     net643[39], net643[40], net643[41], net643[42], net643[43],
     net643[44], net643[45], net643[46], net643[47]}), .bl(bl[107:54]),
     .bot_op_01({slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0], slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0]}), .sp12_h_l_01({net634[0],
     net634[1], net634[2], net634[3], net634[4], net634[5], net634[6],
     net634[7], net634[8], net634[9], net634[10], net634[11],
     net634[12], net634[13], net634[14], net634[15], net634[16],
     net634[17], net634[18], net634[19], net634[20], net634[21],
     net634[22], net634[23]}), .sp12_h_l_02({net633[0], net633[1],
     net633[2], net633[3], net633[4], net633[5], net633[6], net633[7],
     net633[8], net633[9], net633[10], net633[11], net633[12],
     net633[13], net633[14], net633[15], net633[16], net633[17],
     net633[18], net633[19], net633[20], net633[21], net633[22],
     net633[23]}), .sp12_h_l_03({net632[0], net632[1], net632[2],
     net632[3], net632[4], net632[5], net632[6], net632[7], net632[8],
     net632[9], net632[10], net632[11], net632[12], net632[13],
     net632[14], net632[15], net632[16], net632[17], net632[18],
     net632[19], net632[20], net632[21], net632[22], net632[23]}),
     .sp12_h_l_04({net631[0], net631[1], net631[2], net631[3],
     net631[4], net631[5], net631[6], net631[7], net631[8], net631[9],
     net631[10], net631[11], net631[12], net631[13], net631[14],
     net631[15], net631[16], net631[17], net631[18], net631[19],
     net631[20], net631[21], net631[22], net631[23]}),
     .sp4_v_b_04({net636[0], net636[1], net636[2], net636[3],
     net636[4], net636[5], net636[6], net636[7], net636[8], net636[9],
     net636[10], net636[11], net636[12], net636[13], net636[14],
     net636[15], net636[16], net636[17], net636[18], net636[19],
     net636[20], net636[21], net636[22], net636[23], net636[24],
     net636[25], net636[26], net636[27], net636[28], net636[29],
     net636[30], net636[31], net636[32], net636[33], net636[34],
     net636[35], net636[36], net636[37], net636[38], net636[39],
     net636[40], net636[41], net636[42], net636[43], net636[44],
     net636[45], net636[46], net636[47]}), .sp4_v_b_03({net637[0],
     net637[1], net637[2], net637[3], net637[4], net637[5], net637[6],
     net637[7], net637[8], net637[9], net637[10], net637[11],
     net637[12], net637[13], net637[14], net637[15], net637[16],
     net637[17], net637[18], net637[19], net637[20], net637[21],
     net637[22], net637[23], net637[24], net637[25], net637[26],
     net637[27], net637[28], net637[29], net637[30], net637[31],
     net637[32], net637[33], net637[34], net637[35], net637[36],
     net637[37], net637[38], net637[39], net637[40], net637[41],
     net637[42], net637[43], net637[44], net637[45], net637[46],
     net637[47]}), .sp4_v_b_02({net638[0], net638[1], net638[2],
     net638[3], net638[4], net638[5], net638[6], net638[7], net638[8],
     net638[9], net638[10], net638[11], net638[12], net638[13],
     net638[14], net638[15], net638[16], net638[17], net638[18],
     net638[19], net638[20], net638[21], net638[22], net638[23],
     net638[24], net638[25], net638[26], net638[27], net638[28],
     net638[29], net638[30], net638[31], net638[32], net638[33],
     net638[34], net638[35], net638[36], net638[37], net638[38],
     net638[39], net638[40], net638[41], net638[42], net638[43],
     net638[44], net638[45], net638[46], net638[47]}),
     .bnr_op_01({slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0], slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0]}), .top_op_04(top_op_05_04[7:0]),
     .sp12_v_t_04(sp12_v_t_05_04[23:0]), .tnl_op_04(tnl_op_05_04[7:0]),
     .pgate(pgate_r[79:16]), .reset_b(reset_b_r[79:16]),
     .wl(wl_r[79:16]), .tnr_op_04(tnr_op_05_04[7:0]),
     .sp4_v_t_04(sp4_v_t_05_04[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_05_04), .sp12_v_b_01({net478[0], net478[1],
     net478[2], net478[3], net478[4], net478[5], net478[6], net478[7],
     net478[8], net478[9], net478[10], net478[11], net478[12],
     net478[13], net478[14], net478[15], net478[16], net478[17],
     net478[18], net478[19], net478[20], net478[21], net478[22],
     net478[23]}), .glb_netwk(glb_in_5[7:0]));
lt_1x4_bot_ice384 I806 ( .rgt_op_03({slf_op_07_03[3], slf_op_07_03[2],
     slf_op_07_03[1], slf_op_07_03[0], slf_op_07_03[3],
     slf_op_07_03[2], slf_op_07_03[1], slf_op_07_03[0]}),
     .slf_op_02({net500[0], net500[1], net500[2], net500[3], net500[4],
     net500[5], net500[6], net500[7]}), .rgt_op_02({slf_op_07_02[3],
     slf_op_07_02[2], slf_op_07_02[1], slf_op_07_02[0],
     slf_op_07_02[3], slf_op_07_02[2], slf_op_07_02[1],
     slf_op_07_02[0]}), .rgt_op_01({slf_op_07_01[3], slf_op_07_01[2],
     slf_op_07_01[1], slf_op_07_01[0], slf_op_07_01[3],
     slf_op_07_01[2], slf_op_07_01[1], slf_op_07_01[0]}),
     .purst(purst), .prog(prog), .lft_op_04(slf_op_05_04[7:0]),
     .lft_op_03({net612[0], net612[1], net612[2], net612[3], net612[4],
     net612[5], net612[6], net612[7]}), .lft_op_02({net614[0],
     net614[1], net614[2], net614[3], net614[4], net614[5], net614[6],
     net614[7]}), .lft_op_01({net445[0], net445[1], net445[2],
     net445[3], net445[4], net445[5], net445[6], net445[7]}),
     .rgt_op_04({slf_op_07_04[3], slf_op_07_04[2], slf_op_07_04[1],
     slf_op_07_04[0], slf_op_07_04[3], slf_op_07_04[2],
     slf_op_07_04[1], slf_op_07_04[0]}), .carry_in(tiegnd_bl),
     .bnl_op_01({slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0], slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0]}), .slf_op_04(slf_op_06_04[7:0]),
     .slf_op_03({net498[0], net498[1], net498[2], net498[3], net498[4],
     net498[5], net498[6], net498[7]}), .slf_op_01({net451[0],
     net451[1], net451[2], net451[3], net451[4], net451[5], net451[6],
     net451[7]}), .sp4_h_l_04({net526[0], net526[1], net526[2],
     net526[3], net526[4], net526[5], net526[6], net526[7], net526[8],
     net526[9], net526[10], net526[11], net526[12], net526[13],
     net526[14], net526[15], net526[16], net526[17], net526[18],
     net526[19], net526[20], net526[21], net526[22], net526[23],
     net526[24], net526[25], net526[26], net526[27], net526[28],
     net526[29], net526[30], net526[31], net526[32], net526[33],
     net526[34], net526[35], net526[36], net526[37], net526[38],
     net526[39], net526[40], net526[41], net526[42], net526[43],
     net526[44], net526[45], net526[46], net526[47]}),
     .carry_out(carry_out_06_04), .vdd_cntl(vdd_cntl_r[79:16]),
     .sp12_h_r_04({net574[0], net574[1], net574[2], net574[3],
     net574[4], net574[5], net574[6], net574[7], net574[8], net574[9],
     net574[10], net574[11], net574[12], net574[13], net574[14],
     net574[15], net574[16], net574[17], net574[18], net574[19],
     net574[20], net574[21], net574[22], net574[23]}),
     .sp12_h_r_03({net575[0], net575[1], net575[2], net575[3],
     net575[4], net575[5], net575[6], net575[7], net575[8], net575[9],
     net575[10], net575[11], net575[12], net575[13], net575[14],
     net575[15], net575[16], net575[17], net575[18], net575[19],
     net575[20], net575[21], net575[22], net575[23]}),
     .sp12_h_r_02({net576[0], net576[1], net576[2], net576[3],
     net576[4], net576[5], net576[6], net576[7], net576[8], net576[9],
     net576[10], net576[11], net576[12], net576[13], net576[14],
     net576[15], net576[16], net576[17], net576[18], net576[19],
     net576[20], net576[21], net576[22], net576[23]}),
     .sp12_h_r_01({net577[0], net577[1], net577[2], net577[3],
     net577[4], net577[5], net577[6], net577[7], net577[8], net577[9],
     net577[10], net577[11], net577[12], net577[13], net577[14],
     net577[15], net577[16], net577[17], net577[18], net577[19],
     net577[20], net577[21], net577[22], net577[23]}),
     .sp4_v_b_01({net460[0], net460[1], net460[2], net460[3],
     net460[4], net460[5], net460[6], net460[7], net460[8], net460[9],
     net460[10], net460[11], net460[12], net460[13], net460[14],
     net460[15], net460[16], net460[17], net460[18], net460[19],
     net460[20], net460[21], net460[22], net460[23], net460[24],
     net460[25], net460[26], net460[27], net460[28], net460[29],
     net460[30], net460[31], net460[32], net460[33], net460[34],
     net460[35], net460[36], net460[37], net460[38], net460[39],
     net460[40], net460[41], net460[42], net460[43], net460[44],
     net460[45], net460[46], net460[47]}), .sp4_r_v_b_04({net671[0],
     net671[1], net671[2], net671[3], net671[4], net671[5], net671[6],
     net671[7], net671[8], net671[9], net671[10], net671[11],
     net671[12], net671[13], net671[14], net671[15], net671[16],
     net671[17], net671[18], net671[19], net671[20], net671[21],
     net671[22], net671[23], net671[24], net671[25], net671[26],
     net671[27], net671[28], net671[29], net671[30], net671[31],
     net671[32], net671[33], net671[34], net671[35], net671[36],
     net671[37], net671[38], net671[39], net671[40], net671[41],
     net671[42], net671[43], net671[44], net671[45], net671[46],
     net671[47]}), .sp4_r_v_b_03({net672[0], net672[1], net672[2],
     net672[3], net672[4], net672[5], net672[6], net672[7], net672[8],
     net672[9], net672[10], net672[11], net672[12], net672[13],
     net672[14], net672[15], net672[16], net672[17], net672[18],
     net672[19], net672[20], net672[21], net672[22], net672[23],
     net672[24], net672[25], net672[26], net672[27], net672[28],
     net672[29], net672[30], net672[31], net672[32], net672[33],
     net672[34], net672[35], net672[36], net672[37], net672[38],
     net672[39], net672[40], net672[41], net672[42], net672[43],
     net672[44], net672[45], net672[46], net672[47]}),
     .sp4_r_v_b_02({net670[0], net670[1], net670[2], net670[3],
     net670[4], net670[5], net670[6], net670[7], net670[8], net670[9],
     net670[10], net670[11], net670[12], net670[13], net670[14],
     net670[15], net670[16], net670[17], net670[18], net670[19],
     net670[20], net670[21], net670[22], net670[23], net670[24],
     net670[25], net670[26], net670[27], net670[28], net670[29],
     net670[30], net670[31], net670[32], net670[33], net670[34],
     net670[35], net670[36], net670[37], net670[38], net670[39],
     net670[40], net670[41], net670[42], net670[43], net670[44],
     net670[45], net670[46], net670[47]}), .sp4_r_v_b_01({net673[0],
     net673[1], net673[2], net673[3], net673[4], net673[5], net673[6],
     net673[7], net673[8], net673[9], net673[10], net673[11],
     net673[12], net673[13], net673[14], net673[15], net673[16],
     net673[17], net673[18], net673[19], net673[20], net673[21],
     net673[22], net673[23], net673[24], net673[25], net673[26],
     net673[27], net673[28], net673[29], net673[30], net673[31],
     net673[32], net673[33], net673[34], net673[35], net673[36],
     net673[37], net673[38], net673[39], net673[40], net673[41],
     net673[42], net673[43], net673[44], net673[45], net673[46],
     net673[47]}), .sp4_h_r_04({net583[0], net583[1], net583[2],
     net583[3], net583[4], net583[5], net583[6], net583[7], net583[8],
     net583[9], net583[10], net583[11], net583[12], net583[13],
     net583[14], net583[15], net583[16], net583[17], net583[18],
     net583[19], net583[20], net583[21], net583[22], net583[23],
     net583[24], net583[25], net583[26], net583[27], net583[28],
     net583[29], net583[30], net583[31], net583[32], net583[33],
     net583[34], net583[35], net583[36], net583[37], net583[38],
     net583[39], net583[40], net583[41], net583[42], net583[43],
     net583[44], net583[45], net583[46], net583[47]}),
     .sp4_h_r_03({net584[0], net584[1], net584[2], net584[3],
     net584[4], net584[5], net584[6], net584[7], net584[8], net584[9],
     net584[10], net584[11], net584[12], net584[13], net584[14],
     net584[15], net584[16], net584[17], net584[18], net584[19],
     net584[20], net584[21], net584[22], net584[23], net584[24],
     net584[25], net584[26], net584[27], net584[28], net584[29],
     net584[30], net584[31], net584[32], net584[33], net584[34],
     net584[35], net584[36], net584[37], net584[38], net584[39],
     net584[40], net584[41], net584[42], net584[43], net584[44],
     net584[45], net584[46], net584[47]}), .sp4_h_r_02({net585[0],
     net585[1], net585[2], net585[3], net585[4], net585[5], net585[6],
     net585[7], net585[8], net585[9], net585[10], net585[11],
     net585[12], net585[13], net585[14], net585[15], net585[16],
     net585[17], net585[18], net585[19], net585[20], net585[21],
     net585[22], net585[23], net585[24], net585[25], net585[26],
     net585[27], net585[28], net585[29], net585[30], net585[31],
     net585[32], net585[33], net585[34], net585[35], net585[36],
     net585[37], net585[38], net585[39], net585[40], net585[41],
     net585[42], net585[43], net585[44], net585[45], net585[46],
     net585[47]}), .sp4_h_r_01({net586[0], net586[1], net586[2],
     net586[3], net586[4], net586[5], net586[6], net586[7], net586[8],
     net586[9], net586[10], net586[11], net586[12], net586[13],
     net586[14], net586[15], net586[16], net586[17], net586[18],
     net586[19], net586[20], net586[21], net586[22], net586[23],
     net586[24], net586[25], net586[26], net586[27], net586[28],
     net586[29], net586[30], net586[31], net586[32], net586[33],
     net586[34], net586[35], net586[36], net586[37], net586[38],
     net586[39], net586[40], net586[41], net586[42], net586[43],
     net586[44], net586[45], net586[46], net586[47]}),
     .sp4_h_l_03({net527[0], net527[1], net527[2], net527[3],
     net527[4], net527[5], net527[6], net527[7], net527[8], net527[9],
     net527[10], net527[11], net527[12], net527[13], net527[14],
     net527[15], net527[16], net527[17], net527[18], net527[19],
     net527[20], net527[21], net527[22], net527[23], net527[24],
     net527[25], net527[26], net527[27], net527[28], net527[29],
     net527[30], net527[31], net527[32], net527[33], net527[34],
     net527[35], net527[36], net527[37], net527[38], net527[39],
     net527[40], net527[41], net527[42], net527[43], net527[44],
     net527[45], net527[46], net527[47]}), .sp4_h_l_02({net528[0],
     net528[1], net528[2], net528[3], net528[4], net528[5], net528[6],
     net528[7], net528[8], net528[9], net528[10], net528[11],
     net528[12], net528[13], net528[14], net528[15], net528[16],
     net528[17], net528[18], net528[19], net528[20], net528[21],
     net528[22], net528[23], net528[24], net528[25], net528[26],
     net528[27], net528[28], net528[29], net528[30], net528[31],
     net528[32], net528[33], net528[34], net528[35], net528[36],
     net528[37], net528[38], net528[39], net528[40], net528[41],
     net528[42], net528[43], net528[44], net528[45], net528[46],
     net528[47]}), .sp4_h_l_01({net529[0], net529[1], net529[2],
     net529[3], net529[4], net529[5], net529[6], net529[7], net529[8],
     net529[9], net529[10], net529[11], net529[12], net529[13],
     net529[14], net529[15], net529[16], net529[17], net529[18],
     net529[19], net529[20], net529[21], net529[22], net529[23],
     net529[24], net529[25], net529[26], net529[27], net529[28],
     net529[29], net529[30], net529[31], net529[32], net529[33],
     net529[34], net529[35], net529[36], net529[37], net529[38],
     net529[39], net529[40], net529[41], net529[42], net529[43],
     net529[44], net529[45], net529[46], net529[47]}),
     .bl(bl[161:108]), .bot_op_01({slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0], slf_op_06_00[3],
     slf_op_06_00[2], slf_op_06_00[1], slf_op_06_00[0]}),
     .sp12_h_l_01({net520[0], net520[1], net520[2], net520[3],
     net520[4], net520[5], net520[6], net520[7], net520[8], net520[9],
     net520[10], net520[11], net520[12], net520[13], net520[14],
     net520[15], net520[16], net520[17], net520[18], net520[19],
     net520[20], net520[21], net520[22], net520[23]}),
     .sp12_h_l_02({net519[0], net519[1], net519[2], net519[3],
     net519[4], net519[5], net519[6], net519[7], net519[8], net519[9],
     net519[10], net519[11], net519[12], net519[13], net519[14],
     net519[15], net519[16], net519[17], net519[18], net519[19],
     net519[20], net519[21], net519[22], net519[23]}),
     .sp12_h_l_03({net518[0], net518[1], net518[2], net518[3],
     net518[4], net518[5], net518[6], net518[7], net518[8], net518[9],
     net518[10], net518[11], net518[12], net518[13], net518[14],
     net518[15], net518[16], net518[17], net518[18], net518[19],
     net518[20], net518[21], net518[22], net518[23]}),
     .sp12_h_l_04({net517[0], net517[1], net517[2], net517[3],
     net517[4], net517[5], net517[6], net517[7], net517[8], net517[9],
     net517[10], net517[11], net517[12], net517[13], net517[14],
     net517[15], net517[16], net517[17], net517[18], net517[19],
     net517[20], net517[21], net517[22], net517[23]}),
     .sp4_v_b_04({net522[0], net522[1], net522[2], net522[3],
     net522[4], net522[5], net522[6], net522[7], net522[8], net522[9],
     net522[10], net522[11], net522[12], net522[13], net522[14],
     net522[15], net522[16], net522[17], net522[18], net522[19],
     net522[20], net522[21], net522[22], net522[23], net522[24],
     net522[25], net522[26], net522[27], net522[28], net522[29],
     net522[30], net522[31], net522[32], net522[33], net522[34],
     net522[35], net522[36], net522[37], net522[38], net522[39],
     net522[40], net522[41], net522[42], net522[43], net522[44],
     net522[45], net522[46], net522[47]}), .sp4_v_b_03({net523[0],
     net523[1], net523[2], net523[3], net523[4], net523[5], net523[6],
     net523[7], net523[8], net523[9], net523[10], net523[11],
     net523[12], net523[13], net523[14], net523[15], net523[16],
     net523[17], net523[18], net523[19], net523[20], net523[21],
     net523[22], net523[23], net523[24], net523[25], net523[26],
     net523[27], net523[28], net523[29], net523[30], net523[31],
     net523[32], net523[33], net523[34], net523[35], net523[36],
     net523[37], net523[38], net523[39], net523[40], net523[41],
     net523[42], net523[43], net523[44], net523[45], net523[46],
     net523[47]}), .sp4_v_b_02({net524[0], net524[1], net524[2],
     net524[3], net524[4], net524[5], net524[6], net524[7], net524[8],
     net524[9], net524[10], net524[11], net524[12], net524[13],
     net524[14], net524[15], net524[16], net524[17], net524[18],
     net524[19], net524[20], net524[21], net524[22], net524[23],
     net524[24], net524[25], net524[26], net524[27], net524[28],
     net524[29], net524[30], net524[31], net524[32], net524[33],
     net524[34], net524[35], net524[36], net524[37], net524[38],
     net524[39], net524[40], net524[41], net524[42], net524[43],
     net524[44], net524[45], net524[46], net524[47]}),
     .bnr_op_01({tiegnd_bl, tiegnd_bl, tiegnd_bl, tiegnd_bl, tiegnd_bl,
     tiegnd_bl, tiegnd_bl, tiegnd_bl}), .top_op_04(top_op_06_04[7:0]),
     .sp12_v_t_04(sp12_v_t_06_04[23:0]), .tnl_op_04(tnl_op_06_04[7:0]),
     .pgate(pgate_r[79:16]), .reset_b(reset_b_r[79:16]),
     .wl(wl_r[79:16]), .tnr_op_04(tnr_op_06_04[7:0]),
     .sp4_v_t_04(sp4_v_t_06_04[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_06_04), .sp12_v_b_01({net610[0], net610[1],
     net610[2], net610[3], net610[4], net610[5], net610[6], net610[7],
     net610[8], net610[9], net610[10], net610[11], net610[12],
     net610[13], net610[14], net610[15], net610[16], net610[17],
     net610[18], net610[19], net610[20], net610[21], net610[22],
     net610[23]}), .glb_netwk(glb_in_6[7:0]));
lt_1x4_bot_ice384 I804 ( .rgt_op_03({net612[0], net612[1], net612[2],
     net612[3], net612[4], net612[5], net612[6], net612[7]}),
     .slf_op_02(slf_op_04_02[7:0]), .rgt_op_02({net614[0], net614[1],
     net614[2], net614[3], net614[4], net614[5], net614[6],
     net614[7]}), .rgt_op_01({net445[0], net445[1], net445[2],
     net445[3], net445[4], net445[5], net445[6], net445[7]}),
     .purst(purst), .prog(prog), .lft_op_04(lft_op_04_04[7:0]),
     .lft_op_03(lft_op_04_03[7:0]), .lft_op_02(lft_op_04_02[7:0]),
     .lft_op_01(lft_op_04_01[7:0]), .rgt_op_04(slf_op_05_04[7:0]),
     .carry_in(tiegnd_bl), .bnl_op_01({bnl_op_04_01[3],
     bnl_op_04_01[2], bnl_op_04_01[1], bnl_op_04_01[0],
     bnl_op_04_01[3], bnl_op_04_01[2], bnl_op_04_01[1],
     bnl_op_04_01[0]}), .slf_op_04(slf_op_04_04[7:0]),
     .slf_op_03(slf_op_04_03[7:0]), .slf_op_01(slf_op_04_01[7:0]),
     .sp4_h_l_04(sp4_h_l_04_04[47:0]), .carry_out(carry_out_04_04),
     .vdd_cntl(vdd_cntl_r[79:16]), .sp12_h_r_04({net631[0], net631[1],
     net631[2], net631[3], net631[4], net631[5], net631[6], net631[7],
     net631[8], net631[9], net631[10], net631[11], net631[12],
     net631[13], net631[14], net631[15], net631[16], net631[17],
     net631[18], net631[19], net631[20], net631[21], net631[22],
     net631[23]}), .sp12_h_r_03({net632[0], net632[1], net632[2],
     net632[3], net632[4], net632[5], net632[6], net632[7], net632[8],
     net632[9], net632[10], net632[11], net632[12], net632[13],
     net632[14], net632[15], net632[16], net632[17], net632[18],
     net632[19], net632[20], net632[21], net632[22], net632[23]}),
     .sp12_h_r_02({net633[0], net633[1], net633[2], net633[3],
     net633[4], net633[5], net633[6], net633[7], net633[8], net633[9],
     net633[10], net633[11], net633[12], net633[13], net633[14],
     net633[15], net633[16], net633[17], net633[18], net633[19],
     net633[20], net633[21], net633[22], net633[23]}),
     .sp12_h_r_01({net634[0], net634[1], net634[2], net634[3],
     net634[4], net634[5], net634[6], net634[7], net634[8], net634[9],
     net634[10], net634[11], net634[12], net634[13], net634[14],
     net634[15], net634[16], net634[17], net634[18], net634[19],
     net634[20], net634[21], net634[22], net634[23]}),
     .sp4_v_b_01(sp4_v_b_04_01[47:0]), .sp4_r_v_b_04({net636[0],
     net636[1], net636[2], net636[3], net636[4], net636[5], net636[6],
     net636[7], net636[8], net636[9], net636[10], net636[11],
     net636[12], net636[13], net636[14], net636[15], net636[16],
     net636[17], net636[18], net636[19], net636[20], net636[21],
     net636[22], net636[23], net636[24], net636[25], net636[26],
     net636[27], net636[28], net636[29], net636[30], net636[31],
     net636[32], net636[33], net636[34], net636[35], net636[36],
     net636[37], net636[38], net636[39], net636[40], net636[41],
     net636[42], net636[43], net636[44], net636[45], net636[46],
     net636[47]}), .sp4_r_v_b_03({net637[0], net637[1], net637[2],
     net637[3], net637[4], net637[5], net637[6], net637[7], net637[8],
     net637[9], net637[10], net637[11], net637[12], net637[13],
     net637[14], net637[15], net637[16], net637[17], net637[18],
     net637[19], net637[20], net637[21], net637[22], net637[23],
     net637[24], net637[25], net637[26], net637[27], net637[28],
     net637[29], net637[30], net637[31], net637[32], net637[33],
     net637[34], net637[35], net637[36], net637[37], net637[38],
     net637[39], net637[40], net637[41], net637[42], net637[43],
     net637[44], net637[45], net637[46], net637[47]}),
     .sp4_r_v_b_02({net638[0], net638[1], net638[2], net638[3],
     net638[4], net638[5], net638[6], net638[7], net638[8], net638[9],
     net638[10], net638[11], net638[12], net638[13], net638[14],
     net638[15], net638[16], net638[17], net638[18], net638[19],
     net638[20], net638[21], net638[22], net638[23], net638[24],
     net638[25], net638[26], net638[27], net638[28], net638[29],
     net638[30], net638[31], net638[32], net638[33], net638[34],
     net638[35], net638[36], net638[37], net638[38], net638[39],
     net638[40], net638[41], net638[42], net638[43], net638[44],
     net638[45], net638[46], net638[47]}), .sp4_r_v_b_01({net443[0],
     net443[1], net443[2], net443[3], net443[4], net443[5], net443[6],
     net443[7], net443[8], net443[9], net443[10], net443[11],
     net443[12], net443[13], net443[14], net443[15], net443[16],
     net443[17], net443[18], net443[19], net443[20], net443[21],
     net443[22], net443[23], net443[24], net443[25], net443[26],
     net443[27], net443[28], net443[29], net443[30], net443[31],
     net443[32], net443[33], net443[34], net443[35], net443[36],
     net443[37], net443[38], net443[39], net443[40], net443[41],
     net443[42], net443[43], net443[44], net443[45], net443[46],
     net443[47]}), .sp4_h_r_04({net640[0], net640[1], net640[2],
     net640[3], net640[4], net640[5], net640[6], net640[7], net640[8],
     net640[9], net640[10], net640[11], net640[12], net640[13],
     net640[14], net640[15], net640[16], net640[17], net640[18],
     net640[19], net640[20], net640[21], net640[22], net640[23],
     net640[24], net640[25], net640[26], net640[27], net640[28],
     net640[29], net640[30], net640[31], net640[32], net640[33],
     net640[34], net640[35], net640[36], net640[37], net640[38],
     net640[39], net640[40], net640[41], net640[42], net640[43],
     net640[44], net640[45], net640[46], net640[47]}),
     .sp4_h_r_03({net641[0], net641[1], net641[2], net641[3],
     net641[4], net641[5], net641[6], net641[7], net641[8], net641[9],
     net641[10], net641[11], net641[12], net641[13], net641[14],
     net641[15], net641[16], net641[17], net641[18], net641[19],
     net641[20], net641[21], net641[22], net641[23], net641[24],
     net641[25], net641[26], net641[27], net641[28], net641[29],
     net641[30], net641[31], net641[32], net641[33], net641[34],
     net641[35], net641[36], net641[37], net641[38], net641[39],
     net641[40], net641[41], net641[42], net641[43], net641[44],
     net641[45], net641[46], net641[47]}), .sp4_h_r_02({net642[0],
     net642[1], net642[2], net642[3], net642[4], net642[5], net642[6],
     net642[7], net642[8], net642[9], net642[10], net642[11],
     net642[12], net642[13], net642[14], net642[15], net642[16],
     net642[17], net642[18], net642[19], net642[20], net642[21],
     net642[22], net642[23], net642[24], net642[25], net642[26],
     net642[27], net642[28], net642[29], net642[30], net642[31],
     net642[32], net642[33], net642[34], net642[35], net642[36],
     net642[37], net642[38], net642[39], net642[40], net642[41],
     net642[42], net642[43], net642[44], net642[45], net642[46],
     net642[47]}), .sp4_h_r_01({net643[0], net643[1], net643[2],
     net643[3], net643[4], net643[5], net643[6], net643[7], net643[8],
     net643[9], net643[10], net643[11], net643[12], net643[13],
     net643[14], net643[15], net643[16], net643[17], net643[18],
     net643[19], net643[20], net643[21], net643[22], net643[23],
     net643[24], net643[25], net643[26], net643[27], net643[28],
     net643[29], net643[30], net643[31], net643[32], net643[33],
     net643[34], net643[35], net643[36], net643[37], net643[38],
     net643[39], net643[40], net643[41], net643[42], net643[43],
     net643[44], net643[45], net643[46], net643[47]}),
     .sp4_h_l_03(sp4_h_l_04_03[47:0]),
     .sp4_h_l_02(sp4_h_l_04_02[47:0]),
     .sp4_h_l_01(sp4_h_l_04_01[47:0]), .bl(bl[53:0]),
     .bot_op_01({slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0], slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0]}),
     .sp12_h_l_01(sp12_h_l_04_01[23:0]),
     .sp12_h_l_02(sp12_h_l_04_02[23:0]),
     .sp12_h_l_03(sp12_h_l_04_03[23:0]),
     .sp12_h_l_04(sp12_h_l_04_04[23:0]),
     .sp4_v_b_04(sp4_v_b_04_04[47:0]),
     .sp4_v_b_03(sp4_v_b_04_03[47:0]),
     .sp4_v_b_02(sp4_v_b_04_02[47:0]), .bnr_op_01({slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0],
     slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0]}), .top_op_04(top_op_04_04[7:0]),
     .sp12_v_t_04(sp12_v_t_04_04[23:0]), .tnl_op_04(tnl_op_04_04[7:0]),
     .pgate(pgate_r[79:16]), .reset_b(reset_b_r[79:16]),
     .wl(wl_r[79:16]), .tnr_op_04(tnr_op_04_04[7:0]),
     .sp4_v_t_04(sp4_v_t_04_04[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_04_04), .sp12_v_b_01({net463[0], net463[1],
     net463[2], net463[3], net463[4], net463[5], net463[6], net463[7],
     net463[8], net463[9], net463[10], net463[11], net463[12],
     net463[13], net463[14], net463[15], net463[16], net463[17],
     net463[18], net463[19], net463[20], net463[21], net463[22],
     net463[23]}), .glb_netwk(glb_in_4[7:0]));
tielo I450 ( .tielo(tiegnd_bl));
fabric_buf_ice8p I454 ( .f_in(net0668), .f_out(padin_04_00a));
fabric_buf_ice8p I485 ( .f_in(net691), .f_out(padin_07_04b));
pinlatbuf12p_1 I486 ( .pad_in(padin_b_r[6]), .icegate(hold_b_r),
     .cbit(cf_b_r[15]), .cout(net0668), .prog(prog));
pinlatbuf12p_1 I484 ( .pad_in(padin_r[7]), .icegate(hold_r_b),
     .cbit(cf_r[87]), .cout(net691), .prog(prog));

endmodule
// Library - ice384chip, Cell - io_rgt_top_1x4_ice384, View - schematic
// LAST TIME SAVED: Nov 14 19:01:03 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_rgt_top_1x4_ice384 ( cf_r, fabric_out_07_05,
     fabric_out_07_06, padeb, pado, sdo, slf_op_07_05, slf_op_07_06,
     slf_op_07_07, slf_op_07_08, tclk_o, SP4_h_l_07_05, SP4_h_l_07_06,
     SP4_h_l_07_07, SP4_h_l_07_08, SP12_h_l_07_05, SP12_h_l_07_06,
     SP12_h_l_07_07, SP12_h_l_07_08, bl, pgate, reset_b, sp4_v_b_07_05,
     sp4_v_t_07_08, vdd_cntl, wl, bnl_op_07_05, bs_en, ceb, glb_netwk,
     hiz_b, hold, jtag_rowtest_mode_rowu3_b, last_rsr, lft_op_07_05,
     lft_op_07_06, lft_op_07_07, lft_op_07_08, mode, padin, prog, r,
     sdi, shift, tclk, tnl_op_07_08, update );
output  fabric_out_07_05, fabric_out_07_06, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu3_b, mode, prog,
     r, sdi, shift, tclk, update;

output [3:0]  slf_op_07_08;
output [3:0]  slf_op_07_05;
output [3:0]  slf_op_07_07;
output [15:8]  padeb;
output [95:0]  cf_r;
output [15:8]  pado;
output [3:0]  slf_op_07_06;

inout [47:0]  SP4_h_l_07_05;
inout [23:0]  SP12_h_l_07_07;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_07_07;
inout [47:0]  SP4_h_l_07_08;
inout [23:0]  SP12_h_l_07_06;
inout [15:0]  sp4_v_b_07_05;
inout [23:0]  SP12_h_l_07_05;
inout [15:0]  sp4_v_t_07_08;
inout [47:0]  SP4_h_l_07_06;
inout [63:0]  vdd_cntl;
inout [63:0]  pgate;
inout [63:0]  reset_b;
inout [23:0]  SP12_h_l_07_08;
inout [63:0]  wl;

input [7:0]  lft_op_07_06;
input [7:0]  lft_op_07_05;
input [7:0]  glb_netwk;
input [7:0]  tnl_op_07_08;
input [7:0]  lft_op_07_08;
input [7:0]  lft_op_07_07;
input [3:3]  last_rsr;
input [7:0]  bnl_op_07_05;
input [15:8]  padin;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net590;

wire  [15:0]  net514;

wire  [7:0]  net461;

wire  [15:0]  net478;

wire  [15:0]  net550;

wire  [1:0]  net620;

wire  [1:0]  net630;

wire  [7:0]  net0466;

wire  [1:0]  net624;

wire  [7:0]  net497;

wire  [7:0]  net623;



fabric_buf_ice8p I171 ( .f_in(net0350), .f_out(fabric_out_07_06));
fabric_buf_ice8p I166 ( .f_in(net0386), .f_out(fabric_out_07_05));
io_col4_rgt_ice8p_v2 I_io_07_06 ( .cbit_colcntl({net461[0], net461[1],
     net461[2], net461[3], net461[4], net461[5], net461[6],
     net461[7]}), .ceb(ceb), .sdo(net463), .sdi(net499),
     .spiout({tiegnd, last_rsr[3]}),
     .cdone_in(jtag_rowtest_mode_rowu3_b), .spioeb({tievdd, tiegnd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin(padin[11:10]),
     .pado(pado[11:10]), .padeb(padeb[11:10]), .sp4_v_t({net478[0],
     net478[1], net478[2], net478[3], net478[4], net478[5], net478[6],
     net478[7], net478[8], net478[9], net478[10], net478[11],
     net478[12], net478[13], net478[14], net478[15]}),
     .sp4_h_l(SP4_h_l_07_06[47:0]), .sp12_h_l(SP12_h_l_07_06[23:0]),
     .prog(prog), .spi_ss_in_b({net630[0], net630[1]}),
     .tnl_op(lft_op_07_07[7:0]), .lft_op(lft_op_07_06[7:0]),
     .bnl_op(lft_op_07_05[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b({net514[0], net514[1], net514[2],
     net514[3], net514[4], net514[5], net514[6], net514[7], net514[8],
     net514[9], net514[10], net514[11], net514[12], net514[13],
     net514[14], net514[15]}), .wl(wl[31:16]), .cf(cf_r[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_07_06[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(net0350));
io_col4_rgt_ice8p_v2 I_io_07_05 ( .cbit_colcntl({net497[0], net497[1],
     net497[2], net497[3], net497[4], net497[5], net497[6],
     net497[7]}), .ceb(ceb), .sdo(net499), .sdi(sdi), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin(padin[9:8]),
     .pado(pado[9:8]), .padeb(padeb[9:8]), .sp4_v_t({net514[0],
     net514[1], net514[2], net514[3], net514[4], net514[5], net514[6],
     net514[7], net514[8], net514[9], net514[10], net514[11],
     net514[12], net514[13], net514[14], net514[15]}),
     .sp4_h_l(SP4_h_l_07_05[47:0]), .sp12_h_l(SP12_h_l_07_05[23:0]),
     .prog(prog), .spi_ss_in_b({net620[0], net620[1]}),
     .tnl_op(lft_op_07_06[7:0]), .lft_op(lft_op_07_05[7:0]),
     .bnl_op(bnl_op_07_05[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_07_05[15:0]),
     .wl(wl[15:0]), .cf(cf_r[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_07_05[3:0]),
     .glb_netwk(glb_netwk[7:0]), .hold(hold), .fabric_out(net0386));
io_col4_rgt_ice8p_v2 I_io_07_07 ( .cbit_colcntl({net623[0], net623[1],
     net623[2], net623[3], net623[4], net623[5], net623[6],
     net623[7]}), .ceb(ceb), .sdo(net535), .sdi(net463),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[13:12]), .pado(pado[13:12]), .padeb(padeb[13:12]),
     .sp4_v_t({net550[0], net550[1], net550[2], net550[3], net550[4],
     net550[5], net550[6], net550[7], net550[8], net550[9], net550[10],
     net550[11], net550[12], net550[13], net550[14], net550[15]}),
     .sp4_h_l(SP4_h_l_07_07[47:0]), .sp12_h_l(SP12_h_l_07_07[23:0]),
     .prog(prog), .spi_ss_in_b({net624[0], net624[1]}),
     .tnl_op(lft_op_07_08[7:0]), .lft_op(lft_op_07_07[7:0]),
     .bnl_op(lft_op_07_06[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b({net478[0], net478[1], net478[2],
     net478[3], net478[4], net478[5], net478[6], net478[7], net478[8],
     net478[9], net478[10], net478[11], net478[12], net478[13],
     net478[14], net478[15]}), .wl(wl[47:32]), .cf(cf_r[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_07_07[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(net568));
io_col4_rgt_ice8p_v2 I_io_07_08 ( .cbit_colcntl({net0466[0],
     net0466[1], net0466[2], net0466[3], net0466[4], net0466[5],
     net0466[6], net0466[7]}), .ceb(ceb), .sdo(sdo), .sdi(net535),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[15:14]), .pado(pado[15:14]), .padeb(padeb[15:14]),
     .sp4_v_t(sp4_v_t_07_08[15:0]), .sp4_h_l(SP4_h_l_07_08[47:0]),
     .sp12_h_l(SP12_h_l_07_08[23:0]), .prog(prog),
     .spi_ss_in_b({net590[0], net590[1]}), .tnl_op(tnl_op_07_08[7:0]),
     .lft_op(lft_op_07_08[7:0]), .bnl_op(lft_op_07_07[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]), .sp4_v_b({net550[0],
     net550[1], net550[2], net550[3], net550[4], net550[5], net550[6],
     net550[7], net550[8], net550[9], net550[10], net550[11],
     net550[12], net550[13], net550[14], net550[15]}), .wl(wl[63:48]),
     .cf(cf_r[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_07_08[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(net604));
tckbufx32_ice8p I165 ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));

endmodule
// Library - ice8chip, Cell - io_col4_top_ice8p, View - schematic
// LAST TIME SAVED: Aug  3 19:20:04 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_col4_top_ice8p ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [23:0]  cf;
output [1:0]  pado;
output [1:0]  spi_ss_in_b;
output [1:0]  padeb;
output [3:0]  slf_op;

inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [17:0]  bl;

input [1:0]  spioeb;
input [1:0]  padin;
input [7:0]  glb_netwk;
input [15:0]  wl;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [1:0]  spiout;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net0100;

wire  [5:0]  ti;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  om;

wire  [1:0]  oenm;



RM6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
RM6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
RM6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
RM6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
RM6  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
RM6  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
RM6  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
RM6  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
RM6  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
RM6  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
RM6  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
RM6  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
RM6  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
RM6  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
RM6  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
RM6  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
sbox1_colbdlc_v3 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
io_gmux_x16bare_v3 I_io_gmux_x16bare_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .cbitb_colcntl({net0100[0], net0100[1], net0100[2], net0100[3],
     net0100[4], net0100[5], net0100[6], net0100[7]}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));

endmodule
// Library - ice384chip, Cell - io_top_rgt_1x3_ice384, View - schematic
// LAST TIME SAVED: Nov 30 14:39:28 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_top_rgt_1x3_ice384 ( bs_en_o, ceb_o, cf_top_r,
     fabric_out_04_09, fabric_out_05_09, hiz_b_o, mode_o, padeb_t_r,
     pado_t_r, r_o, sdo, shift_o, slf_op_04_09, slf_op_05_09,
     slf_op_06_09, tclk_o, update_o, bl_04, bl_05, bl_06,
     sp4_h_l_04_09, sp4_h_r_06_09, sp4_v_b_04_09, sp4_v_b_05_09,
     sp4_v_b_06_09, sp12_v_b_04_09, sp12_v_b_05_09, sp12_v_b_06_09,
     bnl_op_04_09, bnr_op_06_09, bs_en_i, ceb_i, glb_net_04,
     glb_net_05, glb_net_06, hiz_b_i, hold_t_r, lft_op_04_09,
     lft_op_05_09, lft_op_06_09, mode_i, padin_t_r, pgate_l, prog, r_i,
     reset_l, sdi, shift_i, tclk_i, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_04_09, fabric_out_05_09, hiz_b_o,
     mode_o, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_r, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_04_09;
output [3:0]  slf_op_05_09;
output [3:0]  slf_op_06_09;
output [11:6]  padeb_t_r;
output [71:0]  cf_top_r;
output [11:6]  pado_t_r;

inout [47:0]  sp4_v_b_05_09;
inout [23:0]  sp12_v_b_05_09;
inout [15:0]  sp4_h_r_06_09;
inout [23:0]  sp12_v_b_06_09;
inout [47:0]  sp4_v_b_06_09;
inout [23:0]  sp12_v_b_04_09;
inout [15:0]  sp4_h_l_04_09;
inout [47:0]  sp4_v_b_04_09;
inout [53:0]  bl_06;
inout [53:0]  bl_04;
inout [53:0]  bl_05;

input [7:0]  bnr_op_06_09;
input [15:0]  wl_l;
input [7:0]  glb_net_04;
input [7:0]  bnl_op_04_09;
input [7:0]  lft_op_06_09;
input [7:0]  glb_net_05;
input [15:0]  pgate_l;
input [15:0]  reset_l;
input [7:0]  lft_op_04_09;
input [7:0]  glb_net_06;
input [15:0]  vdd_cntl_l;
input [11:6]  padin_t_r;
input [7:0]  lft_op_05_09;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  net1357;

wire  [15:0]  net1427;

wire  [1:0]  net1312;

wire  [1:0]  net1431;

wire  [1:0]  net1361;



fabric_buf_ice8p I388 ( .f_in(net1445), .f_out(fabric_out_04_09));
fabric_buf_ice8p I347 ( .f_in(net1320), .f_out(fabric_out_05_09));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(net0262), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));
scan_buf_ice8p I345 ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net0262), .shift_o(shift_o),
     .sdo(net1517), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_top_ice8p I_IO_05_09 ( .sdo(net1412), .sdi(net1342),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1427[0], net1427[1], net1427[2],
     net1427[3], net1427[4], net1427[5], net1427[6], net1427[7],
     net1427[8], net1427[9], net1427[10], net1427[11], net1427[12],
     net1427[13], net1427[14], net1427[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_r[9:8]),
     .pado(pado_t_r[9:8]), .padeb(padeb_t_r[9:8]),
     .sp4_v_b({net1357[0], net1357[1], net1357[2], net1357[3],
     net1357[4], net1357[5], net1357[6], net1357[7], net1357[8],
     net1357[9], net1357[10], net1357[11], net1357[12], net1357[13],
     net1357[14], net1357[15]}), .sp4_h_l(sp4_v_b_05_09[47:0]),
     .sp12_h_l(sp12_v_b_05_09[23:0]), .prog(prog),
     .spi_ss_in_b({net1361[0], net1361[1]}),
     .tnl_op(lft_op_04_09[7:0]), .lft_op(lft_op_05_09[7:0]),
     .bnl_op(lft_op_06_09[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_r[47:24]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_09[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_t_r), .fabric_out(net1320));
io_col4_top_ice8p I_IO_04_09 ( .sdo(sdo), .sdi(net1412),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_04_09[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_r[7:6]),
     .pado(pado_t_r[7:6]), .padeb(padeb_t_r[7:6]),
     .sp4_v_b({net1427[0], net1427[1], net1427[2], net1427[3],
     net1427[4], net1427[5], net1427[6], net1427[7], net1427[8],
     net1427[9], net1427[10], net1427[11], net1427[12], net1427[13],
     net1427[14], net1427[15]}), .sp4_h_l(sp4_v_b_04_09[47:0]),
     .sp12_h_l(sp12_v_b_04_09[23:0]), .prog(prog),
     .spi_ss_in_b({net1431[0], net1431[1]}),
     .tnl_op(bnl_op_04_09[7:0]), .lft_op(lft_op_04_09[7:0]),
     .bnl_op(lft_op_05_09[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_r[23:0]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_09[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_t_r), .fabric_out(net1445));
io_col4_top_ice8p I_IO_06_09 ( .sdo(net1342), .sdi(net1517),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1357[0], net1357[1], net1357[2],
     net1357[3], net1357[4], net1357[5], net1357[6], net1357[7],
     net1357[8], net1357[9], net1357[10], net1357[11], net1357[12],
     net1357[13], net1357[14], net1357[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_r[11:10]),
     .pado(pado_t_r[11:10]), .padeb(padeb_t_r[11:10]),
     .sp4_v_b(sp4_h_r_06_09[15:0]), .sp4_h_l(sp4_v_b_06_09[47:0]),
     .sp12_h_l(sp12_v_b_06_09[23:0]), .prog(prog),
     .spi_ss_in_b({net1312[0], net1312[1]}),
     .tnl_op(lft_op_05_09[7:0]), .lft_op(lft_op_06_09[7:0]),
     .bnl_op(bnr_op_06_09[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_06[5], bl_06[4], bl_06[37],
     bl_06[36], bl_06[35], bl_06[34], bl_06[33], bl_06[32], bl_06[14],
     bl_06[20], bl_06[19], bl_06[18], bl_06[17], bl_06[16], bl_06[27],
     bl_06[26], bl_06[25], bl_06[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_r[71:48]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_09[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_t_r), .fabric_out(net0307));

endmodule
// Library - ice384chip, Cell - lt_1x4_top_ice384, View - schematic
// LAST TIME SAVED: Nov  8 15:08:00 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module lt_1x4_top_ice384 ( carry_out, op_vic, slf_op_01, slf_op_02,
     slf_op_03, slf_op_04, bl, glb_netwk, pgate, reset_b, sp4_h_l_01,
     sp4_h_l_02, sp4_h_l_03, sp4_h_l_04, sp4_h_r_01, sp4_h_r_02,
     sp4_h_r_03, sp4_h_r_04, sp4_r_v_b_01, sp4_r_v_b_02, sp4_r_v_b_03,
     sp4_r_v_b_04, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03, sp4_v_b_04,
     sp4_v_t_04, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04,
     sp12_h_r_01, sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_v_b_01,
     sp12_v_t_04, vdd_cntl, wl, bnl_op_01, bnr_op_01, bot_op_01,
     carry_in, lc_bot, lft_op_01, lft_op_02, lft_op_03, lft_op_04,
     prog, purst, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04,
     tnl_op_04, tnr_op_04, top_op_04 );
output  carry_out, op_vic;


input  carry_in, lc_bot, prog, purst;

output [7:0]  slf_op_02;
output [7:0]  slf_op_03;
output [7:0]  slf_op_04;
output [7:0]  slf_op_01;

inout [47:0]  sp4_h_l_02;
inout [53:0]  bl;
inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_h_r_03;
inout [23:0]  sp12_h_l_03;
inout [23:0]  sp12_h_r_04;
inout [47:0]  sp4_v_b_01;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_r_v_b_04;
inout [23:0]  sp12_v_b_01;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_h_r_04;
inout [23:0]  sp12_v_t_04;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_v_t_04;
inout [47:0]  sp4_h_l_04;
inout [47:0]  sp4_v_b_03;
inout [7:0]  glb_netwk;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_r_v_b_02;
inout [63:0]  vdd_cntl;
inout [63:0]  reset_b;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_l_01;
inout [63:0]  wl;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_h_r_01;
inout [63:0]  pgate;
inout [23:0]  sp12_h_l_04;

input [7:0]  lft_op_01;
input [7:0]  lft_op_03;
input [7:0]  tnr_op_04;
input [7:0]  bnr_op_01;
input [7:0]  tnl_op_04;
input [7:0]  rgt_op_01;
input [7:0]  lft_op_04;
input [7:0]  bnl_op_01;
input [7:0]  rgt_op_04;
input [7:0]  top_op_04;
input [7:0]  rgt_op_02;
input [7:0]  bot_op_01;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_02;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net311;

wire  [23:0]  net199;

wire  [7:0]  net280;

wire  [7:0]  net249;

wire  [23:0]  net292;

wire  [7:0]  net187;

wire  [23:0]  net261;



ltile4_ice1f I_LT03 ( .cntl_cbit({net187[0], net187[1], net187[2],
     net187[3], net187[4], net187[5], net187[6], net187[7]}),
     .op_bot(net282), .op_vic(net189), .prog(prog), .carry_out(net191),
     .lft_op(lft_op_03[7:0]), .sp12_h_l(sp12_h_l_03[23:0]),
     .sp4_h_l(sp4_h_l_03[47:0]), .sp4_v_b(sp4_v_b_03[47:0]),
     .sp12_v_b({net292[0], net292[1], net292[2], net292[3], net292[4],
     net292[5], net292[6], net292[7], net292[8], net292[9], net292[10],
     net292[11], net292[12], net292[13], net292[14], net292[15],
     net292[16], net292[17], net292[18], net292[19], net292[20],
     net292[21], net292[22], net292[23]}),
     .sp12_h_r(sp12_h_r_03[23:0]), .sp4_h_r(sp4_h_r_03[47:0]),
     .sp12_v_t({net199[0], net199[1], net199[2], net199[3], net199[4],
     net199[5], net199[6], net199[7], net199[8], net199[9], net199[10],
     net199[11], net199[12], net199[13], net199[14], net199[15],
     net199[16], net199[17], net199[18], net199[19], net199[20],
     net199[21], net199[22], net199[23]}), .sp4_v_t(sp4_v_b_04[47:0]),
     .sp4_r_v_b(sp4_r_v_b_03[47:0]), .wl(wl[47:32]),
     .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net284), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4_ice1f I_LT04 ( .cntl_cbit({net311[0], net311[1], net311[2],
     net311[3], net311[4], net311[5], net311[6], net311[7]}),
     .op_bot(net189), .op_vic(op_vic), .prog(prog),
     .carry_out(carry_out), .lft_op(lft_op_04[7:0]),
     .sp12_h_l(sp12_h_l_04[23:0]), .sp4_h_l(sp4_h_l_04[47:0]),
     .sp4_v_b(sp4_v_b_04[47:0]), .sp12_v_b({net199[0], net199[1],
     net199[2], net199[3], net199[4], net199[5], net199[6], net199[7],
     net199[8], net199[9], net199[10], net199[11], net199[12],
     net199[13], net199[14], net199[15], net199[16], net199[17],
     net199[18], net199[19], net199[20], net199[21], net199[22],
     net199[23]}), .sp12_h_r(sp12_h_r_04[23:0]),
     .sp4_h_r(sp4_h_r_04[47:0]), .sp12_v_t(sp12_v_t_04[23:0]),
     .sp4_v_t(sp4_v_t_04[47:0]), .sp4_r_v_b(sp4_r_v_b_04[47:0]),
     .wl(wl[63:48]), .top_op(top_op_04[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net191), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(tnr_op_04[7:0]),
     .tnl_op(tnl_op_04[7:0]));
ltile4_ice1f I_LT01 ( .cntl_cbit({net249[0], net249[1], net249[2],
     net249[3], net249[4], net249[5], net249[6], net249[7]}),
     .op_bot(lc_bot), .op_vic(net251), .prog(prog), .carry_out(net253),
     .lft_op(lft_op_01[7:0]), .sp12_h_l(sp12_h_l_01[23:0]),
     .sp4_h_l(sp4_h_l_01[47:0]), .sp4_v_b(sp4_v_b_01[47:0]),
     .sp12_v_b(sp12_v_b_01[23:0]), .sp12_h_r(sp12_h_r_01[23:0]),
     .sp4_h_r(sp4_h_r_01[47:0]), .sp12_v_t({net261[0], net261[1],
     net261[2], net261[3], net261[4], net261[5], net261[6], net261[7],
     net261[8], net261[9], net261[10], net261[11], net261[12],
     net261[13], net261[14], net261[15], net261[16], net261[17],
     net261[18], net261[19], net261[20], net261[21], net261[22],
     net261[23]}), .sp4_v_t(sp4_v_b_02[47:0]),
     .sp4_r_v_b(sp4_r_v_b_01[47:0]), .wl(wl[15:0]),
     .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4_ice1f I_LT02 ( .cntl_cbit({net280[0], net280[1], net280[2],
     net280[3], net280[4], net280[5], net280[6], net280[7]}),
     .op_bot(net251), .op_vic(net282), .prog(prog), .carry_out(net284),
     .lft_op(lft_op_02[7:0]), .sp12_h_l(sp12_h_l_02[23:0]),
     .sp4_h_l(sp4_h_l_02[47:0]), .sp4_v_b(sp4_v_b_02[47:0]),
     .sp12_v_b({net261[0], net261[1], net261[2], net261[3], net261[4],
     net261[5], net261[6], net261[7], net261[8], net261[9], net261[10],
     net261[11], net261[12], net261[13], net261[14], net261[15],
     net261[16], net261[17], net261[18], net261[19], net261[20],
     net261[21], net261[22], net261[23]}),
     .sp12_h_r(sp12_h_r_02[23:0]), .sp4_h_r(sp4_h_r_02[47:0]),
     .sp12_v_t({net292[0], net292[1], net292[2], net292[3], net292[4],
     net292[5], net292[6], net292[7], net292[8], net292[9], net292[10],
     net292[11], net292[12], net292[13], net292[14], net292[15],
     net292[16], net292[17], net292[18], net292[19], net292[20],
     net292[21], net292[22], net292[23]}), .sp4_v_t(sp4_v_b_03[47:0]),
     .sp4_r_v_b(sp4_r_v_b_02[47:0]), .wl(wl[31:16]),
     .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net253), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_resbot_40nm, View - schematic
// LAST TIME SAVED: Nov 16 16:07:51 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_sa_resbot_40nm ( bl_in, bl_out, in_dec, sa_ngate );
inout  bl_in, bl_out, in_dec;


input [4:1]  sa_ngate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



RNPPO_LP_pcell2460 R16 ( .B(gnd_), .MINUS(bl_in), .PLUS(bl_in));
RNPPO_LP_pcell2460 R7 ( .B(gnd_), .MINUS(net026), .PLUS(in_dec));
RNPPO_LP_pcell2460 R12 ( .B(gnd_), .MINUS(bl_in), .PLUS(bl_in));
RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(in_dec), .PLUS(bl_in));
RNPPO_LP_pcell2460 R9 ( .B(gnd_), .MINUS(bl_out), .PLUS(net132));
RNPPO_LP_pcell2460 R15 ( .B(gnd_), .MINUS(bl_in), .PLUS(bl_in));
RNPPO_LP_pcell2460 R8 ( .B(gnd_), .MINUS(net072), .PLUS(net026));
RNPPO_LP_pcell2460 R10 ( .B(gnd_), .MINUS(net132), .PLUS(net072));
N_11_LPHVT  M9 ( .D(net026), .B(GND_), .G(sa_ngate[2]), .S(gnd_));
N_11_LPHVT  M20 ( .D(in_dec), .B(GND_), .G(sa_ngate[1]), .S(gnd_));
N_11_LPHVT  M10 ( .D(net072), .B(GND_), .G(sa_ngate[3]), .S(gnd_));
N_11_LPHVT  M11 ( .D(net132), .B(GND_), .G(sa_ngate[4]), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_yp3_x8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:18 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_yp3_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M5_7_ ( .D(bl[7]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M5_6_ ( .D(bl[6]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M5_5_ ( .D(bl[5]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M5_4_ ( .D(bl[4]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M5_3_ ( .D(bl[3]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M5_2_ ( .D(bl[2]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M5_1_ ( .D(bl[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M5_0_ ( .D(bl[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
N_25_LP  M16 ( .D(bl[6]), .B(GND_), .G(yp3_25[6]), .S(bl_out));
N_25_LP  M18 ( .D(bl[4]), .B(GND_), .G(yp3_25[4]), .S(bl_out));
N_25_LP  M19 ( .D(bl[3]), .B(GND_), .G(yp3_25[3]), .S(bl_out));
N_25_LP  M26 ( .D(bl[0]), .B(GND_), .G(yp3_b_25[0]), .S(vblinhi_rde));
N_25_LP  M0 ( .D(bl[1]), .B(GND_), .G(yp3_b_25[1]), .S(vblinhi_rdo));
N_25_LP  M3 ( .D(bl[3]), .B(GND_), .G(yp3_b_25[3]), .S(vblinhi_rdo));
N_25_LP  M2 ( .D(bl[2]), .B(GND_), .G(yp3_b_25[2]), .S(vblinhi_rde));
N_25_LP  M4 ( .D(bl[4]), .B(GND_), .G(yp3_b_25[4]), .S(vblinhi_rde));
N_25_LP  M6 ( .D(bl[5]), .B(GND_), .G(yp3_b_25[5]), .S(vblinhi_rdo));
N_25_LP  M22 ( .D(bl[0]), .B(GND_), .G(yp3_25[0]), .S(bl_out));
N_25_LP  M20 ( .D(bl[2]), .B(GND_), .G(yp3_25[2]), .S(bl_out));
N_25_LP  M21 ( .D(bl[1]), .B(GND_), .G(yp3_25[1]), .S(bl_out));
N_25_LP  M8 ( .D(bl[7]), .B(GND_), .G(yp3_b_25[7]), .S(vblinhi_rdo));
N_25_LP  M17 ( .D(bl[5]), .B(GND_), .G(yp3_25[5]), .S(bl_out));
N_25_LP  M15 ( .D(bl[7]), .B(GND_), .G(yp3_25[7]), .S(bl_out));
N_25_LP  M7 ( .D(bl[6]), .B(GND_), .G(yp3_b_25[6]), .S(vblinhi_rde));

endmodule
// Library - ice384chip, Cell - quad_tr_ice384, View - schematic
// LAST TIME SAVED: Nov 30 14:43:58 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module quad_tr_ice384 ( bs_en_o, ceb_o, cf_r, cf_top_r,
     fabric_out_04_09, fabric_out_05_09, fabric_out_07_05,
     fabric_out_07_06, hiz_b_o, mode_o, padeb_r_t, padeb_t_r,
     padin_04_09a, padin_07_05a, pado_r_t, pado_t_r, r_o, sdo, shift_o,
     slf_op_04_05, slf_op_04_06, slf_op_04_07, slf_op_04_08,
     slf_op_04_09, slf_op_05_05, slf_op_06_05, slf_op_07_05, tclk_o,
     update_o, bl, pgate_r, reset_b_r, sp4_h_l_04_05, sp4_h_l_04_06,
     sp4_h_l_04_07, sp4_h_l_04_08, sp4_h_l_04_09, sp4_h_r_07_05,
     sp4_v_b_04_05, sp4_v_b_04_06, sp4_v_b_04_07, sp4_v_b_04_08,
     sp4_v_b_05_05, sp4_v_b_06_05, sp12_h_l_04_05, sp12_h_l_04_06,
     sp12_h_l_04_07, sp12_h_l_04_08, sp12_v_b_04_05, sp12_v_b_05_05,
     sp12_v_b_06_05, vdd_cntl_r, wl_r, bnl_op_04_05, bnl_op_05_05,
     bnl_op_06_05, bnl_op_07_05, bnr_op_04_05, bnr_op_05_05,
     bnr_op_06_05, bot_op_04_05, bot_op_05_05, bot_op_06_05, bs_en_i,
     carry_in_04_05, carry_in_05_05, carry_in_06_05, ceb_i, glb_in_4,
     glb_in_5, glb_in_6, glb_in_7, hiz_b_i, hold_r_t, hold_t_r,
     jtag_rowtest_mode_rowu3_b, last_rsr, lc_bot_04_05, lc_bot_05_05,
     lc_bot_06_05, lft_op_04_05, lft_op_04_06, lft_op_04_07,
     lft_op_04_08, mode_i, padin_r_t, padin_t_r, prog, purst, r_i, sdi,
     shift_i, tclk_i, tnl_op_04_08, update_i );
output  bs_en_o, ceb_o, fabric_out_04_09, fabric_out_05_09,
     fabric_out_07_05, fabric_out_07_06, hiz_b_o, mode_o, padin_04_09a,
     padin_07_05a, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, carry_in_04_05, carry_in_05_05, carry_in_06_05, ceb_i,
     hiz_b_i, hold_r_t, hold_t_r, jtag_rowtest_mode_rowu3_b,
     lc_bot_04_05, lc_bot_05_05, lc_bot_06_05, mode_i, prog, purst,
     r_i, sdi, shift_i, tclk_i, update_i;

output [15:8]  pado_r_t;
output [7:0]  slf_op_05_05;
output [15:8]  padeb_r_t;
output [7:0]  slf_op_04_05;
output [11:6]  padeb_t_r;
output [7:0]  slf_op_04_07;
output [3:0]  slf_op_04_09;
output [11:6]  pado_t_r;
output [7:0]  slf_op_04_06;
output [71:0]  cf_top_r;
output [7:0]  slf_op_06_05;
output [3:0]  slf_op_07_05;
output [7:0]  slf_op_04_08;
output [95:0]  cf_r;

inout [47:0]  sp4_h_l_04_07;
inout [23:0]  sp12_h_l_04_06;
inout [23:0]  sp12_v_b_05_05;
inout [23:0]  sp12_h_l_04_05;
inout [23:0]  sp12_h_l_04_07;
inout [47:0]  sp4_v_b_06_05;
inout [47:0]  sp4_v_b_05_05;
inout [47:0]  sp4_v_b_04_08;
inout [23:0]  sp12_h_l_04_08;
inout [47:0]  sp4_h_l_04_08;
inout [47:0]  sp4_v_b_04_07;
inout [47:0]  sp4_h_l_04_05;
inout [23:0]  sp12_v_b_06_05;
inout [47:0]  sp4_v_b_04_06;
inout [47:0]  sp4_v_b_04_05;
inout [47:0]  sp4_h_l_04_06;
inout [79:0]  wl_r;
inout [15:0]  sp4_h_l_04_09;
inout [15:0]  sp4_h_r_07_05;
inout [79:0]  pgate_r;
inout [79:0]  reset_b_r;
inout [179:0]  bl;
inout [79:0]  vdd_cntl_r;
inout [23:0]  sp12_v_b_04_05;

input [7:0]  bnr_op_06_05;
input [7:0]  bnr_op_05_05;
input [7:0]  glb_in_4;
input [7:0]  bnl_op_05_05;
input [7:0]  bot_op_06_05;
input [7:0]  bot_op_05_05;
input [7:0]  bnl_op_07_05;
input [7:0]  lft_op_04_06;
input [7:0]  bot_op_04_05;
input [3:3]  last_rsr;
input [7:0]  bnl_op_06_05;
input [7:0]  glb_in_5;
input [7:0]  lft_op_04_05;
input [7:0]  lft_op_04_07;
input [3:0]  tnl_op_04_08;
input [7:0]  bnr_op_04_05;
input [11:6]  padin_t_r;
input [7:0]  bnl_op_04_05;
input [7:0]  lft_op_04_08;
input [7:0]  glb_in_6;
input [15:8]  padin_r_t;
input [7:0]  glb_in_7;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [47:0]  net474;

wire  [23:0]  net469;

wire  [23:0]  net528;

wire  [23:0]  net471;

wire  [47:0]  net580;

wire  [47:0]  net538;

wire  [47:0]  net421;

wire  [47:0]  net475;

wire  [47:0]  net537;

wire  [47:0]  net481;

wire  [47:0]  net419;

wire  [7:0]  net452;

wire  [23:0]  net529;

wire  [23:0]  net414;

wire  [47:0]  net479;

wire  [23:0]  net415;

wire  [47:0]  net577;

wire  [23:0]  net472;

wire  [23:0]  net527;

wire  [7:0]  net393;

wire  [47:0]  net476;

wire  [47:0]  net578;

wire  [7:0]  net450;

wire  [23:0]  net563;

wire  [47:0]  net424;

wire  [7:0]  net403;

wire  [47:0]  net418;

wire  [47:0]  net536;

wire  [23:0]  net526;

wire  [23:0]  net470;

wire  [15:0]  net330;

wire  [47:0]  net562;

wire  [23:0]  net449;

wire  [47:0]  net417;

wire  [7:0]  net395;

wire  [23:0]  net413;

wire  [47:0]  net422;

wire  [47:0]  net505;

wire  [47:0]  net535;

wire  [47:0]  net581;

wire  [47:0]  net480;

wire  [47:0]  net478;

wire  [3:0]  slf_op_07_08;

wire  [23:0]  net412;

wire  [3:0]  slf_op_05_09;

wire  [47:0]  net448;

wire  [3:0]  slf_op_07_06;

wire  [23:0]  net506;

wire  [3:0]  slf_op_06_09;

wire  [7:0]  net460;

wire  [3:0]  slf_op_07_07;

wire  [47:0]  net423;



scan_buf_ice8p I409 ( .update_i(update_i), .tclk_i(net331),
     .shift_i(shift_i), .sdi(net307), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net372), .tclk_o(net373), .shift_o(net374),
     .sdo(net375), .r_o(net377), .mode_o(net380), .hiz_b_o(net381),
     .ceb_o(net392), .bs_en_o(net382));
io_rgt_top_1x4_ice384 I407 ( .shift(shift_i), .bs_en(bs_en_i),
     .mode(mode_i), .sdi(sdi), .hiz_b(hiz_b_i), .prog(prog),
     .hold(hold_r_t), .update(update_i), .r(r_i),
     .slf_op_07_06(slf_op_07_06[3:0]), .glb_netwk(glb_in_7[7:0]),
     .slf_op_07_05(slf_op_07_05[3:0]), .sdo(net307), .bl(bl[179:162]),
     .tclk(tclk_i), .reset_b(reset_b_r[63:0]),
     .tnl_op_07_08({slf_op_06_09[3], slf_op_06_09[2], slf_op_06_09[1],
     slf_op_06_09[0], slf_op_06_09[3], slf_op_06_09[2],
     slf_op_06_09[1], slf_op_06_09[0]}),
     .slf_op_07_07(slf_op_07_07[3:0]),
     .slf_op_07_08(slf_op_07_08[3:0]), .padeb(padeb_r_t[15:8]),
     .SP4_h_l_07_08({net535[0], net535[1], net535[2], net535[3],
     net535[4], net535[5], net535[6], net535[7], net535[8], net535[9],
     net535[10], net535[11], net535[12], net535[13], net535[14],
     net535[15], net535[16], net535[17], net535[18], net535[19],
     net535[20], net535[21], net535[22], net535[23], net535[24],
     net535[25], net535[26], net535[27], net535[28], net535[29],
     net535[30], net535[31], net535[32], net535[33], net535[34],
     net535[35], net535[36], net535[37], net535[38], net535[39],
     net535[40], net535[41], net535[42], net535[43], net535[44],
     net535[45], net535[46], net535[47]}), .SP4_h_l_07_06({net537[0],
     net537[1], net537[2], net537[3], net537[4], net537[5], net537[6],
     net537[7], net537[8], net537[9], net537[10], net537[11],
     net537[12], net537[13], net537[14], net537[15], net537[16],
     net537[17], net537[18], net537[19], net537[20], net537[21],
     net537[22], net537[23], net537[24], net537[25], net537[26],
     net537[27], net537[28], net537[29], net537[30], net537[31],
     net537[32], net537[33], net537[34], net537[35], net537[36],
     net537[37], net537[38], net537[39], net537[40], net537[41],
     net537[42], net537[43], net537[44], net537[45], net537[46],
     net537[47]}), .SP4_h_l_07_07({net536[0], net536[1], net536[2],
     net536[3], net536[4], net536[5], net536[6], net536[7], net536[8],
     net536[9], net536[10], net536[11], net536[12], net536[13],
     net536[14], net536[15], net536[16], net536[17], net536[18],
     net536[19], net536[20], net536[21], net536[22], net536[23],
     net536[24], net536[25], net536[26], net536[27], net536[28],
     net536[29], net536[30], net536[31], net536[32], net536[33],
     net536[34], net536[35], net536[36], net536[37], net536[38],
     net536[39], net536[40], net536[41], net536[42], net536[43],
     net536[44], net536[45], net536[46], net536[47]}),
     .SP4_h_l_07_05({net538[0], net538[1], net538[2], net538[3],
     net538[4], net538[5], net538[6], net538[7], net538[8], net538[9],
     net538[10], net538[11], net538[12], net538[13], net538[14],
     net538[15], net538[16], net538[17], net538[18], net538[19],
     net538[20], net538[21], net538[22], net538[23], net538[24],
     net538[25], net538[26], net538[27], net538[28], net538[29],
     net538[30], net538[31], net538[32], net538[33], net538[34],
     net538[35], net538[36], net538[37], net538[38], net538[39],
     net538[40], net538[41], net538[42], net538[43], net538[44],
     net538[45], net538[46], net538[47]}), .lft_op_07_07({net450[0],
     net450[1], net450[2], net450[3], net450[4], net450[5], net450[6],
     net450[7]}), .lft_op_07_08({net460[0], net460[1], net460[2],
     net460[3], net460[4], net460[5], net460[6], net460[7]}),
     .lft_op_07_05(slf_op_06_05[7:0]), .last_rsr(last_rsr[3]),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .wl(wl_r[63:0]), .cf_r(cf_r[95:0]), .vdd_cntl(vdd_cntl_r[63:0]),
     .pgate(pgate_r[63:0]), .padin(padin_r_t[15:8]),
     .pado(pado_r_t[15:8]), .sp4_v_t_07_08({net330[0], net330[1],
     net330[2], net330[3], net330[4], net330[5], net330[6], net330[7],
     net330[8], net330[9], net330[10], net330[11], net330[12],
     net330[13], net330[14], net330[15]}), .tclk_o(net331),
     .ceb(ceb_i), .fabric_out_07_06(fabric_out_07_06),
     .SP12_h_l_07_07({net527[0], net527[1], net527[2], net527[3],
     net527[4], net527[5], net527[6], net527[7], net527[8], net527[9],
     net527[10], net527[11], net527[12], net527[13], net527[14],
     net527[15], net527[16], net527[17], net527[18], net527[19],
     net527[20], net527[21], net527[22], net527[23]}),
     .SP12_h_l_07_08({net526[0], net526[1], net526[2], net526[3],
     net526[4], net526[5], net526[6], net526[7], net526[8], net526[9],
     net526[10], net526[11], net526[12], net526[13], net526[14],
     net526[15], net526[16], net526[17], net526[18], net526[19],
     net526[20], net526[21], net526[22], net526[23]}),
     .SP12_h_l_07_06({net528[0], net528[1], net528[2], net528[3],
     net528[4], net528[5], net528[6], net528[7], net528[8], net528[9],
     net528[10], net528[11], net528[12], net528[13], net528[14],
     net528[15], net528[16], net528[17], net528[18], net528[19],
     net528[20], net528[21], net528[22], net528[23]}),
     .bnl_op_07_05(bnl_op_07_05[7:0]), .SP12_h_l_07_05({net529[0],
     net529[1], net529[2], net529[3], net529[4], net529[5], net529[6],
     net529[7], net529[8], net529[9], net529[10], net529[11],
     net529[12], net529[13], net529[14], net529[15], net529[16],
     net529[17], net529[18], net529[19], net529[20], net529[21],
     net529[22], net529[23]}), .lft_op_07_06({net452[0], net452[1],
     net452[2], net452[3], net452[4], net452[5], net452[6],
     net452[7]}), .sp4_v_b_07_05(sp4_h_r_07_05[15:0]),
     .fabric_out_07_05(fabric_out_07_05));
io_top_rgt_1x3_ice384 I398 ( .hold_t_r(hold_t_r),
     .sp12_v_b_04_09({net449[0], net449[1], net449[2], net449[3],
     net449[4], net449[5], net449[6], net449[7], net449[8], net449[9],
     net449[10], net449[11], net449[12], net449[13], net449[14],
     net449[15], net449[16], net449[17], net449[18], net449[19],
     net449[20], net449[21], net449[22], net449[23]}),
     .lft_op_05_09({net403[0], net403[1], net403[2], net403[3],
     net403[4], net403[5], net403[6], net403[7]}),
     .sp4_v_b_06_09({net562[0], net562[1], net562[2], net562[3],
     net562[4], net562[5], net562[6], net562[7], net562[8], net562[9],
     net562[10], net562[11], net562[12], net562[13], net562[14],
     net562[15], net562[16], net562[17], net562[18], net562[19],
     net562[20], net562[21], net562[22], net562[23], net562[24],
     net562[25], net562[26], net562[27], net562[28], net562[29],
     net562[30], net562[31], net562[32], net562[33], net562[34],
     net562[35], net562[36], net562[37], net562[38], net562[39],
     net562[40], net562[41], net562[42], net562[43], net562[44],
     net562[45], net562[46], net562[47]}),
     .slf_op_06_09(slf_op_06_09[3:0]), .glb_net_06(glb_in_6[7:0]),
     .sp12_v_b_05_09({net506[0], net506[1], net506[2], net506[3],
     net506[4], net506[5], net506[6], net506[7], net506[8], net506[9],
     net506[10], net506[11], net506[12], net506[13], net506[14],
     net506[15], net506[16], net506[17], net506[18], net506[19],
     net506[20], net506[21], net506[22], net506[23]}),
     .sp4_v_b_04_09({net448[0], net448[1], net448[2], net448[3],
     net448[4], net448[5], net448[6], net448[7], net448[8], net448[9],
     net448[10], net448[11], net448[12], net448[13], net448[14],
     net448[15], net448[16], net448[17], net448[18], net448[19],
     net448[20], net448[21], net448[22], net448[23], net448[24],
     net448[25], net448[26], net448[27], net448[28], net448[29],
     net448[30], net448[31], net448[32], net448[33], net448[34],
     net448[35], net448[36], net448[37], net448[38], net448[39],
     net448[40], net448[41], net448[42], net448[43], net448[44],
     net448[45], net448[46], net448[47]}),
     .fabric_out_04_09(fabric_out_04_09),
     .lft_op_04_09(slf_op_04_08[7:0]),
     .sp4_h_l_04_09(sp4_h_l_04_09[15:0]),
     .bnl_op_04_09(lft_op_04_08[7:0]), .sp4_v_b_05_09({net505[0],
     net505[1], net505[2], net505[3], net505[4], net505[5], net505[6],
     net505[7], net505[8], net505[9], net505[10], net505[11],
     net505[12], net505[13], net505[14], net505[15], net505[16],
     net505[17], net505[18], net505[19], net505[20], net505[21],
     net505[22], net505[23], net505[24], net505[25], net505[26],
     net505[27], net505[28], net505[29], net505[30], net505[31],
     net505[32], net505[33], net505[34], net505[35], net505[36],
     net505[37], net505[38], net505[39], net505[40], net505[41],
     net505[42], net505[43], net505[44], net505[45], net505[46],
     net505[47]}), .glb_net_05(glb_in_5[7:0]),
     .lft_op_06_09({net460[0], net460[1], net460[2], net460[3],
     net460[4], net460[5], net460[6], net460[7]}),
     .glb_net_04(glb_in_4[7:0]), .sp12_v_b_06_09({net563[0], net563[1],
     net563[2], net563[3], net563[4], net563[5], net563[6], net563[7],
     net563[8], net563[9], net563[10], net563[11], net563[12],
     net563[13], net563[14], net563[15], net563[16], net563[17],
     net563[18], net563[19], net563[20], net563[21], net563[22],
     net563[23]}), .slf_op_05_09(slf_op_05_09[3:0]), .bl_04(bl[53:0]),
     .slf_op_04_09(slf_op_04_09[3:0]), .bl_05(bl[107:54]),
     .bl_06(bl[161:108]), .fabric_out_05_09(fabric_out_05_09),
     .cf_top_r(cf_top_r[71:0]), .padeb_t_r(padeb_t_r[11:6]),
     .sp4_h_r_06_09({net330[0], net330[1], net330[2], net330[3],
     net330[4], net330[5], net330[6], net330[7], net330[8], net330[9],
     net330[10], net330[11], net330[12], net330[13], net330[14],
     net330[15]}), .pado_t_r(pado_t_r[11:6]),
     .padin_t_r(padin_t_r[11:6]), .bnr_op_06_09({slf_op_07_08[3],
     slf_op_07_08[2], slf_op_07_08[1], slf_op_07_08[0],
     slf_op_07_08[3], slf_op_07_08[2], slf_op_07_08[1],
     slf_op_07_08[0]}), .wl_l({wl_r[78], wl_r[79], wl_r[77], wl_r[76],
     wl_r[74], wl_r[75], wl_r[73], wl_r[72], wl_r[70], wl_r[71],
     wl_r[69], wl_r[68], wl_r[66], wl_r[67], wl_r[65], wl_r[64]}),
     .vdd_cntl_l({vdd_cntl_r[78], vdd_cntl_r[79], vdd_cntl_r[77],
     vdd_cntl_r[76], vdd_cntl_r[74], vdd_cntl_r[75], vdd_cntl_r[73],
     vdd_cntl_r[72], vdd_cntl_r[70], vdd_cntl_r[71], vdd_cntl_r[69],
     vdd_cntl_r[68], vdd_cntl_r[66], vdd_cntl_r[67], vdd_cntl_r[65],
     vdd_cntl_r[64]}), .update_i(net372), .tclk_i(net373),
     .shift_i(net374), .sdi(net375), .reset_l({reset_b_r[78],
     reset_b_r[79], reset_b_r[77], reset_b_r[76], reset_b_r[74],
     reset_b_r[75], reset_b_r[73], reset_b_r[72], reset_b_r[70],
     reset_b_r[71], reset_b_r[69], reset_b_r[68], reset_b_r[66],
     reset_b_r[67], reset_b_r[65], reset_b_r[64]}), .r_i(net377),
     .prog(prog), .pgate_l({pgate_r[78], pgate_r[79], pgate_r[77],
     pgate_r[76], pgate_r[74], pgate_r[75], pgate_r[73], pgate_r[72],
     pgate_r[70], pgate_r[71], pgate_r[69], pgate_r[68], pgate_r[66],
     pgate_r[67], pgate_r[65], pgate_r[64]}), .mode_i(net380),
     .hiz_b_i(net381), .bs_en_i(net382), .update_o(update_o),
     .tclk_o(tclk_o), .shift_o(shift_o), .sdo(sdo), .r_o(r_o),
     .mode_o(mode_o), .hiz_b_o(hiz_b_o), .bs_en_o(bs_en_o),
     .ceb_o(ceb_o), .ceb_i(net392));
lt_1x4_top_ice384 I394 ( .rgt_op_03({net393[0], net393[1], net393[2],
     net393[3], net393[4], net393[5], net393[6], net393[7]}),
     .slf_op_02(slf_op_04_06[7:0]), .rgt_op_02({net395[0], net395[1],
     net395[2], net395[3], net395[4], net395[5], net395[6],
     net395[7]}), .rgt_op_01(slf_op_05_05[7:0]), .purst(purst),
     .prog(prog), .lft_op_04(lft_op_04_08[7:0]),
     .lft_op_03(lft_op_04_07[7:0]), .lft_op_02(lft_op_04_06[7:0]),
     .lft_op_01(lft_op_04_05[7:0]), .rgt_op_04({net403[0], net403[1],
     net403[2], net403[3], net403[4], net403[5], net403[6],
     net403[7]}), .carry_in(carry_in_04_05),
     .bnl_op_01(bnl_op_04_05[7:0]), .slf_op_04(slf_op_04_08[7:0]),
     .slf_op_03(slf_op_04_07[7:0]), .slf_op_01(slf_op_04_05[7:0]),
     .sp4_h_l_04(sp4_h_l_04_08[47:0]), .carry_out(net410),
     .vdd_cntl(vdd_cntl_r[63:0]), .sp12_h_r_04({net412[0], net412[1],
     net412[2], net412[3], net412[4], net412[5], net412[6], net412[7],
     net412[8], net412[9], net412[10], net412[11], net412[12],
     net412[13], net412[14], net412[15], net412[16], net412[17],
     net412[18], net412[19], net412[20], net412[21], net412[22],
     net412[23]}), .sp12_h_r_03({net413[0], net413[1], net413[2],
     net413[3], net413[4], net413[5], net413[6], net413[7], net413[8],
     net413[9], net413[10], net413[11], net413[12], net413[13],
     net413[14], net413[15], net413[16], net413[17], net413[18],
     net413[19], net413[20], net413[21], net413[22], net413[23]}),
     .sp12_h_r_02({net414[0], net414[1], net414[2], net414[3],
     net414[4], net414[5], net414[6], net414[7], net414[8], net414[9],
     net414[10], net414[11], net414[12], net414[13], net414[14],
     net414[15], net414[16], net414[17], net414[18], net414[19],
     net414[20], net414[21], net414[22], net414[23]}),
     .sp12_h_r_01({net415[0], net415[1], net415[2], net415[3],
     net415[4], net415[5], net415[6], net415[7], net415[8], net415[9],
     net415[10], net415[11], net415[12], net415[13], net415[14],
     net415[15], net415[16], net415[17], net415[18], net415[19],
     net415[20], net415[21], net415[22], net415[23]}),
     .sp4_v_b_01(sp4_v_b_04_05[47:0]), .sp4_r_v_b_04({net417[0],
     net417[1], net417[2], net417[3], net417[4], net417[5], net417[6],
     net417[7], net417[8], net417[9], net417[10], net417[11],
     net417[12], net417[13], net417[14], net417[15], net417[16],
     net417[17], net417[18], net417[19], net417[20], net417[21],
     net417[22], net417[23], net417[24], net417[25], net417[26],
     net417[27], net417[28], net417[29], net417[30], net417[31],
     net417[32], net417[33], net417[34], net417[35], net417[36],
     net417[37], net417[38], net417[39], net417[40], net417[41],
     net417[42], net417[43], net417[44], net417[45], net417[46],
     net417[47]}), .sp4_r_v_b_03({net418[0], net418[1], net418[2],
     net418[3], net418[4], net418[5], net418[6], net418[7], net418[8],
     net418[9], net418[10], net418[11], net418[12], net418[13],
     net418[14], net418[15], net418[16], net418[17], net418[18],
     net418[19], net418[20], net418[21], net418[22], net418[23],
     net418[24], net418[25], net418[26], net418[27], net418[28],
     net418[29], net418[30], net418[31], net418[32], net418[33],
     net418[34], net418[35], net418[36], net418[37], net418[38],
     net418[39], net418[40], net418[41], net418[42], net418[43],
     net418[44], net418[45], net418[46], net418[47]}),
     .sp4_r_v_b_02({net419[0], net419[1], net419[2], net419[3],
     net419[4], net419[5], net419[6], net419[7], net419[8], net419[9],
     net419[10], net419[11], net419[12], net419[13], net419[14],
     net419[15], net419[16], net419[17], net419[18], net419[19],
     net419[20], net419[21], net419[22], net419[23], net419[24],
     net419[25], net419[26], net419[27], net419[28], net419[29],
     net419[30], net419[31], net419[32], net419[33], net419[34],
     net419[35], net419[36], net419[37], net419[38], net419[39],
     net419[40], net419[41], net419[42], net419[43], net419[44],
     net419[45], net419[46], net419[47]}),
     .sp4_r_v_b_01(sp4_v_b_05_05[47:0]), .sp4_h_r_04({net421[0],
     net421[1], net421[2], net421[3], net421[4], net421[5], net421[6],
     net421[7], net421[8], net421[9], net421[10], net421[11],
     net421[12], net421[13], net421[14], net421[15], net421[16],
     net421[17], net421[18], net421[19], net421[20], net421[21],
     net421[22], net421[23], net421[24], net421[25], net421[26],
     net421[27], net421[28], net421[29], net421[30], net421[31],
     net421[32], net421[33], net421[34], net421[35], net421[36],
     net421[37], net421[38], net421[39], net421[40], net421[41],
     net421[42], net421[43], net421[44], net421[45], net421[46],
     net421[47]}), .sp4_h_r_03({net422[0], net422[1], net422[2],
     net422[3], net422[4], net422[5], net422[6], net422[7], net422[8],
     net422[9], net422[10], net422[11], net422[12], net422[13],
     net422[14], net422[15], net422[16], net422[17], net422[18],
     net422[19], net422[20], net422[21], net422[22], net422[23],
     net422[24], net422[25], net422[26], net422[27], net422[28],
     net422[29], net422[30], net422[31], net422[32], net422[33],
     net422[34], net422[35], net422[36], net422[37], net422[38],
     net422[39], net422[40], net422[41], net422[42], net422[43],
     net422[44], net422[45], net422[46], net422[47]}),
     .sp4_h_r_02({net423[0], net423[1], net423[2], net423[3],
     net423[4], net423[5], net423[6], net423[7], net423[8], net423[9],
     net423[10], net423[11], net423[12], net423[13], net423[14],
     net423[15], net423[16], net423[17], net423[18], net423[19],
     net423[20], net423[21], net423[22], net423[23], net423[24],
     net423[25], net423[26], net423[27], net423[28], net423[29],
     net423[30], net423[31], net423[32], net423[33], net423[34],
     net423[35], net423[36], net423[37], net423[38], net423[39],
     net423[40], net423[41], net423[42], net423[43], net423[44],
     net423[45], net423[46], net423[47]}), .sp4_h_r_01({net424[0],
     net424[1], net424[2], net424[3], net424[4], net424[5], net424[6],
     net424[7], net424[8], net424[9], net424[10], net424[11],
     net424[12], net424[13], net424[14], net424[15], net424[16],
     net424[17], net424[18], net424[19], net424[20], net424[21],
     net424[22], net424[23], net424[24], net424[25], net424[26],
     net424[27], net424[28], net424[29], net424[30], net424[31],
     net424[32], net424[33], net424[34], net424[35], net424[36],
     net424[37], net424[38], net424[39], net424[40], net424[41],
     net424[42], net424[43], net424[44], net424[45], net424[46],
     net424[47]}), .sp4_h_l_03(sp4_h_l_04_07[47:0]),
     .sp4_h_l_02(sp4_h_l_04_06[47:0]),
     .sp4_h_l_01(sp4_h_l_04_05[47:0]), .bl(bl[53:0]),
     .bot_op_01(bot_op_04_05[7:0]), .sp12_h_l_01(sp12_h_l_04_05[23:0]),
     .sp12_h_l_02(sp12_h_l_04_06[23:0]),
     .sp12_h_l_03(sp12_h_l_04_07[23:0]),
     .sp12_h_l_04(sp12_h_l_04_08[23:0]),
     .sp4_v_b_04(sp4_v_b_04_08[47:0]),
     .sp4_v_b_03(sp4_v_b_04_07[47:0]),
     .sp4_v_b_02(sp4_v_b_04_06[47:0]), .bnr_op_01(bnr_op_04_05[7:0]),
     .tnr_op_04({slf_op_05_09[3], slf_op_05_09[2], slf_op_05_09[1],
     slf_op_05_09[0], slf_op_05_09[3], slf_op_05_09[2],
     slf_op_05_09[1], slf_op_05_09[0]}), .glb_netwk(glb_in_4[7:0]),
     .tnl_op_04({tnl_op_04_08[3], tnl_op_04_08[2], tnl_op_04_08[1],
     tnl_op_04_08[0], tnl_op_04_08[3], tnl_op_04_08[2],
     tnl_op_04_08[1], tnl_op_04_08[0]}), .pgate(pgate_r[63:0]),
     .reset_b(reset_b_r[63:0]), .wl(wl_r[63:0]),
     .top_op_04({slf_op_04_09[3], slf_op_04_09[2], slf_op_04_09[1],
     slf_op_04_09[0], slf_op_04_09[3], slf_op_04_09[2],
     slf_op_04_09[1], slf_op_04_09[0]}), .lc_bot(lc_bot_04_05),
     .op_vic(net446), .sp12_v_b_01(sp12_v_b_04_05[23:0]),
     .sp4_v_t_04({net448[0], net448[1], net448[2], net448[3],
     net448[4], net448[5], net448[6], net448[7], net448[8], net448[9],
     net448[10], net448[11], net448[12], net448[13], net448[14],
     net448[15], net448[16], net448[17], net448[18], net448[19],
     net448[20], net448[21], net448[22], net448[23], net448[24],
     net448[25], net448[26], net448[27], net448[28], net448[29],
     net448[30], net448[31], net448[32], net448[33], net448[34],
     net448[35], net448[36], net448[37], net448[38], net448[39],
     net448[40], net448[41], net448[42], net448[43], net448[44],
     net448[45], net448[46], net448[47]}), .sp12_v_t_04({net449[0],
     net449[1], net449[2], net449[3], net449[4], net449[5], net449[6],
     net449[7], net449[8], net449[9], net449[10], net449[11],
     net449[12], net449[13], net449[14], net449[15], net449[16],
     net449[17], net449[18], net449[19], net449[20], net449[21],
     net449[22], net449[23]}));
lt_1x4_top_ice384 I399 ( .rgt_op_03({net450[0], net450[1], net450[2],
     net450[3], net450[4], net450[5], net450[6], net450[7]}),
     .slf_op_02({net395[0], net395[1], net395[2], net395[3], net395[4],
     net395[5], net395[6], net395[7]}), .rgt_op_02({net452[0],
     net452[1], net452[2], net452[3], net452[4], net452[5], net452[6],
     net452[7]}), .rgt_op_01(slf_op_06_05[7:0]), .purst(purst),
     .prog(prog), .lft_op_04(slf_op_04_08[7:0]),
     .lft_op_03(slf_op_04_07[7:0]), .lft_op_02(slf_op_04_06[7:0]),
     .lft_op_01(slf_op_04_05[7:0]), .rgt_op_04({net460[0], net460[1],
     net460[2], net460[3], net460[4], net460[5], net460[6],
     net460[7]}), .carry_in(carry_in_05_05),
     .bnl_op_01(bnl_op_05_05[7:0]), .slf_op_04({net403[0], net403[1],
     net403[2], net403[3], net403[4], net403[5], net403[6],
     net403[7]}), .slf_op_03({net393[0], net393[1], net393[2],
     net393[3], net393[4], net393[5], net393[6], net393[7]}),
     .slf_op_01(slf_op_05_05[7:0]), .sp4_h_l_04({net421[0], net421[1],
     net421[2], net421[3], net421[4], net421[5], net421[6], net421[7],
     net421[8], net421[9], net421[10], net421[11], net421[12],
     net421[13], net421[14], net421[15], net421[16], net421[17],
     net421[18], net421[19], net421[20], net421[21], net421[22],
     net421[23], net421[24], net421[25], net421[26], net421[27],
     net421[28], net421[29], net421[30], net421[31], net421[32],
     net421[33], net421[34], net421[35], net421[36], net421[37],
     net421[38], net421[39], net421[40], net421[41], net421[42],
     net421[43], net421[44], net421[45], net421[46], net421[47]}),
     .carry_out(net467), .vdd_cntl(vdd_cntl_r[63:0]),
     .sp12_h_r_04({net469[0], net469[1], net469[2], net469[3],
     net469[4], net469[5], net469[6], net469[7], net469[8], net469[9],
     net469[10], net469[11], net469[12], net469[13], net469[14],
     net469[15], net469[16], net469[17], net469[18], net469[19],
     net469[20], net469[21], net469[22], net469[23]}),
     .sp12_h_r_03({net470[0], net470[1], net470[2], net470[3],
     net470[4], net470[5], net470[6], net470[7], net470[8], net470[9],
     net470[10], net470[11], net470[12], net470[13], net470[14],
     net470[15], net470[16], net470[17], net470[18], net470[19],
     net470[20], net470[21], net470[22], net470[23]}),
     .sp12_h_r_02({net471[0], net471[1], net471[2], net471[3],
     net471[4], net471[5], net471[6], net471[7], net471[8], net471[9],
     net471[10], net471[11], net471[12], net471[13], net471[14],
     net471[15], net471[16], net471[17], net471[18], net471[19],
     net471[20], net471[21], net471[22], net471[23]}),
     .sp12_h_r_01({net472[0], net472[1], net472[2], net472[3],
     net472[4], net472[5], net472[6], net472[7], net472[8], net472[9],
     net472[10], net472[11], net472[12], net472[13], net472[14],
     net472[15], net472[16], net472[17], net472[18], net472[19],
     net472[20], net472[21], net472[22], net472[23]}),
     .sp4_v_b_01(sp4_v_b_05_05[47:0]), .sp4_r_v_b_04({net474[0],
     net474[1], net474[2], net474[3], net474[4], net474[5], net474[6],
     net474[7], net474[8], net474[9], net474[10], net474[11],
     net474[12], net474[13], net474[14], net474[15], net474[16],
     net474[17], net474[18], net474[19], net474[20], net474[21],
     net474[22], net474[23], net474[24], net474[25], net474[26],
     net474[27], net474[28], net474[29], net474[30], net474[31],
     net474[32], net474[33], net474[34], net474[35], net474[36],
     net474[37], net474[38], net474[39], net474[40], net474[41],
     net474[42], net474[43], net474[44], net474[45], net474[46],
     net474[47]}), .sp4_r_v_b_03({net475[0], net475[1], net475[2],
     net475[3], net475[4], net475[5], net475[6], net475[7], net475[8],
     net475[9], net475[10], net475[11], net475[12], net475[13],
     net475[14], net475[15], net475[16], net475[17], net475[18],
     net475[19], net475[20], net475[21], net475[22], net475[23],
     net475[24], net475[25], net475[26], net475[27], net475[28],
     net475[29], net475[30], net475[31], net475[32], net475[33],
     net475[34], net475[35], net475[36], net475[37], net475[38],
     net475[39], net475[40], net475[41], net475[42], net475[43],
     net475[44], net475[45], net475[46], net475[47]}),
     .sp4_r_v_b_02({net476[0], net476[1], net476[2], net476[3],
     net476[4], net476[5], net476[6], net476[7], net476[8], net476[9],
     net476[10], net476[11], net476[12], net476[13], net476[14],
     net476[15], net476[16], net476[17], net476[18], net476[19],
     net476[20], net476[21], net476[22], net476[23], net476[24],
     net476[25], net476[26], net476[27], net476[28], net476[29],
     net476[30], net476[31], net476[32], net476[33], net476[34],
     net476[35], net476[36], net476[37], net476[38], net476[39],
     net476[40], net476[41], net476[42], net476[43], net476[44],
     net476[45], net476[46], net476[47]}),
     .sp4_r_v_b_01(sp4_v_b_06_05[47:0]), .sp4_h_r_04({net478[0],
     net478[1], net478[2], net478[3], net478[4], net478[5], net478[6],
     net478[7], net478[8], net478[9], net478[10], net478[11],
     net478[12], net478[13], net478[14], net478[15], net478[16],
     net478[17], net478[18], net478[19], net478[20], net478[21],
     net478[22], net478[23], net478[24], net478[25], net478[26],
     net478[27], net478[28], net478[29], net478[30], net478[31],
     net478[32], net478[33], net478[34], net478[35], net478[36],
     net478[37], net478[38], net478[39], net478[40], net478[41],
     net478[42], net478[43], net478[44], net478[45], net478[46],
     net478[47]}), .sp4_h_r_03({net479[0], net479[1], net479[2],
     net479[3], net479[4], net479[5], net479[6], net479[7], net479[8],
     net479[9], net479[10], net479[11], net479[12], net479[13],
     net479[14], net479[15], net479[16], net479[17], net479[18],
     net479[19], net479[20], net479[21], net479[22], net479[23],
     net479[24], net479[25], net479[26], net479[27], net479[28],
     net479[29], net479[30], net479[31], net479[32], net479[33],
     net479[34], net479[35], net479[36], net479[37], net479[38],
     net479[39], net479[40], net479[41], net479[42], net479[43],
     net479[44], net479[45], net479[46], net479[47]}),
     .sp4_h_r_02({net480[0], net480[1], net480[2], net480[3],
     net480[4], net480[5], net480[6], net480[7], net480[8], net480[9],
     net480[10], net480[11], net480[12], net480[13], net480[14],
     net480[15], net480[16], net480[17], net480[18], net480[19],
     net480[20], net480[21], net480[22], net480[23], net480[24],
     net480[25], net480[26], net480[27], net480[28], net480[29],
     net480[30], net480[31], net480[32], net480[33], net480[34],
     net480[35], net480[36], net480[37], net480[38], net480[39],
     net480[40], net480[41], net480[42], net480[43], net480[44],
     net480[45], net480[46], net480[47]}), .sp4_h_r_01({net481[0],
     net481[1], net481[2], net481[3], net481[4], net481[5], net481[6],
     net481[7], net481[8], net481[9], net481[10], net481[11],
     net481[12], net481[13], net481[14], net481[15], net481[16],
     net481[17], net481[18], net481[19], net481[20], net481[21],
     net481[22], net481[23], net481[24], net481[25], net481[26],
     net481[27], net481[28], net481[29], net481[30], net481[31],
     net481[32], net481[33], net481[34], net481[35], net481[36],
     net481[37], net481[38], net481[39], net481[40], net481[41],
     net481[42], net481[43], net481[44], net481[45], net481[46],
     net481[47]}), .sp4_h_l_03({net422[0], net422[1], net422[2],
     net422[3], net422[4], net422[5], net422[6], net422[7], net422[8],
     net422[9], net422[10], net422[11], net422[12], net422[13],
     net422[14], net422[15], net422[16], net422[17], net422[18],
     net422[19], net422[20], net422[21], net422[22], net422[23],
     net422[24], net422[25], net422[26], net422[27], net422[28],
     net422[29], net422[30], net422[31], net422[32], net422[33],
     net422[34], net422[35], net422[36], net422[37], net422[38],
     net422[39], net422[40], net422[41], net422[42], net422[43],
     net422[44], net422[45], net422[46], net422[47]}),
     .sp4_h_l_02({net423[0], net423[1], net423[2], net423[3],
     net423[4], net423[5], net423[6], net423[7], net423[8], net423[9],
     net423[10], net423[11], net423[12], net423[13], net423[14],
     net423[15], net423[16], net423[17], net423[18], net423[19],
     net423[20], net423[21], net423[22], net423[23], net423[24],
     net423[25], net423[26], net423[27], net423[28], net423[29],
     net423[30], net423[31], net423[32], net423[33], net423[34],
     net423[35], net423[36], net423[37], net423[38], net423[39],
     net423[40], net423[41], net423[42], net423[43], net423[44],
     net423[45], net423[46], net423[47]}), .sp4_h_l_01({net424[0],
     net424[1], net424[2], net424[3], net424[4], net424[5], net424[6],
     net424[7], net424[8], net424[9], net424[10], net424[11],
     net424[12], net424[13], net424[14], net424[15], net424[16],
     net424[17], net424[18], net424[19], net424[20], net424[21],
     net424[22], net424[23], net424[24], net424[25], net424[26],
     net424[27], net424[28], net424[29], net424[30], net424[31],
     net424[32], net424[33], net424[34], net424[35], net424[36],
     net424[37], net424[38], net424[39], net424[40], net424[41],
     net424[42], net424[43], net424[44], net424[45], net424[46],
     net424[47]}), .bl(bl[107:54]), .bot_op_01(bot_op_05_05[7:0]),
     .sp12_h_l_01({net415[0], net415[1], net415[2], net415[3],
     net415[4], net415[5], net415[6], net415[7], net415[8], net415[9],
     net415[10], net415[11], net415[12], net415[13], net415[14],
     net415[15], net415[16], net415[17], net415[18], net415[19],
     net415[20], net415[21], net415[22], net415[23]}),
     .sp12_h_l_02({net414[0], net414[1], net414[2], net414[3],
     net414[4], net414[5], net414[6], net414[7], net414[8], net414[9],
     net414[10], net414[11], net414[12], net414[13], net414[14],
     net414[15], net414[16], net414[17], net414[18], net414[19],
     net414[20], net414[21], net414[22], net414[23]}),
     .sp12_h_l_03({net413[0], net413[1], net413[2], net413[3],
     net413[4], net413[5], net413[6], net413[7], net413[8], net413[9],
     net413[10], net413[11], net413[12], net413[13], net413[14],
     net413[15], net413[16], net413[17], net413[18], net413[19],
     net413[20], net413[21], net413[22], net413[23]}),
     .sp12_h_l_04({net412[0], net412[1], net412[2], net412[3],
     net412[4], net412[5], net412[6], net412[7], net412[8], net412[9],
     net412[10], net412[11], net412[12], net412[13], net412[14],
     net412[15], net412[16], net412[17], net412[18], net412[19],
     net412[20], net412[21], net412[22], net412[23]}),
     .sp4_v_b_04({net417[0], net417[1], net417[2], net417[3],
     net417[4], net417[5], net417[6], net417[7], net417[8], net417[9],
     net417[10], net417[11], net417[12], net417[13], net417[14],
     net417[15], net417[16], net417[17], net417[18], net417[19],
     net417[20], net417[21], net417[22], net417[23], net417[24],
     net417[25], net417[26], net417[27], net417[28], net417[29],
     net417[30], net417[31], net417[32], net417[33], net417[34],
     net417[35], net417[36], net417[37], net417[38], net417[39],
     net417[40], net417[41], net417[42], net417[43], net417[44],
     net417[45], net417[46], net417[47]}), .sp4_v_b_03({net418[0],
     net418[1], net418[2], net418[3], net418[4], net418[5], net418[6],
     net418[7], net418[8], net418[9], net418[10], net418[11],
     net418[12], net418[13], net418[14], net418[15], net418[16],
     net418[17], net418[18], net418[19], net418[20], net418[21],
     net418[22], net418[23], net418[24], net418[25], net418[26],
     net418[27], net418[28], net418[29], net418[30], net418[31],
     net418[32], net418[33], net418[34], net418[35], net418[36],
     net418[37], net418[38], net418[39], net418[40], net418[41],
     net418[42], net418[43], net418[44], net418[45], net418[46],
     net418[47]}), .sp4_v_b_02({net419[0], net419[1], net419[2],
     net419[3], net419[4], net419[5], net419[6], net419[7], net419[8],
     net419[9], net419[10], net419[11], net419[12], net419[13],
     net419[14], net419[15], net419[16], net419[17], net419[18],
     net419[19], net419[20], net419[21], net419[22], net419[23],
     net419[24], net419[25], net419[26], net419[27], net419[28],
     net419[29], net419[30], net419[31], net419[32], net419[33],
     net419[34], net419[35], net419[36], net419[37], net419[38],
     net419[39], net419[40], net419[41], net419[42], net419[43],
     net419[44], net419[45], net419[46], net419[47]}),
     .bnr_op_01(bnr_op_05_05[7:0]), .tnr_op_04({slf_op_06_09[3],
     slf_op_06_09[2], slf_op_06_09[1], slf_op_06_09[0],
     slf_op_06_09[3], slf_op_06_09[2], slf_op_06_09[1],
     slf_op_06_09[0]}), .glb_netwk(glb_in_5[7:0]),
     .tnl_op_04({slf_op_04_09[3], slf_op_04_09[2], slf_op_04_09[1],
     slf_op_04_09[0], slf_op_04_09[3], slf_op_04_09[2],
     slf_op_04_09[1], slf_op_04_09[0]}), .pgate(pgate_r[63:0]),
     .reset_b(reset_b_r[63:0]), .wl(wl_r[63:0]),
     .top_op_04({slf_op_05_09[3], slf_op_05_09[2], slf_op_05_09[1],
     slf_op_05_09[0], slf_op_05_09[3], slf_op_05_09[2],
     slf_op_05_09[1], slf_op_05_09[0]}), .lc_bot(lc_bot_05_05),
     .op_vic(net583), .sp12_v_b_01(sp12_v_b_05_05[23:0]),
     .sp4_v_t_04({net505[0], net505[1], net505[2], net505[3],
     net505[4], net505[5], net505[6], net505[7], net505[8], net505[9],
     net505[10], net505[11], net505[12], net505[13], net505[14],
     net505[15], net505[16], net505[17], net505[18], net505[19],
     net505[20], net505[21], net505[22], net505[23], net505[24],
     net505[25], net505[26], net505[27], net505[28], net505[29],
     net505[30], net505[31], net505[32], net505[33], net505[34],
     net505[35], net505[36], net505[37], net505[38], net505[39],
     net505[40], net505[41], net505[42], net505[43], net505[44],
     net505[45], net505[46], net505[47]}), .sp12_v_t_04({net506[0],
     net506[1], net506[2], net506[3], net506[4], net506[5], net506[6],
     net506[7], net506[8], net506[9], net506[10], net506[11],
     net506[12], net506[13], net506[14], net506[15], net506[16],
     net506[17], net506[18], net506[19], net506[20], net506[21],
     net506[22], net506[23]}));
lt_1x4_top_ice384 I400 ( .rgt_op_03({slf_op_07_07[3], slf_op_07_07[2],
     slf_op_07_07[1], slf_op_07_07[0], slf_op_07_07[3],
     slf_op_07_07[2], slf_op_07_07[1], slf_op_07_07[0]}),
     .slf_op_02({net452[0], net452[1], net452[2], net452[3], net452[4],
     net452[5], net452[6], net452[7]}), .rgt_op_02({slf_op_07_06[3],
     slf_op_07_06[2], slf_op_07_06[1], slf_op_07_06[0],
     slf_op_07_06[3], slf_op_07_06[2], slf_op_07_06[1],
     slf_op_07_06[0]}), .rgt_op_01({slf_op_07_05[3], slf_op_07_05[2],
     slf_op_07_05[1], slf_op_07_05[0], slf_op_07_05[3],
     slf_op_07_05[2], slf_op_07_05[1], slf_op_07_05[0]}),
     .purst(purst), .prog(prog), .lft_op_04({net403[0], net403[1],
     net403[2], net403[3], net403[4], net403[5], net403[6],
     net403[7]}), .lft_op_03({net393[0], net393[1], net393[2],
     net393[3], net393[4], net393[5], net393[6], net393[7]}),
     .lft_op_02({net395[0], net395[1], net395[2], net395[3], net395[4],
     net395[5], net395[6], net395[7]}), .lft_op_01(slf_op_05_05[7:0]),
     .rgt_op_04({slf_op_07_08[3], slf_op_07_08[2], slf_op_07_08[1],
     slf_op_07_08[0], slf_op_07_08[3], slf_op_07_08[2],
     slf_op_07_08[1], slf_op_07_08[0]}), .carry_in(carry_in_06_05),
     .bnl_op_01(bnl_op_06_05[7:0]), .slf_op_04({net460[0], net460[1],
     net460[2], net460[3], net460[4], net460[5], net460[6],
     net460[7]}), .slf_op_03({net450[0], net450[1], net450[2],
     net450[3], net450[4], net450[5], net450[6], net450[7]}),
     .slf_op_01(slf_op_06_05[7:0]), .sp4_h_l_04({net478[0], net478[1],
     net478[2], net478[3], net478[4], net478[5], net478[6], net478[7],
     net478[8], net478[9], net478[10], net478[11], net478[12],
     net478[13], net478[14], net478[15], net478[16], net478[17],
     net478[18], net478[19], net478[20], net478[21], net478[22],
     net478[23], net478[24], net478[25], net478[26], net478[27],
     net478[28], net478[29], net478[30], net478[31], net478[32],
     net478[33], net478[34], net478[35], net478[36], net478[37],
     net478[38], net478[39], net478[40], net478[41], net478[42],
     net478[43], net478[44], net478[45], net478[46], net478[47]}),
     .carry_out(net524), .vdd_cntl(vdd_cntl_r[63:0]),
     .sp12_h_r_04({net526[0], net526[1], net526[2], net526[3],
     net526[4], net526[5], net526[6], net526[7], net526[8], net526[9],
     net526[10], net526[11], net526[12], net526[13], net526[14],
     net526[15], net526[16], net526[17], net526[18], net526[19],
     net526[20], net526[21], net526[22], net526[23]}),
     .sp12_h_r_03({net527[0], net527[1], net527[2], net527[3],
     net527[4], net527[5], net527[6], net527[7], net527[8], net527[9],
     net527[10], net527[11], net527[12], net527[13], net527[14],
     net527[15], net527[16], net527[17], net527[18], net527[19],
     net527[20], net527[21], net527[22], net527[23]}),
     .sp12_h_r_02({net528[0], net528[1], net528[2], net528[3],
     net528[4], net528[5], net528[6], net528[7], net528[8], net528[9],
     net528[10], net528[11], net528[12], net528[13], net528[14],
     net528[15], net528[16], net528[17], net528[18], net528[19],
     net528[20], net528[21], net528[22], net528[23]}),
     .sp12_h_r_01({net529[0], net529[1], net529[2], net529[3],
     net529[4], net529[5], net529[6], net529[7], net529[8], net529[9],
     net529[10], net529[11], net529[12], net529[13], net529[14],
     net529[15], net529[16], net529[17], net529[18], net529[19],
     net529[20], net529[21], net529[22], net529[23]}),
     .sp4_v_b_01(sp4_v_b_06_05[47:0]), .sp4_r_v_b_04({net578[0],
     net578[1], net578[2], net578[3], net578[4], net578[5], net578[6],
     net578[7], net578[8], net578[9], net578[10], net578[11],
     net578[12], net578[13], net578[14], net578[15], net578[16],
     net578[17], net578[18], net578[19], net578[20], net578[21],
     net578[22], net578[23], net578[24], net578[25], net578[26],
     net578[27], net578[28], net578[29], net578[30], net578[31],
     net578[32], net578[33], net578[34], net578[35], net578[36],
     net578[37], net578[38], net578[39], net578[40], net578[41],
     net578[42], net578[43], net578[44], net578[45], net578[46],
     net578[47]}), .sp4_r_v_b_03({net580[0], net580[1], net580[2],
     net580[3], net580[4], net580[5], net580[6], net580[7], net580[8],
     net580[9], net580[10], net580[11], net580[12], net580[13],
     net580[14], net580[15], net580[16], net580[17], net580[18],
     net580[19], net580[20], net580[21], net580[22], net580[23],
     net580[24], net580[25], net580[26], net580[27], net580[28],
     net580[29], net580[30], net580[31], net580[32], net580[33],
     net580[34], net580[35], net580[36], net580[37], net580[38],
     net580[39], net580[40], net580[41], net580[42], net580[43],
     net580[44], net580[45], net580[46], net580[47]}),
     .sp4_r_v_b_02({net581[0], net581[1], net581[2], net581[3],
     net581[4], net581[5], net581[6], net581[7], net581[8], net581[9],
     net581[10], net581[11], net581[12], net581[13], net581[14],
     net581[15], net581[16], net581[17], net581[18], net581[19],
     net581[20], net581[21], net581[22], net581[23], net581[24],
     net581[25], net581[26], net581[27], net581[28], net581[29],
     net581[30], net581[31], net581[32], net581[33], net581[34],
     net581[35], net581[36], net581[37], net581[38], net581[39],
     net581[40], net581[41], net581[42], net581[43], net581[44],
     net581[45], net581[46], net581[47]}), .sp4_r_v_b_01({net577[0],
     net577[1], net577[2], net577[3], net577[4], net577[5], net577[6],
     net577[7], net577[8], net577[9], net577[10], net577[11],
     net577[12], net577[13], net577[14], net577[15], net577[16],
     net577[17], net577[18], net577[19], net577[20], net577[21],
     net577[22], net577[23], net577[24], net577[25], net577[26],
     net577[27], net577[28], net577[29], net577[30], net577[31],
     net577[32], net577[33], net577[34], net577[35], net577[36],
     net577[37], net577[38], net577[39], net577[40], net577[41],
     net577[42], net577[43], net577[44], net577[45], net577[46],
     net577[47]}), .sp4_h_r_04({net535[0], net535[1], net535[2],
     net535[3], net535[4], net535[5], net535[6], net535[7], net535[8],
     net535[9], net535[10], net535[11], net535[12], net535[13],
     net535[14], net535[15], net535[16], net535[17], net535[18],
     net535[19], net535[20], net535[21], net535[22], net535[23],
     net535[24], net535[25], net535[26], net535[27], net535[28],
     net535[29], net535[30], net535[31], net535[32], net535[33],
     net535[34], net535[35], net535[36], net535[37], net535[38],
     net535[39], net535[40], net535[41], net535[42], net535[43],
     net535[44], net535[45], net535[46], net535[47]}),
     .sp4_h_r_03({net536[0], net536[1], net536[2], net536[3],
     net536[4], net536[5], net536[6], net536[7], net536[8], net536[9],
     net536[10], net536[11], net536[12], net536[13], net536[14],
     net536[15], net536[16], net536[17], net536[18], net536[19],
     net536[20], net536[21], net536[22], net536[23], net536[24],
     net536[25], net536[26], net536[27], net536[28], net536[29],
     net536[30], net536[31], net536[32], net536[33], net536[34],
     net536[35], net536[36], net536[37], net536[38], net536[39],
     net536[40], net536[41], net536[42], net536[43], net536[44],
     net536[45], net536[46], net536[47]}), .sp4_h_r_02({net537[0],
     net537[1], net537[2], net537[3], net537[4], net537[5], net537[6],
     net537[7], net537[8], net537[9], net537[10], net537[11],
     net537[12], net537[13], net537[14], net537[15], net537[16],
     net537[17], net537[18], net537[19], net537[20], net537[21],
     net537[22], net537[23], net537[24], net537[25], net537[26],
     net537[27], net537[28], net537[29], net537[30], net537[31],
     net537[32], net537[33], net537[34], net537[35], net537[36],
     net537[37], net537[38], net537[39], net537[40], net537[41],
     net537[42], net537[43], net537[44], net537[45], net537[46],
     net537[47]}), .sp4_h_r_01({net538[0], net538[1], net538[2],
     net538[3], net538[4], net538[5], net538[6], net538[7], net538[8],
     net538[9], net538[10], net538[11], net538[12], net538[13],
     net538[14], net538[15], net538[16], net538[17], net538[18],
     net538[19], net538[20], net538[21], net538[22], net538[23],
     net538[24], net538[25], net538[26], net538[27], net538[28],
     net538[29], net538[30], net538[31], net538[32], net538[33],
     net538[34], net538[35], net538[36], net538[37], net538[38],
     net538[39], net538[40], net538[41], net538[42], net538[43],
     net538[44], net538[45], net538[46], net538[47]}),
     .sp4_h_l_03({net479[0], net479[1], net479[2], net479[3],
     net479[4], net479[5], net479[6], net479[7], net479[8], net479[9],
     net479[10], net479[11], net479[12], net479[13], net479[14],
     net479[15], net479[16], net479[17], net479[18], net479[19],
     net479[20], net479[21], net479[22], net479[23], net479[24],
     net479[25], net479[26], net479[27], net479[28], net479[29],
     net479[30], net479[31], net479[32], net479[33], net479[34],
     net479[35], net479[36], net479[37], net479[38], net479[39],
     net479[40], net479[41], net479[42], net479[43], net479[44],
     net479[45], net479[46], net479[47]}), .sp4_h_l_02({net480[0],
     net480[1], net480[2], net480[3], net480[4], net480[5], net480[6],
     net480[7], net480[8], net480[9], net480[10], net480[11],
     net480[12], net480[13], net480[14], net480[15], net480[16],
     net480[17], net480[18], net480[19], net480[20], net480[21],
     net480[22], net480[23], net480[24], net480[25], net480[26],
     net480[27], net480[28], net480[29], net480[30], net480[31],
     net480[32], net480[33], net480[34], net480[35], net480[36],
     net480[37], net480[38], net480[39], net480[40], net480[41],
     net480[42], net480[43], net480[44], net480[45], net480[46],
     net480[47]}), .sp4_h_l_01({net481[0], net481[1], net481[2],
     net481[3], net481[4], net481[5], net481[6], net481[7], net481[8],
     net481[9], net481[10], net481[11], net481[12], net481[13],
     net481[14], net481[15], net481[16], net481[17], net481[18],
     net481[19], net481[20], net481[21], net481[22], net481[23],
     net481[24], net481[25], net481[26], net481[27], net481[28],
     net481[29], net481[30], net481[31], net481[32], net481[33],
     net481[34], net481[35], net481[36], net481[37], net481[38],
     net481[39], net481[40], net481[41], net481[42], net481[43],
     net481[44], net481[45], net481[46], net481[47]}),
     .bl(bl[161:108]), .bot_op_01(bot_op_06_05[7:0]),
     .sp12_h_l_01({net472[0], net472[1], net472[2], net472[3],
     net472[4], net472[5], net472[6], net472[7], net472[8], net472[9],
     net472[10], net472[11], net472[12], net472[13], net472[14],
     net472[15], net472[16], net472[17], net472[18], net472[19],
     net472[20], net472[21], net472[22], net472[23]}),
     .sp12_h_l_02({net471[0], net471[1], net471[2], net471[3],
     net471[4], net471[5], net471[6], net471[7], net471[8], net471[9],
     net471[10], net471[11], net471[12], net471[13], net471[14],
     net471[15], net471[16], net471[17], net471[18], net471[19],
     net471[20], net471[21], net471[22], net471[23]}),
     .sp12_h_l_03({net470[0], net470[1], net470[2], net470[3],
     net470[4], net470[5], net470[6], net470[7], net470[8], net470[9],
     net470[10], net470[11], net470[12], net470[13], net470[14],
     net470[15], net470[16], net470[17], net470[18], net470[19],
     net470[20], net470[21], net470[22], net470[23]}),
     .sp12_h_l_04({net469[0], net469[1], net469[2], net469[3],
     net469[4], net469[5], net469[6], net469[7], net469[8], net469[9],
     net469[10], net469[11], net469[12], net469[13], net469[14],
     net469[15], net469[16], net469[17], net469[18], net469[19],
     net469[20], net469[21], net469[22], net469[23]}),
     .sp4_v_b_04({net474[0], net474[1], net474[2], net474[3],
     net474[4], net474[5], net474[6], net474[7], net474[8], net474[9],
     net474[10], net474[11], net474[12], net474[13], net474[14],
     net474[15], net474[16], net474[17], net474[18], net474[19],
     net474[20], net474[21], net474[22], net474[23], net474[24],
     net474[25], net474[26], net474[27], net474[28], net474[29],
     net474[30], net474[31], net474[32], net474[33], net474[34],
     net474[35], net474[36], net474[37], net474[38], net474[39],
     net474[40], net474[41], net474[42], net474[43], net474[44],
     net474[45], net474[46], net474[47]}), .sp4_v_b_03({net475[0],
     net475[1], net475[2], net475[3], net475[4], net475[5], net475[6],
     net475[7], net475[8], net475[9], net475[10], net475[11],
     net475[12], net475[13], net475[14], net475[15], net475[16],
     net475[17], net475[18], net475[19], net475[20], net475[21],
     net475[22], net475[23], net475[24], net475[25], net475[26],
     net475[27], net475[28], net475[29], net475[30], net475[31],
     net475[32], net475[33], net475[34], net475[35], net475[36],
     net475[37], net475[38], net475[39], net475[40], net475[41],
     net475[42], net475[43], net475[44], net475[45], net475[46],
     net475[47]}), .sp4_v_b_02({net476[0], net476[1], net476[2],
     net476[3], net476[4], net476[5], net476[6], net476[7], net476[8],
     net476[9], net476[10], net476[11], net476[12], net476[13],
     net476[14], net476[15], net476[16], net476[17], net476[18],
     net476[19], net476[20], net476[21], net476[22], net476[23],
     net476[24], net476[25], net476[26], net476[27], net476[28],
     net476[29], net476[30], net476[31], net476[32], net476[33],
     net476[34], net476[35], net476[36], net476[37], net476[38],
     net476[39], net476[40], net476[41], net476[42], net476[43],
     net476[44], net476[45], net476[46], net476[47]}),
     .bnr_op_01(bnr_op_06_05[7:0]), .tnr_op_04({net569, net569, net569,
     net569, net569, net569, net569, net569}),
     .glb_netwk(glb_in_6[7:0]), .tnl_op_04({slf_op_05_09[3],
     slf_op_05_09[2], slf_op_05_09[1], slf_op_05_09[0],
     slf_op_05_09[3], slf_op_05_09[2], slf_op_05_09[1],
     slf_op_05_09[0]}), .pgate(pgate_r[63:0]),
     .reset_b(reset_b_r[63:0]), .wl(wl_r[63:0]),
     .top_op_04({slf_op_06_09[3], slf_op_06_09[2], slf_op_06_09[1],
     slf_op_06_09[0], slf_op_06_09[3], slf_op_06_09[2],
     slf_op_06_09[1], slf_op_06_09[0]}), .lc_bot(lc_bot_06_05),
     .op_vic(net560), .sp12_v_b_01(sp12_v_b_06_05[23:0]),
     .sp4_v_t_04({net562[0], net562[1], net562[2], net562[3],
     net562[4], net562[5], net562[6], net562[7], net562[8], net562[9],
     net562[10], net562[11], net562[12], net562[13], net562[14],
     net562[15], net562[16], net562[17], net562[18], net562[19],
     net562[20], net562[21], net562[22], net562[23], net562[24],
     net562[25], net562[26], net562[27], net562[28], net562[29],
     net562[30], net562[31], net562[32], net562[33], net562[34],
     net562[35], net562[36], net562[37], net562[38], net562[39],
     net562[40], net562[41], net562[42], net562[43], net562[44],
     net562[45], net562[46], net562[47]}), .sp12_v_t_04({net563[0],
     net563[1], net563[2], net563[3], net563[4], net563[5], net563[6],
     net563[7], net563[8], net563[9], net563[10], net563[11],
     net563[12], net563[13], net563[14], net563[15], net563[16],
     net563[17], net563[18], net563[19], net563[20], net563[21],
     net563[22], net563[23]}));
pinlatbuf12p I_pinlatbuf12p_r ( .pad_in(padin_r_t[8]),
     .icegate(hold_r_t), .cbit(cf_r[15]), .cout(net0599), .prog(prog));
pinlatbuf12p I389 ( .pad_in(padin_t_r[6]), .icegate(hold_t_r),
     .cbit(cf_top_r[15]), .cout(net567), .prog(prog));
tielo I450 ( .tielo(net569));
fabric_buf_ice8p I390 ( .f_in(net567), .f_out(padin_04_09a));
fabric_buf_ice8p I461 ( .f_in(net0599), .f_out(padin_07_05a));

endmodule
// Library - ice384chip, Cell - io_lft_top_1x4_ice384, View - schematic
// LAST TIME SAVED: Nov 11 16:28:40 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_lft_top_1x4_ice384 ( cf_l, fabric_out_05, padeb, pado, sdo,
     slf_op_01, slf_op_02, slf_op_03, slf_op_04, tclk_o, SP4_h_l_01,
     SP4_h_l_02, SP4_h_l_03, SP4_h_l_04, SP12_h_l_01, SP12_h_l_02,
     SP12_h_l_03, SP12_h_l_04, bl, glb_netwk, pgate, reset_b,
     sp4_v_b_00_05, sp4_v_t_04, vdd_cntl, wl, bnr_op_00_05, bs_en, ceb,
     hiz_b, hold, jtag_rowtest_mode_rowu1_b, last_rsr, mode, padin,
     prog, r, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04, sdi, shift,
     tclk, tnr_op_04, update );
output  fabric_out_05, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu1_b, mode, prog,
     r, sdi, shift, tclk, update;

output [3:0]  slf_op_01;
output [3:0]  slf_op_03;
output [3:0]  slf_op_02;
output [95:0]  cf_l;
output [3:0]  slf_op_04;
output [15:8]  padeb;
output [15:8]  pado;

inout [47:0]  SP4_h_l_01;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_02;
inout [15:0]  sp4_v_t_04;
inout [47:0]  SP4_h_l_04;
inout [23:0]  SP12_h_l_01;
inout [23:0]  SP12_h_l_04;
inout [23:0]  SP12_h_l_02;
inout [7:0]  glb_netwk;
inout [23:0]  SP12_h_l_03;
inout [63:0]  wl;
inout [63:0]  vdd_cntl;
inout [63:0]  reset_b;
inout [63:0]  pgate;
inout [47:0]  SP4_h_l_03;
inout [15:0]  sp4_v_b_00_05;

input [7:0]  rgt_op_02;
input [7:0]  rgt_op_01;
input [7:0]  tnr_op_04;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_04;
input [7:0]  bnr_op_00_05;
input [15:8]  padin;
input [1:1]  last_rsr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net1009;

wire  [15:0]  net901;

wire  [7:0]  net1007;

wire  [15:0]  net937;

wire  [15:0]  net865;

wire  [1:0]  net1005;

wire  [7:0]  net1008;

wire  [1:0]  net1002;

wire  [7:0]  net884;

wire  [1:0]  net1014;

wire  [7:0]  net0429;



fabric_buf_ice8p I385 ( .f_in(net0263), .f_out(fabric_out_05));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
io_col4_lft_ice8p_v2 I_io_00_02 ( .cbit_colcntl({net1007[0],
     net1007[1], net1007[2], net1007[3], net1007[4], net1007[5],
     net1007[6], net1007[7]}), .ceb(ceb), .sdo(net887), .sdi(net851),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[11:10]), .pado(pado[11:10]), .padeb(padeb[11:10]),
     .sp4_v_t({net865[0], net865[1], net865[2], net865[3], net865[4],
     net865[5], net865[6], net865[7], net865[8], net865[9], net865[10],
     net865[11], net865[12], net865[13], net865[14], net865[15]}),
     .sp4_h_l(SP4_h_l_02[47:0]), .sp12_h_l(SP12_h_l_02[23:0]),
     .prog(prog), .spi_ss_in_b({net1014[0], net1014[1]}),
     .tnl_op(rgt_op_03[7:0]), .lft_op(rgt_op_02[7:0]),
     .bnl_op(rgt_op_01[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15]}), .wl(wl[31:16]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(net0229));
io_col4_lft_ice8p_v2 I_io_00_01 ( .cbit_colcntl({net884[0], net884[1],
     net884[2], net884[3], net884[4], net884[5], net884[6],
     net884[7]}), .ceb(ceb), .sdo(sdo), .sdi(net887), .spiout({tiegnd,
     last_rsr[1]}), .cdone_in(jtag_rowtest_mode_rowu1_b),
     .spioeb({tievdd, tiegnd}), .mode(mode), .shift(shift),
     .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[9:8]), .pado(pado[9:8]),
     .padeb(padeb[9:8]), .sp4_v_t({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15]}), .sp4_h_l(SP4_h_l_01[47:0]),
     .sp12_h_l(SP12_h_l_01[23:0]), .prog(prog),
     .spi_ss_in_b({net1005[0], net1005[1]}), .tnl_op(rgt_op_02[7:0]),
     .lft_op(rgt_op_01[7:0]), .bnl_op(bnr_op_00_05[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_v_b_00_05[15:0]), .wl(wl[15:0]), .cf(cf_l[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk[7:0]), .hold(hold), .fabric_out(net0263));
io_col4_lft_ice8p_v2 I_io_00_03 ( .cbit_colcntl({net1008[0],
     net1008[1], net1008[2], net1008[3], net1008[4], net1008[5],
     net1008[6], net1008[7]}), .ceb(ceb), .sdo(net851), .sdi(net923),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[13:12]), .pado(pado[13:12]), .padeb(padeb[13:12]),
     .sp4_v_t({net937[0], net937[1], net937[2], net937[3], net937[4],
     net937[5], net937[6], net937[7], net937[8], net937[9], net937[10],
     net937[11], net937[12], net937[13], net937[14], net937[15]}),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b({net1009[0], net1009[1]}),
     .tnl_op(rgt_op_04[7:0]), .lft_op(rgt_op_03[7:0]),
     .bnl_op(rgt_op_02[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b({net865[0], net865[1], net865[2],
     net865[3], net865[4], net865[5], net865[6], net865[7], net865[8],
     net865[9], net865[10], net865[11], net865[12], net865[13],
     net865[14], net865[15]}), .wl(wl[47:32]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(net0301));
io_col4_lft_ice8p_v2 I_io_00_04 ( .cbit_colcntl({net0429[0],
     net0429[1], net0429[2], net0429[3], net0429[4], net0429[5],
     net0429[6], net0429[7]}), .ceb(ceb), .sdo(net923), .sdi(sdi),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[15:14]), .pado(pado[15:14]), .padeb(padeb[15:14]),
     .sp4_v_t(sp4_v_t_04[15:0]), .sp4_h_l(SP4_h_l_04[47:0]),
     .sp12_h_l(SP12_h_l_04[23:0]), .prog(prog),
     .spi_ss_in_b({net1002[0], net1002[1]}), .tnl_op(tnr_op_04[7:0]),
     .lft_op(rgt_op_04[7:0]), .bnl_op(rgt_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]), .sp4_v_b({net937[0],
     net937[1], net937[2], net937[3], net937[4], net937[5], net937[6],
     net937[7], net937[8], net937[9], net937[10], net937[11],
     net937[12], net937[13], net937[14], net937[15]}), .wl(wl[63:48]),
     .cf(cf_l[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(net0337));

endmodule
// Library - ice384chip, Cell - io_top_lft_1x3_ice384, View - schematic
// LAST TIME SAVED: Nov 11 16:27:57 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module io_top_lft_1x3_ice384 ( bs_en_o, ceb_o, cf_top_l,
     fabric_out_03_09, hiz_b_o, mode_o, padeb_t_l, pado_t_l, r_o, sdo,
     shift_o, slf_op_01_09, slf_op_02_09, slf_op_03_09, tclk_o,
     update_o, bl_01, bl_02, bl_03, sp4_h_l_01_09, sp4_h_r_03_09,
     sp4_v_b_01_09, sp4_v_b_02_09, sp4_v_b_03_09, sp12_v_b_01_09,
     sp12_v_b_02_09, sp12_v_b_03_09, bnl_op_01_09, bnr_op_03_09,
     bs_en_i, ceb_i, glb_net_01, glb_net_02, glb_net_03, hiz_b_i,
     hold_t_l, lft_op_01_09, lft_op_02_09, lft_op_03_09, mode_i,
     padin_t_l, pgate_l, prog, r_i, reset_l, sdi, shift_i, tclk_i,
     update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_03_09, hiz_b_o, mode_o, r_o, sdo,
     shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_02_09;
output [3:0]  slf_op_01_09;
output [3:0]  slf_op_03_09;
output [71:0]  cf_top_l;
output [5:0]  pado_t_l;
output [5:0]  padeb_t_l;

inout [23:0]  sp12_v_b_01_09;
inout [23:0]  sp12_v_b_03_09;
inout [47:0]  sp4_v_b_03_09;
inout [23:0]  sp12_v_b_02_09;
inout [47:0]  sp4_v_b_01_09;
inout [15:0]  sp4_h_r_03_09;
inout [47:0]  sp4_v_b_02_09;
inout [15:0]  sp4_h_l_01_09;
inout [53:0]  bl_02;
inout [53:0]  bl_03;
inout [53:0]  bl_01;

input [15:0]  reset_l;
input [7:0]  glb_net_03;
input [7:0]  bnl_op_01_09;
input [7:0]  bnr_op_03_09;
input [7:0]  lft_op_01_09;
input [7:0]  lft_op_03_09;
input [15:0]  pgate_l;
input [15:0]  wl_l;
input [7:0]  lft_op_02_09;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_02;
input [5:0]  padin_t_l;
input [7:0]  glb_net_01;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  net1427;

wire  [15:0]  net1357;

wire  [1:0]  net1431;

wire  [1:0]  net1361;

wire  [1:0]  net1312;



fabric_buf_ice8p I388 ( .f_in(net0307), .f_out(fabric_out_03_09));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(net0262), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));
scan_buf_ice8p I345 ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net0262), .shift_o(shift_o),
     .sdo(net1517), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_top_ice8p I_IO_02_09 ( .sdo(net1412), .sdi(net1342),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1427[0], net1427[1], net1427[2],
     net1427[3], net1427[4], net1427[5], net1427[6], net1427[7],
     net1427[8], net1427[9], net1427[10], net1427[11], net1427[12],
     net1427[13], net1427[14], net1427[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[3:2]),
     .pado(pado_t_l[3:2]), .padeb(padeb_t_l[3:2]),
     .sp4_v_b({net1357[0], net1357[1], net1357[2], net1357[3],
     net1357[4], net1357[5], net1357[6], net1357[7], net1357[8],
     net1357[9], net1357[10], net1357[11], net1357[12], net1357[13],
     net1357[14], net1357[15]}), .sp4_h_l(sp4_v_b_02_09[47:0]),
     .sp12_h_l(sp12_v_b_02_09[23:0]), .prog(prog),
     .spi_ss_in_b({net1361[0], net1361[1]}),
     .tnl_op(lft_op_01_09[7:0]), .lft_op(lft_op_02_09[7:0]),
     .bnl_op(lft_op_03_09[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[47:24]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_09[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_t_l), .fabric_out(net1320));
io_col4_top_ice8p I_IO_01_09 ( .sdo(sdo), .sdi(net1412),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_01_09[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[1:0]),
     .pado(pado_t_l[1:0]), .padeb(padeb_t_l[1:0]),
     .sp4_v_b({net1427[0], net1427[1], net1427[2], net1427[3],
     net1427[4], net1427[5], net1427[6], net1427[7], net1427[8],
     net1427[9], net1427[10], net1427[11], net1427[12], net1427[13],
     net1427[14], net1427[15]}), .sp4_h_l(sp4_v_b_01_09[47:0]),
     .sp12_h_l(sp12_v_b_01_09[23:0]), .prog(prog),
     .spi_ss_in_b({net1431[0], net1431[1]}),
     .tnl_op(bnl_op_01_09[7:0]), .lft_op(lft_op_01_09[7:0]),
     .bnl_op(lft_op_02_09[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[23:0]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_09[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_t_l), .fabric_out(net1445));
io_col4_top_ice8p I_IO_03_09 ( .sdo(net1342), .sdi(net1517),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1357[0], net1357[1], net1357[2],
     net1357[3], net1357[4], net1357[5], net1357[6], net1357[7],
     net1357[8], net1357[9], net1357[10], net1357[11], net1357[12],
     net1357[13], net1357[14], net1357[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[5:4]),
     .pado(pado_t_l[5:4]), .padeb(padeb_t_l[5:4]),
     .sp4_v_b(sp4_h_r_03_09[15:0]), .sp4_h_l(sp4_v_b_03_09[47:0]),
     .sp12_h_l(sp12_v_b_03_09[23:0]), .prog(prog),
     .spi_ss_in_b({net1312[0], net1312[1]}),
     .tnl_op(lft_op_02_09[7:0]), .lft_op(lft_op_03_09[7:0]),
     .bnl_op(bnr_op_03_09[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[71:48]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_09[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_t_l), .fabric_out(net0307));

endmodule
// Library - ice384chip, Cell - quad_tl_ice384, View - schematic
// LAST TIME SAVED: Nov 23 12:21:17 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module quad_tl_ice384 ( bs_en_o, ceb_o, cf_l, cf_top_l,
     fabric_out_00_05, fabric_out_03_09, hiz_b_o, mode_o, padeb_l_t,
     padeb_t_l, padin_00_05a, padin_03_09b, pado_l_t, pado_t_l, r_o,
     sdo, shift_o, slf_op_00_05, slf_op_01_05, slf_op_02_05,
     slf_op_03_05, slf_op_03_06, slf_op_03_07, slf_op_03_08,
     slf_op_03_09, tclk_o, update_o, bl, pgate_l, reset_b_l,
     sp4_h_r_03_05, sp4_h_r_03_06, sp4_h_r_03_07, sp4_h_r_03_08,
     sp4_h_r_03_09, sp4_r_v_b_03_05, sp4_r_v_b_03_06, sp4_r_v_b_03_07,
     sp4_r_v_b_03_08, sp4_v_b_00_05, sp4_v_b_01_05, sp4_v_b_02_05,
     sp4_v_b_03_05, sp12_h_r_03_05, sp12_h_r_03_06, sp12_h_r_03_07,
     sp12_h_r_03_08, sp12_v_b_01_05, sp12_v_b_02_05, sp12_v_b_03_05,
     vdd_cntl_l, wl_l, bnl_op_01_05, bnl_op_02_05, bnl_op_03_05,
     bnr_op_00_05, bnr_op_01_05, bnr_op_02_05, bnr_op_03_05,
     bot_op_01_05, bot_op_02_05, bot_op_03_05, bs_en_i, carry_in_01_05,
     carry_in_02_05, carry_in_03_05, ceb_i, glb_in_0, glb_in_1,
     glb_in_2, glb_in_3, hiz_b_i, hold_l_t, hold_t_l,
     jtag_rowtest_mode_rowu1_b, last_rsr, lc_bot_01_05, lc_bot_02_05,
     lc_bot_03_05, mode_i, padin_l_t, padin_t_l, prog, purst, r_i,
     rgt_op_03_05, rgt_op_03_06, rgt_op_03_07, rgt_op_03_08, sdi,
     shift_i, tclk_i, tnr_op_03_08, update_i );
output  bs_en_o, ceb_o, fabric_out_00_05, fabric_out_03_09, hiz_b_o,
     mode_o, padin_00_05a, padin_03_09b, r_o, sdo, shift_o, tclk_o,
     update_o;


input  bs_en_i, carry_in_01_05, carry_in_02_05, carry_in_03_05, ceb_i,
     hiz_b_i, hold_l_t, hold_t_l, jtag_rowtest_mode_rowu1_b,
     lc_bot_01_05, lc_bot_02_05, lc_bot_03_05, mode_i, prog, purst,
     r_i, sdi, shift_i, tclk_i, update_i;

output [7:0]  slf_op_03_06;
output [15:8]  pado_l_t;
output [7:0]  slf_op_03_05;
output [7:0]  slf_op_03_08;
output [5:0]  padeb_t_l;
output [7:0]  slf_op_02_05;
output [7:0]  slf_op_01_05;
output [95:0]  cf_l;
output [5:0]  pado_t_l;
output [3:0]  slf_op_00_05;
output [3:0]  slf_op_03_09;
output [71:0]  cf_top_l;
output [15:8]  padeb_l_t;
output [7:0]  slf_op_03_07;

inout [47:0]  sp4_r_v_b_03_08;
inout [47:0]  sp4_h_r_03_08;
inout [47:0]  sp4_v_b_01_05;
inout [15:0]  sp4_v_b_00_05;
inout [23:0]  sp12_h_r_03_07;
inout [47:0]  sp4_r_v_b_03_07;
inout [23:0]  sp12_v_b_01_05;
inout [47:0]  sp4_h_r_03_05;
inout [23:0]  sp12_h_r_03_08;
inout [15:0]  sp4_h_r_03_09;
inout [23:0]  sp12_v_b_03_05;
inout [23:0]  sp12_h_r_03_06;
inout [47:0]  sp4_v_b_03_05;
inout [47:0]  sp4_v_b_02_05;
inout [23:0]  sp12_h_r_03_05;
inout [23:0]  sp12_v_b_02_05;
inout [79:0]  pgate_l;
inout [79:0]  reset_b_l;
inout [79:0]  vdd_cntl_l;
inout [47:0]  sp4_h_r_03_07;
inout [179:0]  bl;
inout [47:0]  sp4_h_r_03_06;
inout [79:0]  wl_l;
inout [47:0]  sp4_r_v_b_03_05;
inout [47:0]  sp4_r_v_b_03_06;

input [7:0]  bnr_op_01_05;
input [7:0]  rgt_op_03_05;
input [7:0]  bnr_op_02_05;
input [7:0]  bnl_op_03_05;
input [7:0]  bnr_op_00_05;
input [7:0]  glb_in_2;
input [7:0]  glb_in_0;
input [1:1]  last_rsr;
input [7:0]  bnl_op_01_05;
input [7:0]  bnl_op_02_05;
input [7:0]  rgt_op_03_07;
input [7:0]  rgt_op_03_08;
input [7:0]  bot_op_02_05;
input [15:8]  padin_l_t;
input [5:0]  padin_t_l;
input [7:0]  glb_in_3;
input [7:0]  glb_in_1;
input [3:0]  tnr_op_03_08;
input [7:0]  rgt_op_03_06;
input [7:0]  bot_op_03_05;
input [7:0]  bot_op_01_05;
input [7:0]  bnr_op_03_05;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [47:0]  net496;

wire  [23:0]  net352;

wire  [23:0]  net580;

wire  [23:0]  net351;

wire  [3:0]  slf_op_02_09;

wire  [3:0]  slf_op_01_09;

wire  [3:0]  slf_op_00_07;

wire  [3:0]  slf_op_00_06;

wire  [3:0]  slf_op_00_08;

wire  [47:0]  net498;

wire  [7:0]  net410;

wire  [47:0]  net435;

wire  [47:0]  net434;

wire  [23:0]  net523;

wire  [47:0]  net441;

wire  [23:0]  net432;

wire  [7:0]  net357;

wire  [47:0]  net493;

wire  [23:0]  net487;

wire  [47:0]  net334;

wire  [23:0]  net466;

wire  [47:0]  net492;

wire  [47:0]  net491;

wire  [7:0]  net337;

wire  [23:0]  net430;

wire  [7:0]  net330;

wire  [47:0]  net335;

wire  [47:0]  net336;

wire  [47:0]  net452;

wire  [47:0]  net453;

wire  [7:0]  net420;

wire  [23:0]  net488;

wire  [15:0]  net358;

wire  [23:0]  net354;

wire  [7:0]  net412;

wire  [23:0]  net353;

wire  [47:0]  net522;

wire  [23:0]  net489;

wire  [47:0]  net465;

wire  [47:0]  net451;

wire  [47:0]  net495;

wire  [47:0]  net497;

wire  [47:0]  net579;

wire  [47:0]  net333;

wire  [47:0]  net439;

wire  [23:0]  net486;

wire  [47:0]  net436;

wire  [23:0]  net429;

wire  [23:0]  net431;

wire  [47:0]  net438;

wire  [47:0]  net440;



io_lft_top_1x4_ice384 I396 ( .shift(shift_o), .bs_en(bs_en_o),
     .mode(mode_o), .sdi(net316), .hiz_b(hiz_b_o), .prog(prog),
     .hold(hold_l_t), .update(update_o), .r(r_o),
     .glb_netwk(glb_in_0[7:0]), .slf_op_01(slf_op_00_05[3:0]),
     .slf_op_02(slf_op_00_06[3:0]), .sdo(sdo), .bl({bl[0], bl[1],
     bl[2], bl[3], bl[4], bl[5], bl[6], bl[7], bl[8], bl[9], bl[10],
     bl[11], bl[12], bl[13], bl[14], bl[15], bl[16], bl[17]}),
     .sp4_v_b_00_05(sp4_v_b_00_05[15:0]), .tclk(net328),
     .reset_b(reset_b_l[63:0]), .rgt_op_02({net330[0], net330[1],
     net330[2], net330[3], net330[4], net330[5], net330[6],
     net330[7]}), .slf_op_04(slf_op_00_08[3:0]),
     .slf_op_03(slf_op_00_07[3:0]), .SP4_h_l_03({net333[0], net333[1],
     net333[2], net333[3], net333[4], net333[5], net333[6], net333[7],
     net333[8], net333[9], net333[10], net333[11], net333[12],
     net333[13], net333[14], net333[15], net333[16], net333[17],
     net333[18], net333[19], net333[20], net333[21], net333[22],
     net333[23], net333[24], net333[25], net333[26], net333[27],
     net333[28], net333[29], net333[30], net333[31], net333[32],
     net333[33], net333[34], net333[35], net333[36], net333[37],
     net333[38], net333[39], net333[40], net333[41], net333[42],
     net333[43], net333[44], net333[45], net333[46], net333[47]}),
     .SP4_h_l_04({net334[0], net334[1], net334[2], net334[3],
     net334[4], net334[5], net334[6], net334[7], net334[8], net334[9],
     net334[10], net334[11], net334[12], net334[13], net334[14],
     net334[15], net334[16], net334[17], net334[18], net334[19],
     net334[20], net334[21], net334[22], net334[23], net334[24],
     net334[25], net334[26], net334[27], net334[28], net334[29],
     net334[30], net334[31], net334[32], net334[33], net334[34],
     net334[35], net334[36], net334[37], net334[38], net334[39],
     net334[40], net334[41], net334[42], net334[43], net334[44],
     net334[45], net334[46], net334[47]}), .SP4_h_l_02({net335[0],
     net335[1], net335[2], net335[3], net335[4], net335[5], net335[6],
     net335[7], net335[8], net335[9], net335[10], net335[11],
     net335[12], net335[13], net335[14], net335[15], net335[16],
     net335[17], net335[18], net335[19], net335[20], net335[21],
     net335[22], net335[23], net335[24], net335[25], net335[26],
     net335[27], net335[28], net335[29], net335[30], net335[31],
     net335[32], net335[33], net335[34], net335[35], net335[36],
     net335[37], net335[38], net335[39], net335[40], net335[41],
     net335[42], net335[43], net335[44], net335[45], net335[46],
     net335[47]}), .SP4_h_l_01({net336[0], net336[1], net336[2],
     net336[3], net336[4], net336[5], net336[6], net336[7], net336[8],
     net336[9], net336[10], net336[11], net336[12], net336[13],
     net336[14], net336[15], net336[16], net336[17], net336[18],
     net336[19], net336[20], net336[21], net336[22], net336[23],
     net336[24], net336[25], net336[26], net336[27], net336[28],
     net336[29], net336[30], net336[31], net336[32], net336[33],
     net336[34], net336[35], net336[36], net336[37], net336[38],
     net336[39], net336[40], net336[41], net336[42], net336[43],
     net336[44], net336[45], net336[46], net336[47]}),
     .rgt_op_03({net337[0], net337[1], net337[2], net337[3], net337[4],
     net337[5], net337[6], net337[7]}), .rgt_op_01(slf_op_01_05[7:0]),
     .vdd_cntl(vdd_cntl_l[63:0]), .last_rsr(last_rsr[1]),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .tnr_op_04({slf_op_01_09[3], slf_op_01_09[2], slf_op_01_09[1],
     slf_op_01_09[0], slf_op_01_09[3], slf_op_01_09[2],
     slf_op_01_09[1], slf_op_01_09[0]}), .padin(padin_l_t[15:8]),
     .bnr_op_00_05(bnr_op_00_05[7:0]), .pado(pado_l_t[15:8]),
     .padeb(padeb_l_t[15:8]), .wl(wl_l[63:0]), .cf_l(cf_l[95:0]),
     .tclk_o(tclk_o), .ceb(ceb_o), .SP12_h_l_02({net351[0], net351[1],
     net351[2], net351[3], net351[4], net351[5], net351[6], net351[7],
     net351[8], net351[9], net351[10], net351[11], net351[12],
     net351[13], net351[14], net351[15], net351[16], net351[17],
     net351[18], net351[19], net351[20], net351[21], net351[22],
     net351[23]}), .SP12_h_l_04({net352[0], net352[1], net352[2],
     net352[3], net352[4], net352[5], net352[6], net352[7], net352[8],
     net352[9], net352[10], net352[11], net352[12], net352[13],
     net352[14], net352[15], net352[16], net352[17], net352[18],
     net352[19], net352[20], net352[21], net352[22], net352[23]}),
     .SP12_h_l_01({net353[0], net353[1], net353[2], net353[3],
     net353[4], net353[5], net353[6], net353[7], net353[8], net353[9],
     net353[10], net353[11], net353[12], net353[13], net353[14],
     net353[15], net353[16], net353[17], net353[18], net353[19],
     net353[20], net353[21], net353[22], net353[23]}),
     .SP12_h_l_03({net354[0], net354[1], net354[2], net354[3],
     net354[4], net354[5], net354[6], net354[7], net354[8], net354[9],
     net354[10], net354[11], net354[12], net354[13], net354[14],
     net354[15], net354[16], net354[17], net354[18], net354[19],
     net354[20], net354[21], net354[22], net354[23]}),
     .pgate(pgate_l[63:0]), .fabric_out_05(fabric_out_00_05),
     .rgt_op_04({net357[0], net357[1], net357[2], net357[3], net357[4],
     net357[5], net357[6], net357[7]}), .sp4_v_t_04({net358[0],
     net358[1], net358[2], net358[3], net358[4], net358[5], net358[6],
     net358[7], net358[8], net358[9], net358[10], net358[11],
     net358[12], net358[13], net358[14], net358[15]}));
io_top_lft_1x3_ice384 I398 ( .wl_l({wl_l[78], wl_l[79], wl_l[77],
     wl_l[76], wl_l[74], wl_l[75], wl_l[73], wl_l[72], wl_l[70],
     wl_l[71], wl_l[69], wl_l[68], wl_l[66], wl_l[67], wl_l[65],
     wl_l[64]}), .sp12_v_b_01_09({net466[0], net466[1], net466[2],
     net466[3], net466[4], net466[5], net466[6], net466[7], net466[8],
     net466[9], net466[10], net466[11], net466[12], net466[13],
     net466[14], net466[15], net466[16], net466[17], net466[18],
     net466[19], net466[20], net466[21], net466[22], net466[23]}),
     .vdd_cntl_l({vdd_cntl_l[78], vdd_cntl_l[79], vdd_cntl_l[77],
     vdd_cntl_l[76], vdd_cntl_l[74], vdd_cntl_l[75], vdd_cntl_l[73],
     vdd_cntl_l[72], vdd_cntl_l[70], vdd_cntl_l[71], vdd_cntl_l[69],
     vdd_cntl_l[68], vdd_cntl_l[66], vdd_cntl_l[67], vdd_cntl_l[65],
     vdd_cntl_l[64]}), .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .reset_l({reset_b_l[78],
     reset_b_l[79], reset_b_l[77], reset_b_l[76], reset_b_l[74],
     reset_b_l[75], reset_b_l[73], reset_b_l[72], reset_b_l[70],
     reset_b_l[71], reset_b_l[69], reset_b_l[68], reset_b_l[66],
     reset_b_l[67], reset_b_l[65], reset_b_l[64]}), .r_i(r_i),
     .prog(prog), .pgate_l({pgate_l[78], pgate_l[79], pgate_l[77],
     pgate_l[76], pgate_l[74], pgate_l[75], pgate_l[73], pgate_l[72],
     pgate_l[70], pgate_l[71], pgate_l[69], pgate_l[68], pgate_l[66],
     pgate_l[67], pgate_l[65], pgate_l[64]}), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .bs_en_i(bs_en_i), .update_o(net592),
     .tclk_o(net593), .shift_o(net594), .sdo(net595), .r_o(net596),
     .mode_o(net597), .hiz_b_o(net598), .glb_net_02(glb_in_2[7:0]),
     .glb_net_01(glb_in_1[7:0]), .bs_en_o(net600), .bl_03(bl[179:126]),
     .sp4_v_b_03_09({net579[0], net579[1], net579[2], net579[3],
     net579[4], net579[5], net579[6], net579[7], net579[8], net579[9],
     net579[10], net579[11], net579[12], net579[13], net579[14],
     net579[15], net579[16], net579[17], net579[18], net579[19],
     net579[20], net579[21], net579[22], net579[23], net579[24],
     net579[25], net579[26], net579[27], net579[28], net579[29],
     net579[30], net579[31], net579[32], net579[33], net579[34],
     net579[35], net579[36], net579[37], net579[38], net579[39],
     net579[40], net579[41], net579[42], net579[43], net579[44],
     net579[45], net579[46], net579[47]}),
     .bnr_op_03_09(rgt_op_03_08[7:0]), .bl_02(bl[125:72]),
     .bl_01(bl[71:18]), .fabric_out_03_09(fabric_out_03_09),
     .cf_top_l(cf_top_l[71:0]), .bnl_op_01_09({slf_op_00_08[3],
     slf_op_00_08[2], slf_op_00_08[1], slf_op_00_08[0],
     slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0]}), .sp4_v_b_01_09({net465[0], net465[1],
     net465[2], net465[3], net465[4], net465[5], net465[6], net465[7],
     net465[8], net465[9], net465[10], net465[11], net465[12],
     net465[13], net465[14], net465[15], net465[16], net465[17],
     net465[18], net465[19], net465[20], net465[21], net465[22],
     net465[23], net465[24], net465[25], net465[26], net465[27],
     net465[28], net465[29], net465[30], net465[31], net465[32],
     net465[33], net465[34], net465[35], net465[36], net465[37],
     net465[38], net465[39], net465[40], net465[41], net465[42],
     net465[43], net465[44], net465[45], net465[46], net465[47]}),
     .padin_t_l(padin_t_l[5:0]), .slf_op_02_09(slf_op_02_09[3:0]),
     .slf_op_03_09(slf_op_03_09[3:0]),
     .lft_op_03_09(slf_op_03_08[7:0]), .sp12_v_b_02_09({net523[0],
     net523[1], net523[2], net523[3], net523[4], net523[5], net523[6],
     net523[7], net523[8], net523[9], net523[10], net523[11],
     net523[12], net523[13], net523[14], net523[15], net523[16],
     net523[17], net523[18], net523[19], net523[20], net523[21],
     net523[22], net523[23]}), .glb_net_03(glb_in_3[7:0]),
     .lft_op_01_09({net357[0], net357[1], net357[2], net357[3],
     net357[4], net357[5], net357[6], net357[7]}),
     .slf_op_01_09(slf_op_01_09[3:0]),
     .sp4_h_r_03_09(sp4_h_r_03_09[15:0]), .sp4_v_b_02_09({net522[0],
     net522[1], net522[2], net522[3], net522[4], net522[5], net522[6],
     net522[7], net522[8], net522[9], net522[10], net522[11],
     net522[12], net522[13], net522[14], net522[15], net522[16],
     net522[17], net522[18], net522[19], net522[20], net522[21],
     net522[22], net522[23], net522[24], net522[25], net522[26],
     net522[27], net522[28], net522[29], net522[30], net522[31],
     net522[32], net522[33], net522[34], net522[35], net522[36],
     net522[37], net522[38], net522[39], net522[40], net522[41],
     net522[42], net522[43], net522[44], net522[45], net522[46],
     net522[47]}), .lft_op_02_09({net420[0], net420[1], net420[2],
     net420[3], net420[4], net420[5], net420[6], net420[7]}),
     .padeb_t_l(padeb_t_l[5:0]), .ceb_o(net599),
     .pado_t_l(pado_t_l[5:0]), .sp12_v_b_03_09({net580[0], net580[1],
     net580[2], net580[3], net580[4], net580[5], net580[6], net580[7],
     net580[8], net580[9], net580[10], net580[11], net580[12],
     net580[13], net580[14], net580[15], net580[16], net580[17],
     net580[18], net580[19], net580[20], net580[21], net580[22],
     net580[23]}), .hold_t_l(hold_t_l), .sp4_h_l_01_09({net358[0],
     net358[1], net358[2], net358[3], net358[4], net358[5], net358[6],
     net358[7], net358[8], net358[9], net358[10], net358[11],
     net358[12], net358[13], net358[14], net358[15]}), .ceb_i(ceb_i));
lt_1x4_top_ice384 I394 ( .rgt_op_03({net410[0], net410[1], net410[2],
     net410[3], net410[4], net410[5], net410[6], net410[7]}),
     .slf_op_02({net330[0], net330[1], net330[2], net330[3], net330[4],
     net330[5], net330[6], net330[7]}), .rgt_op_02({net412[0],
     net412[1], net412[2], net412[3], net412[4], net412[5], net412[6],
     net412[7]}), .rgt_op_01(slf_op_02_05[7:0]), .purst(purst),
     .prog(prog), .lft_op_04({slf_op_00_08[3], slf_op_00_08[2],
     slf_op_00_08[1], slf_op_00_08[0], slf_op_00_08[3],
     slf_op_00_08[2], slf_op_00_08[1], slf_op_00_08[0]}),
     .lft_op_03({slf_op_00_07[3], slf_op_00_07[2], slf_op_00_07[1],
     slf_op_00_07[0], slf_op_00_07[3], slf_op_00_07[2],
     slf_op_00_07[1], slf_op_00_07[0]}), .lft_op_02({slf_op_00_06[3],
     slf_op_00_06[2], slf_op_00_06[1], slf_op_00_06[0],
     slf_op_00_06[3], slf_op_00_06[2], slf_op_00_06[1],
     slf_op_00_06[0]}), .lft_op_01({slf_op_00_05[3], slf_op_00_05[2],
     slf_op_00_05[1], slf_op_00_05[0], slf_op_00_05[3],
     slf_op_00_05[2], slf_op_00_05[1], slf_op_00_05[0]}),
     .rgt_op_04({net420[0], net420[1], net420[2], net420[3], net420[4],
     net420[5], net420[6], net420[7]}), .carry_in(carry_in_01_05),
     .bnl_op_01(bnl_op_01_05[7:0]), .slf_op_04({net357[0], net357[1],
     net357[2], net357[3], net357[4], net357[5], net357[6],
     net357[7]}), .slf_op_03({net337[0], net337[1], net337[2],
     net337[3], net337[4], net337[5], net337[6], net337[7]}),
     .slf_op_01(slf_op_01_05[7:0]), .sp4_h_l_04({net334[0], net334[1],
     net334[2], net334[3], net334[4], net334[5], net334[6], net334[7],
     net334[8], net334[9], net334[10], net334[11], net334[12],
     net334[13], net334[14], net334[15], net334[16], net334[17],
     net334[18], net334[19], net334[20], net334[21], net334[22],
     net334[23], net334[24], net334[25], net334[26], net334[27],
     net334[28], net334[29], net334[30], net334[31], net334[32],
     net334[33], net334[34], net334[35], net334[36], net334[37],
     net334[38], net334[39], net334[40], net334[41], net334[42],
     net334[43], net334[44], net334[45], net334[46], net334[47]}),
     .carry_out(net427), .vdd_cntl(vdd_cntl_l[63:0]),
     .sp12_h_r_04({net429[0], net429[1], net429[2], net429[3],
     net429[4], net429[5], net429[6], net429[7], net429[8], net429[9],
     net429[10], net429[11], net429[12], net429[13], net429[14],
     net429[15], net429[16], net429[17], net429[18], net429[19],
     net429[20], net429[21], net429[22], net429[23]}),
     .sp12_h_r_03({net430[0], net430[1], net430[2], net430[3],
     net430[4], net430[5], net430[6], net430[7], net430[8], net430[9],
     net430[10], net430[11], net430[12], net430[13], net430[14],
     net430[15], net430[16], net430[17], net430[18], net430[19],
     net430[20], net430[21], net430[22], net430[23]}),
     .sp12_h_r_02({net431[0], net431[1], net431[2], net431[3],
     net431[4], net431[5], net431[6], net431[7], net431[8], net431[9],
     net431[10], net431[11], net431[12], net431[13], net431[14],
     net431[15], net431[16], net431[17], net431[18], net431[19],
     net431[20], net431[21], net431[22], net431[23]}),
     .sp12_h_r_01({net432[0], net432[1], net432[2], net432[3],
     net432[4], net432[5], net432[6], net432[7], net432[8], net432[9],
     net432[10], net432[11], net432[12], net432[13], net432[14],
     net432[15], net432[16], net432[17], net432[18], net432[19],
     net432[20], net432[21], net432[22], net432[23]}),
     .sp4_v_b_01(sp4_v_b_01_05[47:0]), .sp4_r_v_b_04({net434[0],
     net434[1], net434[2], net434[3], net434[4], net434[5], net434[6],
     net434[7], net434[8], net434[9], net434[10], net434[11],
     net434[12], net434[13], net434[14], net434[15], net434[16],
     net434[17], net434[18], net434[19], net434[20], net434[21],
     net434[22], net434[23], net434[24], net434[25], net434[26],
     net434[27], net434[28], net434[29], net434[30], net434[31],
     net434[32], net434[33], net434[34], net434[35], net434[36],
     net434[37], net434[38], net434[39], net434[40], net434[41],
     net434[42], net434[43], net434[44], net434[45], net434[46],
     net434[47]}), .sp4_r_v_b_03({net435[0], net435[1], net435[2],
     net435[3], net435[4], net435[5], net435[6], net435[7], net435[8],
     net435[9], net435[10], net435[11], net435[12], net435[13],
     net435[14], net435[15], net435[16], net435[17], net435[18],
     net435[19], net435[20], net435[21], net435[22], net435[23],
     net435[24], net435[25], net435[26], net435[27], net435[28],
     net435[29], net435[30], net435[31], net435[32], net435[33],
     net435[34], net435[35], net435[36], net435[37], net435[38],
     net435[39], net435[40], net435[41], net435[42], net435[43],
     net435[44], net435[45], net435[46], net435[47]}),
     .sp4_r_v_b_02({net436[0], net436[1], net436[2], net436[3],
     net436[4], net436[5], net436[6], net436[7], net436[8], net436[9],
     net436[10], net436[11], net436[12], net436[13], net436[14],
     net436[15], net436[16], net436[17], net436[18], net436[19],
     net436[20], net436[21], net436[22], net436[23], net436[24],
     net436[25], net436[26], net436[27], net436[28], net436[29],
     net436[30], net436[31], net436[32], net436[33], net436[34],
     net436[35], net436[36], net436[37], net436[38], net436[39],
     net436[40], net436[41], net436[42], net436[43], net436[44],
     net436[45], net436[46], net436[47]}),
     .sp4_r_v_b_01(sp4_v_b_02_05[47:0]), .sp4_h_r_04({net438[0],
     net438[1], net438[2], net438[3], net438[4], net438[5], net438[6],
     net438[7], net438[8], net438[9], net438[10], net438[11],
     net438[12], net438[13], net438[14], net438[15], net438[16],
     net438[17], net438[18], net438[19], net438[20], net438[21],
     net438[22], net438[23], net438[24], net438[25], net438[26],
     net438[27], net438[28], net438[29], net438[30], net438[31],
     net438[32], net438[33], net438[34], net438[35], net438[36],
     net438[37], net438[38], net438[39], net438[40], net438[41],
     net438[42], net438[43], net438[44], net438[45], net438[46],
     net438[47]}), .sp4_h_r_03({net439[0], net439[1], net439[2],
     net439[3], net439[4], net439[5], net439[6], net439[7], net439[8],
     net439[9], net439[10], net439[11], net439[12], net439[13],
     net439[14], net439[15], net439[16], net439[17], net439[18],
     net439[19], net439[20], net439[21], net439[22], net439[23],
     net439[24], net439[25], net439[26], net439[27], net439[28],
     net439[29], net439[30], net439[31], net439[32], net439[33],
     net439[34], net439[35], net439[36], net439[37], net439[38],
     net439[39], net439[40], net439[41], net439[42], net439[43],
     net439[44], net439[45], net439[46], net439[47]}),
     .sp4_h_r_02({net440[0], net440[1], net440[2], net440[3],
     net440[4], net440[5], net440[6], net440[7], net440[8], net440[9],
     net440[10], net440[11], net440[12], net440[13], net440[14],
     net440[15], net440[16], net440[17], net440[18], net440[19],
     net440[20], net440[21], net440[22], net440[23], net440[24],
     net440[25], net440[26], net440[27], net440[28], net440[29],
     net440[30], net440[31], net440[32], net440[33], net440[34],
     net440[35], net440[36], net440[37], net440[38], net440[39],
     net440[40], net440[41], net440[42], net440[43], net440[44],
     net440[45], net440[46], net440[47]}), .sp4_h_r_01({net441[0],
     net441[1], net441[2], net441[3], net441[4], net441[5], net441[6],
     net441[7], net441[8], net441[9], net441[10], net441[11],
     net441[12], net441[13], net441[14], net441[15], net441[16],
     net441[17], net441[18], net441[19], net441[20], net441[21],
     net441[22], net441[23], net441[24], net441[25], net441[26],
     net441[27], net441[28], net441[29], net441[30], net441[31],
     net441[32], net441[33], net441[34], net441[35], net441[36],
     net441[37], net441[38], net441[39], net441[40], net441[41],
     net441[42], net441[43], net441[44], net441[45], net441[46],
     net441[47]}), .sp4_h_l_03({net333[0], net333[1], net333[2],
     net333[3], net333[4], net333[5], net333[6], net333[7], net333[8],
     net333[9], net333[10], net333[11], net333[12], net333[13],
     net333[14], net333[15], net333[16], net333[17], net333[18],
     net333[19], net333[20], net333[21], net333[22], net333[23],
     net333[24], net333[25], net333[26], net333[27], net333[28],
     net333[29], net333[30], net333[31], net333[32], net333[33],
     net333[34], net333[35], net333[36], net333[37], net333[38],
     net333[39], net333[40], net333[41], net333[42], net333[43],
     net333[44], net333[45], net333[46], net333[47]}),
     .sp4_h_l_02({net335[0], net335[1], net335[2], net335[3],
     net335[4], net335[5], net335[6], net335[7], net335[8], net335[9],
     net335[10], net335[11], net335[12], net335[13], net335[14],
     net335[15], net335[16], net335[17], net335[18], net335[19],
     net335[20], net335[21], net335[22], net335[23], net335[24],
     net335[25], net335[26], net335[27], net335[28], net335[29],
     net335[30], net335[31], net335[32], net335[33], net335[34],
     net335[35], net335[36], net335[37], net335[38], net335[39],
     net335[40], net335[41], net335[42], net335[43], net335[44],
     net335[45], net335[46], net335[47]}), .sp4_h_l_01({net336[0],
     net336[1], net336[2], net336[3], net336[4], net336[5], net336[6],
     net336[7], net336[8], net336[9], net336[10], net336[11],
     net336[12], net336[13], net336[14], net336[15], net336[16],
     net336[17], net336[18], net336[19], net336[20], net336[21],
     net336[22], net336[23], net336[24], net336[25], net336[26],
     net336[27], net336[28], net336[29], net336[30], net336[31],
     net336[32], net336[33], net336[34], net336[35], net336[36],
     net336[37], net336[38], net336[39], net336[40], net336[41],
     net336[42], net336[43], net336[44], net336[45], net336[46],
     net336[47]}), .bl(bl[71:18]), .bot_op_01(bot_op_01_05[7:0]),
     .sp12_h_l_01({net353[0], net353[1], net353[2], net353[3],
     net353[4], net353[5], net353[6], net353[7], net353[8], net353[9],
     net353[10], net353[11], net353[12], net353[13], net353[14],
     net353[15], net353[16], net353[17], net353[18], net353[19],
     net353[20], net353[21], net353[22], net353[23]}),
     .sp12_h_l_02({net351[0], net351[1], net351[2], net351[3],
     net351[4], net351[5], net351[6], net351[7], net351[8], net351[9],
     net351[10], net351[11], net351[12], net351[13], net351[14],
     net351[15], net351[16], net351[17], net351[18], net351[19],
     net351[20], net351[21], net351[22], net351[23]}),
     .sp12_h_l_03({net354[0], net354[1], net354[2], net354[3],
     net354[4], net354[5], net354[6], net354[7], net354[8], net354[9],
     net354[10], net354[11], net354[12], net354[13], net354[14],
     net354[15], net354[16], net354[17], net354[18], net354[19],
     net354[20], net354[21], net354[22], net354[23]}),
     .sp12_h_l_04({net352[0], net352[1], net352[2], net352[3],
     net352[4], net352[5], net352[6], net352[7], net352[8], net352[9],
     net352[10], net352[11], net352[12], net352[13], net352[14],
     net352[15], net352[16], net352[17], net352[18], net352[19],
     net352[20], net352[21], net352[22], net352[23]}),
     .sp4_v_b_04({net451[0], net451[1], net451[2], net451[3],
     net451[4], net451[5], net451[6], net451[7], net451[8], net451[9],
     net451[10], net451[11], net451[12], net451[13], net451[14],
     net451[15], net451[16], net451[17], net451[18], net451[19],
     net451[20], net451[21], net451[22], net451[23], net451[24],
     net451[25], net451[26], net451[27], net451[28], net451[29],
     net451[30], net451[31], net451[32], net451[33], net451[34],
     net451[35], net451[36], net451[37], net451[38], net451[39],
     net451[40], net451[41], net451[42], net451[43], net451[44],
     net451[45], net451[46], net451[47]}), .sp4_v_b_03({net452[0],
     net452[1], net452[2], net452[3], net452[4], net452[5], net452[6],
     net452[7], net452[8], net452[9], net452[10], net452[11],
     net452[12], net452[13], net452[14], net452[15], net452[16],
     net452[17], net452[18], net452[19], net452[20], net452[21],
     net452[22], net452[23], net452[24], net452[25], net452[26],
     net452[27], net452[28], net452[29], net452[30], net452[31],
     net452[32], net452[33], net452[34], net452[35], net452[36],
     net452[37], net452[38], net452[39], net452[40], net452[41],
     net452[42], net452[43], net452[44], net452[45], net452[46],
     net452[47]}), .sp4_v_b_02({net453[0], net453[1], net453[2],
     net453[3], net453[4], net453[5], net453[6], net453[7], net453[8],
     net453[9], net453[10], net453[11], net453[12], net453[13],
     net453[14], net453[15], net453[16], net453[17], net453[18],
     net453[19], net453[20], net453[21], net453[22], net453[23],
     net453[24], net453[25], net453[26], net453[27], net453[28],
     net453[29], net453[30], net453[31], net453[32], net453[33],
     net453[34], net453[35], net453[36], net453[37], net453[38],
     net453[39], net453[40], net453[41], net453[42], net453[43],
     net453[44], net453[45], net453[46], net453[47]}),
     .bnr_op_01(bnr_op_01_05[7:0]), .tnr_op_04({slf_op_02_09[3],
     slf_op_02_09[2], slf_op_02_09[1], slf_op_02_09[0],
     slf_op_02_09[3], slf_op_02_09[2], slf_op_02_09[1],
     slf_op_02_09[0]}), .glb_netwk(glb_in_1[7:0]),
     .tnl_op_04({tiegnd_qtl, tiegnd_qtl, tiegnd_qtl, tiegnd_qtl,
     tiegnd_qtl, tiegnd_qtl, tiegnd_qtl, tiegnd_qtl}),
     .pgate(pgate_l[63:0]), .reset_b(reset_b_l[63:0]), .wl(wl_l[63:0]),
     .top_op_04({slf_op_01_09[3], slf_op_01_09[2], slf_op_01_09[1],
     slf_op_01_09[0], slf_op_01_09[3], slf_op_01_09[2],
     slf_op_01_09[1], slf_op_01_09[0]}), .lc_bot(lc_bot_01_05),
     .op_vic(net463), .sp12_v_b_01(sp12_v_b_01_05[23:0]),
     .sp4_v_t_04({net465[0], net465[1], net465[2], net465[3],
     net465[4], net465[5], net465[6], net465[7], net465[8], net465[9],
     net465[10], net465[11], net465[12], net465[13], net465[14],
     net465[15], net465[16], net465[17], net465[18], net465[19],
     net465[20], net465[21], net465[22], net465[23], net465[24],
     net465[25], net465[26], net465[27], net465[28], net465[29],
     net465[30], net465[31], net465[32], net465[33], net465[34],
     net465[35], net465[36], net465[37], net465[38], net465[39],
     net465[40], net465[41], net465[42], net465[43], net465[44],
     net465[45], net465[46], net465[47]}), .sp12_v_t_04({net466[0],
     net466[1], net466[2], net466[3], net466[4], net466[5], net466[6],
     net466[7], net466[8], net466[9], net466[10], net466[11],
     net466[12], net466[13], net466[14], net466[15], net466[16],
     net466[17], net466[18], net466[19], net466[20], net466[21],
     net466[22], net466[23]}));
lt_1x4_top_ice384 I399 ( .rgt_op_03(slf_op_03_07[7:0]),
     .slf_op_02({net412[0], net412[1], net412[2], net412[3], net412[4],
     net412[5], net412[6], net412[7]}), .rgt_op_02(slf_op_03_06[7:0]),
     .rgt_op_01(slf_op_03_05[7:0]), .purst(purst), .prog(prog),
     .lft_op_04({net357[0], net357[1], net357[2], net357[3], net357[4],
     net357[5], net357[6], net357[7]}), .lft_op_03({net337[0],
     net337[1], net337[2], net337[3], net337[4], net337[5], net337[6],
     net337[7]}), .lft_op_02({net330[0], net330[1], net330[2],
     net330[3], net330[4], net330[5], net330[6], net330[7]}),
     .lft_op_01(slf_op_01_05[7:0]), .rgt_op_04(slf_op_03_08[7:0]),
     .carry_in(carry_in_02_05), .bnl_op_01(bnl_op_02_05[7:0]),
     .slf_op_04({net420[0], net420[1], net420[2], net420[3], net420[4],
     net420[5], net420[6], net420[7]}), .slf_op_03({net410[0],
     net410[1], net410[2], net410[3], net410[4], net410[5], net410[6],
     net410[7]}), .slf_op_01(slf_op_02_05[7:0]),
     .sp4_h_l_04({net438[0], net438[1], net438[2], net438[3],
     net438[4], net438[5], net438[6], net438[7], net438[8], net438[9],
     net438[10], net438[11], net438[12], net438[13], net438[14],
     net438[15], net438[16], net438[17], net438[18], net438[19],
     net438[20], net438[21], net438[22], net438[23], net438[24],
     net438[25], net438[26], net438[27], net438[28], net438[29],
     net438[30], net438[31], net438[32], net438[33], net438[34],
     net438[35], net438[36], net438[37], net438[38], net438[39],
     net438[40], net438[41], net438[42], net438[43], net438[44],
     net438[45], net438[46], net438[47]}), .carry_out(net484),
     .vdd_cntl(vdd_cntl_l[63:0]), .sp12_h_r_04({net486[0], net486[1],
     net486[2], net486[3], net486[4], net486[5], net486[6], net486[7],
     net486[8], net486[9], net486[10], net486[11], net486[12],
     net486[13], net486[14], net486[15], net486[16], net486[17],
     net486[18], net486[19], net486[20], net486[21], net486[22],
     net486[23]}), .sp12_h_r_03({net487[0], net487[1], net487[2],
     net487[3], net487[4], net487[5], net487[6], net487[7], net487[8],
     net487[9], net487[10], net487[11], net487[12], net487[13],
     net487[14], net487[15], net487[16], net487[17], net487[18],
     net487[19], net487[20], net487[21], net487[22], net487[23]}),
     .sp12_h_r_02({net488[0], net488[1], net488[2], net488[3],
     net488[4], net488[5], net488[6], net488[7], net488[8], net488[9],
     net488[10], net488[11], net488[12], net488[13], net488[14],
     net488[15], net488[16], net488[17], net488[18], net488[19],
     net488[20], net488[21], net488[22], net488[23]}),
     .sp12_h_r_01({net489[0], net489[1], net489[2], net489[3],
     net489[4], net489[5], net489[6], net489[7], net489[8], net489[9],
     net489[10], net489[11], net489[12], net489[13], net489[14],
     net489[15], net489[16], net489[17], net489[18], net489[19],
     net489[20], net489[21], net489[22], net489[23]}),
     .sp4_v_b_01(sp4_v_b_02_05[47:0]), .sp4_r_v_b_04({net491[0],
     net491[1], net491[2], net491[3], net491[4], net491[5], net491[6],
     net491[7], net491[8], net491[9], net491[10], net491[11],
     net491[12], net491[13], net491[14], net491[15], net491[16],
     net491[17], net491[18], net491[19], net491[20], net491[21],
     net491[22], net491[23], net491[24], net491[25], net491[26],
     net491[27], net491[28], net491[29], net491[30], net491[31],
     net491[32], net491[33], net491[34], net491[35], net491[36],
     net491[37], net491[38], net491[39], net491[40], net491[41],
     net491[42], net491[43], net491[44], net491[45], net491[46],
     net491[47]}), .sp4_r_v_b_03({net492[0], net492[1], net492[2],
     net492[3], net492[4], net492[5], net492[6], net492[7], net492[8],
     net492[9], net492[10], net492[11], net492[12], net492[13],
     net492[14], net492[15], net492[16], net492[17], net492[18],
     net492[19], net492[20], net492[21], net492[22], net492[23],
     net492[24], net492[25], net492[26], net492[27], net492[28],
     net492[29], net492[30], net492[31], net492[32], net492[33],
     net492[34], net492[35], net492[36], net492[37], net492[38],
     net492[39], net492[40], net492[41], net492[42], net492[43],
     net492[44], net492[45], net492[46], net492[47]}),
     .sp4_r_v_b_02({net493[0], net493[1], net493[2], net493[3],
     net493[4], net493[5], net493[6], net493[7], net493[8], net493[9],
     net493[10], net493[11], net493[12], net493[13], net493[14],
     net493[15], net493[16], net493[17], net493[18], net493[19],
     net493[20], net493[21], net493[22], net493[23], net493[24],
     net493[25], net493[26], net493[27], net493[28], net493[29],
     net493[30], net493[31], net493[32], net493[33], net493[34],
     net493[35], net493[36], net493[37], net493[38], net493[39],
     net493[40], net493[41], net493[42], net493[43], net493[44],
     net493[45], net493[46], net493[47]}),
     .sp4_r_v_b_01(sp4_v_b_03_05[47:0]), .sp4_h_r_04({net495[0],
     net495[1], net495[2], net495[3], net495[4], net495[5], net495[6],
     net495[7], net495[8], net495[9], net495[10], net495[11],
     net495[12], net495[13], net495[14], net495[15], net495[16],
     net495[17], net495[18], net495[19], net495[20], net495[21],
     net495[22], net495[23], net495[24], net495[25], net495[26],
     net495[27], net495[28], net495[29], net495[30], net495[31],
     net495[32], net495[33], net495[34], net495[35], net495[36],
     net495[37], net495[38], net495[39], net495[40], net495[41],
     net495[42], net495[43], net495[44], net495[45], net495[46],
     net495[47]}), .sp4_h_r_03({net496[0], net496[1], net496[2],
     net496[3], net496[4], net496[5], net496[6], net496[7], net496[8],
     net496[9], net496[10], net496[11], net496[12], net496[13],
     net496[14], net496[15], net496[16], net496[17], net496[18],
     net496[19], net496[20], net496[21], net496[22], net496[23],
     net496[24], net496[25], net496[26], net496[27], net496[28],
     net496[29], net496[30], net496[31], net496[32], net496[33],
     net496[34], net496[35], net496[36], net496[37], net496[38],
     net496[39], net496[40], net496[41], net496[42], net496[43],
     net496[44], net496[45], net496[46], net496[47]}),
     .sp4_h_r_02({net497[0], net497[1], net497[2], net497[3],
     net497[4], net497[5], net497[6], net497[7], net497[8], net497[9],
     net497[10], net497[11], net497[12], net497[13], net497[14],
     net497[15], net497[16], net497[17], net497[18], net497[19],
     net497[20], net497[21], net497[22], net497[23], net497[24],
     net497[25], net497[26], net497[27], net497[28], net497[29],
     net497[30], net497[31], net497[32], net497[33], net497[34],
     net497[35], net497[36], net497[37], net497[38], net497[39],
     net497[40], net497[41], net497[42], net497[43], net497[44],
     net497[45], net497[46], net497[47]}), .sp4_h_r_01({net498[0],
     net498[1], net498[2], net498[3], net498[4], net498[5], net498[6],
     net498[7], net498[8], net498[9], net498[10], net498[11],
     net498[12], net498[13], net498[14], net498[15], net498[16],
     net498[17], net498[18], net498[19], net498[20], net498[21],
     net498[22], net498[23], net498[24], net498[25], net498[26],
     net498[27], net498[28], net498[29], net498[30], net498[31],
     net498[32], net498[33], net498[34], net498[35], net498[36],
     net498[37], net498[38], net498[39], net498[40], net498[41],
     net498[42], net498[43], net498[44], net498[45], net498[46],
     net498[47]}), .sp4_h_l_03({net439[0], net439[1], net439[2],
     net439[3], net439[4], net439[5], net439[6], net439[7], net439[8],
     net439[9], net439[10], net439[11], net439[12], net439[13],
     net439[14], net439[15], net439[16], net439[17], net439[18],
     net439[19], net439[20], net439[21], net439[22], net439[23],
     net439[24], net439[25], net439[26], net439[27], net439[28],
     net439[29], net439[30], net439[31], net439[32], net439[33],
     net439[34], net439[35], net439[36], net439[37], net439[38],
     net439[39], net439[40], net439[41], net439[42], net439[43],
     net439[44], net439[45], net439[46], net439[47]}),
     .sp4_h_l_02({net440[0], net440[1], net440[2], net440[3],
     net440[4], net440[5], net440[6], net440[7], net440[8], net440[9],
     net440[10], net440[11], net440[12], net440[13], net440[14],
     net440[15], net440[16], net440[17], net440[18], net440[19],
     net440[20], net440[21], net440[22], net440[23], net440[24],
     net440[25], net440[26], net440[27], net440[28], net440[29],
     net440[30], net440[31], net440[32], net440[33], net440[34],
     net440[35], net440[36], net440[37], net440[38], net440[39],
     net440[40], net440[41], net440[42], net440[43], net440[44],
     net440[45], net440[46], net440[47]}), .sp4_h_l_01({net441[0],
     net441[1], net441[2], net441[3], net441[4], net441[5], net441[6],
     net441[7], net441[8], net441[9], net441[10], net441[11],
     net441[12], net441[13], net441[14], net441[15], net441[16],
     net441[17], net441[18], net441[19], net441[20], net441[21],
     net441[22], net441[23], net441[24], net441[25], net441[26],
     net441[27], net441[28], net441[29], net441[30], net441[31],
     net441[32], net441[33], net441[34], net441[35], net441[36],
     net441[37], net441[38], net441[39], net441[40], net441[41],
     net441[42], net441[43], net441[44], net441[45], net441[46],
     net441[47]}), .bl(bl[125:72]), .bot_op_01(bot_op_02_05[7:0]),
     .sp12_h_l_01({net432[0], net432[1], net432[2], net432[3],
     net432[4], net432[5], net432[6], net432[7], net432[8], net432[9],
     net432[10], net432[11], net432[12], net432[13], net432[14],
     net432[15], net432[16], net432[17], net432[18], net432[19],
     net432[20], net432[21], net432[22], net432[23]}),
     .sp12_h_l_02({net431[0], net431[1], net431[2], net431[3],
     net431[4], net431[5], net431[6], net431[7], net431[8], net431[9],
     net431[10], net431[11], net431[12], net431[13], net431[14],
     net431[15], net431[16], net431[17], net431[18], net431[19],
     net431[20], net431[21], net431[22], net431[23]}),
     .sp12_h_l_03({net430[0], net430[1], net430[2], net430[3],
     net430[4], net430[5], net430[6], net430[7], net430[8], net430[9],
     net430[10], net430[11], net430[12], net430[13], net430[14],
     net430[15], net430[16], net430[17], net430[18], net430[19],
     net430[20], net430[21], net430[22], net430[23]}),
     .sp12_h_l_04({net429[0], net429[1], net429[2], net429[3],
     net429[4], net429[5], net429[6], net429[7], net429[8], net429[9],
     net429[10], net429[11], net429[12], net429[13], net429[14],
     net429[15], net429[16], net429[17], net429[18], net429[19],
     net429[20], net429[21], net429[22], net429[23]}),
     .sp4_v_b_04({net434[0], net434[1], net434[2], net434[3],
     net434[4], net434[5], net434[6], net434[7], net434[8], net434[9],
     net434[10], net434[11], net434[12], net434[13], net434[14],
     net434[15], net434[16], net434[17], net434[18], net434[19],
     net434[20], net434[21], net434[22], net434[23], net434[24],
     net434[25], net434[26], net434[27], net434[28], net434[29],
     net434[30], net434[31], net434[32], net434[33], net434[34],
     net434[35], net434[36], net434[37], net434[38], net434[39],
     net434[40], net434[41], net434[42], net434[43], net434[44],
     net434[45], net434[46], net434[47]}), .sp4_v_b_03({net435[0],
     net435[1], net435[2], net435[3], net435[4], net435[5], net435[6],
     net435[7], net435[8], net435[9], net435[10], net435[11],
     net435[12], net435[13], net435[14], net435[15], net435[16],
     net435[17], net435[18], net435[19], net435[20], net435[21],
     net435[22], net435[23], net435[24], net435[25], net435[26],
     net435[27], net435[28], net435[29], net435[30], net435[31],
     net435[32], net435[33], net435[34], net435[35], net435[36],
     net435[37], net435[38], net435[39], net435[40], net435[41],
     net435[42], net435[43], net435[44], net435[45], net435[46],
     net435[47]}), .sp4_v_b_02({net436[0], net436[1], net436[2],
     net436[3], net436[4], net436[5], net436[6], net436[7], net436[8],
     net436[9], net436[10], net436[11], net436[12], net436[13],
     net436[14], net436[15], net436[16], net436[17], net436[18],
     net436[19], net436[20], net436[21], net436[22], net436[23],
     net436[24], net436[25], net436[26], net436[27], net436[28],
     net436[29], net436[30], net436[31], net436[32], net436[33],
     net436[34], net436[35], net436[36], net436[37], net436[38],
     net436[39], net436[40], net436[41], net436[42], net436[43],
     net436[44], net436[45], net436[46], net436[47]}),
     .bnr_op_01(bnr_op_02_05[7:0]), .tnr_op_04({slf_op_03_09[3],
     slf_op_03_09[2], slf_op_03_09[1], slf_op_03_09[0],
     slf_op_03_09[3], slf_op_03_09[2], slf_op_03_09[1],
     slf_op_03_09[0]}), .glb_netwk(glb_in_2[7:0]),
     .tnl_op_04({slf_op_01_09[3], slf_op_01_09[2], slf_op_01_09[1],
     slf_op_01_09[0], slf_op_01_09[3], slf_op_01_09[2],
     slf_op_01_09[1], slf_op_01_09[0]}), .pgate(pgate_l[63:0]),
     .reset_b(reset_b_l[63:0]), .wl(wl_l[63:0]),
     .top_op_04({slf_op_02_09[3], slf_op_02_09[2], slf_op_02_09[1],
     slf_op_02_09[0], slf_op_02_09[3], slf_op_02_09[2],
     slf_op_02_09[1], slf_op_02_09[0]}), .lc_bot(lc_bot_02_05),
     .op_vic(net520), .sp12_v_b_01(sp12_v_b_02_05[23:0]),
     .sp4_v_t_04({net522[0], net522[1], net522[2], net522[3],
     net522[4], net522[5], net522[6], net522[7], net522[8], net522[9],
     net522[10], net522[11], net522[12], net522[13], net522[14],
     net522[15], net522[16], net522[17], net522[18], net522[19],
     net522[20], net522[21], net522[22], net522[23], net522[24],
     net522[25], net522[26], net522[27], net522[28], net522[29],
     net522[30], net522[31], net522[32], net522[33], net522[34],
     net522[35], net522[36], net522[37], net522[38], net522[39],
     net522[40], net522[41], net522[42], net522[43], net522[44],
     net522[45], net522[46], net522[47]}), .sp12_v_t_04({net523[0],
     net523[1], net523[2], net523[3], net523[4], net523[5], net523[6],
     net523[7], net523[8], net523[9], net523[10], net523[11],
     net523[12], net523[13], net523[14], net523[15], net523[16],
     net523[17], net523[18], net523[19], net523[20], net523[21],
     net523[22], net523[23]}));
lt_1x4_top_ice384 I400 ( .rgt_op_03(rgt_op_03_07[7:0]),
     .slf_op_02(slf_op_03_06[7:0]), .rgt_op_02(rgt_op_03_06[7:0]),
     .rgt_op_01(rgt_op_03_05[7:0]), .purst(purst), .prog(prog),
     .lft_op_04({net420[0], net420[1], net420[2], net420[3], net420[4],
     net420[5], net420[6], net420[7]}), .lft_op_03({net410[0],
     net410[1], net410[2], net410[3], net410[4], net410[5], net410[6],
     net410[7]}), .lft_op_02({net412[0], net412[1], net412[2],
     net412[3], net412[4], net412[5], net412[6], net412[7]}),
     .lft_op_01(slf_op_02_05[7:0]), .rgt_op_04(rgt_op_03_08[7:0]),
     .carry_in(carry_in_03_05), .bnl_op_01(bnl_op_03_05[7:0]),
     .slf_op_04(slf_op_03_08[7:0]), .slf_op_03(slf_op_03_07[7:0]),
     .slf_op_01(slf_op_03_05[7:0]), .sp4_h_l_04({net495[0], net495[1],
     net495[2], net495[3], net495[4], net495[5], net495[6], net495[7],
     net495[8], net495[9], net495[10], net495[11], net495[12],
     net495[13], net495[14], net495[15], net495[16], net495[17],
     net495[18], net495[19], net495[20], net495[21], net495[22],
     net495[23], net495[24], net495[25], net495[26], net495[27],
     net495[28], net495[29], net495[30], net495[31], net495[32],
     net495[33], net495[34], net495[35], net495[36], net495[37],
     net495[38], net495[39], net495[40], net495[41], net495[42],
     net495[43], net495[44], net495[45], net495[46], net495[47]}),
     .carry_out(net541), .vdd_cntl(vdd_cntl_l[63:0]),
     .sp12_h_r_04(sp12_h_r_03_08[23:0]),
     .sp12_h_r_03(sp12_h_r_03_07[23:0]),
     .sp12_h_r_02(sp12_h_r_03_06[23:0]),
     .sp12_h_r_01(sp12_h_r_03_05[23:0]),
     .sp4_v_b_01(sp4_v_b_03_05[47:0]),
     .sp4_r_v_b_04(sp4_r_v_b_03_08[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_03_07[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_03_06[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_03_05[47:0]),
     .sp4_h_r_04(sp4_h_r_03_08[47:0]),
     .sp4_h_r_03(sp4_h_r_03_07[47:0]),
     .sp4_h_r_02(sp4_h_r_03_06[47:0]),
     .sp4_h_r_01(sp4_h_r_03_05[47:0]), .sp4_h_l_03({net496[0],
     net496[1], net496[2], net496[3], net496[4], net496[5], net496[6],
     net496[7], net496[8], net496[9], net496[10], net496[11],
     net496[12], net496[13], net496[14], net496[15], net496[16],
     net496[17], net496[18], net496[19], net496[20], net496[21],
     net496[22], net496[23], net496[24], net496[25], net496[26],
     net496[27], net496[28], net496[29], net496[30], net496[31],
     net496[32], net496[33], net496[34], net496[35], net496[36],
     net496[37], net496[38], net496[39], net496[40], net496[41],
     net496[42], net496[43], net496[44], net496[45], net496[46],
     net496[47]}), .sp4_h_l_02({net497[0], net497[1], net497[2],
     net497[3], net497[4], net497[5], net497[6], net497[7], net497[8],
     net497[9], net497[10], net497[11], net497[12], net497[13],
     net497[14], net497[15], net497[16], net497[17], net497[18],
     net497[19], net497[20], net497[21], net497[22], net497[23],
     net497[24], net497[25], net497[26], net497[27], net497[28],
     net497[29], net497[30], net497[31], net497[32], net497[33],
     net497[34], net497[35], net497[36], net497[37], net497[38],
     net497[39], net497[40], net497[41], net497[42], net497[43],
     net497[44], net497[45], net497[46], net497[47]}),
     .sp4_h_l_01({net498[0], net498[1], net498[2], net498[3],
     net498[4], net498[5], net498[6], net498[7], net498[8], net498[9],
     net498[10], net498[11], net498[12], net498[13], net498[14],
     net498[15], net498[16], net498[17], net498[18], net498[19],
     net498[20], net498[21], net498[22], net498[23], net498[24],
     net498[25], net498[26], net498[27], net498[28], net498[29],
     net498[30], net498[31], net498[32], net498[33], net498[34],
     net498[35], net498[36], net498[37], net498[38], net498[39],
     net498[40], net498[41], net498[42], net498[43], net498[44],
     net498[45], net498[46], net498[47]}), .bl(bl[179:126]),
     .bot_op_01(bot_op_03_05[7:0]), .sp12_h_l_01({net489[0], net489[1],
     net489[2], net489[3], net489[4], net489[5], net489[6], net489[7],
     net489[8], net489[9], net489[10], net489[11], net489[12],
     net489[13], net489[14], net489[15], net489[16], net489[17],
     net489[18], net489[19], net489[20], net489[21], net489[22],
     net489[23]}), .sp12_h_l_02({net488[0], net488[1], net488[2],
     net488[3], net488[4], net488[5], net488[6], net488[7], net488[8],
     net488[9], net488[10], net488[11], net488[12], net488[13],
     net488[14], net488[15], net488[16], net488[17], net488[18],
     net488[19], net488[20], net488[21], net488[22], net488[23]}),
     .sp12_h_l_03({net487[0], net487[1], net487[2], net487[3],
     net487[4], net487[5], net487[6], net487[7], net487[8], net487[9],
     net487[10], net487[11], net487[12], net487[13], net487[14],
     net487[15], net487[16], net487[17], net487[18], net487[19],
     net487[20], net487[21], net487[22], net487[23]}),
     .sp12_h_l_04({net486[0], net486[1], net486[2], net486[3],
     net486[4], net486[5], net486[6], net486[7], net486[8], net486[9],
     net486[10], net486[11], net486[12], net486[13], net486[14],
     net486[15], net486[16], net486[17], net486[18], net486[19],
     net486[20], net486[21], net486[22], net486[23]}),
     .sp4_v_b_04({net491[0], net491[1], net491[2], net491[3],
     net491[4], net491[5], net491[6], net491[7], net491[8], net491[9],
     net491[10], net491[11], net491[12], net491[13], net491[14],
     net491[15], net491[16], net491[17], net491[18], net491[19],
     net491[20], net491[21], net491[22], net491[23], net491[24],
     net491[25], net491[26], net491[27], net491[28], net491[29],
     net491[30], net491[31], net491[32], net491[33], net491[34],
     net491[35], net491[36], net491[37], net491[38], net491[39],
     net491[40], net491[41], net491[42], net491[43], net491[44],
     net491[45], net491[46], net491[47]}), .sp4_v_b_03({net492[0],
     net492[1], net492[2], net492[3], net492[4], net492[5], net492[6],
     net492[7], net492[8], net492[9], net492[10], net492[11],
     net492[12], net492[13], net492[14], net492[15], net492[16],
     net492[17], net492[18], net492[19], net492[20], net492[21],
     net492[22], net492[23], net492[24], net492[25], net492[26],
     net492[27], net492[28], net492[29], net492[30], net492[31],
     net492[32], net492[33], net492[34], net492[35], net492[36],
     net492[37], net492[38], net492[39], net492[40], net492[41],
     net492[42], net492[43], net492[44], net492[45], net492[46],
     net492[47]}), .sp4_v_b_02({net493[0], net493[1], net493[2],
     net493[3], net493[4], net493[5], net493[6], net493[7], net493[8],
     net493[9], net493[10], net493[11], net493[12], net493[13],
     net493[14], net493[15], net493[16], net493[17], net493[18],
     net493[19], net493[20], net493[21], net493[22], net493[23],
     net493[24], net493[25], net493[26], net493[27], net493[28],
     net493[29], net493[30], net493[31], net493[32], net493[33],
     net493[34], net493[35], net493[36], net493[37], net493[38],
     net493[39], net493[40], net493[41], net493[42], net493[43],
     net493[44], net493[45], net493[46], net493[47]}),
     .bnr_op_01(bnr_op_03_05[7:0]), .tnr_op_04({tnr_op_03_08[3],
     tnr_op_03_08[2], tnr_op_03_08[1], tnr_op_03_08[0],
     tnr_op_03_08[3], tnr_op_03_08[2], tnr_op_03_08[1],
     tnr_op_03_08[0]}), .glb_netwk(glb_in_3[7:0]),
     .tnl_op_04({slf_op_02_09[3], slf_op_02_09[2], slf_op_02_09[1],
     slf_op_02_09[0], slf_op_02_09[3], slf_op_02_09[2],
     slf_op_02_09[1], slf_op_02_09[0]}), .pgate(pgate_l[63:0]),
     .reset_b(reset_b_l[63:0]), .wl(wl_l[63:0]),
     .top_op_04({slf_op_03_09[3], slf_op_03_09[2], slf_op_03_09[1],
     slf_op_03_09[0], slf_op_03_09[3], slf_op_03_09[2],
     slf_op_03_09[1], slf_op_03_09[0]}), .lc_bot(lc_bot_03_05),
     .op_vic(net577), .sp12_v_b_01(sp12_v_b_03_05[23:0]),
     .sp4_v_t_04({net579[0], net579[1], net579[2], net579[3],
     net579[4], net579[5], net579[6], net579[7], net579[8], net579[9],
     net579[10], net579[11], net579[12], net579[13], net579[14],
     net579[15], net579[16], net579[17], net579[18], net579[19],
     net579[20], net579[21], net579[22], net579[23], net579[24],
     net579[25], net579[26], net579[27], net579[28], net579[29],
     net579[30], net579[31], net579[32], net579[33], net579[34],
     net579[35], net579[36], net579[37], net579[38], net579[39],
     net579[40], net579[41], net579[42], net579[43], net579[44],
     net579[45], net579[46], net579[47]}), .sp12_v_t_04({net580[0],
     net580[1], net580[2], net580[3], net580[4], net580[5], net580[6],
     net580[7], net580[8], net580[9], net580[10], net580[11],
     net580[12], net580[13], net580[14], net580[15], net580[16],
     net580[17], net580[18], net580[19], net580[20], net580[21],
     net580[22], net580[23]}));
pinlatbuf12p I389 ( .pad_in(padin_t_l[5]), .icegate(hold_t_l),
     .cbit(cf_top_l[63]), .cout(net584), .prog(prog));
pinlatbuf12p I_pinlatbuf12p_l ( .pad_in(padin_l_t[8]),
     .icegate(hold_l_t), .cbit(cf_l[15]), .cout(net614), .prog(prog));
tielo I369 ( .tielo(tiegnd_qtl));
scan_buf_ice8p I_scanbuf_8p_tl ( .update_i(net592), .tclk_i(net593),
     .shift_i(net594), .sdi(net595), .r_i(net596), .mode_i(net597),
     .hiz_b_i(net598), .ceb_i(net599), .bs_en_i(net600),
     .update_o(update_o), .tclk_o(net328), .shift_o(shift_o),
     .sdo(net316), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
fabric_buf_ice8p I390 ( .f_in(net584), .f_out(padin_03_09b));
fabric_buf_ice8p I391 ( .f_in(net614), .f_out(padin_00_05a));

endmodule
// Library - ice8chip, Cell - clk_mux_2to1_ice8p, View - schematic
// LAST TIME SAVED: Jul 30 23:15:00 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module clk_mux_2to1_ice8p ( clk, cbit, cbitb, min, prog );
output  clk;

input  cbit, cbitb, prog;

input [1:0]  min;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I_inv0 ( .A(prog), .Y(net030));
nand2_lvt I_nand2_1 ( .A(st2), .Y(clkb), .B(net030));
inv_lvt I_inv2 ( .A(clkb), .Y(clk));
txgate_lvt I_txgate_hvt0 ( .in(min[0]), .out(st2), .pp(cbit),
     .nn(cbitb));
txgate_lvt I_txgate_hvt1 ( .in(min[1]), .out(st2), .pp(cbitb),
     .nn(cbit));

endmodule
// Library - ice8chip, Cell - clk_mux2to1_ice8p, View - schematic
// LAST TIME SAVED: Aug  3 19:20:01 2011
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module clk_mux2to1_ice8p ( gnet, bl, min0, min1, min2, min3, pgate_l,
     pgate_r, prog, reset_l, reset_r, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r );


input  prog;

output [3:0]  gnet;

inout [3:0]  bl;

input [1:0]  wl_r;
input [1:0]  min1;
input [1:0]  pgate_l;
input [1:0]  min0;
input [1:0]  reset_r;
input [1:0]  wl_l;
input [1:0]  reset_l;
input [1:0]  vdd_cntl_l;
input [1:0]  vdd_cntl_r;
input [1:0]  pgate_r;
input [1:0]  min2;
input [1:0]  min3;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  l_vdd;

wire  [1:0]  r_vdd;

wire  [7:0]  cbitb;

wire  [7:0]  cbit;



P_11_LPHVT  I_pch_hvt_l_1_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl_l[1]),
     .D(l_vdd[0]));
P_11_LPHVT  I_pch_hvt_l_0_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl_l[0]),
     .D(l_vdd[1]));
P_11_LPHVT  M0_1_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl_r[1]),
     .D(r_vdd[1]));
P_11_LPHVT  M0_0_ ( .S(vdd_), .B(vdd_), .G(vdd_cntl_r[0]),
     .D(r_vdd[0]));
clk_mux_2to1_ice8p I_clkmux3 ( .prog(prog), .cbit(cbit[3]),
     .cbitb(cbitb[3]), .min(min3[1:0]), .clk(gnet[3]));
clk_mux_2to1_ice8p I_clkmux1 ( .prog(prog), .cbit(cbit[1]),
     .cbitb(cbitb[1]), .min(min1[1:0]), .clk(gnet[1]));
clk_mux_2to1_ice8p I_clkmux2 ( .prog(prog), .cbit(cbit[2]),
     .cbitb(cbitb[2]), .min(min2[1:0]), .clk(gnet[2]));
clk_mux_2to1_ice8p I_clkmux0 ( .prog(prog), .cbit(cbit[0]),
     .cbitb(cbitb[0]), .min(min0[1:0]), .clk(gnet[0]));
cram2x2 I_cram2x2_lft ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset_l[1:0]), .q(cbit[3:0]), .wl(wl_l[1:0]),
     .r_vdd({l_vdd[0], l_vdd[1]}), .pgate(pgate_l[1:0]));
cram2x2 I_cram2x2_rgt ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset_r[1:0]), .q(cbit[7:4]), .wl(wl_r[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate_r[1:0]));

endmodule
// Library - ice384chip, Cell - quad_x4_ice384, View - schematic
// LAST TIME SAVED: Jan 13 16:44:53 2012
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module quad_x4_ice384 ( cf_b[143:0], cf_l[191:0], cf_r[191:0],
     cf_t[143:0], padeb_b[11:0], padeb_l[15:0], padeb_r[15:0],
     padeb_t[11:0], pado_b[11:0], pado_l[15:0], pado_r[15:0],
     pado_t[11:0], sdo_pad, spi_ss_in_bbank[4:0], tck_pad, tdi_pad,
     tms_pad, bl_bot[363:0], bl_top[363:0], bs_en, ceb, end_of_startup,
     hiz_b, jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[0],
     last_rsr[1], last_rsr[2], last_rsr[3], md_spi_b, mode,
     mux_jtag_sel_b, padin_b[11:0], padin_l[15:0], padin_r[15:0],
     padin_t[11:0], pgate_l[159:0], pgate_r[159:0], prog, purst, r,
     reset_b_l[159:0], reset_b_r[159:0], sdi_pad, sdo_enable, shift,
     spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out, tclk, totdopad,
     trstb_pad, update, vdd_cntl_l[159:0], vdd_cntl_r[159:0],
     wl_l[159:0], wl_r[159:0] );
output  sdo_pad, tck_pad, tdi_pad, tms_pad;


input  bs_en, ceb, end_of_startup, hiz_b, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, md_spi_b, mode, mux_jtag_sel_b, prog,
     purst, r, sdi_pad, sdo_enable, shift, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk, totdopad, trstb_pad, update;

output [4:0]  spi_ss_in_bbank;
output [15:0]  pado_r;
output [11:0]  pado_t;
output [191:0]  cf_l;
output [15:0]  pado_l;
output [191:0]  cf_r;
output [15:0]  padeb_l;
output [11:0]  padeb_t;
output [15:0]  padeb_r;
output [143:0]  cf_t;
output [11:0]  padeb_b;
output [11:0]  pado_b;
output [143:0]  cf_b;

inout [363:0]  bl_top;
inout [363:0]  bl_bot;

input [11:0]  padin_t;
input [159:0]  vdd_cntl_l;
input [15:0]  padin_r;
input [11:0]  padin_b;
input [159:0]  pgate_l;
input [159:0]  wl_l;
input [15:0]  padin_l;
input [3:0]  last_rsr;
input [159:0]  pgate_r;
input [159:0]  reset_b_r;
input [159:0]  vdd_cntl_r;
input [159:0]  reset_b_l;
input [159:0]  wl_r;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [47:0]  net492;

wire  [7:0]  net454;

wire  [7:0]  net589;

wire  [7:0]  net713;

wire  [3:0]  slf_op_01_04;

wire  [7:0]  gclk;

wire  [47:0]  net795;

wire  [23:0]  net794;

wire  [7:0]  net579;

wire  [3:0]  net790;

wire  [7:0]  net484;

wire  [23:0]  net487;

wire  [23:0]  net496;

wire  [47:0]  net602;

wire  [7:0]  net599;

wire  [7:0]  net483;

wire  [47:0]  net810;

wire  [15:0]  net513;

wire  [7:0]  net0471;

wire  [47:0]  net489;

wire  [7:0]  net767;

wire  [7:0]  net766;

wire  [47:0]  net498;

wire  [23:0]  net595;

wire  [7:0]  net481;

wire  [7:0]  net469;

wire  [47:0]  net467;

wire  [7:0]  net430;

wire  [47:0]  net499;

wire  [47:0]  net465;

wire  [7:0]  net580;

wire  [3:0]  net470;

wire  [23:0]  net451;

wire  [23:0]  net812;

wire  [3:0]  net461;

wire  [7:0]  net802;

wire  [23:0]  net488;

wire  [7:0]  net0504;

wire  [7:0]  net471;

wire  [7:0]  net764;

wire  [7:0]  net801;

wire  [7:0]  net608;

wire  [7:0]  net466;

wire  [7:0]  net468;

wire  [47:0]  net808;

wire  [7:0]  net472;

wire  [7:0]  net800;

wire  [23:0]  net477;

wire  [15:0]  net814;

wire  [15:0]  net505;

wire  [23:0]  net815;

wire  [3:0]  slf_op_07_05;

wire  [7:0]  net459;

wire  [47:0]  net494;

wire  [23:0]  net813;

wire  [7:0]  net598;

wire  [23:0]  net596;

wire  [47:0]  net781;

wire  [47:0]  net485;

wire  [47:0]  net601;

wire  [23:0]  net597;

wire  [3:0]  net826;

wire  [3:0]  slf_op_00_04;

wire  [47:0]  net779;

wire  [47:0]  net809;

wire  [7:0]  net460;

wire  [7:0]  net607;

wire  [23:0]  net503;

wire  [15:0]  net603;

wire  [47:0]  net588;

wire  [7:0]  net765;

wire  [7:0]  net455;

wire  [47:0]  net495;

wire  [47:0]  net811;

wire  [47:0]  net456;

wire  [23:0]  net486;

wire  [7:0]  net491;

wire  [47:0]  net497;

wire  [3:0]  slf_op_07_04;

wire  [7:0]  net478;



quad_clk_drv_l Iquad_clk_drv__lleft ( .gclk(gclk[7:0]),
     .glb_in_2({net0504[0], net0504[1], net0504[2], net0504[3],
     net0504[4], net0504[5], net0504[6], net0504[7]}),
     .glb_in_3({net481[0], net481[1], net481[2], net481[3], net481[4],
     net481[5], net481[6], net481[7]}), .glb_in_1({net0471[0],
     net0471[1], net0471[2], net0471[3], net0471[4], net0471[5],
     net0471[6], net0471[7]}), .glb_in_0({net491[0], net491[1],
     net491[2], net491[3], net491[4], net491[5], net491[6],
     net491[7]}));
quad_clk_drv Iquad_clk_drv_rgt ( .gclk(gclk[7:0]),
     .glb_in_2({net580[0], net580[1], net580[2], net580[3], net580[4],
     net580[5], net580[6], net580[7]}), .glb_in_3({net579[0],
     net579[1], net579[2], net579[3], net579[4], net579[5], net579[6],
     net579[7]}), .glb_in_1({net713[0], net713[1], net713[2],
     net713[3], net713[4], net713[5], net713[6], net713[7]}),
     .glb_in_0({net430[0], net430[1], net430[2], net430[3], net430[4],
     net430[5], net430[6], net430[7]}));
ice384_cram_row78col4 Icram_row78col4_bot ( .wl_r(wl_r[77:0]),
     .vdd_cntl_r(vdd_cntl_r[77:0]), .reset_r(reset_b_r[77:0]),
     .pgate_r(pgate_r[77:0]), .pgate_l(pgate_l[77:0]),
     .wl_l(wl_l[77:0]), .vdd_cntl_l(vdd_cntl_l[77:0]),
     .reset_l(reset_b_l[77:0]), .bl(bl_bot[183:180]));
ice384_cram_row78col4 Icram_row78col4_top ( .wl_r(wl_r[159:82]),
     .vdd_cntl_r(vdd_cntl_r[159:82]), .reset_r(reset_b_r[159:82]),
     .pgate_r(pgate_r[159:82]), .pgate_l(pgate_l[159:82]),
     .wl_l(wl_l[159:82]), .vdd_cntl_l(vdd_cntl_l[159:82]),
     .reset_l(reset_b_l[159:82]), .bl(bl_top[183:180]));
quad_bl_ice384 i_bl_quad ( .padin_03_00b(padin_03_00b),
     .padin_00_04b(padin_00_04b), .sp12_v_t_03_04({net451[0],
     net451[1], net451[2], net451[3], net451[4], net451[5], net451[6],
     net451[7], net451[8], net451[9], net451[10], net451[11],
     net451[12], net451[13], net451[14], net451[15], net451[16],
     net451[17], net451[18], net451[19], net451[20], net451[21],
     net451[22], net451[23]}), .top_op_02_04({net455[0], net455[1],
     net455[2], net455[3], net455[4], net455[5], net455[6],
     net455[7]}), .top_op_01_04({net466[0], net466[1], net466[2],
     net466[3], net466[4], net466[5], net466[6], net466[7]}),
     .tnr_op_02_04({net454[0], net454[1], net454[2], net454[3],
     net454[4], net454[5], net454[6], net454[7]}),
     .tnr_op_01_04({net455[0], net455[1], net455[2], net455[3],
     net455[4], net455[5], net455[6], net455[7]}),
     .sp4_v_t_03_04({net456[0], net456[1], net456[2], net456[3],
     net456[4], net456[5], net456[6], net456[7], net456[8], net456[9],
     net456[10], net456[11], net456[12], net456[13], net456[14],
     net456[15], net456[16], net456[17], net456[18], net456[19],
     net456[20], net456[21], net456[22], net456[23], net456[24],
     net456[25], net456[26], net456[27], net456[28], net456[29],
     net456[30], net456[31], net456[32], net456[33], net456[34],
     net456[35], net456[36], net456[37], net456[38], net456[39],
     net456[40], net456[41], net456[42], net456[43], net456[44],
     net456[45], net456[46], net456[47]}), .glb_in_1({net0471[0],
     net0471[1], net0471[2], net0471[3], net0471[4], net0471[5],
     net0471[6], net0471[7]}), .tnl_op_02_04({net466[0], net466[1],
     net466[2], net466[3], net466[4], net466[5], net466[6],
     net466[7]}), .rgt_op_03_03({net459[0], net459[1], net459[2],
     net459[3], net459[4], net459[5], net459[6], net459[7]}),
     .rgt_op_03_02({net460[0], net460[1], net460[2], net460[3],
     net460[4], net460[5], net460[6], net460[7]}),
     .bnr_op_03_01({net461[0], net461[1], net461[2], net461[3]}),
     .rgt_op_03_04({net766[0], net766[1], net766[2], net766[3],
     net766[4], net766[5], net766[6], net766[7]}),
     .pado_b_l(pado_b[5:0]), .padin_l_b(padin_l[7:0]),
     .sp4_v_t_01_04({net465[0], net465[1], net465[2], net465[3],
     net465[4], net465[5], net465[6], net465[7], net465[8], net465[9],
     net465[10], net465[11], net465[12], net465[13], net465[14],
     net465[15], net465[16], net465[17], net465[18], net465[19],
     net465[20], net465[21], net465[22], net465[23], net465[24],
     net465[25], net465[26], net465[27], net465[28], net465[29],
     net465[30], net465[31], net465[32], net465[33], net465[34],
     net465[35], net465[36], net465[37], net465[38], net465[39],
     net465[40], net465[41], net465[42], net465[43], net465[44],
     net465[45], net465[46], net465[47]}), .tnr_op_00_04({net466[0],
     net466[1], net466[2], net466[3], net466[4], net466[5], net466[6],
     net466[7]}), .sp4_h_r_03_04({net467[0], net467[1], net467[2],
     net467[3], net467[4], net467[5], net467[6], net467[7], net467[8],
     net467[9], net467[10], net467[11], net467[12], net467[13],
     net467[14], net467[15], net467[16], net467[17], net467[18],
     net467[19], net467[20], net467[21], net467[22], net467[23],
     net467[24], net467[25], net467[26], net467[27], net467[28],
     net467[29], net467[30], net467[31], net467[32], net467[33],
     net467[34], net467[35], net467[36], net467[37], net467[38],
     net467[39], net467[40], net467[41], net467[42], net467[43],
     net467[44], net467[45], net467[46], net467[47]}),
     .slf_op_03_03({net468[0], net468[1], net468[2], net468[3],
     net468[4], net468[5], net468[6], net468[7]}),
     .slf_op_03_02({net469[0], net469[1], net469[2], net469[3],
     net469[4], net469[5], net469[6], net469[7]}),
     .slf_op_03_00({net470[0], net470[1], net470[2], net470[3]}),
     .slf_op_03_04({net471[0], net471[1], net471[2], net471[3],
     net471[4], net471[5], net471[6], net471[7]}),
     .slf_op_02_04({net472[0], net472[1], net472[2], net472[3],
     net472[4], net472[5], net472[6], net472[7]}),
     .padeb_b_l(padeb_b[5:0]), .padin_b_l(padin_b[5:0]),
     .padeb_l_b(padeb_l[7:0]), .fabric_out_00_04(fabric_out_00_04),
     .sp12_v_t_01_04({net477[0], net477[1], net477[2], net477[3],
     net477[4], net477[5], net477[6], net477[7], net477[8], net477[9],
     net477[10], net477[11], net477[12], net477[13], net477[14],
     net477[15], net477[16], net477[17], net477[18], net477[19],
     net477[20], net477[21], net477[22], net477[23]}),
     .slf_op_01_04({net478[0], net478[1], net478[2], net478[3],
     net478[4], net478[5], net478[6], net478[7]}),
     .carry_out_01_04(net479), .carry_out_03_04(net480),
     .glb_in_0({net491[0], net491[1], net491[2], net491[3], net491[4],
     net491[5], net491[6], net491[7]}), .vdd_cntl_l(vdd_cntl_l[79:0]),
     .rgt_op_03_01({net483[0], net483[1], net483[2], net483[3],
     net483[4], net483[5], net483[6], net483[7]}),
     .slf_op_03_01({net484[0], net484[1], net484[2], net484[3],
     net484[4], net484[5], net484[6], net484[7]}),
     .sp4_r_v_b_03_01({net485[0], net485[1], net485[2], net485[3],
     net485[4], net485[5], net485[6], net485[7], net485[8], net485[9],
     net485[10], net485[11], net485[12], net485[13], net485[14],
     net485[15], net485[16], net485[17], net485[18], net485[19],
     net485[20], net485[21], net485[22], net485[23], net485[24],
     net485[25], net485[26], net485[27], net485[28], net485[29],
     net485[30], net485[31], net485[32], net485[33], net485[34],
     net485[35], net485[36], net485[37], net485[38], net485[39],
     net485[40], net485[41], net485[42], net485[43], net485[44],
     net485[45], net485[46], net485[47]}), .sp12_h_r_03_03({net486[0],
     net486[1], net486[2], net486[3], net486[4], net486[5], net486[6],
     net486[7], net486[8], net486[9], net486[10], net486[11],
     net486[12], net486[13], net486[14], net486[15], net486[16],
     net486[17], net486[18], net486[19], net486[20], net486[21],
     net486[22], net486[23]}), .sp12_h_r_03_02({net487[0], net487[1],
     net487[2], net487[3], net487[4], net487[5], net487[6], net487[7],
     net487[8], net487[9], net487[10], net487[11], net487[12],
     net487[13], net487[14], net487[15], net487[16], net487[17],
     net487[18], net487[19], net487[20], net487[21], net487[22],
     net487[23]}), .sp12_h_r_03_01({net488[0], net488[1], net488[2],
     net488[3], net488[4], net488[5], net488[6], net488[7], net488[8],
     net488[9], net488[10], net488[11], net488[12], net488[13],
     net488[14], net488[15], net488[16], net488[17], net488[18],
     net488[19], net488[20], net488[21], net488[22], net488[23]}),
     .sp4_r_v_b_03_04({net489[0], net489[1], net489[2], net489[3],
     net489[4], net489[5], net489[6], net489[7], net489[8], net489[9],
     net489[10], net489[11], net489[12], net489[13], net489[14],
     net489[15], net489[16], net489[17], net489[18], net489[19],
     net489[20], net489[21], net489[22], net489[23], net489[24],
     net489[25], net489[26], net489[27], net489[28], net489[29],
     net489[30], net489[31], net489[32], net489[33], net489[34],
     net489[35], net489[36], net489[37], net489[38], net489[39],
     net489[40], net489[41], net489[42], net489[43], net489[44],
     net489[45], net489[46], net489[47]}), .glb_in_2({net0504[0],
     net0504[1], net0504[2], net0504[3], net0504[4], net0504[5],
     net0504[6], net0504[7]}), .glb_in_3({net481[0], net481[1],
     net481[2], net481[3], net481[4], net481[5], net481[6],
     net481[7]}), .sp4_v_t_02_04({net492[0], net492[1], net492[2],
     net492[3], net492[4], net492[5], net492[6], net492[7], net492[8],
     net492[9], net492[10], net492[11], net492[12], net492[13],
     net492[14], net492[15], net492[16], net492[17], net492[18],
     net492[19], net492[20], net492[21], net492[22], net492[23],
     net492[24], net492[25], net492[26], net492[27], net492[28],
     net492[29], net492[30], net492[31], net492[32], net492[33],
     net492[34], net492[35], net492[36], net492[37], net492[38],
     net492[39], net492[40], net492[41], net492[42], net492[43],
     net492[44], net492[45], net492[46], net492[47]}),
     .tnl_op_01_04({slf_op_01_04[3], slf_op_01_04[2], slf_op_01_04[1],
     slf_op_01_04[0], slf_op_01_04[3], slf_op_01_04[2],
     slf_op_01_04[1], slf_op_01_04[0]}), .sp4_r_v_b_03_03({net494[0],
     net494[1], net494[2], net494[3], net494[4], net494[5], net494[6],
     net494[7], net494[8], net494[9], net494[10], net494[11],
     net494[12], net494[13], net494[14], net494[15], net494[16],
     net494[17], net494[18], net494[19], net494[20], net494[21],
     net494[22], net494[23], net494[24], net494[25], net494[26],
     net494[27], net494[28], net494[29], net494[30], net494[31],
     net494[32], net494[33], net494[34], net494[35], net494[36],
     net494[37], net494[38], net494[39], net494[40], net494[41],
     net494[42], net494[43], net494[44], net494[45], net494[46],
     net494[47]}), .sp4_r_v_b_03_02({net495[0], net495[1], net495[2],
     net495[3], net495[4], net495[5], net495[6], net495[7], net495[8],
     net495[9], net495[10], net495[11], net495[12], net495[13],
     net495[14], net495[15], net495[16], net495[17], net495[18],
     net495[19], net495[20], net495[21], net495[22], net495[23],
     net495[24], net495[25], net495[26], net495[27], net495[28],
     net495[29], net495[30], net495[31], net495[32], net495[33],
     net495[34], net495[35], net495[36], net495[37], net495[38],
     net495[39], net495[40], net495[41], net495[42], net495[43],
     net495[44], net495[45], net495[46], net495[47]}),
     .sp12_h_r_03_04({net496[0], net496[1], net496[2], net496[3],
     net496[4], net496[5], net496[6], net496[7], net496[8], net496[9],
     net496[10], net496[11], net496[12], net496[13], net496[14],
     net496[15], net496[16], net496[17], net496[18], net496[19],
     net496[20], net496[21], net496[22], net496[23]}),
     .sp4_h_r_03_03({net497[0], net497[1], net497[2], net497[3],
     net497[4], net497[5], net497[6], net497[7], net497[8], net497[9],
     net497[10], net497[11], net497[12], net497[13], net497[14],
     net497[15], net497[16], net497[17], net497[18], net497[19],
     net497[20], net497[21], net497[22], net497[23], net497[24],
     net497[25], net497[26], net497[27], net497[28], net497[29],
     net497[30], net497[31], net497[32], net497[33], net497[34],
     net497[35], net497[36], net497[37], net497[38], net497[39],
     net497[40], net497[41], net497[42], net497[43], net497[44],
     net497[45], net497[46], net497[47]}), .sp4_h_r_03_02({net498[0],
     net498[1], net498[2], net498[3], net498[4], net498[5], net498[6],
     net498[7], net498[8], net498[9], net498[10], net498[11],
     net498[12], net498[13], net498[14], net498[15], net498[16],
     net498[17], net498[18], net498[19], net498[20], net498[21],
     net498[22], net498[23], net498[24], net498[25], net498[26],
     net498[27], net498[28], net498[29], net498[30], net498[31],
     net498[32], net498[33], net498[34], net498[35], net498[36],
     net498[37], net498[38], net498[39], net498[40], net498[41],
     net498[42], net498[43], net498[44], net498[45], net498[46],
     net498[47]}), .sp4_h_r_03_01({net499[0], net499[1], net499[2],
     net499[3], net499[4], net499[5], net499[6], net499[7], net499[8],
     net499[9], net499[10], net499[11], net499[12], net499[13],
     net499[14], net499[15], net499[16], net499[17], net499[18],
     net499[19], net499[20], net499[21], net499[22], net499[23],
     net499[24], net499[25], net499[26], net499[27], net499[28],
     net499[29], net499[30], net499[31], net499[32], net499[33],
     net499[34], net499[35], net499[36], net499[37], net499[38],
     net499[39], net499[40], net499[41], net499[42], net499[43],
     net499[44], net499[45], net499[46], net499[47]}),
     .tnr_op_03_04({net589[0], net589[1], net589[2], net589[3],
     net589[4], net589[5], net589[6], net589[7]}),
     .reset_b_l(reset_b_l[79:0]), .pgate_l(pgate_l[79:0]),
     .sp12_v_t_02_04({net503[0], net503[1], net503[2], net503[3],
     net503[4], net503[5], net503[6], net503[7], net503[8], net503[9],
     net503[10], net503[11], net503[12], net503[13], net503[14],
     net503[15], net503[16], net503[17], net503[18], net503[19],
     net503[20], net503[21], net503[22], net503[23]}),
     .bl(bl_bot[179:0]), .sp4_v_t_00_04({net505[0], net505[1],
     net505[2], net505[3], net505[4], net505[5], net505[6], net505[7],
     net505[8], net505[9], net505[10], net505[11], net505[12],
     net505[13], net505[14], net505[15]}), .pado_l_b(pado_l[7:0]),
     .fabric_out_03_00(fabric_out_03_00), .op_vic_03_04(op_vic_03),
     .op_vic_02_04(op_vic_02),
     .fabric_out_02_00(fabric_out_02_00_bicegate),
     .op_vic_01_04(op_vic_01), .carry_out_02_04(net512),
     .sp4_h_r_03_00({net513[0], net513[1], net513[2], net513[3],
     net513[4], net513[5], net513[6], net513[7], net513[8], net513[9],
     net513[10], net513[11], net513[12], net513[13], net513[14],
     net513[15]}), .fabric_out_00_03(fabric_out_00_03_licegate),
     .tnl_op_03_04({net455[0], net455[1], net455[2], net455[3],
     net455[4], net455[5], net455[6], net455[7]}),
     .top_op_03_04({net454[0], net454[1], net454[2], net454[3],
     net454[4], net454[5], net454[6], net454[7]}),
     .slf_op_00_04(slf_op_00_04[3:0]), .cf_b_l(cf_b[71:0]),
     .wl_l(wl_l[79:0]), .cf_l(cf_l[95:0]), .update_i(net521),
     .last_rsr(last_rsr[0]),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .tclk_i(tclkio_ml), .shift_i(net525), .sdi(sdio_ml), .r_i(net527),
     .purst(purst), .prog(prog), .mode_i(net530), .hiz_b_i(net531),
     .ceb_i(net532), .bs_en_i(net533), .update_o(net534),
     .tclk_o(tclkio_mb), .shift_o(net536), .sdo(sdio_mb), .r_o(net538),
     .mode_o(net539), .hiz_b_o(net540),
     .hold_b_l(fabric_out_02_00_bicegate),
     .hold_l_b(fabric_out_00_03_licegate), .ceb_o(net543),
     .bs_en_o(net544));
quad_br_ice384 i_br_quad ( .padin_07_04b(padin_07_04b),
     .slf_op_04_00({net461[0], net461[1], net461[2], net461[3]}),
     .slf_op_07_04(slf_op_07_04[3:0]), .padeb_b_r(padeb_b[11:6]),
     .op_vic_06_04(op_vic_06), .slf_op_04_02({net460[0], net460[1],
     net460[2], net460[3], net460[4], net460[5], net460[6],
     net460[7]}), .slf_op_04_01({net483[0], net483[1], net483[2],
     net483[3], net483[4], net483[5], net483[6], net483[7]}),
     .slf_op_04_03({net459[0], net459[1], net459[2], net459[3],
     net459[4], net459[5], net459[6], net459[7]}),
     .pado_b_r(pado_b[11:6]), .pado_r(pado_r[7:0]),
     .pgate_r(pgate_r[79:0]), .op_vic_05_04(op_vic_05),
     .sp12_h_l_04_01({net488[0], net488[1], net488[2], net488[3],
     net488[4], net488[5], net488[6], net488[7], net488[8], net488[9],
     net488[10], net488[11], net488[12], net488[13], net488[14],
     net488[15], net488[16], net488[17], net488[18], net488[19],
     net488[20], net488[21], net488[22], net488[23]}),
     .sp12_h_l_04_03({net486[0], net486[1], net486[2], net486[3],
     net486[4], net486[5], net486[6], net486[7], net486[8], net486[9],
     net486[10], net486[11], net486[12], net486[13], net486[14],
     net486[15], net486[16], net486[17], net486[18], net486[19],
     net486[20], net486[21], net486[22], net486[23]}),
     .sp12_h_l_04_02({net487[0], net487[1], net487[2], net487[3],
     net487[4], net487[5], net487[6], net487[7], net487[8], net487[9],
     net487[10], net487[11], net487[12], net487[13], net487[14],
     net487[15], net487[16], net487[17], net487[18], net487[19],
     net487[20], net487[21], net487[22], net487[23]}),
     .sp4_v_b_04_04({net489[0], net489[1], net489[2], net489[3],
     net489[4], net489[5], net489[6], net489[7], net489[8], net489[9],
     net489[10], net489[11], net489[12], net489[13], net489[14],
     net489[15], net489[16], net489[17], net489[18], net489[19],
     net489[20], net489[21], net489[22], net489[23], net489[24],
     net489[25], net489[26], net489[27], net489[28], net489[29],
     net489[30], net489[31], net489[32], net489[33], net489[34],
     net489[35], net489[36], net489[37], net489[38], net489[39],
     net489[40], net489[41], net489[42], net489[43], net489[44],
     net489[45], net489[46], net489[47]}), .slf_op_04_04({net766[0],
     net766[1], net766[2], net766[3], net766[4], net766[5], net766[6],
     net766[7]}), .sp4_v_b_04_03({net494[0], net494[1], net494[2],
     net494[3], net494[4], net494[5], net494[6], net494[7], net494[8],
     net494[9], net494[10], net494[11], net494[12], net494[13],
     net494[14], net494[15], net494[16], net494[17], net494[18],
     net494[19], net494[20], net494[21], net494[22], net494[23],
     net494[24], net494[25], net494[26], net494[27], net494[28],
     net494[29], net494[30], net494[31], net494[32], net494[33],
     net494[34], net494[35], net494[36], net494[37], net494[38],
     net494[39], net494[40], net494[41], net494[42], net494[43],
     net494[44], net494[45], net494[46], net494[47]}),
     .sp4_v_b_04_02({net495[0], net495[1], net495[2], net495[3],
     net495[4], net495[5], net495[6], net495[7], net495[8], net495[9],
     net495[10], net495[11], net495[12], net495[13], net495[14],
     net495[15], net495[16], net495[17], net495[18], net495[19],
     net495[20], net495[21], net495[22], net495[23], net495[24],
     net495[25], net495[26], net495[27], net495[28], net495[29],
     net495[30], net495[31], net495[32], net495[33], net495[34],
     net495[35], net495[36], net495[37], net495[38], net495[39],
     net495[40], net495[41], net495[42], net495[43], net495[44],
     net495[45], net495[46], net495[47]}), .sp4_v_b_04_01({net485[0],
     net485[1], net485[2], net485[3], net485[4], net485[5], net485[6],
     net485[7], net485[8], net485[9], net485[10], net485[11],
     net485[12], net485[13], net485[14], net485[15], net485[16],
     net485[17], net485[18], net485[19], net485[20], net485[21],
     net485[22], net485[23], net485[24], net485[25], net485[26],
     net485[27], net485[28], net485[29], net485[30], net485[31],
     net485[32], net485[33], net485[34], net485[35], net485[36],
     net485[37], net485[38], net485[39], net485[40], net485[41],
     net485[42], net485[43], net485[44], net485[45], net485[46],
     net485[47]}), .sp12_h_l_04_04({net496[0], net496[1], net496[2],
     net496[3], net496[4], net496[5], net496[6], net496[7], net496[8],
     net496[9], net496[10], net496[11], net496[12], net496[13],
     net496[14], net496[15], net496[16], net496[17], net496[18],
     net496[19], net496[20], net496[21], net496[22], net496[23]}),
     .sp4_h_l_04_01({net499[0], net499[1], net499[2], net499[3],
     net499[4], net499[5], net499[6], net499[7], net499[8], net499[9],
     net499[10], net499[11], net499[12], net499[13], net499[14],
     net499[15], net499[16], net499[17], net499[18], net499[19],
     net499[20], net499[21], net499[22], net499[23], net499[24],
     net499[25], net499[26], net499[27], net499[28], net499[29],
     net499[30], net499[31], net499[32], net499[33], net499[34],
     net499[35], net499[36], net499[37], net499[38], net499[39],
     net499[40], net499[41], net499[42], net499[43], net499[44],
     net499[45], net499[46], net499[47]}), .sp4_h_l_04_03({net497[0],
     net497[1], net497[2], net497[3], net497[4], net497[5], net497[6],
     net497[7], net497[8], net497[9], net497[10], net497[11],
     net497[12], net497[13], net497[14], net497[15], net497[16],
     net497[17], net497[18], net497[19], net497[20], net497[21],
     net497[22], net497[23], net497[24], net497[25], net497[26],
     net497[27], net497[28], net497[29], net497[30], net497[31],
     net497[32], net497[33], net497[34], net497[35], net497[36],
     net497[37], net497[38], net497[39], net497[40], net497[41],
     net497[42], net497[43], net497[44], net497[45], net497[46],
     net497[47]}), .sp4_h_l_04_02({net498[0], net498[1], net498[2],
     net498[3], net498[4], net498[5], net498[6], net498[7], net498[8],
     net498[9], net498[10], net498[11], net498[12], net498[13],
     net498[14], net498[15], net498[16], net498[17], net498[18],
     net498[19], net498[20], net498[21], net498[22], net498[23],
     net498[24], net498[25], net498[26], net498[27], net498[28],
     net498[29], net498[30], net498[31], net498[32], net498[33],
     net498[34], net498[35], net498[36], net498[37], net498[38],
     net498[39], net498[40], net498[41], net498[42], net498[43],
     net498[44], net498[45], net498[46], net498[47]}),
     .sp4_h_l_04_04({net467[0], net467[1], net467[2], net467[3],
     net467[4], net467[5], net467[6], net467[7], net467[8], net467[9],
     net467[10], net467[11], net467[12], net467[13], net467[14],
     net467[15], net467[16], net467[17], net467[18], net467[19],
     net467[20], net467[21], net467[22], net467[23], net467[24],
     net467[25], net467[26], net467[27], net467[28], net467[29],
     net467[30], net467[31], net467[32], net467[33], net467[34],
     net467[35], net467[36], net467[37], net467[38], net467[39],
     net467[40], net467[41], net467[42], net467[43], net467[44],
     net467[45], net467[46], net467[47]}), .tnl_op_04_04({net454[0],
     net454[1], net454[2], net454[3], net454[4], net454[5], net454[6],
     net454[7]}), .vdd_cntl_r(vdd_cntl_r[79:0]),
     .reset_b_r(reset_b_r[79:0]), .lft_op_04_02({net469[0], net469[1],
     net469[2], net469[3], net469[4], net469[5], net469[6],
     net469[7]}), .bnl_op_04_01({net470[0], net470[1], net470[2],
     net470[3]}), .lft_op_04_04({net471[0], net471[1], net471[2],
     net471[3], net471[4], net471[5], net471[6], net471[7]}),
     .op_vic_04_04(op_vic_04), .lft_op_04_03({net468[0], net468[1],
     net468[2], net468[3], net468[4], net468[5], net468[6],
     net468[7]}), .bl(bl_bot[363:184]), .wl_r(wl_r[79:0]),
     .glb_in_7({net579[0], net579[1], net579[2], net579[3], net579[4],
     net579[5], net579[6], net579[7]}), .glb_in_6({net580[0],
     net580[1], net580[2], net580[3], net580[4], net580[5], net580[6],
     net580[7]}), .glb_in_5({net713[0], net713[1], net713[2],
     net713[3], net713[4], net713[5], net713[6], net713[7]}),
     .glb_in_4({net430[0], net430[1], net430[2], net430[3], net430[4],
     net430[5], net430[6], net430[7]}), .padin_b_r(padin_b[11:6]),
     .cf_b_r(cf_b[143:72]), .padin_r(padin_r[7:0]),
     .padeb_r(padeb_r[7:0]), .lft_op_04_01({net484[0], net484[1],
     net484[2], net484[3], net484[4], net484[5], net484[6],
     net484[7]}), .sp4_v_t_04_04({net588[0], net588[1], net588[2],
     net588[3], net588[4], net588[5], net588[6], net588[7], net588[8],
     net588[9], net588[10], net588[11], net588[12], net588[13],
     net588[14], net588[15], net588[16], net588[17], net588[18],
     net588[19], net588[20], net588[21], net588[22], net588[23],
     net588[24], net588[25], net588[26], net588[27], net588[28],
     net588[29], net588[30], net588[31], net588[32], net588[33],
     net588[34], net588[35], net588[36], net588[37], net588[38],
     net588[39], net588[40], net588[41], net588[42], net588[43],
     net588[44], net588[45], net588[46], net588[47]}),
     .top_op_04_04({net589[0], net589[1], net589[2], net589[3],
     net589[4], net589[5], net589[6], net589[7]}),
     .top_op_05_04({net598[0], net598[1], net598[2], net598[3],
     net598[4], net598[5], net598[6], net598[7]}),
     .top_op_06_04({net599[0], net599[1], net599[2], net599[3],
     net599[4], net599[5], net599[6], net599[7]}),
     .carry_out_04_04(net592), .carry_out_05_04(net593),
     .carry_out_06_04(net594), .sp12_v_t_04_04({net595[0], net595[1],
     net595[2], net595[3], net595[4], net595[5], net595[6], net595[7],
     net595[8], net595[9], net595[10], net595[11], net595[12],
     net595[13], net595[14], net595[15], net595[16], net595[17],
     net595[18], net595[19], net595[20], net595[21], net595[22],
     net595[23]}), .sp12_v_t_05_04({net596[0], net596[1], net596[2],
     net596[3], net596[4], net596[5], net596[6], net596[7], net596[8],
     net596[9], net596[10], net596[11], net596[12], net596[13],
     net596[14], net596[15], net596[16], net596[17], net596[18],
     net596[19], net596[20], net596[21], net596[22], net596[23]}),
     .sp12_v_t_06_04({net597[0], net597[1], net597[2], net597[3],
     net597[4], net597[5], net597[6], net597[7], net597[8], net597[9],
     net597[10], net597[11], net597[12], net597[13], net597[14],
     net597[15], net597[16], net597[17], net597[18], net597[19],
     net597[20], net597[21], net597[22], net597[23]}),
     .tnr_op_04_04({net598[0], net598[1], net598[2], net598[3],
     net598[4], net598[5], net598[6], net598[7]}),
     .tnr_op_05_04({net599[0], net599[1], net599[2], net599[3],
     net599[4], net599[5], net599[6], net599[7]}),
     .tnr_op_06_04({slf_op_07_05[3], slf_op_07_05[2], slf_op_07_05[1],
     slf_op_07_05[0], slf_op_07_05[3], slf_op_07_05[2],
     slf_op_07_05[1], slf_op_07_05[0]}), .sp4_v_t_05_04({net601[0],
     net601[1], net601[2], net601[3], net601[4], net601[5], net601[6],
     net601[7], net601[8], net601[9], net601[10], net601[11],
     net601[12], net601[13], net601[14], net601[15], net601[16],
     net601[17], net601[18], net601[19], net601[20], net601[21],
     net601[22], net601[23], net601[24], net601[25], net601[26],
     net601[27], net601[28], net601[29], net601[30], net601[31],
     net601[32], net601[33], net601[34], net601[35], net601[36],
     net601[37], net601[38], net601[39], net601[40], net601[41],
     net601[42], net601[43], net601[44], net601[45], net601[46],
     net601[47]}), .sp4_v_t_06_04({net602[0], net602[1], net602[2],
     net602[3], net602[4], net602[5], net602[6], net602[7], net602[8],
     net602[9], net602[10], net602[11], net602[12], net602[13],
     net602[14], net602[15], net602[16], net602[17], net602[18],
     net602[19], net602[20], net602[21], net602[22], net602[23],
     net602[24], net602[25], net602[26], net602[27], net602[28],
     net602[29], net602[30], net602[31], net602[32], net602[33],
     net602[34], net602[35], net602[36], net602[37], net602[38],
     net602[39], net602[40], net602[41], net602[42], net602[43],
     net602[44], net602[45], net602[46], net602[47]}),
     .sp4_v_t_07_04({net603[0], net603[1], net603[2], net603[3],
     net603[4], net603[5], net603[6], net603[7], net603[8], net603[9],
     net603[10], net603[11], net603[12], net603[13], net603[14],
     net603[15]}), .tnl_op_07_04({net599[0], net599[1], net599[2],
     net599[3], net599[4], net599[5], net599[6], net599[7]}),
     .tnl_op_05_04({net589[0], net589[1], net589[2], net589[3],
     net589[4], net589[5], net589[6], net589[7]}),
     .tnl_op_06_04({net598[0], net598[1], net598[2], net598[3],
     net598[4], net598[5], net598[6], net598[7]}),
     .slf_op_05_04({net607[0], net607[1], net607[2], net607[3],
     net607[4], net607[5], net607[6], net607[7]}),
     .slf_op_06_04({net608[0], net608[1], net608[2], net608[3],
     net608[4], net608[5], net608[6], net608[7]}),
     .sp4_h_l_04_00({net513[0], net513[1], net513[2], net513[3],
     net513[4], net513[5], net513[6], net513[7], net513[8], net513[9],
     net513[10], net513[11], net513[12], net513[13], net513[14],
     net513[15]}), .cf_r(cf_r[95:0]),
     .fabric_out_04_00(fabric_out_04_00), .padin_04_00a(padin_04_00a),
     .fabric_out_07_04(fabric_out_07_04), .trstb_pad(trstb_pad),
     .sdo_pad(sdo_pad), .update_mi(update), .update_i(net534),
     .tclk_mi(tclk), .tclk_i(tclkio_mb), .shift_mi(shift),
     .shift_i(net536), .sdi_pad(sdi_pad), .sdi(sdio_mb), .r_mi(r),
     .r_i(net538), .purst(purst), .prog(prog), .mode_mi(mode),
     .mode_i(net539), .hold_r_b(fabric_out_07_06_ricegate),
     .hold_b_r(fabric_out_02_00_bicegate), .hiz_b_mi(hiz_b),
     .hiz_b_i(net540), .ceb_mi(ceb), .ceb_i(net543), .bs_en_mi(bs_en),
     .bs_en_i(net544), .update_o(net639), .tclk_o(tclkio_mr),
     .shift_o(net641), .sdo(sdio_mr), .r_o(net643), .mode_o(net644),
     .hiz_b_o(net645), .ceb_o(net646), .bs_en_o(net647),
     .last_rsr(last_rsr[2]), .spi_clk_out(spi_clk_out),
     .spi_ss_out(spi_ss_out), .spi_ss_in_bbank(spi_ss_in_bbank[4:0]),
     .spi_sdo(spi_sdo), .spi_sdo_oe_b(spi_sdo_oe_b),
     .md_spi_b(md_spi_b), .end_of_startup(end_of_startup),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .mux_jtag_sel_b(mux_jtag_sel_b), .tms_pad(tms_pad),
     .tdi_pad(tdi_pad), .tck_pad(tck_pad), .totdopad(totdopad),
     .sdo_enable(sdo_enable));
quad_tr_ice384 i_tr_quad ( .padin_04_09a(padin_04_09a),
     .slf_op_07_05(slf_op_07_05[3:0]), .sp4_v_b_04_05({net588[0],
     net588[1], net588[2], net588[3], net588[4], net588[5], net588[6],
     net588[7], net588[8], net588[9], net588[10], net588[11],
     net588[12], net588[13], net588[14], net588[15], net588[16],
     net588[17], net588[18], net588[19], net588[20], net588[21],
     net588[22], net588[23], net588[24], net588[25], net588[26],
     net588[27], net588[28], net588[29], net588[30], net588[31],
     net588[32], net588[33], net588[34], net588[35], net588[36],
     net588[37], net588[38], net588[39], net588[40], net588[41],
     net588[42], net588[43], net588[44], net588[45], net588[46],
     net588[47]}), .fabric_out_07_05(fabric_out_07_05),
     .tnl_op_04_08({net790[0], net790[1], net790[2], net790[3]}),
     .carry_in_04_05(net592), .carry_in_06_05(net594),
     .sp4_v_b_06_05({net602[0], net602[1], net602[2], net602[3],
     net602[4], net602[5], net602[6], net602[7], net602[8], net602[9],
     net602[10], net602[11], net602[12], net602[13], net602[14],
     net602[15], net602[16], net602[17], net602[18], net602[19],
     net602[20], net602[21], net602[22], net602[23], net602[24],
     net602[25], net602[26], net602[27], net602[28], net602[29],
     net602[30], net602[31], net602[32], net602[33], net602[34],
     net602[35], net602[36], net602[37], net602[38], net602[39],
     net602[40], net602[41], net602[42], net602[43], net602[44],
     net602[45], net602[46], net602[47]}), .bnl_op_07_05({net608[0],
     net608[1], net608[2], net608[3], net608[4], net608[5], net608[6],
     net608[7]}), .bnl_op_06_05({net607[0], net607[1], net607[2],
     net607[3], net607[4], net607[5], net607[6], net607[7]}),
     .bot_op_04_05({net766[0], net766[1], net766[2], net766[3],
     net766[4], net766[5], net766[6], net766[7]}),
     .bot_op_06_05({net608[0], net608[1], net608[2], net608[3],
     net608[4], net608[5], net608[6], net608[7]}),
     .bot_op_05_05({net607[0], net607[1], net607[2], net607[3],
     net607[4], net607[5], net607[6], net607[7]}),
     .lft_op_04_06({net802[0], net802[1], net802[2], net802[3],
     net802[4], net802[5], net802[6], net802[7]}),
     .carry_in_05_05(net593), .sp4_h_r_07_05({net603[0], net603[1],
     net603[2], net603[3], net603[4], net603[5], net603[6], net603[7],
     net603[8], net603[9], net603[10], net603[11], net603[12],
     net603[13], net603[14], net603[15]}), .sp12_h_l_04_05({net812[0],
     net812[1], net812[2], net812[3], net812[4], net812[5], net812[6],
     net812[7], net812[8], net812[9], net812[10], net812[11],
     net812[12], net812[13], net812[14], net812[15], net812[16],
     net812[17], net812[18], net812[19], net812[20], net812[21],
     net812[22], net812[23]}), .sp12_h_l_04_08({net794[0], net794[1],
     net794[2], net794[3], net794[4], net794[5], net794[6], net794[7],
     net794[8], net794[9], net794[10], net794[11], net794[12],
     net794[13], net794[14], net794[15], net794[16], net794[17],
     net794[18], net794[19], net794[20], net794[21], net794[22],
     net794[23]}), .sp12_h_l_04_07({net815[0], net815[1], net815[2],
     net815[3], net815[4], net815[5], net815[6], net815[7], net815[8],
     net815[9], net815[10], net815[11], net815[12], net815[13],
     net815[14], net815[15], net815[16], net815[17], net815[18],
     net815[19], net815[20], net815[21], net815[22], net815[23]}),
     .sp12_v_b_05_05({net596[0], net596[1], net596[2], net596[3],
     net596[4], net596[5], net596[6], net596[7], net596[8], net596[9],
     net596[10], net596[11], net596[12], net596[13], net596[14],
     net596[15], net596[16], net596[17], net596[18], net596[19],
     net596[20], net596[21], net596[22], net596[23]}),
     .padin_07_05a(padin_07_05a),
     .fabric_out_05_09(fabric_out_05_09_ticegate), .wl_r(wl_r[159:80]),
     .bnr_op_04_05({net607[0], net607[1], net607[2], net607[3],
     net607[4], net607[5], net607[6], net607[7]}),
     .bnr_op_06_05({slf_op_07_04[3], slf_op_07_04[2], slf_op_07_04[1],
     slf_op_07_04[0], slf_op_07_04[3], slf_op_07_04[2],
     slf_op_07_04[1], slf_op_07_04[0]}), .bnr_op_05_05({net608[0],
     net608[1], net608[2], net608[3], net608[4], net608[5], net608[6],
     net608[7]}), .last_rsr(last_rsr[3]), .sp4_h_l_04_09({net814[0],
     net814[1], net814[2], net814[3], net814[4], net814[5], net814[6],
     net814[7], net814[8], net814[9], net814[10], net814[11],
     net814[12], net814[13], net814[14], net814[15]}),
     .sp4_v_b_04_06({net795[0], net795[1], net795[2], net795[3],
     net795[4], net795[5], net795[6], net795[7], net795[8], net795[9],
     net795[10], net795[11], net795[12], net795[13], net795[14],
     net795[15], net795[16], net795[17], net795[18], net795[19],
     net795[20], net795[21], net795[22], net795[23], net795[24],
     net795[25], net795[26], net795[27], net795[28], net795[29],
     net795[30], net795[31], net795[32], net795[33], net795[34],
     net795[35], net795[36], net795[37], net795[38], net795[39],
     net795[40], net795[41], net795[42], net795[43], net795[44],
     net795[45], net795[46], net795[47]}), .sp4_v_b_04_08({net779[0],
     net779[1], net779[2], net779[3], net779[4], net779[5], net779[6],
     net779[7], net779[8], net779[9], net779[10], net779[11],
     net779[12], net779[13], net779[14], net779[15], net779[16],
     net779[17], net779[18], net779[19], net779[20], net779[21],
     net779[22], net779[23], net779[24], net779[25], net779[26],
     net779[27], net779[28], net779[29], net779[30], net779[31],
     net779[32], net779[33], net779[34], net779[35], net779[36],
     net779[37], net779[38], net779[39], net779[40], net779[41],
     net779[42], net779[43], net779[44], net779[45], net779[46],
     net779[47]}), .sp4_v_b_04_07({net781[0], net781[1], net781[2],
     net781[3], net781[4], net781[5], net781[6], net781[7], net781[8],
     net781[9], net781[10], net781[11], net781[12], net781[13],
     net781[14], net781[15], net781[16], net781[17], net781[18],
     net781[19], net781[20], net781[21], net781[22], net781[23],
     net781[24], net781[25], net781[26], net781[27], net781[28],
     net781[29], net781[30], net781[31], net781[32], net781[33],
     net781[34], net781[35], net781[36], net781[37], net781[38],
     net781[39], net781[40], net781[41], net781[42], net781[43],
     net781[44], net781[45], net781[46], net781[47]}),
     .sp4_v_b_05_05({net601[0], net601[1], net601[2], net601[3],
     net601[4], net601[5], net601[6], net601[7], net601[8], net601[9],
     net601[10], net601[11], net601[12], net601[13], net601[14],
     net601[15], net601[16], net601[17], net601[18], net601[19],
     net601[20], net601[21], net601[22], net601[23], net601[24],
     net601[25], net601[26], net601[27], net601[28], net601[29],
     net601[30], net601[31], net601[32], net601[33], net601[34],
     net601[35], net601[36], net601[37], net601[38], net601[39],
     net601[40], net601[41], net601[42], net601[43], net601[44],
     net601[45], net601[46], net601[47]}),
     .fabric_out_07_06(fabric_out_07_06_ricegate),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .sp12_v_b_04_05({net595[0], net595[1], net595[2], net595[3],
     net595[4], net595[5], net595[6], net595[7], net595[8], net595[9],
     net595[10], net595[11], net595[12], net595[13], net595[14],
     net595[15], net595[16], net595[17], net595[18], net595[19],
     net595[20], net595[21], net595[22], net595[23]}),
     .sp12_v_b_06_05({net597[0], net597[1], net597[2], net597[3],
     net597[4], net597[5], net597[6], net597[7], net597[8], net597[9],
     net597[10], net597[11], net597[12], net597[13], net597[14],
     net597[15], net597[16], net597[17], net597[18], net597[19],
     net597[20], net597[21], net597[22], net597[23]}),
     .padin_t_r(padin_t[11:6]), .sp4_h_l_04_05({net811[0], net811[1],
     net811[2], net811[3], net811[4], net811[5], net811[6], net811[7],
     net811[8], net811[9], net811[10], net811[11], net811[12],
     net811[13], net811[14], net811[15], net811[16], net811[17],
     net811[18], net811[19], net811[20], net811[21], net811[22],
     net811[23], net811[24], net811[25], net811[26], net811[27],
     net811[28], net811[29], net811[30], net811[31], net811[32],
     net811[33], net811[34], net811[35], net811[36], net811[37],
     net811[38], net811[39], net811[40], net811[41], net811[42],
     net811[43], net811[44], net811[45], net811[46], net811[47]}),
     .bnl_op_04_05({net471[0], net471[1], net471[2], net471[3],
     net471[4], net471[5], net471[6], net471[7]}),
     .sp4_h_l_04_08({net810[0], net810[1], net810[2], net810[3],
     net810[4], net810[5], net810[6], net810[7], net810[8], net810[9],
     net810[10], net810[11], net810[12], net810[13], net810[14],
     net810[15], net810[16], net810[17], net810[18], net810[19],
     net810[20], net810[21], net810[22], net810[23], net810[24],
     net810[25], net810[26], net810[27], net810[28], net810[29],
     net810[30], net810[31], net810[32], net810[33], net810[34],
     net810[35], net810[36], net810[37], net810[38], net810[39],
     net810[40], net810[41], net810[42], net810[43], net810[44],
     net810[45], net810[46], net810[47]}), .sp4_h_l_04_07({net809[0],
     net809[1], net809[2], net809[3], net809[4], net809[5], net809[6],
     net809[7], net809[8], net809[9], net809[10], net809[11],
     net809[12], net809[13], net809[14], net809[15], net809[16],
     net809[17], net809[18], net809[19], net809[20], net809[21],
     net809[22], net809[23], net809[24], net809[25], net809[26],
     net809[27], net809[28], net809[29], net809[30], net809[31],
     net809[32], net809[33], net809[34], net809[35], net809[36],
     net809[37], net809[38], net809[39], net809[40], net809[41],
     net809[42], net809[43], net809[44], net809[45], net809[46],
     net809[47]}), .bnl_op_05_05({net766[0], net766[1], net766[2],
     net766[3], net766[4], net766[5], net766[6], net766[7]}),
     .lft_op_04_05({net454[0], net454[1], net454[2], net454[3],
     net454[4], net454[5], net454[6], net454[7]}),
     .lft_op_04_08({net764[0], net764[1], net764[2], net764[3],
     net764[4], net764[5], net764[6], net764[7]}),
     .lft_op_04_07({net801[0], net801[1], net801[2], net801[3],
     net801[4], net801[5], net801[6], net801[7]}),
     .vdd_cntl_r(vdd_cntl_r[159:80]), .bl(bl_top[363:184]),
     .glb_in_7({net579[0], net579[1], net579[2], net579[3], net579[4],
     net579[5], net579[6], net579[7]}), .glb_in_6({net580[0],
     net580[1], net580[2], net580[3], net580[4], net580[5], net580[6],
     net580[7]}), .reset_b_r(reset_b_r[159:80]), .glb_in_5({net713[0],
     net713[1], net713[2], net713[3], net713[4], net713[5], net713[6],
     net713[7]}), .glb_in_4({net430[0], net430[1], net430[2],
     net430[3], net430[4], net430[5], net430[6], net430[7]}),
     .sp4_h_l_04_06({net808[0], net808[1], net808[2], net808[3],
     net808[4], net808[5], net808[6], net808[7], net808[8], net808[9],
     net808[10], net808[11], net808[12], net808[13], net808[14],
     net808[15], net808[16], net808[17], net808[18], net808[19],
     net808[20], net808[21], net808[22], net808[23], net808[24],
     net808[25], net808[26], net808[27], net808[28], net808[29],
     net808[30], net808[31], net808[32], net808[33], net808[34],
     net808[35], net808[36], net808[37], net808[38], net808[39],
     net808[40], net808[41], net808[42], net808[43], net808[44],
     net808[45], net808[46], net808[47]}), .sp12_h_l_04_06({net813[0],
     net813[1], net813[2], net813[3], net813[4], net813[5], net813[6],
     net813[7], net813[8], net813[9], net813[10], net813[11],
     net813[12], net813[13], net813[14], net813[15], net813[16],
     net813[17], net813[18], net813[19], net813[20], net813[21],
     net813[22], net813[23]}), .lc_bot_04_05(op_vic_04),
     .cf_top_r(cf_t[143:72]), .padin_r_t(padin_r[15:8]),
     .pgate_r(pgate_r[159:80]), .cf_r(cf_r[191:96]),
     .lc_bot_06_05(op_vic_06), .lc_bot_05_05(op_vic_05),
     .pado_t_r(pado_t[11:6]), .fabric_out_04_09(fabric_out_04_09),
     .slf_op_05_05({net598[0], net598[1], net598[2], net598[3],
     net598[4], net598[5], net598[6], net598[7]}),
     .slf_op_06_05({net599[0], net599[1], net599[2], net599[3],
     net599[4], net599[5], net599[6], net599[7]}),
     .padeb_t_r(padeb_t[11:6]), .slf_op_04_09({net826[0], net826[1],
     net826[2], net826[3]}), .slf_op_04_06({net767[0], net767[1],
     net767[2], net767[3], net767[4], net767[5], net767[6],
     net767[7]}), .slf_op_04_07({net765[0], net765[1], net765[2],
     net765[3], net765[4], net765[5], net765[6], net765[7]}),
     .slf_op_04_05({net589[0], net589[1], net589[2], net589[3],
     net589[4], net589[5], net589[6], net589[7]}),
     .slf_op_04_08({net800[0], net800[1], net800[2], net800[3],
     net800[4], net800[5], net800[6], net800[7]}),
     .padeb_r_t(padeb_r[15:8]), .pado_r_t(pado_r[15:8]),
     .update_i(net639), .tclk_i(tclkio_mr), .shift_i(net641),
     .sdi(sdio_mr), .r_i(net643), .purst(purst), .prog(prog),
     .mode_i(net644), .hold_t_r(fabric_out_05_09_ticegate),
     .hold_r_t(fabric_out_07_06_ricegate), .hiz_b_i(net645),
     .ceb_i(net646), .bs_en_i(net647), .update_o(net840),
     .tclk_o(tclkio_mt), .shift_o(net842), .sdo(sdio_mt), .r_o(net844),
     .mode_o(net847), .hiz_b_o(net850), .ceb_o(net839),
     .bs_en_o(net851));
quad_tl_ice384 i_tl_quad ( .fabric_out_00_05(fabric_out_00_05),
     .padin_l_t(padin_l[15:8]), .pado_l_t(pado_l[15:8]),
     .padin_03_09b(padin_03_09b), .cf_l(cf_l[191:96]),
     .fabric_out_03_09(fabric_out_03_09), .slf_op_03_08({net764[0],
     net764[1], net764[2], net764[3], net764[4], net764[5], net764[6],
     net764[7]}), .rgt_op_03_07({net765[0], net765[1], net765[2],
     net765[3], net765[4], net765[5], net765[6], net765[7]}),
     .bnr_op_03_05({net766[0], net766[1], net766[2], net766[3],
     net766[4], net766[5], net766[6], net766[7]}),
     .rgt_op_03_06({net767[0], net767[1], net767[2], net767[3],
     net767[4], net767[5], net767[6], net767[7]}),
     .rgt_op_03_05({net589[0], net589[1], net589[2], net589[3],
     net589[4], net589[5], net589[6], net589[7]}),
     .vdd_cntl_l(vdd_cntl_l[159:80]), .sp4_v_b_00_05({net505[0],
     net505[1], net505[2], net505[3], net505[4], net505[5], net505[6],
     net505[7], net505[8], net505[9], net505[10], net505[11],
     net505[12], net505[13], net505[14], net505[15]}),
     .sp12_v_b_02_05({net503[0], net503[1], net503[2], net503[3],
     net503[4], net503[5], net503[6], net503[7], net503[8], net503[9],
     net503[10], net503[11], net503[12], net503[13], net503[14],
     net503[15], net503[16], net503[17], net503[18], net503[19],
     net503[20], net503[21], net503[22], net503[23]}),
     .sp12_v_b_03_05({net451[0], net451[1], net451[2], net451[3],
     net451[4], net451[5], net451[6], net451[7], net451[8], net451[9],
     net451[10], net451[11], net451[12], net451[13], net451[14],
     net451[15], net451[16], net451[17], net451[18], net451[19],
     net451[20], net451[21], net451[22], net451[23]}),
     .sp4_v_b_02_05({net492[0], net492[1], net492[2], net492[3],
     net492[4], net492[5], net492[6], net492[7], net492[8], net492[9],
     net492[10], net492[11], net492[12], net492[13], net492[14],
     net492[15], net492[16], net492[17], net492[18], net492[19],
     net492[20], net492[21], net492[22], net492[23], net492[24],
     net492[25], net492[26], net492[27], net492[28], net492[29],
     net492[30], net492[31], net492[32], net492[33], net492[34],
     net492[35], net492[36], net492[37], net492[38], net492[39],
     net492[40], net492[41], net492[42], net492[43], net492[44],
     net492[45], net492[46], net492[47]}), .slf_op_01_05({net466[0],
     net466[1], net466[2], net466[3], net466[4], net466[5], net466[6],
     net466[7]}), .slf_op_00_05(slf_op_01_04[3:0]),
     .sp12_v_b_01_05({net477[0], net477[1], net477[2], net477[3],
     net477[4], net477[5], net477[6], net477[7], net477[8], net477[9],
     net477[10], net477[11], net477[12], net477[13], net477[14],
     net477[15], net477[16], net477[17], net477[18], net477[19],
     net477[20], net477[21], net477[22], net477[23]}),
     .sp4_v_b_01_05({net465[0], net465[1], net465[2], net465[3],
     net465[4], net465[5], net465[6], net465[7], net465[8], net465[9],
     net465[10], net465[11], net465[12], net465[13], net465[14],
     net465[15], net465[16], net465[17], net465[18], net465[19],
     net465[20], net465[21], net465[22], net465[23], net465[24],
     net465[25], net465[26], net465[27], net465[28], net465[29],
     net465[30], net465[31], net465[32], net465[33], net465[34],
     net465[35], net465[36], net465[37], net465[38], net465[39],
     net465[40], net465[41], net465[42], net465[43], net465[44],
     net465[45], net465[46], net465[47]}), .sp4_v_b_03_05({net456[0],
     net456[1], net456[2], net456[3], net456[4], net456[5], net456[6],
     net456[7], net456[8], net456[9], net456[10], net456[11],
     net456[12], net456[13], net456[14], net456[15], net456[16],
     net456[17], net456[18], net456[19], net456[20], net456[21],
     net456[22], net456[23], net456[24], net456[25], net456[26],
     net456[27], net456[28], net456[29], net456[30], net456[31],
     net456[32], net456[33], net456[34], net456[35], net456[36],
     net456[37], net456[38], net456[39], net456[40], net456[41],
     net456[42], net456[43], net456[44], net456[45], net456[46],
     net456[47]}), .sp4_r_v_b_03_08({net779[0], net779[1], net779[2],
     net779[3], net779[4], net779[5], net779[6], net779[7], net779[8],
     net779[9], net779[10], net779[11], net779[12], net779[13],
     net779[14], net779[15], net779[16], net779[17], net779[18],
     net779[19], net779[20], net779[21], net779[22], net779[23],
     net779[24], net779[25], net779[26], net779[27], net779[28],
     net779[29], net779[30], net779[31], net779[32], net779[33],
     net779[34], net779[35], net779[36], net779[37], net779[38],
     net779[39], net779[40], net779[41], net779[42], net779[43],
     net779[44], net779[45], net779[46], net779[47]}),
     .sp4_r_v_b_03_05({net588[0], net588[1], net588[2], net588[3],
     net588[4], net588[5], net588[6], net588[7], net588[8], net588[9],
     net588[10], net588[11], net588[12], net588[13], net588[14],
     net588[15], net588[16], net588[17], net588[18], net588[19],
     net588[20], net588[21], net588[22], net588[23], net588[24],
     net588[25], net588[26], net588[27], net588[28], net588[29],
     net588[30], net588[31], net588[32], net588[33], net588[34],
     net588[35], net588[36], net588[37], net588[38], net588[39],
     net588[40], net588[41], net588[42], net588[43], net588[44],
     net588[45], net588[46], net588[47]}), .sp4_r_v_b_03_07({net781[0],
     net781[1], net781[2], net781[3], net781[4], net781[5], net781[6],
     net781[7], net781[8], net781[9], net781[10], net781[11],
     net781[12], net781[13], net781[14], net781[15], net781[16],
     net781[17], net781[18], net781[19], net781[20], net781[21],
     net781[22], net781[23], net781[24], net781[25], net781[26],
     net781[27], net781[28], net781[29], net781[30], net781[31],
     net781[32], net781[33], net781[34], net781[35], net781[36],
     net781[37], net781[38], net781[39], net781[40], net781[41],
     net781[42], net781[43], net781[44], net781[45], net781[46],
     net781[47]}), .bl(bl_top[179:0]), .bot_op_03_05({net471[0],
     net471[1], net471[2], net471[3], net471[4], net471[5], net471[6],
     net471[7]}), .bnl_op_02_05({net478[0], net478[1], net478[2],
     net478[3], net478[4], net478[5], net478[6], net478[7]}),
     .bnl_op_03_05({net472[0], net472[1], net472[2], net472[3],
     net472[4], net472[5], net472[6], net472[7]}),
     .slf_op_02_05({net455[0], net455[1], net455[2], net455[3],
     net455[4], net455[5], net455[6], net455[7]}),
     .lc_bot_01_05(op_vic_01), .bnr_op_01_05({net472[0], net472[1],
     net472[2], net472[3], net472[4], net472[5], net472[6],
     net472[7]}), .bnr_op_02_05({net471[0], net471[1], net471[2],
     net471[3], net471[4], net471[5], net471[6], net471[7]}),
     .slf_op_03_09({net790[0], net790[1], net790[2], net790[3]}),
     .bnr_op_00_05({net478[0], net478[1], net478[2], net478[3],
     net478[4], net478[5], net478[6], net478[7]}),
     .pgate_l(pgate_l[159:80]), .reset_b_l(reset_b_l[159:80]),
     .sp12_h_r_03_08({net794[0], net794[1], net794[2], net794[3],
     net794[4], net794[5], net794[6], net794[7], net794[8], net794[9],
     net794[10], net794[11], net794[12], net794[13], net794[14],
     net794[15], net794[16], net794[17], net794[18], net794[19],
     net794[20], net794[21], net794[22], net794[23]}),
     .sp4_r_v_b_03_06({net795[0], net795[1], net795[2], net795[3],
     net795[4], net795[5], net795[6], net795[7], net795[8], net795[9],
     net795[10], net795[11], net795[12], net795[13], net795[14],
     net795[15], net795[16], net795[17], net795[18], net795[19],
     net795[20], net795[21], net795[22], net795[23], net795[24],
     net795[25], net795[26], net795[27], net795[28], net795[29],
     net795[30], net795[31], net795[32], net795[33], net795[34],
     net795[35], net795[36], net795[37], net795[38], net795[39],
     net795[40], net795[41], net795[42], net795[43], net795[44],
     net795[45], net795[46], net795[47]}), .carry_in_01_05(net479),
     .carry_in_02_05(net512), .bot_op_01_05({net478[0], net478[1],
     net478[2], net478[3], net478[4], net478[5], net478[6],
     net478[7]}), .bot_op_02_05({net472[0], net472[1], net472[2],
     net472[3], net472[4], net472[5], net472[6], net472[7]}),
     .rgt_op_03_08({net800[0], net800[1], net800[2], net800[3],
     net800[4], net800[5], net800[6], net800[7]}),
     .slf_op_03_07({net801[0], net801[1], net801[2], net801[3],
     net801[4], net801[5], net801[6], net801[7]}),
     .slf_op_03_06({net802[0], net802[1], net802[2], net802[3],
     net802[4], net802[5], net802[6], net802[7]}),
     .slf_op_03_05({net454[0], net454[1], net454[2], net454[3],
     net454[4], net454[5], net454[6], net454[7]}),
     .lc_bot_02_05(op_vic_02), .lc_bot_03_05(op_vic_03),
     .carry_in_03_05(net480), .padin_00_05a(padin_00_05a),
     .sp4_h_r_03_06({net808[0], net808[1], net808[2], net808[3],
     net808[4], net808[5], net808[6], net808[7], net808[8], net808[9],
     net808[10], net808[11], net808[12], net808[13], net808[14],
     net808[15], net808[16], net808[17], net808[18], net808[19],
     net808[20], net808[21], net808[22], net808[23], net808[24],
     net808[25], net808[26], net808[27], net808[28], net808[29],
     net808[30], net808[31], net808[32], net808[33], net808[34],
     net808[35], net808[36], net808[37], net808[38], net808[39],
     net808[40], net808[41], net808[42], net808[43], net808[44],
     net808[45], net808[46], net808[47]}), .sp4_h_r_03_07({net809[0],
     net809[1], net809[2], net809[3], net809[4], net809[5], net809[6],
     net809[7], net809[8], net809[9], net809[10], net809[11],
     net809[12], net809[13], net809[14], net809[15], net809[16],
     net809[17], net809[18], net809[19], net809[20], net809[21],
     net809[22], net809[23], net809[24], net809[25], net809[26],
     net809[27], net809[28], net809[29], net809[30], net809[31],
     net809[32], net809[33], net809[34], net809[35], net809[36],
     net809[37], net809[38], net809[39], net809[40], net809[41],
     net809[42], net809[43], net809[44], net809[45], net809[46],
     net809[47]}), .sp4_h_r_03_08({net810[0], net810[1], net810[2],
     net810[3], net810[4], net810[5], net810[6], net810[7], net810[8],
     net810[9], net810[10], net810[11], net810[12], net810[13],
     net810[14], net810[15], net810[16], net810[17], net810[18],
     net810[19], net810[20], net810[21], net810[22], net810[23],
     net810[24], net810[25], net810[26], net810[27], net810[28],
     net810[29], net810[30], net810[31], net810[32], net810[33],
     net810[34], net810[35], net810[36], net810[37], net810[38],
     net810[39], net810[40], net810[41], net810[42], net810[43],
     net810[44], net810[45], net810[46], net810[47]}),
     .sp4_h_r_03_05({net811[0], net811[1], net811[2], net811[3],
     net811[4], net811[5], net811[6], net811[7], net811[8], net811[9],
     net811[10], net811[11], net811[12], net811[13], net811[14],
     net811[15], net811[16], net811[17], net811[18], net811[19],
     net811[20], net811[21], net811[22], net811[23], net811[24],
     net811[25], net811[26], net811[27], net811[28], net811[29],
     net811[30], net811[31], net811[32], net811[33], net811[34],
     net811[35], net811[36], net811[37], net811[38], net811[39],
     net811[40], net811[41], net811[42], net811[43], net811[44],
     net811[45], net811[46], net811[47]}), .sp12_h_r_03_05({net812[0],
     net812[1], net812[2], net812[3], net812[4], net812[5], net812[6],
     net812[7], net812[8], net812[9], net812[10], net812[11],
     net812[12], net812[13], net812[14], net812[15], net812[16],
     net812[17], net812[18], net812[19], net812[20], net812[21],
     net812[22], net812[23]}), .sp12_h_r_03_06({net813[0], net813[1],
     net813[2], net813[3], net813[4], net813[5], net813[6], net813[7],
     net813[8], net813[9], net813[10], net813[11], net813[12],
     net813[13], net813[14], net813[15], net813[16], net813[17],
     net813[18], net813[19], net813[20], net813[21], net813[22],
     net813[23]}), .sp4_h_r_03_09({net814[0], net814[1], net814[2],
     net814[3], net814[4], net814[5], net814[6], net814[7], net814[8],
     net814[9], net814[10], net814[11], net814[12], net814[13],
     net814[14], net814[15]}), .sp12_h_r_03_07({net815[0], net815[1],
     net815[2], net815[3], net815[4], net815[5], net815[6], net815[7],
     net815[8], net815[9], net815[10], net815[11], net815[12],
     net815[13], net815[14], net815[15], net815[16], net815[17],
     net815[18], net815[19], net815[20], net815[21], net815[22],
     net815[23]}), .cf_top_l(cf_t[71:0]), .padeb_t_l(padeb_t[5:0]),
     .pado_t_l(pado_t[5:0]), .padin_t_l(padin_t[5:0]),
     .padeb_l_t(padeb_l[15:8]), .bnl_op_01_05({slf_op_00_04[3],
     slf_op_00_04[2], slf_op_00_04[1], slf_op_00_04[0],
     slf_op_00_04[3], slf_op_00_04[2], slf_op_00_04[1],
     slf_op_00_04[0]}), .glb_in_3({net481[0], net481[1], net481[2],
     net481[3], net481[4], net481[5], net481[6], net481[7]}),
     .glb_in_2({net0504[0], net0504[1], net0504[2], net0504[3],
     net0504[4], net0504[5], net0504[6], net0504[7]}),
     .glb_in_1({net0471[0], net0471[1], net0471[2], net0471[3],
     net0471[4], net0471[5], net0471[6], net0471[7]}),
     .glb_in_0({net491[0], net491[1], net491[2], net491[3], net491[4],
     net491[5], net491[6], net491[7]}), .tnr_op_03_08({net826[0],
     net826[1], net826[2], net826[3]}), .wl_l(wl_l[159:80]),
     .mode_o(net530), .hiz_b_o(net531), .ceb_o(net532),
     .bs_en_o(net533), .tclk_o(tclkio_ml), .update_o(net521),
     .shift_o(net525), .sdo(sdio_ml), .r_o(net527),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .last_rsr(last_rsr[1]), .ceb_i(net839), .update_i(net840),
     .tclk_i(tclkio_mt), .shift_i(net842), .sdi(sdio_mt), .r_i(net844),
     .purst(purst), .prog(prog), .mode_i(net847),
     .hold_t_l(fabric_out_05_09_ticegate),
     .hold_l_t(fabric_out_00_03_licegate), .hiz_b_i(net850),
     .bs_en_i(net851));
clk_mux2to1_ice8p I_glb_ck_tree_top5432 ( .bl(bl_top[183:180]),
     .gnet(gclk[5:2]), .reset_r(reset_b_r[81:80]), .min0({padin_04_09a,
     fabric_out_07_05}), .min1({padin_04_00a, fabric_out_00_05}),
     .min2({padin_00_05a, fabric_out_03_09}), .min3({padin_07_05a,
     fabric_out_03_00}), .pgate_l(pgate_l[81:80]), .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[81:80]), .reset_l(reset_b_l[81:80]),
     .wl_l(wl_l[81:80]), .wl_r(wl_r[81:80]), .pgate_r(pgate_r[81:80]),
     .vdd_cntl_r(vdd_cntl_r[81:80]));
clk_mux2to1_ice8p I_glb_ck_tree_bot7610 ( .bl(bl_bot[183:180]),
     .gnet({gclk[7], gclk[6], gclk[1], gclk[0]}),
     .reset_r(reset_b_r[79:78]), .min0({padin_07_04b,
     fabric_out_04_00}), .min1({padin_00_04b, fabric_out_04_09}),
     .min2({padin_03_00b, fabric_out_00_04}), .min3({padin_03_09b,
     fabric_out_07_04}), .pgate_l(pgate_l[79:78]), .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[79:78]), .reset_l(reset_b_l[79:78]),
     .wl_l(wl_l[79:78]), .wl_r(wl_r[79:78]), .pgate_r(pgate_r[79:78]),
     .vdd_cntl_r(vdd_cntl_r[79:78]));

endmodule
// Library - ice384chip, Cell - chip_ice384, View - schematic
// LAST TIME SAVED: Jan 12 11:50:55 2012
// NETLIST TIME: Jan 18 18:48:21 2012
`timescale 1ns / 1ns 

module chip_ice384 ( cdone, pad_b, pad_l, pad_r, pad_t, vpp, creset_b,
     trstb );

inout  cdone, vpp;

input  creset_b, trstb;

inout [15:0]  pad_l;
inout [11:0]  pad_b;
inout [15:0]  pad_r;
inout [11:0]  pad_t;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  pado_r;

wire  [4:0]  spi_ss_in_bbank;

wire  [15:0]  padin_l;

wire  [159:0]  wl_l;

wire  [159:0]  pgate_l;

wire  [159:0]  vdd_cntl_l;

wire  [363:0]  bl_bot;

wire  [159:0]  reset_l;

wire  [15:0]  pado_l;

wire  [11:0]  padeb_t;

wire  [15:0]  padeb_r;

wire  [15:0]  padeb_l;

wire  [11:0]  pado_t;

wire  [363:0]  bl_top;

wire  [11:0]  padeb_b;

wire  [159:0]  vdd_cntl_r;

wire  [11:0]  padin_b;

wire  [159:0]  pgate_r;

wire  [15:0]  padin_r;

wire  [3:0]  last_rsr;

wire  [143:0]  cf_bank_t;

wire  [11:0]  padin_t;

wire  [159:0]  wl_r;

wire  [191:0]  cf_bank_l;

wire  [191:0]  cf_bank_r;

wire  [159:0]  reset_r;

wire  [143:0]  cf_bank_b;

wire  [11:0]  pado_b;



ring_route_ice384 Iring_route ( bs_en0, ceb, end_of_startup, gint_hz,
     gsr, hiz_b0, j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr[1], last_rsr[0], last_rsr[3],
     last_rsr[2], md_spi_b, mode0, mux_jtag_sel_b, padin_b[11:0],
     padin_l[15:0], padin_r[15:0], padin_t[11:0], pgate_l[159:0],
     pgate_r[159:0], reset_l[159:0], reset_r[159:0], sdo_enable,
     shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out, totdopad,
     trstb_pad, update0, vdd_cntl_l[159:0], vdd_cntl_r[159:0],
     wl_l[159:0], wl_r[159:0], bl_bot[363:0], bl_top[363:0], cdone,
     pad_b[11:0], pad_l[15:0], pad_r[15:0], pad_t[11:0], vpp, creset_b,
     fromsdo, {cf_bank_b[132], cf_bank_b[131], cf_bank_b[108],
     cf_bank_b[107], cf_bank_b[84], cf_bank_b[83], cf_bank_b[60],
     cf_bank_b[59], cf_bank_b[36], cf_bank_b[35], cf_bank_b[12],
     cf_bank_b[11]}, {cf_bank_l[180], cf_bank_l[179], cf_bank_l[156],
     cf_bank_l[155], cf_bank_l[132], cf_bank_l[131], cf_bank_l[108],
     cf_bank_l[107], cf_bank_l[84], cf_bank_l[83], cf_bank_l[60],
     cf_bank_l[59], cf_bank_l[36], cf_bank_l[35], cf_bank_l[12],
     cf_bank_l[11]}, {cf_bank_r[180], cf_bank_r[179], cf_bank_r[156],
     cf_bank_r[155], cf_bank_r[132], cf_bank_r[131], cf_bank_r[108],
     cf_bank_r[107], cf_bank_r[84], cf_bank_r[83], cf_bank_r[60],
     cf_bank_r[59], cf_bank_r[36], cf_bank_r[35], cf_bank_r[12],
     cf_bank_r[11]}, {cf_bank_t[132], cf_bank_t[131], cf_bank_t[108],
     cf_bank_t[107], cf_bank_t[84], cf_bank_t[83], cf_bank_t[60],
     cf_bank_t[59], cf_bank_t[36], cf_bank_t[35], cf_bank_t[12],
     cf_bank_t[11]}, {cf_bank_l[181], cf_bank_l[157], cf_bank_l[133],
     cf_bank_l[109], cf_bank_l[85], cf_bank_l[61], cf_bank_l[37],
     cf_bank_l[13]}, padeb_b[11:0], padeb_l[15:0], padeb_r[15:0],
     padeb_t[11:0], pado_b[11:0], pado_l[15:0], pado_r[15:0],
     pado_t[11:0], {cf_bank_b[130], cf_bank_b[120], cf_bank_b[106],
     cf_bank_b[96], cf_bank_b[82], cf_bank_b[72], cf_bank_b[58],
     cf_bank_b[48], cf_bank_b[34], cf_bank_b[24], cf_bank_b[10],
     cf_bank_b[0]}, {cf_bank_l[178], cf_bank_l[168], cf_bank_l[154],
     cf_bank_l[144], cf_bank_l[130], cf_bank_l[120], cf_bank_l[106],
     cf_bank_l[96], cf_bank_l[82], cf_bank_l[72], cf_bank_l[58],
     cf_bank_l[48], cf_bank_l[34], cf_bank_l[24], cf_bank_l[10],
     cf_bank_l[0]}, {cf_bank_r[38], cf_bank_r[178], cf_bank_r[168],
     cf_bank_r[154], cf_bank_r[144], cf_bank_r[130], cf_bank_r[120],
     cf_bank_r[106], cf_bank_r[96], cf_bank_r[82], cf_bank_r[72],
     cf_bank_r[58], cf_bank_r[48], cf_bank_r[34], cf_bank_r[24],
     cf_bank_r[10], cf_bank_r[0]}, {cf_bank_t[130], cf_bank_t[120],
     cf_bank_t[106], cf_bank_t[96], cf_bank_t[82], cf_bank_t[72],
     cf_bank_t[58], cf_bank_t[48], cf_bank_t[34], cf_bank_t[24],
     cf_bank_t[10], cf_bank_t[0]}, spi_ss_in_bbank[4:0], tck_pad,
     tdi_pad, tms_pad, trstb);
quad_x4_ice384 quad_x4_ice384 ( cf_bank_b[143:0], cf_bank_l[191:0],
     cf_bank_r[191:0], cf_bank_t[143:0], padeb_b[11:0], padeb_l[15:0],
     padeb_r[15:0], padeb_t[11:0], pado_b[11:0], pado_l[15:0],
     pado_r[15:0], pado_t[11:0], fromsdo, spi_ss_in_bbank[4:0],
     tck_pad, tdi_pad, tms_pad, bl_bot[363:0], bl_top[363:0], bs_en0,
     ceb, end_of_startup, hiz_b0, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr[0], last_rsr[1], last_rsr[2],
     last_rsr[3], md_spi_b, mode0, mux_jtag_sel_b, padin_b[11:0],
     padin_l[15:0], padin_r[15:0], padin_t[11:0], pgate_l[159:0],
     pgate_r[159:0], gint_hz, gsr, gsr, reset_l[159:0], reset_r[159:0],
     j_tdi, sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, j_tck, totdopad, trstb_pad, update0,
     vdd_cntl_l[159:0], vdd_cntl_r[159:0], wl_l[159:0], wl_r[159:0]);

endmodule
// Library - sbtlibn65lp, Cell - vdd_tielow, View - schematic
// LAST TIME SAVED: Aug  3 19:21:57 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module vdd_tielow ( gnd_tiel );
inout  gnd_tiel;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M3 ( .D(net9), .B(vdd_), .G(net9), .S(vdd_));
N_11_LPHVT  M2 ( .D(gnd_tiel), .B(GND_), .G(net9), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_gwlgnd_nor2, View - schematic
// LAST TIME SAVED: Aug  3 19:29:08 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_rock_gwlgnd_nor2 ( gwl_gnd_25, gwl_b_sup_25, gwl_b_25,
     gwl_b_gnden_25 );
output  gwl_gnd_25;

inout  gwl_b_sup_25;

input  gwl_b_25, gwl_b_gnden_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M2 ( .D(gwl_gnd_25), .B(gwl_b_sup_25), .G(gwl_b_25),
     .S(gwl_b_sup_25));
N_25_LP  M5 ( .D(net14), .B(GND_), .G(gwl_b_gnden_25), .S(GND_));
N_25_LP  M0 ( .D(gwl_gnd_25), .B(GND_), .G(gwl_b_25), .S(net14));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp, View - schematic
// LAST TIME SAVED: Aug  3 19:29:09 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp ( wp, gwl_gnd_rp_25, ngate_25, gwl_b_25,
     gwl_gnd_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv );
output  wp;

inout  gwl_gnd_rp_25, ngate_25;

input  gwl_b_25, gwl_gnd_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M6 ( .D(wp), .B(gwp_hv), .G(s_b_hv), .S(gwp_hv));
P_25_LP  M0 ( .D(gwl_gnd_rp_25), .B(gwp_hv), .G(s_rd_b_hv), .S(wp));
N_25_LP  M11 ( .D(net18), .B(GND_), .G(s_b_25), .S(gwl_gnd_25));
N_25_LP  M12 ( .D(wp), .B(GND_), .G(ngate_25), .S(net18));
N_25_LP  M10 ( .D(net18), .B(GND_), .G(gwl_b_25), .S(gwl_gnd_25));

endmodule
// Library - sbtlibn65lp, Cell - nand2_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:55 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nand2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M2 ( .D(Y), .B(Pb), .G(B), .S(P));
P_25_LP  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
N_25_LP  M0 ( .D(Y), .B(Gb), .G(A), .S(net16));
N_25_LP  M3 ( .D(net16), .B(Gb), .G(B), .S(G));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp, View - schematic
// LAST TIME SAVED: Aug  3 19:28:59 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_sa_comp ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_b_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M3 ( .D(out_ref), .B(vddp_), .G(in_ref), .S(net65));
P_25_LP  M4_1_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
P_25_LP  M4_0_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
P_25_LP  M6 ( .D(out_div), .B(vddp_), .G(in_div), .S(net65));
N_25_LP  M2 ( .D(out_div), .B(GND_), .G(out_ref), .S(gnd_));
N_25_LP  M8 ( .D(out_ref), .B(GND_), .G(saen_b_25), .S(gnd_));
N_25_LP  M1 ( .D(out_ref), .B(GND_), .G(out_ref), .S(gnd_));
N_25_LP  M5 ( .D(out_div), .B(GND_), .G(saen_b_25), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_top, View - schematic
// LAST TIME SAVED: Nov 16 16:08:22 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_sa_comp_top ( sa_out, vdd_tieh, in_div, in_ref, saen_25
     );
output  sa_out;

inout  vdd_tieh;

input  in_div, in_ref, saen_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M43 ( .D(sa_bias), .B(vddp_), .G(saen_25), .S(vddp_));
P_25_LP  M4_1_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
P_25_LP  M4_0_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
P_25_LP  M7 ( .D(sa_out_b_25), .B(vddp_), .G(out_div2), .S(net089));
P_25_LP  M3 ( .D(net089), .B(vddp_), .G(sa_bias), .S(vddp_));
RNPPO_LP_pcell2460 R1 ( .B(gnd_), .MINUS(net053), .PLUS(net039));
RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(net039), .PLUS(net45));
N_25_LP  M6 ( .D(sa_out_b_25), .B(gnd_), .G(saen_b_25), .S(gnd_));
N_25_LP  M0 ( .D(net053), .B(gnd_), .G(saen_25), .S(gnd_));
N_25_LP  M5 ( .D(sa_out_b_25), .B(gnd_), .G(out_div2), .S(gnd_));
N_25_LP  M1 ( .D(sa_bias), .B(gnd_), .G(vdd_tieh), .S(net45));
nand2_25 I80 ( .G(gnd_), .Pb(vdd_), .A(net051), .Y(net038), .P(vdd_),
     .B(saen_25), .Gb(gnd_));
inv_25 I89 ( .IN(sa_out_b_25), .OUT(net051), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I91 ( .IN(saen_25), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net038), .OUT(sa_out), .P(vdd_), .Pb(vdd_), .G(gnd_),
     .Gb(gnd_));
ml_core_sa_comp Icore_sa_comp0 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp Icore_sa_comp1 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref2), .in_div(in_div2),
     .out_ref(out_ref), .out_div(out_div2));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa, View - schematic
// LAST TIME SAVED: Sep 24 16:16:00 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_sa ( nv_dataout, blsa, vdd_tieh, vddp_tieh, vpxa,
     dec_ok, dec_trim, fsm_rst_b, fsm_sample, fsm_tm_ref,
     fsm_tm_testdec, sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, tm_testdec_wr );
output  nv_dataout;

inout  blsa, vdd_tieh, vddp_tieh, vpxa;

input  dec_ok, fsm_rst_b, fsm_sample, fsm_tm_testdec, saen_25,
     saen_b_vpxa, saprd_b_vpxa, testdec_en_b, tm_testdec_wr;

input [1:0]  fsm_tm_ref;
input [4:1]  sa_ngate;
input [7:5]  dec_trim;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  ref;



N_25_LP  M22 ( .D(net167), .B(GND_), .G(vddp_tieh), .S(net228));
N_11_LPHVT  M23 ( .D(net220), .B(GND_), .G(dec_trim[7]), .S(gnd_));
N_11_LPHVT  M31 ( .D(gnd_), .B(GND_), .G(net226), .S(net0131));
N_11_LPHVT  M16 ( .D(net175), .B(GND_), .G(net226), .S(gnd_));
N_11_LPHVT  M13 ( .D(net228), .B(GND_), .G(vdd_tieh), .S(net240));
N_11_LPHVT  M18 ( .D(net151), .B(GND_), .G(vdd_tieh), .S(net142));
N_11_LPHVT  M25 ( .D(gnd_), .B(GND_), .G(sa_ngate[2]), .S(net0117));
N_11_LPHVT  M29 ( .D(gnd_), .B(GND_), .G(dec_trim[6]), .S(net0160));
N_11_LPHVT  M24 ( .D(gnd_), .B(GND_), .G(sa_ngate[1]), .S(net0150));
N_11_LPHVT  M21 ( .D(net0137), .B(GND_), .G(dec_trim[6]), .S(gnd_));
N_11_LPHVT  M28 ( .D(gnd_), .B(GND_), .G(dec_trim[5]), .S(net0210));
N_11_LPHVT  M19 ( .D(net236), .B(GND_), .G(vdd_tieh), .S(gnd_));
N_11_LPHVT  M26 ( .D(gnd_), .B(GND_), .G(sa_ngate[3]), .S(net0134));
N_11_LPHVT  M20 ( .D(net171), .B(GND_), .G(dec_trim[5]), .S(gnd_));
N_11_LPHVT  M30 ( .D(gnd_), .B(GND_), .G(dec_trim[7]), .S(gnd_));
N_11_LPHVT  M27 ( .D(gnd_), .B(GND_), .G(sa_ngate[4]), .S(net0152));
N_11_LPHVT  M12 ( .D(net240), .B(GND_), .G(vdd_tieh), .S(net151));
P_11_LPRVT  M0 ( .D(net167), .B(vdd_), .G(testdec_en_b), .S(vdd_));
RNPPO_LP_pcell2460 R6 ( .B(GND_), .MINUS(net0150), .PLUS(net0155));
RNPPO_LP_pcell2460 R9 ( .B(gnd_), .MINUS(net171), .PLUS(net175));
RNPPO_LP_pcell2460 R18 ( .B(GND_), .MINUS(net0160), .PLUS(net0210));
RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(net0137), .PLUS(net171));
RNPPO_LP_pcell2460 R1 ( .B(gnd_), .MINUS(net220), .PLUS(net0137));
RNPPO_LP_pcell2460 R16 ( .B(GND_), .MINUS(net0155), .PLUS(blsa));
RNPPO_LP_pcell2460 R11 ( .B(GND_), .MINUS(net0210), .PLUS(net0131));
RNPPO_LP_pcell2460 R7 ( .B(GND_), .MINUS(net0117), .PLUS(net0150));
RNPPO_LP_pcell2460 R10 ( .B(GND_), .MINUS(net0152), .PLUS(net0134));
RNPPO_LP_pcell2460 R17 ( .B(GND_), .MINUS(net0134), .PLUS(net0117));
RNPPO_LP_pcell2460 R19 ( .B(GND_), .MINUS(net0131), .PLUS(net0152));
RNPPO_LP_pcell2460 R13 ( .B(GND_), .MINUS(gnd_), .PLUS(net0160));
N_11_LPRVT  WR_CELL ( .D(net0159), .B(GND_), .G(testdec_b),
     .S(net167));
NCAP_25_LP  C0 ( .MINUS(GND_), .PLUS(in_ref));
ml_dff_nvcm I132 ( .R(net273), .D(net274), .CLK(fsm_sample),
     .QN(net276), .Q(nv_dataout));
ml_core_sa_resref_40nm Irref_bot ( .bl_in(net142), .bl_out(net236),
     .ref(ref[3:0]));
ml_core_sa_restop_40nm Irref_top ( .bl_top(net0221), .bl_bot(net0159));
ml_core_sa_resbot_40nm Irsen_bot ( .bl_in(net0141), .bl_out(net175),
     .sa_ngate(sa_ngate[4:1]), .in_dec(net0247));
nor2_hvt I214 ( .B(high_res_b), .Y(net214), .A(fsm_tm_testdec));
nor3_hvt I102 ( .B(dec_trim[6]), .Y(high_res_b), .A(dec_trim[5]),
     .C(dec_trim[7]));
mux2_hvt I206 ( .in1(blsa), .in0(net0150), .out(in_div),
     .sel(testdec_b));
mux2_hvt I270 ( .in1(ref[1]), .in0(ref[0]), .out(net185),
     .sel(fsm_tm_ref[0]));
mux2_hvt I271 ( .in1(ref[3]), .in0(ref[2]), .out(net184),
     .sel(fsm_tm_ref[0]));
mux2_hvt I279 ( .in1(net0195), .in0(ref[2]), .out(in_ref),
     .sel(testdec_b));
mux2_hvt I234 ( .in1(dec_ok), .in0(sa_out), .out(net274),
     .sel(tm_testdec_wr));
mux2_hvt I272 ( .in1(net184), .in0(net185), .out(net0195),
     .sel(fsm_tm_ref[1]));
inv_hvt I247 ( .A(fsm_rst_b), .Y(net273));
inv_hvt I208 ( .A(fsm_tm_testdec), .Y(testdec_b));
inv_hvt I248 ( .A(net214), .Y(net226));
vdd_tielow I204 ( .gnd_tiel(gnd_tlow));
ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 ( .gwl_b_gnden_25(vddp_tieh),
     .gwl_b_sup_25(vpxa), .gwl_b_25(saen_b_vpxa),
     .gwl_gnd_25(gwl_gnd_25_ref));
ml_rock_lwldrv_wp Irock_lwldrv_wp ( .gwl_gnd_rp_25(gwl_gnd_25_ref),
     .s_rd_b_hv(saprd_b_vpxa), .gwl_gnd_25(gwl_gnd_25_ref),
     .s_b_hv(gwl_gnd_25_ref), .gwp_hv(gwl_gnd_25_ref),
     .gwl_b_25(gnd_tlow), .ngate_25(vpxa), .s_b_25(saprd_b_vpxa),
     .wp(net0221));
ml_core_sa_comp_top Icore_sa_comp_top ( .vdd_tieh(vdd_tieh),
     .saen_25(saen_25), .in_ref(in_ref), .in_div(in_div),
     .sa_out(sa_out));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_top, View - schematic
// LAST TIME SAVED: Aug  3 19:29:00 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_sa_top ( nv_dataout, bl_out, bl_pgm_glb, vdd_tieh,
     vddp_tieh, vpxa, dec_ok, dec_trim, fsm_rst_b, fsm_sample,
     fsm_tm_ref, fsm_tm_testdec, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     tm_dma, tm_testdec_wr );
output  nv_dataout;

inout  bl_out, bl_pgm_glb, vdd_tieh, vddp_tieh, vpxa;

input  dec_ok, fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, tm_dma, tm_testdec_wr;

input [1:0]  fsm_tm_ref;
input [7:5]  dec_trim;
input [4:1]  sa_ngate;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_11_LPHVT  M1 ( .D(bl_out), .B(GND_), .G(sa_bl_to_pgm_glb),
     .S(bl_pgm_glb));
N_11_LPHVT  M4 ( .D(net71), .B(GND_), .G(tm_dma), .S(gnd_));
N_11_LPHVT  M2 ( .D(bl_out), .B(GND_), .G(sa_bl_to_blsa), .S(net71));
inv_hvt I131 ( .A(net073), .Y(net048));
inv_hvt I45 ( .A(net048), .Y(nv_dataout));
ml_core_sa Iml_core_sa ( .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .vddp_tieh(vddp_tieh),
     .vdd_tieh(vdd_tieh), .sa_ngate(sa_ngate[4:1]), .dec_ok(dec_ok),
     .testdec_en_b(testdec_en_b), .tm_testdec_wr(tm_testdec_wr),
     .fsm_tm_testdec(fsm_tm_testdec), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .dec_trim(dec_trim[7:5]), .nv_dataout(net073), .vpxa(vpxa),
     .blsa(net71));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_core_40nm, View - schematic
// LAST TIME SAVED: Aug  3 19:29:04 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_hv_ls_inv_core_40nm ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M15 ( .D(net37), .B(GND_), .G(sel_b_25), .S(gnd_));
N_25_LP  M10 ( .D(out_b_hv), .B(GND_), .G(vddp_tieh), .S(net29));
N_25_LP  M14 ( .D(net29), .B(GND_), .G(sel_25), .S(gnd_));
N_25_LP  M12 ( .D(net19), .B(GND_), .G(vddp_tieh), .S(net37));
P_25_LP  M2 ( .D(out_b_hv), .B(net26), .G(sel_25), .S(net26));
P_25_LP  M5 ( .D(net19), .B(net22), .G(sel_b_25), .S(net22));
P_25_LP  M7 ( .D(net26), .B(in_hv), .G(net19), .S(in_hv));
P_25_LP  M6 ( .D(net22), .B(in_hv), .G(out_b_hv), .S(in_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_s_b_hv_sw, View - schematic
// LAST TIME SAVED: Aug  3 19:29:10 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_s_b_hv_sw ( sbout_hv, ssup_hv, sbout_gnd_25, sbout_high_25,
     vddp_tieh );
inout  sbout_hv, ssup_hv;

input  sbout_gnd_25, sbout_high_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(net46), .B(ssup_hv), .G(sbout_hv_b), .S(ssup_hv));
P_25_LP  M2 ( .D(sbout_hv), .B(net46), .G(sbout_gnd_25), .S(net46));
N_25_LP  M23 ( .D(sbout_hv), .B(GND_), .G(vddp_tieh), .S(net34));
N_25_LP  M7 ( .D(net34), .B(GND_), .G(sbout_gnd_25), .S(gnd_));
ml_hv_ls_inv_core_40nm Iml_hv_ls_inv_core_40nm ( .sel_b_25(net62),
     .sel_25(sbout_high_25), .out_b_hv(sbout_hv_b), .in_hv(ssup_hv),
     .vddp_tieh(vddp_tieh));
inv_25 I114 ( .IN(sbout_high_25), .OUT(net62), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:15 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_bls_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_wp_ctrl, View - schematic
// LAST TIME SAVED: Aug  3 19:29:14 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_wp_ctrl ( s_b_25, s_b_hv, sb25sup_25, sbhvsup_hv, vddp_tieh,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25 );
inout  sb25sup_25, sbhvsup_hv, vddp_tieh;


inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [3:0]  sb25_high_25;
input [3:0]  sb25_gnd_25;
input [3:0]  sbhv_high_25;
input [3:0]  sbhv_gnd_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_s_b_hv_sw Iml_s_b_25_sw_3_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[3]),
     .sbout_hv(s_b_25[3]), .sbout_high_25(sb25_high_25[3]));
ml_s_b_hv_sw Iml_s_b_25_sw_2_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[2]),
     .sbout_hv(s_b_25[2]), .sbout_high_25(sb25_high_25[2]));
ml_s_b_hv_sw Iml_s_b_25_sw_1_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[1]),
     .sbout_hv(s_b_25[1]), .sbout_high_25(sb25_high_25[1]));
ml_s_b_hv_sw Iml_s_b_25_sw_0_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[0]),
     .sbout_hv(s_b_25[0]), .sbout_high_25(sb25_high_25[0]));
ml_s_b_hv_sw Iml_s_b_hv_sw_3_ ( .sbout_high_25(sbhv_high_25[3]),
     .sbout_hv(s_b_hv[3]), .sbout_gnd_25(sbhv_gnd_25[3]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_2_ ( .sbout_high_25(sbhv_high_25[2]),
     .sbout_hv(s_b_hv[2]), .sbout_gnd_25(sbhv_gnd_25[2]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_1_ ( .sbout_high_25(sbhv_high_25[1]),
     .sbout_hv(s_b_hv[1]), .sbout_gnd_25(sbhv_gnd_25[1]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_0_ ( .sbout_high_25(sbhv_high_25[0]),
     .sbout_hv(s_b_hv[0]), .sbout_gnd_25(sbhv_gnd_25[0]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_top_1f, View - schematic
// LAST TIME SAVED: Aug  3 19:28:58 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_ctrl_top_1f ( gwl_b_gnden_25, nv_dataout, s_rd, yp1,
     yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25, yp_test, yp_test_25,
     yp_test_b_25, bl_out, bl_pgm_glb, s_b_25, s_b_hv, sb25sup_25,
     sbhvsup_hv, vblinhi_pgm_25, vdd_tieh, vpxa, ysup_25, dec_ok,
     fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, testdec_en_b, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );
output  gwl_b_gnden_25, nv_dataout;

inout  bl_out, bl_pgm_glb, sb25sup_25, sbhvsup_hv, vblinhi_pgm_25,
     vdd_tieh, vpxa, ysup_25;

input  dec_ok, fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [3:0]  s_rd;
output [5:0]  yp1_b_25;
output [1:0]  yp_test_b_25;
output [5:0]  yp1;
output [7:0]  yp2_b_25;
output [7:0]  yp2;
output [7:0]  yp3_b_25;
output [7:0]  yp3_25;
output [1:0]  yp_test_25;
output [1:0]  yp_test;

inout [3:0]  s_b_25;
inout [3:0]  s_b_hv;

input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
input [4:1]  sa_ngate;
input [1:0]  fsm_tm_ref;
input [3:0]  fsm_blkadd;
input [9:0]  fsm_coladd;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp3_sel;

wire  [7:5]  dec_trim;

wire  [3:0]  sb25_high_25;

wire  [5:0]  yp1_sel;

wire  [3:0]  sbhv_high_25;

wire  [3:0]  sb25_gnd_25;

wire  [7:0]  yp2_sel;

wire  [3:0]  sbhv_gnd_25;



N_11_LPHVT  M3 ( .D(net223), .B(GND_), .G(net223), .S(gnd_));
P_25_LP  M4 ( .D(vddp_tieh), .B(vddp_), .G(net223), .S(vddp_));
P_11_LPHVT  M0 ( .D(vdd_tieh), .B(vdd_), .G(net223), .S(vdd_));
ml_ymux_ctrl_1f Iml_ymux_ctrl_1f ( .yp1_b_25(yp1_b_25[5:0]),
     .yp1(yp1[5:0]), .yp1_sel(yp1_sel[5:0]), .yp2(yp2[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2_sel(yp2_sel[7:0]),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_sel(yp3_sel[7:0]), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test(yp_test[1:0]),
     .yp2_b_low_b(yp21_b_low_b), .yp1_b_low_b(yp21_b_low_b),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .yp_test_25(yp_test_25[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_core_ctrl_logic_1f Icore_ctrl_logic_1f (
     .fsm_coladd(fsm_coladd[9:0]), .yp1_sel(yp1_sel[5:0]),
     .vdd_tieh(vdd_tieh), .fsm_tm_rprd(fsm_tm_rprd), .s_rd(s_rd[3:0]),
     .tm_allbank_sel(tm_allbank_sel), .yp2_sel(yp2_sel[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_tm_allwl_l(tm_allwl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25), .tm_tcol(tm_tcol),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_allbl_l(tm_allbl_l), .fsm_pgm(fsm_pgm),
     .fsm_tm_allbl_h(tm_allbl_h), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_nvcmen(fsm_nvcmen), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_blkadd(fsm_blkadd[3:0]),
     .yp_test(yp_test[1:0]), .yp21_b_low_b(yp21_b_low_b),
     .yp3_sel(yp3_sel[7:0]), .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .sbhv_high_25(sbhv_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sb25_gnd_25(sb25_gnd_25[3:0]),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .dec_trim(dec_trim[7:5]));
inv_25 I38 ( .IN(net240), .OUT(gwl_b_gnden_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I30 ( .IN(fsm_gwlbdis_b_25), .OUT(net240), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_core_sa_top Icore_sa_top ( .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .vddp_tieh(vddp_tieh),
     .vdd_tieh(vdd_tieh), .sa_ngate(sa_ngate[4:1]), .dec_ok(dec_ok),
     .testdec_en_b(testdec_en_b), .tm_dma(tm_dma),
     .fsm_tm_testdec(fsm_tm_testdec), .tm_testdec_wr(tm_testdec_wr),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .dec_trim(dec_trim[7:5]), .nv_dataout(nv_dataout), .vpxa(vpxa),
     .bl_pgm_glb(bl_pgm_glb), .bl_out(bl_out));
ml_wp_ctrl Iml_wp_ctrl ( .vddp_tieh(vddp_tieh),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .sbhv_high_25(sbhv_high_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_gnd_25(sb25_gnd_25[3:0]), .s_b_25(s_b_25[3:0]),
     .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM_40nm, Cell - cell_1x1, View - schematic
// LAST TIME SAVED: Nov 17 16:24:23 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module cell_1x1 ( bl, wp, wr );
inout  bl;

input  wp, wr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_11_LPRVT  WR_CELL ( .D(net08), .B(gnd_), .G(wr), .S(bl));
N_11_LPRVT  WP_CELL ( .D(net011), .B(gnd_), .G(wp), .S(net08));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_1x8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:19 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_1x8 ( bl, wp, wr );

input  wp, wr;

inout [7:0]  bl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



cell_1x1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
cell_1x1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));
cell_1x1 m2 ( .wp(wp), .wr(wr), .bl(bl[2]));
cell_1x1 m3 ( .wp(wp), .wr(wr), .bl(bl[3]));
cell_1x1 m4 ( .wp(wp), .wr(wr), .bl(bl[4]));
cell_1x1 m5 ( .wp(wp), .wr(wr), .bl(bl[5]));
cell_1x1 m6 ( .wp(wp), .wr(wr), .bl(bl[6]));
cell_1x1 m7 ( .wp(wp), .wr(wr), .bl(bl[7]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_8x4, View - schematic
// LAST TIME SAVED: Jan 18 16:57:38 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_8x4 ( bl, wp, wr );


inout [7:0]  bl;

input [3:0]  wp;
input [3:0]  wr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 m0 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 m1 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 m2 ( .bl(bl[7:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_1x8 m3 ( .bl(bl[7:0]), .wr(wr[3]), .wp(wp[3]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_16x4, View - schematic
// LAST TIME SAVED: Jan 18 17:00:49 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_16x4 ( bl, wp, wr );


inout [15:0]  bl;

input [3:0]  wr;
input [3:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_8x4 m0 ( .wr(wr[3:0]), .wp(wp[3:0]), .bl(bl[7:0]));
nvcm_cell_8x4 m1 ( .wr(wr[3:0]), .wp(wp[3:0]), .bl(bl[15:8]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x1, View - schematic
// LAST TIME SAVED: Aug  3 19:29:19 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_2x1 ( bl, wp, wr );

input  wp, wr;

inout [1:0]  bl;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



cell_1x1 I11 ( .wp(wp), .wr(wr), .bl(bl[0]));
cell_1x1 I12 ( .wp(wp), .wr(wr), .bl(bl[1]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x4, View - schematic
// LAST TIME SAVED: Jan 18 17:00:42 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_2x4 ( bl, wp, wr );


inout [1:0]  bl;

input [3:0]  wr;
input [3:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m3 ( .bl(bl[1:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_2x1 m2 ( .bl(bl[1:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_336x4, View - schematic
// LAST TIME SAVED: Jan 18 17:00:53 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_336x4 ( bl, bl_dummyl, bl_dummyr, bl_test, wp, wr );


inout [327:0]  bl;
inout [5:0]  bl_dummyr;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;

input [3:0]  wr;
input [3:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_16x4 Invcm_cell_16x4_19_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[319:304]));
nvcm_cell_16x4 Invcm_cell_16x4_18_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[303:288]));
nvcm_cell_16x4 Invcm_cell_16x4_17_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[287:272]));
nvcm_cell_16x4 Invcm_cell_16x4_16_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[271:256]));
nvcm_cell_16x4 Invcm_cell_16x4_15_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[255:240]));
nvcm_cell_16x4 Invcm_cell_16x4_14_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[239:224]));
nvcm_cell_16x4 Invcm_cell_16x4_13_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[223:208]));
nvcm_cell_16x4 Invcm_cell_16x4_12_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[207:192]));
nvcm_cell_16x4 Invcm_cell_16x4_11_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[191:176]));
nvcm_cell_16x4 Invcm_cell_16x4_10_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[175:160]));
nvcm_cell_16x4 Invcm_cell_16x4_9_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[159:144]));
nvcm_cell_16x4 Invcm_cell_16x4_8_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[143:128]));
nvcm_cell_16x4 Invcm_cell_16x4_7_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[127:112]));
nvcm_cell_16x4 Invcm_cell_16x4_6_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[111:96]));
nvcm_cell_16x4 Invcm_cell_16x4_5_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[95:80]));
nvcm_cell_16x4 Invcm_cell_16x4_4_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[79:64]));
nvcm_cell_16x4 Invcm_cell_16x4_3_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[63:48]));
nvcm_cell_16x4 Invcm_cell_16x4_2_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[47:32]));
nvcm_cell_16x4 Invcm_cell_16x4_1_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[31:16]));
nvcm_cell_16x4 Invcm_cell_16x4_0_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl(bl[15:0]));
nvcm_cell_16x4 Invcm_cell_16x4_20_ ( .wp(wp[3:0]), .wr(wr[3:0]),
     .bl({bl_dummyr[5:0], bl_test[1:0], bl[327:320]}));
nvcm_cell_2x4 Invcm_cell_2x4 ( .bl(bl_dummyl[1:0]), .wr(wr[3:0]),
     .wp(wp[3:0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x2, View - schematic
// LAST TIME SAVED: Oct 24 17:12:35 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_2x2 ( bl, wp, wr );


inout [1:0]  bl;

input [1:0]  wr;
input [1:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_dummy, View - schematic
// LAST TIME SAVED: Aug  3 19:29:14 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_bls_dummy ( bl_dummyr, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, pgminhi_dmmy_b_25, vdd_tieh );
inout  vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo;

input  pgminhi_dmmy_b_25, vdd_tieh;

inout [1:0]  bl_dummyr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(bl_dummyr[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M8 ( .D(bl_dummyr[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
N_25_LP  M1 ( .D(bl_dummyr[1]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rdo));
N_25_LP  M2 ( .D(bl_dummyr[0]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rde));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_16x2, View - schematic
// LAST TIME SAVED: Oct 26 17:14:50 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_16x2 ( bl, wp, wr );


inout [15:0]  bl;

input [1:0]  wr;
input [1:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 Inst_0 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 Inst_1 ( .bl(bl[15:8]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 Inst_2 ( .bl(bl[15:8]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 Inst_3 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_336x2, View - schematic
// LAST TIME SAVED: Oct 24 17:12:38 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_336x2 ( bl, bl_dummyl, bl_dummyr, bl_test, wp, wr );


inout [327:0]  bl;
inout [1:0]  bl_test;
inout [5:0]  bl_dummyr;
inout [1:0]  bl_dummyl;

input [1:0]  wp;
input [1:0]  wr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x2 Invcm_cell_2x8 ( .wr(wr[1:0]), .wp(wp[1:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_16x2 Invcm_cell_16x2_19_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[319:304]));
nvcm_cell_16x2 Invcm_cell_16x2_18_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[303:288]));
nvcm_cell_16x2 Invcm_cell_16x2_17_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[287:272]));
nvcm_cell_16x2 Invcm_cell_16x2_16_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[271:256]));
nvcm_cell_16x2 Invcm_cell_16x2_15_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[255:240]));
nvcm_cell_16x2 Invcm_cell_16x2_14_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[239:224]));
nvcm_cell_16x2 Invcm_cell_16x2_13_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[223:208]));
nvcm_cell_16x2 Invcm_cell_16x2_12_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[207:192]));
nvcm_cell_16x2 Invcm_cell_16x2_11_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[191:176]));
nvcm_cell_16x2 Invcm_cell_16x2_10_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[175:160]));
nvcm_cell_16x2 Invcm_cell_16x2_9_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[159:144]));
nvcm_cell_16x2 Invcm_cell_16x2_8_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[143:128]));
nvcm_cell_16x2 Invcm_cell_16x2_7_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[127:112]));
nvcm_cell_16x2 Invcm_cell_16x2_6_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[111:96]));
nvcm_cell_16x2 Invcm_cell_16x2_5_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[95:80]));
nvcm_cell_16x2 Invcm_cell_16x2_4_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[79:64]));
nvcm_cell_16x2 Invcm_cell_16x2_3_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[63:48]));
nvcm_cell_16x2 Invcm_cell_16x2_2_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[47:32]));
nvcm_cell_16x2 Invcm_cell_16x2_1_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[31:16]));
nvcm_cell_16x2 Invcm_cell_16x2_0_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl(bl[15:0]));
nvcm_cell_16x2 Invcm_cell_16x8_20_ ( .wp(wp[1:0]), .wr(wr[1:0]),
     .bl({bl_dummyr[5:0], bl_test[1:0], bl[327:320]}));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:19 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_2x8 ( bl, wp, wr );


inout [1:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m7 ( .bl(bl[1:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_2x1 m6 ( .bl(bl[1:0]), .wr(wr[6]), .wp(wp[6]));
nvcm_cell_2x1 m5 ( .bl(bl[1:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_2x1 m4 ( .bl(bl[1:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_2x1 m3 ( .bl(bl[1:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_2x1 m2 ( .bl(bl[1:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_8x8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:23 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_8x8 ( bl, wp, wr );


inout [7:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 m0 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 m1 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 m2 ( .bl(bl[7:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_1x8 m3 ( .bl(bl[7:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_1x8 m7 ( .bl(bl[7:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_1x8 m4 ( .bl(bl[7:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_1x8 m5 ( .bl(bl[7:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_1x8 m6 ( .bl(bl[7:0]), .wr(wr[6]), .wp(wp[6]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_16x8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:19 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_16x8 ( bl, wp, wr );


inout [15:0]  bl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_8x8 m0 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[7:0]));
nvcm_cell_8x8 m1 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[15:8]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_336x8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:21 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_336x8 ( bl, bl_dummyl, bl_dummyr, bl_test, wp, wr );


inout [1:0]  bl_test;
inout [5:0]  bl_dummyr;
inout [327:0]  bl;
inout [1:0]  bl_dummyl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x8 Invcm_cell_2x8 ( .wp(wp[7:0]), .wr(wr[7:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_16x8 Invcm_cell_16x8_19_ ( .wp(wp[7:0]), .bl(bl[319:304]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_18_ ( .wp(wp[7:0]), .bl(bl[303:288]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_17_ ( .wp(wp[7:0]), .bl(bl[287:272]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_16_ ( .wp(wp[7:0]), .bl(bl[271:256]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_15_ ( .wp(wp[7:0]), .bl(bl[255:240]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_14_ ( .wp(wp[7:0]), .bl(bl[239:224]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_13_ ( .wp(wp[7:0]), .bl(bl[223:208]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_12_ ( .wp(wp[7:0]), .bl(bl[207:192]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_11_ ( .wp(wp[7:0]), .bl(bl[191:176]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_10_ ( .wp(wp[7:0]), .bl(bl[175:160]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_9_ ( .wp(wp[7:0]), .bl(bl[159:144]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_8_ ( .wp(wp[7:0]), .bl(bl[143:128]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_7_ ( .wp(wp[7:0]), .bl(bl[127:112]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_6_ ( .wp(wp[7:0]), .bl(bl[111:96]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_5_ ( .wp(wp[7:0]), .bl(bl[95:80]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_4_ ( .wp(wp[7:0]), .bl(bl[79:64]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_3_ ( .wp(wp[7:0]), .bl(bl[63:48]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_2_ ( .wp(wp[7:0]), .bl(bl[47:32]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_1_ ( .wp(wp[7:0]), .bl(bl[31:16]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_0_ ( .wp(wp[7:0]), .bl(bl[15:0]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_20_ ( .wp(wp[7:0]), .bl({bl_dummyr[5:0],
     bl_test[1:0], bl[327:320]}), .wr(wr[7:0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_338x24_384, View - schematic
// LAST TIME SAVED: Jan 18 18:04:07 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nvcm_cell_338x24_384 ( bl, bl_dummyl, bl_dummyr, bl_test, wp,
     wp_dummyb, wp_dummyt, wr, wr_dummyb, wr_dummyt );


inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [1:0]  bl_dummyr;
inout [327:0]  bl;

input [1:0]  wp_dummyt;
input [1:0]  wp_dummyb;
input [1:0]  wr_dummyb;
input [1:0]  wr_dummyt;
input [27:0]  wr;
input [27:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_336x4 Invcm_cell_336x4 ( .wr(wr[27:24]), .wp(wp[27:24]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x2 Invcm_cell_336x2_t ( .wr(wr_dummyt[1:0]),
     .wp(wp_dummyt[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x2 Invcm_cell_336x2_b ( .wr(wr_dummyb[1:0]),
     .wp(wp_dummyb[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_2_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[23:16]), .wp(wp[23:16]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_1_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[15:8]), .wp(wp[15:8]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_0_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[7:0]), .wp(wp[7:0]), .bl_dummyl(bl_dummyl[1:0]));

endmodule
// Library - sbtlibn65lp, Cell - vddp_tiehigh, View - schematic
// LAST TIME SAVED: Oct  4 11:04:43 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module vddp_tiehigh ( vddp_tieh );
inout  vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M9 ( .D(vddp_tieh), .B(vddp_), .G(net9), .S(vddp_));
N_25_LP  M8 ( .D(net9), .B(gnd_), .G(net9), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_rows, View - schematic
// LAST TIME SAVED: Aug  3 19:29:11 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_testdec_rows ( dec_bias, dec_det, vddp_tieh, wp, wr );
inout  dec_bias, dec_det;

input  vddp_tieh, wp, wr;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M12 ( .D(net20), .B(gnd_), .G(vddp_tieh), .S(wp));
N_11_LPRVT  M8 ( .D(dec_det), .B(GND_), .G(wr), .S(gnd_));
N_11_LPRVT  M6 ( .D(dec_det), .B(GND_), .G(net20), .S(gnd_));
N_11_LPRVT  M5 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(net20));
N_11_LPRVT  M7 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(wr));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_rowsx108_384, View -
//schematic
// LAST TIME SAVED: Jan 18 18:04:16 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_testdec_rowsx108_384 ( dec_det_buf, dec_bias, dec_det, wp, wr
     );
output  dec_det_buf;

inout  dec_bias, dec_det;


input [27:0]  wr;
input [27:0]  wp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(dec_det), .Y(net18));
inv_hvt I27 ( .A(net18), .Y(dec_det_buf));
vddp_tiehigh I25 ( .vddp_tieh(vddp_tiel));
ml_testdec_rows Itestdec_rows_27_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[27]), .wp(wp[27]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_26_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[26]), .wp(wp[26]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_25_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[25]), .wp(wp[25]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_24_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[24]), .wp(wp[24]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_23_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[23]), .wp(wp[23]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_22_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[22]), .wp(wp[22]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_21_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[21]), .wp(wp[21]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_20_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[20]), .wp(wp[20]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_19_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[19]), .wp(wp[19]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_18_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[18]), .wp(wp[18]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_17_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[17]), .wp(wp[17]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_16_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[16]), .wp(wp[16]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_15_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[15]), .wp(wp[15]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_14_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[14]), .wp(wp[14]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_13_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[13]), .wp(wp[13]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_12_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[12]), .wp(wp[12]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_11_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[11]), .wp(wp[11]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_10_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[10]), .wp(wp[10]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_9_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[9]), .wp(wp[9]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_8_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[8]), .wp(wp[8]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_7_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[7]), .wp(wp[7]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_6_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[6]), .wp(wp[6]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_5_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[5]), .wp(wp[5]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_4_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[4]), .wp(wp[4]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_3_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[3]), .wp(wp[3]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_2_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[2]), .wp(wp[2]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_1_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[1]), .wp(wp[1]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_0_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[0]), .wp(wp[0]),
     .dec_bias(dec_bias));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_yp2_8, View - schematic
// LAST TIME SAVED: Aug  3 19:29:18 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_yp2_8 ( bl, bl_out, vblinhi_rde, vblinhi_rdo, yp2,
     yp2_b_25 );
inout  bl_out, vblinhi_rde, vblinhi_rdo;


inout [7:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M13 ( .D(bl[6]), .B(GND_), .G(yp2_b_25[6]), .S(vblinhi_rde));
N_25_LP  M8 ( .D(bl[1]), .B(GND_), .G(yp2_b_25[1]), .S(vblinhi_rdo));
N_25_LP  M20 ( .D(bl[0]), .B(GND_), .G(yp2_b_25[0]), .S(vblinhi_rde));
N_25_LP  M12 ( .D(bl[5]), .B(GND_), .G(yp2_b_25[5]), .S(vblinhi_rdo));
N_25_LP  M11 ( .D(bl[4]), .B(GND_), .G(yp2_b_25[4]), .S(vblinhi_rde));
N_25_LP  M10 ( .D(bl[3]), .B(GND_), .G(yp2_b_25[3]), .S(vblinhi_rdo));
N_25_LP  M9 ( .D(bl[2]), .B(GND_), .G(yp2_b_25[2]), .S(vblinhi_rde));
N_25_LP  M14 ( .D(bl[7]), .B(GND_), .G(yp2_b_25[7]), .S(vblinhi_rdo));
N_11_LPHVT  M7 ( .D(bl[7]), .B(GND_), .G(yp2[7]), .S(bl_out));
N_11_LPHVT  M0 ( .D(bl[1]), .B(GND_), .G(yp2[1]), .S(bl_out));
N_11_LPHVT  M6 ( .D(bl[6]), .B(GND_), .G(yp2[6]), .S(bl_out));
N_11_LPHVT  M5 ( .D(bl[5]), .B(GND_), .G(yp2[5]), .S(bl_out));
N_11_LPHVT  M4 ( .D(bl[4]), .B(GND_), .G(yp2[4]), .S(bl_out));
N_11_LPHVT  M3 ( .D(bl[3]), .B(GND_), .G(yp2[3]), .S(bl_out));
N_11_LPHVT  M2 ( .D(bl[0]), .B(GND_), .G(yp2[0]), .S(bl_out));
N_11_LPHVT  M1 ( .D(bl[2]), .B(GND_), .G(yp2[2]), .S(bl_out));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp_x4, View - schematic
// LAST TIME SAVED: Aug  3 19:29:09 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x4 ( wp, gwl_b_sup_25, ngate_25, gwl_b_25,
     gwl_b_gnden_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_25, gwl_b_gnden_25, gwp_hv;

output [3:0]  wp;

input [3:0]  s_b_25;
input [3:0]  s_b_hv;
input [3:0]  s_rd_b_hv;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwl_b_25(gwl_b_25), .gwl_gnd_25(gwl_gnd_25));
ml_rock_lwldrv_wp Iml_lwldrv_1 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[1]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[1]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[1]), .wp(wp[1]));
ml_rock_lwldrv_wp Iml_lwldrv_2 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[2]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[2]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[2]), .wp(wp[2]));
ml_rock_lwldrv_wp Iml_lwldrv_3 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[3]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[3]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3]), .wp(wp[3]));
ml_rock_lwldrv_wp Iml_lwldrv_0 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[0]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[0]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp_x24, View - schematic
// LAST TIME SAVED: Jan 18 18:04:00 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x24 ( wp, gwl_b_sup_25, ngate_25, s_b_25,
     s_b_hv, gwl_b_25, gwl_b_gnden_25, gwp_hv, s_rd_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_gnden_25;

output [27:0]  wp;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [6:0]  gwp_hv;
input [6:0]  gwl_b_25;
input [3:0]  s_rd_b_hv;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_6_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[6]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[27:24]),
     .gwl_b_25(gwl_b_25[6]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_5_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[5]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[23:20]),
     .gwl_b_25(gwl_b_25[5]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_4_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[4]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[19:16]),
     .gwl_b_25(gwl_b_25[4]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_3_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[3]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[15:12]),
     .gwl_b_25(gwl_b_25[3]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_2_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[2]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[11:8]),
     .gwl_b_25(gwl_b_25[2]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_1_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[1]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[7:4]),
     .gwl_b_25(gwl_b_25[1]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_0_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[0]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[3:0]),
     .gwl_b_25(gwl_b_25[0]), .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_328x24_top_384, View - schematic
// LAST TIME SAVED: Jan 18 18:04:21 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_328x24_top_384 ( nv_dataout, s_rd, bl_pgm_glb,
     gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde,
     vblinhi_rdo, vpxa, ysup_25, fsm_blkadd, fsm_coladd,
     fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25,
     s_rd_b_hv, sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );
output  nv_dataout;

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  s_rd;

input [3:0]  fsm_blkadd;
input [3:0]  s_rd_b_hv;
input [2:0]  fsm_trim_rrefrd;
input [1:0]  fsm_rowadd;
input [27:0]  wr;
input [6:0]  gwl_b_25;
input [4:1]  sa_ngate;
input [2:0]  fsm_trim_rrefpgm;
input [6:0]  gwp_hv;
input [9:0]  fsm_coladd;
input [1:0]  fsm_tm_ref;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp3;

wire  [1:0]  yp_test_b_25;

wire  [1:0]  yp_test_25;

wire  [27:0]  wp;

wire  [7:0]  yp2;

wire  [3:0]  s_b_25;

wire  [7:0]  yp3_b_25;

wire  [1:0]  yp_test;

wire  [7:0]  yp2_b_25;

wire  [1:0]  bl_test;

wire  [5:0]  yp1_b_25;

wire  [1:0]  bl_dummyr;

wire  [327:0]  bl;

wire  [5:0]  yp1;

wire  [3:0]  s_b_hv;

wire  [1:0]  bl_dummyl;



ml_testdec_bgen Itestdec_bgen ( .dec_ok(dec_ok_l),
     .testdec_en_b(testdec_en_b), .testdec_prec_b(testdec_prec_b),
     .dec_bias(dec_bias), .dec_det(dec_det));
ml_ymux_bls_x328_1f Iml_ymux_bls_x328_1f (
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_25(yp_test_25[1:0]),
     .yp_test(yp_test[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .yp2_b_25(yp2_b_25[7:0]),
     .vblinhi_rdo(vblinhi_rdo), .bl_dummyr(bl_dummyr[1:0]),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyl(bl_dummyl[1:0]), .bl_test(bl_test[1:0]),
     .bl_out(bl_out), .bl(bl[327:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vdd_tieh(vdd_tieh),
     .yp1(yp1[5:0]), .yp2(yp2[7:0]), .yp1_b_25(yp1_b_25[5:0]));
ml_core_ctrl_top_1f Icore_ctrl_top_1f ( .yp1(yp1[5:0]),
     .yp1_b_25(yp1_b_25[5:0]), .dec_ok(dec_ok_l),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .s_rd(s_rd[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .sa_ngate(sa_ngate[4:1]), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .fsm_coladd(fsm_coladd[9:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .gwl_b_gnden_25(gwl_b_gnden_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .vdd_tieh(vdd_tieh), .tm_testdec_wr(tm_testdec_wr),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_blkadd(fsm_blkadd[3:0]), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .nv_dataout(nv_dataout), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_pgm_25(vblinhi_pgm_25),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .bl_out(bl_out),
     .yp_test(yp_test[1:0]));
nvcm_cell_338x24_384 Invcm_cell_338x24_384 ( .wp(wp[27:0]),
     .wr(wr[27:0]), .wr_dummyt({net247, net247}), .wr_dummyb({net247,
     net247}), .wp_dummyt({net247, net247}), .wp_dummyb({net247,
     net247}), .bl_test(bl_test[1:0]), .bl_dummyr(bl_dummyr[1:0]),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
ml_testdec_rowsx108_384 Iml_testdec_rowsx108_384 ( .wr(wr[27:0]),
     .wp(wp[27:0]), .dec_det_buf(dec_det_buf), .dec_bias(dec_bias),
     .dec_det(dec_det));
ml_rock_lwldrv_wp_x24 Iml_rock_lwldrv_wp_x24 ( .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .wp(wp[27:0]), .s_b_hv(s_b_hv[3:0]),
     .s_b_25(s_b_25[3:0]), .ngate_25(ngate_25),
     .gwl_b_sup_25(gwl_b_sup_25), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .gwl_b_gnden_25(gwl_b_gnden_25));
vdd_tielow I47 ( .gnd_tiel(net247));

endmodule
// Library - NVCM_40nm, Cell - ml_core_bank_0_384, View - schematic
// LAST TIME SAVED: Jan 18 17:21:42 2012
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_core_bank_0_384 ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  nv_dataout;

input [3:0]  s_rd_b_hv;
input [27:0]  wr;
input [9:0]  fsm_coladd;
input [4:1]  sa_ngate;
input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
input [1:0]  fsm_tm_ref;
input [3:0]  fsm_blkadd_b;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [6:0]  gwl_b_25;
input [6:0]  gwp_hv;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net380;

wire  [3:0]  net435;

wire  [3:0]  net433;

wire  [3:0]  net434;



ml_core_328x24_top_384 Iblk_2 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net433[0], net433[1], net433[2], net433[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[2]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_328x24_top_384 blk_1 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net434[0], net434[1], net434[2], net434[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[1]),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_tm_trow(fsm_tm_trow),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_rd(fsm_rd),
     .bl_pgm_glb(bl_pgm_glb), .fsm_rowadd(fsm_rowadd[1:0]),
     .gwl_b_sup_25(gwl_b_sup_25), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .ngate_25(ngate_25), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .saen_25(saen_25), .vblinhi_rdo(vblinhi_rdo),
     .saen_b_vpxa(saen_b_vpxa), .testdec_even_b_25(testdec_even_b_25),
     .vpxa(vpxa), .testdec_odd_b_25(testdec_odd_b_25),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ysup_25(ysup_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd[0]}), .tm_testdec_wr(tm_testdec_wr),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_328x24_top_384 Iblk_0 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net435[0], net435[1], net435[2], net435[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[0]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_328x24_top_384 Iblk_3 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net380[0], net380[1], net380[2], net380[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd[1], fsm_blkadd[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[3]),
     .fsm_coladd(fsm_coladd[9:0]));

endmodule
// Library - sbtlibn65lp, Cell - nor3_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:56 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nor3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M1 ( .D(net12), .B(Pb), .G(A), .S(P));
P_25_LP  M2 ( .D(Y), .B(Pb), .G(C), .S(net16));
P_25_LP  M0 ( .D(net16), .B(Pb), .G(B), .S(net12));
N_25_LP  M3 ( .D(Y), .B(Gb), .G(B), .S(G));
N_25_LP  M5 ( .D(Y), .B(Gb), .G(C), .S(G));
N_25_LP  M4 ( .D(Y), .B(Gb), .G(A), .S(G));

endmodule
// Library - sbtlibn65lp, Cell - nand3_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:55 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module nand3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(Y), .B(Pb), .G(B), .S(P));
P_25_LP  M2 ( .D(Y), .B(Pb), .G(C), .S(P));
P_25_LP  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
N_25_LP  M5 ( .D(net21), .B(Gb), .G(C), .S(G));
N_25_LP  M3 ( .D(Y), .B(Gb), .G(A), .S(net25));
N_25_LP  M4 ( .D(net25), .B(Gb), .G(B), .S(net21));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vddp2vpxa, View - schematic
// LAST TIME SAVED: Aug  3 19:29:06 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ls_vddp2vpxa ( out_33, out_b_33, sup, in_25, in_b_25 );
output  out_33, out_b_33;

inout  sup;

input  in_25, in_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M1 ( .D(out_b_33), .B(sup), .G(in_25), .S(net60));
P_25_LP  M2 ( .D(out_33), .B(sup), .G(in_b_25), .S(net56));
P_25_LP  M3 ( .D(net56), .B(sup), .G(out_b_33), .S(sup));
P_25_LP  M5 ( .D(net60), .B(sup), .G(out_33), .S(sup));
N_25_LP  M0 ( .D(out_33), .B(gnd_), .G(in_b_25), .S(gnd_));
N_25_LP  M7 ( .D(out_b_33), .B(gnd_), .G(in_25), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_gwhv, View - schematic
// LAST TIME SAVED: Aug  3 19:29:08 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_rock_lwldrv_gwhv ( gwp_hv, gwp_sup_hv, gwl_25, gwl_25_b,
     vddp_tieh );
output  gwp_hv;

inout  gwp_sup_hv;

input  gwl_25, gwl_25_b, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M16 ( .D(gwp_hv), .B(net067), .G(gwl_25_b), .S(net067));
P_25_LP  M5 ( .D(net054), .B(net087), .G(gwl_25), .S(net087));
P_25_LP  M8 ( .D(net087), .B(gwp_sup_hv), .G(net0129), .S(gwp_sup_hv));
P_25_LP  M9 ( .D(net091), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
P_25_LP  M7 ( .D(net0129), .B(net091), .G(gwl_25_b), .S(net091));
P_25_LP  M6 ( .D(net067), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
N_25_LP  M10 ( .D(net0129), .B(gnd_), .G(vddp_tieh), .S(net050));
N_25_LP  M12 ( .D(gwp_hv), .B(gnd_), .G(vddp_tieh), .S(net034));
N_25_LP  M11 ( .D(net034), .B(gnd_), .G(gwl_25_b), .S(gnd_));
N_25_LP  M13 ( .D(net050), .B(gnd_), .G(gwl_25_b), .S(gnd_));
N_25_LP  M14 ( .D(net054), .B(gnd_), .G(vddp_tieh), .S(net058));
N_25_LP  M15 ( .D(net058), .B(gnd_), .G(gwl_25), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_gwl_drv, View - schematic
// LAST TIME SAVED: Aug  3 19:29:00 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwl_drv ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25,
     radd_1_25, radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );
output  gwl_b_25, gwl_wr_25, gwp_hv;

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25, radd_1_25,
     radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_25 I133 ( .IN(gwl_wp_25), .OUT(gwl_wp_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I100 ( .IN(out_33), .OUT(gwl_b_25), .P(gwl_b_sup_25),
     .Pb(gwl_b_sup_25), .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(gwlb_25), .OUT(gwlb_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nor3_25 I123 ( .B(net76), .A(net68), .C(net84), .Y(dec_sel_25),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nand3_25 I44 ( .B(radd_4_25), .A(radd_5_25), .Y(net76), .C(radd_3_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I122 ( .B(radd_1_25), .A(radd_2_25), .Y(net84), .C(radd_0_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I121 ( .B(gwlgrpsel_25), .A(gwlgrpsel_25), .Y(net68),
     .C(radd_6_25), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nor2_25 I128 ( .A(wr_frcen_25), .Y(net056), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(dec_sel_25));
nor2_25 I127 ( .A(wr_dis_25), .Y(gwl_wr_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(net056));
nor2_25 I129 ( .A(dec_sel_25), .Y(net096), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_en_25));
nor2_25 I130 ( .A(net096), .Y(gwlb_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_dis_25));
nor2_25 I131 ( .A(dec_sel_25), .Y(net058), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_frcen_25));
nor2_25 I132 ( .A(net058), .Y(gwl_wp_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_dis_25));
ml_ls_vddp2vpxa I99 ( .in_25(gwlb_25), .sup(gwl_b_sup_25),
     .in_b_25(gwlb_b_25), .out_33(out_33), .out_b_33(net053));
ml_rock_lwldrv_gwhv Iml_rock_lwldrv_gwhv ( .gwp_sup_hv(gwp_sup_hv),
     .vddp_tieh(vddp_tieh), .gwp_hv(gwp_hv), .gwl_25(gwl_wp_25),
     .gwl_25_b(gwl_wp_b_25));

endmodule
// Library - NVCM_40nm, Cell - ml_gwl_drv_x5_384, View - schematic
// LAST TIME SAVED: Jan 18 18:03:17 2012
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwl_drv_x5_384 ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25,
     gnv2_b_25, gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25,
     gnv5_b_25, gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1,
     gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25, gnv2_b_25,
     gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25, gnv5_b_25,
     gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1, gwl_misc_25,
     gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

output [6:0]  gwl_b_25;
output [6:0]  gwp_hv;
output [6:0]  gwl_wr_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_gwl_drv Igwl_drv_misc_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[5]),
     .radd_0_25(vddp_tieh), .radd_1_25(vddp_tieh),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_misc_25),
     .gwp_hv(gwp_hv[5]), .gwl_wr_25(gwl_wr_25[5]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_5_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[6]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[6]),
     .gwl_wr_25(gwl_wr_25[6]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_4_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[4]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[4]),
     .gwl_wr_25(gwl_wr_25[4]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[3]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[3]),
     .gwl_wr_25(gwl_wr_25[3]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[2]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[2]),
     .gwl_wr_25(gwl_wr_25[2]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[1]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[1]),
     .gwl_wr_25(gwl_wr_25[1]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[0]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25),
     .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[0]), .gwl_wr_25(gwl_wr_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x64, View - schematic
// LAST TIME SAVED: Aug  3 19:29:15 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_bls_x64 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp2, yp2_b_25, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [63:0]  bl;

input [7:0]  yp2;
input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
input [7:0]  yp2_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  bl_med;



ml_ymux_yp2_8 Iml_ymux_yp2_x8 ( .bl(bl_med[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[0]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_2 ( .vdd_tieh(vdd_tieh), .bl(bl[23:16]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[2]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_3 ( .vdd_tieh(vdd_tieh), .bl(bl[31:24]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[3]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_6 ( .vdd_tieh(vdd_tieh), .bl(bl[55:48]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[6]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_7 ( .vdd_tieh(vdd_tieh), .bl(bl[63:56]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[7]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_5 ( .vdd_tieh(vdd_tieh), .bl(bl[47:40]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[5]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_4 ( .vdd_tieh(vdd_tieh), .bl(bl[39:32]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[4]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_1 ( .vdd_tieh(vdd_tieh), .bl(bl[15:8]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[1]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr, View - schematic
// LAST TIME SAVED: Aug  3 19:29:09 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr ( wr, gwl_wr_25, s_25, wr_sup_25 );
output  wr;

input  gwl_wr_25, s_25, wr_sup_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



nand2_25 I59 ( .A(gwl_wr_25), .Y(net27), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(s_25));
inv_25 I38 ( .IN(net27), .OUT(wr), .P(wr_sup_25), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr_x4, View - schematic
// LAST TIME SAVED: Aug  3 19:29:10 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x4 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  gwl_wr_25, wr_sup_25;

output [3:0]  wr;

input [3:0]  s_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr Iml_lwldrv_2 ( .gwl_wr_25(gwl_wr_25), .wr(wr[2]),
     .s_25(s_25[2]), .wr_sup_25(wr_sup_25));
ml_rock_lwldrv_wr Iml_lwldrv_1 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[1]), .wr(wr[1]));
ml_rock_lwldrv_wr Iml_lwldrv_3 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3]), .wr(wr[3]));
ml_rock_lwldrv_wr Iml_lwldrv_0 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[0]), .wr(wr[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr_x24_384, View -
//schematic
// LAST TIME SAVED: Jan 18 17:28:31 2012
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x24_384 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  wr_sup_25;

output [27:0]  wr;

input [3:0]  s_25;
input [6:0]  gwl_wr_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_6_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[27:24]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[6]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_5_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[23:20]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[5]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_4_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[19:16]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[4]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_3_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[15:12]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[3]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_2_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[11:8]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[2]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_1_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[7:4]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[1]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_0_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[3:0]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_384, View - schematic
// LAST TIME SAVED: Jan 18 18:03:20 2012
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_384 ( gwl_b_25, gwp_hv, wr, gwl_b_sup_25, gwp_sup_hv,
     gnv_25, gnv_b_25, gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25,
     gwl_red_25, gwlb_dis_25, gwlb_en_25, s_25, vddp_tieh, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, wr_sup_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wr_sup_25;

output [6:0]  gwp_hv;
output [6:0]  gwl_b_25;
output [27:0]  wr;

input [3:0]  s_25;
input [5:0]  gnv_25;
input [1:0]  gred_b_25;
input [5:0]  gnv_b_25;
input [1:0]  gred_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [6:0]  gwl_wr_25;



ml_gwl_drv_x5_384 Igwl_drv_x5 ( .gwp_hv(gwp_hv[6:0]),
     .gwl_wr_25(gwl_wr_25[6:0]), .gwl_b_25(gwl_b_25[6:0]),
     .gwlb_en_25(gwlb_en_25), .gwlb_dis_25(gwlb_dis_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25_1(gred_b_25[1]), .gred_b_25_0(gred_b_25[0]),
     .gred_25_1(gred_25[1]), .gred_25_0(gred_25[0]),
     .gnv5_b_25(gnv_b_25[5]), .gnv5_25(gnv_25[5]),
     .gnv4_b_25(gnv_b_25[4]), .gnv4_25(gnv_25[4]),
     .gnv3_b_25(gnv_b_25[3]), .gnv3_25(gnv_25[3]),
     .gnv2_b_25(gnv_b_25[2]), .gnv2_25(gnv_25[2]),
     .gnv1_b_25(gnv_b_25[1]), .gnv1_25(gnv_25[1]),
     .gnv0_b_25(gnv_b_25[0]), .gnv0_25(gnv_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));
ml_rock_lwldrv_wr_x24_384 Iml_rock_lwldrv_wr_x24_384 (
     .gwl_wr_25(gwl_wr_25[6:0]), .wr(wr[27:0]), .wr_sup_25(wr_sup_25),
     .s_25(s_25[3:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rdhv_inv, View - schematic
// LAST TIME SAVED: Aug  3 19:29:08 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_rdhv_inv ( s_rd_b_hv, srdsup_hv, s_rdin_hv, vddp_tieh );
output  s_rd_b_hv;

inout  srdsup_hv;

input  s_rdin_hv, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M21 ( .D(s_rd_b_hv), .B(GND_), .G(vddp_tieh), .S(net19));
N_25_LP  M29 ( .D(net19), .B(GND_), .G(rd_in_25), .S(gnd_));
P_25_LP  M3 ( .D(s_rd_b_hv), .B(net12), .G(rd_in_25), .S(net12));
P_25_LP  M0 ( .D(net12), .B(srdsup_hv), .G(s_rdin_hv), .S(srdsup_hv));
N_25_LPNVT  M1 ( .D(rd_in_25), .B(GND_), .G(vddp_tieh), .S(s_rdin_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_invx3_enhance, View - schematic
// LAST TIME SAVED: Aug  3 19:29:04 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv_invx3_enhance ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh
     );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
P_25_LP  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
N_25_LP  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
N_25_LP  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM_40nm, Cell - ml_lshv_6v_switch_enhance, View -
//schematic
// LAST TIME SAVED: Aug  3 19:29:07 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_lshv_6v_switch_enhance ( out_b_hv, out_hv, in_hv, sel_25,
     sel_b_25, vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
P_25_LP  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
P_25_LP  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
P_25_LP  M1 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
N_25_LP  M0 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
N_25_LP  M3 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));
N_25_LP  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
N_25_LP  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_hotsw_enhance, View -
//schematic
// LAST TIME SAVED: Aug  3 19:29:04 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw_enhance ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3_enhance Ihv_invx3 ( .vddp_tieh(vddp_tieh),
     .out_b_hv(out_b_hv), .sel_25(sel_25), .in_hv(in_hv),
     .sel_hv(sel_hv));
ml_lshv_6v_switch_enhance Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_hotswitch_enhance, View -
//schematic
// LAST TIME SAVED: Aug  3 19:29:03 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv_hotswitch_enhance ( hv_in_hv, hv_out_hv, selhv_25,
     vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
P_25_LP  M6 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
N_25_LP  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net042));
N_25_LP  M2 ( .D(net031), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
N_25_LP  M4 ( .D(net031), .B(GND_), .G(selhv_25), .S(net042));
inv_25 I112 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_hotswitch_enhance, View -
//schematic
// LAST TIME SAVED: Aug  3 19:29:05 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch_enhance ( hvin_a_hv, hvin_b_hv, out_hv,
     sel_hv_a_25, sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch_enhance Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x328_1f, View - schematic
// LAST TIME SAVED: Aug  3 19:29:14 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module ml_ymux_bls_x328_1f ( bl, bl_dummyl, bl_dummyr, bl_out, bl_test,
     vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh,
     pgminhi_dmmy_b_25, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test, yp_test_25, yp_test_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25;

inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;
inout [327:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp2;
input [7:0]  yp3_25;
input [7:0]  yp2_b_25;
input [1:0]  yp_test_25;
input [1:0]  yp_test;
input [1:0]  yp_test_b_25;
input [5:0]  yp1;
input [5:0]  yp1_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:5]  blx8_out;

wire  [4:0]  blx64_out;



N_25_LP  M26 ( .D(vblinhi_rdo), .B(GND_), .G(yp_test_b_25[1]),
     .S(bl_test[1]));
N_25_LP  M25 ( .D(bl_test[1]), .B(GND_), .G(yp_test_25[1]),
     .S(net228));
N_25_LP  M18 ( .D(vblinhi_rde), .B(GND_), .G(yp_test_b_25[0]),
     .S(bl_test[0]));
N_25_LP  M1 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[0]),
     .S(blx64_out[0]));
N_25_LP  M11 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[5]),
     .S(blx8_out[5]));
N_25_LP  M17 ( .D(bl_test[0]), .B(GND_), .G(yp_test_25[0]),
     .S(net244));
N_25_LP  M6 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[2]),
     .S(blx64_out[2]));
N_25_LP  M5 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[1]),
     .S(blx64_out[1]));
N_25_LP  M10 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[4]),
     .S(blx64_out[4]));
N_25_LP  M9 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[3]),
     .S(blx64_out[3]));
P_25_LP  M8 ( .D(bl_test[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
P_25_LP  M7 ( .D(bl_test[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
N_11_LPHVT  M21 ( .D(net224), .B(GND_), .G(yp_test[1]), .S(bl_out));
N_11_LPHVT  M19 ( .D(net228), .B(GND_), .G(yp_test[1]), .S(net224));
N_11_LPHVT  M23 ( .D(net232), .B(GND_), .G(yp_test[0]), .S(bl_out));
N_11_LPHVT  M28 ( .D(net236), .B(GND_), .G(yp1[5]), .S(bl_out));
N_11_LPHVT  M0 ( .D(blx64_out[2]), .B(GND_), .G(yp1[2]), .S(bl_out));
N_11_LPHVT  M22 ( .D(net244), .B(GND_), .G(yp_test[0]), .S(net232));
N_11_LPHVT  M24 ( .D(blx64_out[0]), .B(GND_), .G(yp1[0]), .S(bl_out));
N_11_LPHVT  M30 ( .D(blx8_out[5]), .B(GND_), .G(yp1[5]), .S(net236));
N_11_LPHVT  M3 ( .D(blx64_out[4]), .B(GND_), .G(yp1[4]), .S(bl_out));
N_11_LPHVT  M4 ( .D(blx64_out[3]), .B(GND_), .G(yp1[3]), .S(bl_out));
N_11_LPHVT  M2 ( .D(blx64_out[1]), .B(GND_), .G(yp1[1]), .S(bl_out));
ml_ymux_bls_x8 Iml_ymux_bls_x8 ( .bl_out(blx8_out[5]),
     .bl(bl[327:320]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_r ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyr[1:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_l ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyl[1:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_0 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[0]), .bl(bl[63:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_2 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[2]), .bl(bl[191:128]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_4 ( .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]), .bl(bl[319:256]),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .bl_out(blx64_out[4]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo));
ml_ymux_bls_x64 Iml_ymux_bls_x64_1 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[1]), .bl(bl[127:64]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_3 ( .yp2(yp2[7:0]), .bl_out(blx64_out[3]),
     .bl(bl[255:192]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .yp2_b_25(yp2_b_25[7:0]), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tiehigh, View - schematic
// LAST TIME SAVED: Aug  3 19:21:57 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module vdd_tiehigh ( vdd_tieh );
inout  vdd_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_11_LPHVT  M3 ( .D(vdd_tieh), .B(vdd_), .G(net9), .S(vdd_));
N_11_LPHVT  M2 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_logic, View - schematic
// LAST TIME SAVED: Aug  3 19:29:02 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_logic ( gnv, gred, gwl_misc, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, s, sa_trim, saen, testdec_en_b, testdec_even_b,
     testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd, fsm_coladd, fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rprd, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr );
output  gwl_misc, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, saen, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [5:0]  gnv;
output [1:0]  gred;
output [3:0]  s;
output [2:0]  sa_trim;

input [0:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefpgm;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_b;

wire  [5:0]  gnv_b;

wire  [2:0]  sa_trim_b;

wire  [1:0]  xadd_b;

wire  [1:0]  gred_b;

wire  [1:0]  xadd;

wire  [2:0]  net390;

wire  [1:0]  net386;



anor21_hvt I109_1_ ( .A(net386[0]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I109_0_ ( .A(net386[1]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
nor4_hvt I287 ( .B(fsm_nvcmen_b), .Y(net216), .D(testdec_wp),
     .A(fsm_wren_b), .C(net331));
nor4_hvt I286 ( .B(fsm_pgmvfy), .Y(net211), .D(fsm_tm_allwl_h),
     .A(fsm_pgmvfy), .C(fsm_rd));
nor4_hvt I282 ( .B(fsm_tm_allbl_l), .Y(net0258), .D(net282),
     .A(fsm_tm_allbl_l), .C(fsm_nvcmen_b));
nor4_hvt I284 ( .B(pgm_hvpulse), .Y(wrsup_2vdd), .D(fsm_nvcmen_b),
     .A(pgm_hvpulse), .C(testdec_wr));
nor4_hvt I285 ( .B(fsm_nvcmen_b), .Y(net226), .D(fsm_wpen_b),
     .A(testdec_wr), .C(fsm_tm_allwl_l));
nand2_hvt I302 ( .A(net0341), .Y(net307), .B(tm_testdec));
nand2_hvt I297 ( .A(tm_testdec_wr), .Y(testwr_wpgnd_b),
     .B(tm_testdec));
nand2_hvt I269 ( .A(net355), .Y(testdec_even_b), .B(testdec_en));
nand2_hvt I268 ( .A(testdec_en), .Y(testdec_odd_b), .B(fsm_coladd[0]));
nand2_hvt I267 ( .A(fsm_rd), .Y(net0266), .B(tm_testdec));
nand3_hvt I298 ( .Y(net282), .B(net341), .C(fsm_lshven), .A(fsm_pgm));
nand3_hvt I299 ( .Y(net0278), .B(fsm_rd), .C(fsm_ymuxdis),
     .A(tm_testdec));
nand3_hvt I293 ( .Y(net286), .B(fsm_pgm), .C(fsm_tm_allwl_h),
     .A(fsm_wren));
nand3_hvt I288 ( .Y(net274), .B(fsm_tm_allwl_h), .C(fsm_tm_allwl_h),
     .A(stress2));
nand3_hvt I292 ( .Y(net292), .B(tm_allwl_l_b), .C(net307),
     .A(fsm_nvcmen));
nand3_hvt I303 ( .Y(gwlb_dis), .B(fsm_nvcmen), .C(testwr_wpgnd_b),
     .A(net0332));
inv_hvt I307_5_ ( .A(fsm_rowadd[7]), .Y(gnv_b[5]));
inv_hvt I307_4_ ( .A(fsm_rowadd[6]), .Y(gnv_b[4]));
inv_hvt I307_3_ ( .A(fsm_rowadd[5]), .Y(gnv_b[3]));
inv_hvt I307_2_ ( .A(fsm_rowadd[4]), .Y(gnv_b[2]));
inv_hvt I307_1_ ( .A(fsm_rowadd[3]), .Y(gnv_b[1]));
inv_hvt I307_0_ ( .A(fsm_rowadd[2]), .Y(gnv_b[0]));
inv_hvt I238 ( .A(net0274), .Y(gwl_misc));
inv_hvt I234 ( .A(testdec_en), .Y(testdec_en_b));
inv_hvt I240 ( .A(gwlbsup_vddp), .Y(net202));
inv_hvt I236 ( .A(net0300), .Y(testdec_prec_b));
inv_hvt I305_1_ ( .A(gred_b[1]), .Y(gred[1]));
inv_hvt I305_0_ ( .A(gred_b[0]), .Y(gred[0]));
inv_hvt I314_2_ ( .A(sa_trim_b[2]), .Y(sa_trim[2]));
inv_hvt I314_1_ ( .A(sa_trim_b[1]), .Y(sa_trim[1]));
inv_hvt I314_0_ ( .A(sa_trim_b[0]), .Y(sa_trim[0]));
inv_hvt I315_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I315_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I306_5_ ( .A(gnv_b[5]), .Y(gnv[5]));
inv_hvt I306_4_ ( .A(gnv_b[4]), .Y(gnv[4]));
inv_hvt I306_3_ ( .A(gnv_b[3]), .Y(gnv[3]));
inv_hvt I306_2_ ( .A(gnv_b[2]), .Y(gnv[2]));
inv_hvt I306_1_ ( .A(gnv_b[1]), .Y(gnv[1]));
inv_hvt I306_0_ ( .A(gnv_b[0]), .Y(gnv[0]));
inv_hvt I261 ( .A(pgm_hvpulse), .Y(net0390));
inv_hvt I291 ( .A(net0428), .Y(net331));
inv_hvt I263 ( .A(net282), .Y(pgm_hvpulse));
inv_hvt I250 ( .A(fsm_coladd[0]), .Y(net355));
inv_hvt I255 ( .A(net307), .Y(testdec_wp));
inv_hvt I248 ( .A(net246), .Y(net359));
inv_hvt I252 ( .A(fsm_wren), .Y(fsm_wren_b));
inv_hvt I241 ( .A(gwlbsup_vpxa), .Y(net204));
inv_hvt I244 ( .A(net0278), .Y(net0300));
inv_hvt I264 ( .A(fsm_pgmvfy), .Y(net341));
inv_hvt I246_2_ ( .A(net390[0]), .Y(sa_trim_b[2]));
inv_hvt I246_1_ ( .A(net390[1]), .Y(sa_trim_b[1]));
inv_hvt I246_0_ ( .A(net390[2]), .Y(sa_trim_b[0]));
inv_hvt I254 ( .A(net292), .Y(net365));
inv_hvt I242 ( .A(gwphv_vddp), .Y(net206));
inv_hvt I249 ( .A(net0266), .Y(testdec_en));
inv_hvt I266 ( .A(net0388), .Y(net0327));
inv_hvt I243 ( .A(gwphv_vppint), .Y(net200));
inv_hvt I256 ( .A(net286), .Y(net0343));
inv_hvt I258 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I257 ( .A(tm_testdec_wr), .Y(net0341));
inv_hvt I259 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I304_1_ ( .A(fsm_rowadd[3]), .Y(gred_b[1]));
inv_hvt I304_0_ ( .A(fsm_rowadd[2]), .Y(gred_b[0]));
inv_hvt I253 ( .A(net196), .Y(net351));
inv_hvt I251 ( .A(fsm_wpen), .Y(fsm_wpen_b));
inv_hvt I262 ( .A(fsm_pgm), .Y(fsm_pgm_b));
inv_hvt I309 ( .A(net211), .Y(wp_frcen));
inv_hvt I310 ( .A(net216), .Y(wr_dis));
inv_hvt I308 ( .A(net226), .Y(wp_dis));
inv_hvt I311 ( .A(net274), .Y(wr_frcen));
inv_hvt I312 ( .A(testwr_wpgnd_b), .Y(testdec_wr));
inv_hvt I147_3_ ( .A(s_b[3]), .Y(s[3]));
inv_hvt I147_2_ ( .A(s_b[2]), .Y(s[2]));
inv_hvt I147_1_ ( .A(s_b[1]), .Y(s[1]));
inv_hvt I147_0_ ( .A(s_b[0]), .Y(s[0]));
nor2_hvt I272 ( .A(net0258), .B(tm_testdec), .Y(pgminhi_dmmy_b));
nor2_hvt I279 ( .A(fsm_pgm), .B(fsm_pgmvfy), .Y(net0388));
nor2_hvt I313 ( .A(net0288), .B(net0390), .Y(gwlb_en));
nor2_hvt I274 ( .A(net359), .B(net201), .Y(gwphv_vddp));
nor2_hvt I273 ( .A(fsm_nvcmen_b), .B(tm_dma), .Y(saen));
nor2_hvt I278 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I300 ( .A(fsm_pgmdisc), .B(fsm_pgmhv), .Y(net0231));
nor2_hvt I316 ( .A(net207), .B(net246), .Y(gwphv_vppint));
nor2_hvt I275 ( .A(net0232), .B(fsm_nvcmen_b), .Y(net246));
nor2_hvt I276 ( .A(net203), .B(net351), .Y(gwlbsup_vpxa));
nor2_hvt I296 ( .A(fsm_pgmvfy), .B(fsm_pgm_b), .Y(stress2));
nor2_hvt I277 ( .A(net196), .B(net205), .Y(gwlbsup_vddp));
nor3_hvt I290 ( .B(fsm_tm_allwl_l), .Y(net0428), .A(fsm_tm_allwl_l),
     .C(fsm_tm_allwl_l));
nor3_hvt I324 ( .B(fsm_tm_allwl_h), .Y(net0288), .A(fsm_tm_allwl_h),
     .C(fsm_tm_allwl_h));
nor3_hvt I295 ( .B(fsm_tm_trow), .Y(net0274), .A(fsm_nv_rri_trim),
     .C(fsm_nv_sisi_ui));
nor3_hvt I294 ( .B(fsm_tm_rprd), .Y(net196), .A(fsm_tm_rprd),
     .C(fsm_tm_rprd));
mux2_hvt I180_1_ ( .in1(fsm_rowadd[1]), .in0(fsm_rowadd[1]),
     .out(net386[0]), .sel(fsm_nv_rrow));
mux2_hvt I180_0_ ( .in1(fsm_rowadd[0]), .in0(fsm_rowadd[0]),
     .out(net386[1]), .sel(fsm_nv_rrow));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net390[0]), .sel(net0327));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net390[1]), .sel(net0327));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net390[2]), .sel(net0327));
mux2_hvt I221 ( .in1(fsm_wpen), .in0(fsm_wgnden), .out(net0332),
     .sel(pgm_hvpulse));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_pump_a_clkdly I230 ( .in(net0231), .out(net0232));
ml_pump_a_clkdly I208 ( .in(net200), .out(net201));
ml_pump_a_clkdly I202 ( .in(net202), .out(net203));
ml_pump_a_clkdly I198 ( .in(net204), .out(net205));
ml_pump_a_clkdly I207 ( .in(net206), .out(net207));
anor31_hvt I121_3_ ( .A(net365), .D(net0343), .B(xadd[1]), .Y(s_b[3]),
     .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net365), .D(net0343), .B(xadd[1]), .Y(s_b[2]),
     .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net365), .D(net0343), .B(xadd_b[1]),
     .Y(s_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net365), .D(net0343), .B(xadd_b[1]),
     .Y(s_b[0]), .C(xadd_b[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_invx3, View - schematic
// LAST TIME SAVED: Aug  3 19:29:04 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv_invx3 ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
P_25_LP  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
N_25_LP  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
N_25_LP  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM_40nm, Cell - ml_lshv_6v_switch, View - schematic
// LAST TIME SAVED: Aug  3 19:29:07 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_lshv_6v_switch ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
P_25_LP  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
P_25_LP  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
P_25_LP  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
N_25_LP  M3 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));
N_25_LP  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
N_25_LP  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
N_25_LP  M0 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_hotsw, View - schematic
// LAST TIME SAVED: Aug  3 19:29:04 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3 Ihv_invx3 ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));
ml_lshv_6v_switch Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_hotswitch, View - schematic
// LAST TIME SAVED: Aug  3 19:29:03 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hv_hotswitch ( hv_in_hv, hv_out_hv, selhv_25, vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LP  M4 ( .D(net15), .B(GND_), .G(selhv_25), .S(net12));
N_25_LP  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
N_25_LP  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
P_25_LP  M3 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
P_25_LP  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_hotswitch, View - schematic
// LAST TIME SAVED: Aug  3 19:29:05 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch ( hvin_a_hv, hvin_b_hv, out_hv, sel_hv_a_25,
     sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_bldrv, View - schematic
// LAST TIME SAVED: Oct 13 15:09:26 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_bldrv ( bgr, bl_pgm_glb, bl_frc_gnd, fsm_din, fsm_pgm,
     fsm_pgmien, fsm_trim_ipp, tm_dma );
inout  bgr, bl_pgm_glb;

input  bl_frc_gnd, fsm_din, fsm_pgm, fsm_pgmien, tm_dma;

input [3:0]  fsm_trim_ipp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net0115;

wire  [1:0]  net0160;

wire  [7:0]  net0152;

wire  [3:0]  net0172;

wire  [3:0]  net0156;

wire  [1:0]  net0180;



P_25_LP  M14_1_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
P_25_LP  M14_0_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
P_25_LP  M5 ( .D(net0164), .B(vddp_), .G(dec_bias_p), .S(net0241));
P_25_LP  M7_1_ ( .D(net0241), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
P_25_LP  M7_0_ ( .D(net0241), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
P_25_LP  M4 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p), .S(net0241));
P_25_LP  M11 ( .D(pgm_inhi_bias), .B(vddp_), .G(vdd_tieh),
     .S(net0259));
N_11_LPHVT  M37 ( .D(net0107), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
N_11_LPHVT  M31_7_ ( .D(net0115[0]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[0]));
N_11_LPHVT  M31_6_ ( .D(net0115[1]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[1]));
N_11_LPHVT  M31_5_ ( .D(net0115[2]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[2]));
N_11_LPHVT  M31_4_ ( .D(net0115[3]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[3]));
N_11_LPHVT  M31_3_ ( .D(net0115[4]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[4]));
N_11_LPHVT  M31_2_ ( .D(net0115[5]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[5]));
N_11_LPHVT  M31_1_ ( .D(net0115[6]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[6]));
N_11_LPHVT  M31_0_ ( .D(net0115[7]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[7]));
N_11_LPHVT  M19 ( .D(net0135), .B(GND_), .G(fsm_trim_ipp[0]),
     .S(net0131));
N_11_LPHVT  M38_7_ ( .D(net0152[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M38_6_ ( .D(net0152[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M38_5_ ( .D(net0152[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M38_4_ ( .D(net0152[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M38_3_ ( .D(net0152[4]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M38_2_ ( .D(net0152[5]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M38_1_ ( .D(net0152[6]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M38_0_ ( .D(net0152[7]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M39_3_ ( .D(net0156[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M39_2_ ( .D(net0156[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M39_1_ ( .D(net0156[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M39_0_ ( .D(net0156[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M40_1_ ( .D(net0160[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M40_0_ ( .D(net0160[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
N_11_LPHVT  M26 ( .D(net0131), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
N_11_LPHVT  M33 ( .D(bl_pgm_glb), .B(GND_), .G(net0187), .S(gnd_));
N_11_LPHVT  M30_3_ ( .D(net0172[0]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[0]));
N_11_LPHVT  M30_2_ ( .D(net0172[1]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[1]));
N_11_LPHVT  M30_1_ ( .D(net0172[2]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[2]));
N_11_LPHVT  M30_0_ ( .D(net0172[3]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[3]));
N_11_LPHVT  M36 ( .D(net0173), .B(GND_), .G(pgm_trim0_en),
     .S(net0107));
N_11_LPHVT  M34 ( .D(net089), .B(GND_), .G(pgm_trim0_en), .S(gnd_));
N_11_LPHVT  M27_1_ ( .D(net0180[0]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[0]));
N_11_LPHVT  M27_0_ ( .D(net0180[1]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[1]));
N_25_LP  M21 ( .D(pgm_inhi_bias), .B(GND_), .G(pgm_inhi_bias),
     .S(gnd_));
N_25_LP  M12_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[0]));
N_25_LP  M12_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[1]));
N_25_LP  M13_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[0]));
N_25_LP  M13_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[1]));
N_25_LP  M13_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[2]));
N_25_LP  M13_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[3]));
N_25_LP  M6 ( .D(net0164), .B(GND_), .G(net0164), .S(gnd_));
N_25_LP  M3 ( .D(dec_bias_p), .B(GND_), .G(bgr), .S(net0141));
N_25_LP  M20 ( .D(net0173), .B(GND_), .G(pgm_inhi_bias),
     .S(bl_pgm_glb));
N_25_LP  M10 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net089));
N_25_LP  M18_7_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[0]));
N_25_LP  M18_6_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[1]));
N_25_LP  M18_5_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[2]));
N_25_LP  M18_4_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[3]));
N_25_LP  M18_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[4]));
N_25_LP  M18_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[5]));
N_25_LP  M18_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[6]));
N_25_LP  M18_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[7]));
N_25_LP  M9 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net0135));
N_25_LP  M8 ( .D(net0164), .B(GND_), .G(pgmen_b_25), .S(gnd_));
RNPPO_LP_pcell2460 R1 ( .B(GND_), .MINUS(gnd_), .PLUS(gnd_));
RNPPO_LP_pcell2460 R2 ( .B(GND_), .MINUS(gnd_), .PLUS(gnd_));
RNPPO_LP_pcell2460 R0 ( .B(GND_), .MINUS(gnd_), .PLUS(net0141));
nor2_hvt I121 ( .A(net086), .B(fsm_pgmien_b_buf), .Y(pgm_trim0_en));
nor2_hvt I114 ( .B(tm_dma), .Y(net0116), .A(tm_dma));
nor4_hvt I105 ( .D(fsm_trim_ipp[0]), .B(fsm_trim_ipp[2]), .Y(net086),
     .A(fsm_trim_ipp[3]), .C(fsm_trim_ipp[1]));
nand2_hvt I71 ( .B(fsm_din), .A(fsm_pgmien), .Y(fsm_pgmien_b_buf));
inv_hvt I115 ( .A(net0116), .Y(net0187));
inv_hvt I58 ( .A(pgmen_b), .Y(pgmen));
inv_hvt I131 ( .A(fsm_pgm), .Y(pgmen_b));
inv_hvt I72 ( .A(fsm_pgmien_b_buf), .Y(fsm_pgmien_buf));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_ls_vdd2vdd25 I56 ( .in(pgmen), .sup(vddp_),
     .out_vddio_b(pgmen_b_25), .out_vddio(pgmen_25), .in_b(pgmen_b));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_wr_sup, View - schematic
// LAST TIME SAVED: Aug  3 19:29:02 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_wr_sup ( wr_sup_25, wrsup_2vdd, wrsup_2vdd_25 );
inout  wr_sup_25;

input  wrsup_2vdd, wrsup_2vdd_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



N_25_LPNVT  M13 ( .D(vdd_), .B(GND_), .G(wrsup_2vdd_25),
     .S(wr_sup_25));
P_25_LP  M5 ( .D(net17), .B(vddp_), .G(wrsup_2vdd_25), .S(vddp_));
P_25_LP  M0 ( .D(net17), .B(wr_sup_25), .G(wrsup_2vdd), .S(wr_sup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_ls25_1b, View - schematic
// LAST TIME SAVED: Aug  3 19:29:02 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25_1b ( out_25, in );
output  out_25;

input  in;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I145 ( .A(in), .Y(net45));
inv_25 I153 ( .IN(out_b_25), .OUT(out_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I112 ( .in(in), .sup(vddp_), .out_vddio_b(out_b_25),
     .out_vddio(net025), .in_b(net45));

endmodule
// Library - sbtlibn65lp, Cell - inv_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:54 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module inv_25 ( OUT, G, Gb, IN, P, Pb );
output  OUT;

input  G, Gb, IN, P, Pb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M1 ( .D(OUT), .B(Pb), .G(IN), .S(P));
N_25_LP  M0 ( .D(OUT), .B(Gb), .G(IN), .S(G));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_ls25, View - schematic
// LAST TIME SAVED: Aug  3 19:29:02 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25 ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25,
     gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25, s_25,
     testdec_even_b_25, testdec_odd_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, wrsup_2vdd_25, fsm_gwlbdis, gnv, gred,
     gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en, gwlbsup_vddp,
     gwlbsup_vpxa, gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, s,
     testdec_even_b, testdec_odd_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25,
     testdec_even_b_25, testdec_odd_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, wrsup_2vdd_25;

input  fsm_gwlbdis, gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, testdec_even_b, testdec_odd_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

output [3:0]  s_25;
output [1:0]  gred_25;
output [5:0]  gnv_b_25;
output [5:0]  gnv_25;
output [1:0]  gred_b_25;

input [5:0]  gnv;
input [3:0]  s;
input [1:0]  gred;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



inv_25 I_1_ ( .IN(gred_25[1]), .OUT(gred_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I_0_ ( .IN(gred_25[0]), .OUT(gred_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_5_ ( .IN(gnv_25[5]), .OUT(gnv_b_25[5]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_4_ ( .IN(gnv_25[4]), .OUT(gnv_b_25[4]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_3_ ( .IN(gnv_25[3]), .OUT(gnv_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_2_ ( .IN(gnv_25[2]), .OUT(gnv_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_1_ ( .IN(gnv_25[1]), .OUT(gnv_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_0_ ( .IN(gnv_25[0]), .OUT(gnv_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I143 ( .IN(net101), .OUT(fsm_gwlbdis_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_gwlwr_ctrl_ls25_1b I139 ( .in(gwlb_dis), .out_25(gwlb_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_frcen ( .in(wr_frcen),
     .out_25(wr_frcen_25));
ml_gwlwr_ctrl_ls25_1b I144 ( .in(gwlb_en), .out_25(gwlb_en_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vpp ( .in(gwphv_vppint),
     .out_25(gwphv_vppint_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwlb_vddp ( .in(gwlbsup_vddp),
     .out_25(gwlbsup_vddp_25));
ml_gwlwr_ctrl_ls25_1b ls25_gwlb_vpp ( .in(gwlbsup_vpxa),
     .out_25(gwlbsup_vpxa_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_vdd ( .in(wrsup_2vdd),
     .out_25(wrsup_2vdd_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_dis ( .in(wr_dis), .out_25(wr_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vddp ( .in(gwphv_vddp),
     .out_25(gwphv_vddp_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_frcen ( .in(wp_frcen),
     .out_25(wp_frcen_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_dis ( .in(wp_dis), .out_25(wp_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwl_red ( .in(gwl_red),
     .out_25(gwl_red_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_nvcm ( .in(gwl_nvcm),
     .out_25(gwl_nvcm_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_misc ( .in(gwl_misc),
     .out_25(gwl_misc_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_1_ ( .in(gred[1]),
     .out_25(gred_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_0_ ( .in(gred[0]),
     .out_25(gred_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_5_ ( .in(gnv[5]), .out_25(gnv_25[5]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_4_ ( .in(gnv[4]), .out_25(gnv_25[4]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_3_ ( .in(gnv[3]), .out_25(gnv_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_2_ ( .in(gnv[2]), .out_25(gnv_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_1_ ( .in(gnv[1]), .out_25(gnv_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_0_ ( .in(gnv[0]), .out_25(gnv_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_3_ ( .in(s[3]), .out_25(s_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_2_ ( .in(s[2]), .out_25(s_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_1_ ( .in(s[1]), .out_25(s_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_0_ ( .in(s[0]), .out_25(s_25[0]));
ml_gwlwr_ctrl_ls25_1b I136 ( .in(pgminhi_dmmy_b),
     .out_25(pgminhi_dmmy_b_25));
ml_gwlwr_ctrl_ls25_1b I140 ( .in(fsm_gwlbdis), .out_25(net101));
ml_gwlwr_ctrl_ls25_1b I137 ( .in(testdec_even_b),
     .out_25(testdec_even_b_25));
ml_gwlwr_ctrl_ls25_1b I138 ( .in(testdec_odd_b),
     .out_25(testdec_odd_b_25));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_npgate_gen, View - schematic
// LAST TIME SAVED: Aug  3 19:28:59 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_core_sa_npgate_gen ( sa_ngate, saen_25, saen_b_vpxa,
     saprd_b_vpxa, sdiode_en_vpxa, vpxa, fsm_tm_rprd, fsm_tm_sdiode,
     fsm_tm_testdec, saen, satrim, vddp_tieh );
output  saen_25, saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa;

inout  vpxa;

input  fsm_tm_rprd, fsm_tm_sdiode, fsm_tm_testdec, saen, vddp_tieh;

output [4:1]  sa_ngate;

input [2:0]  satrim;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  dec_trim_b;

wire  [4:1]  trim;

wire  [3:0]  net48;

wire  [7:0]  dec_trim;

wire  [2:0]  ydec;

wire  [2:0]  ydec_b;



nand2_hvt I183 ( .Y(net037), .B(fsm_tm_rprd), .A(net078));
inv_25 I149 ( .IN(net052), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nor4_hvt I102 ( .D(fsm_tm_testdec), .C(dec_trim[7]), .A(dec_trim[5]),
     .B(dec_trim[6]), .Y(net47));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_4_ ( .Y(dec_trim_b[4]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_3_ ( .Y(dec_trim_b[3]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_2_ ( .Y(dec_trim_b[2]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nand3_hvt I37_1_ ( .Y(dec_trim_b[1]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_0_ ( .Y(dec_trim_b[0]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nor2_hvt I75_4_ ( .Y(net48[0]), .B(dec_trim[4]), .A(sa_high_res));
nor2_hvt I75_3_ ( .Y(net48[1]), .B(dec_trim[3]), .A(trim[4]));
nor2_hvt I75_2_ ( .Y(net48[2]), .B(dec_trim[2]), .A(trim[3]));
nor2_hvt I75_1_ ( .Y(net48[3]), .B(dec_trim[1]), .A(trim[2]));
inv_hvt I158_2_ ( .A(satrim[2]), .Y(ydec_b[2]));
inv_hvt I158_1_ ( .A(satrim[1]), .Y(ydec_b[1]));
inv_hvt I158_0_ ( .A(satrim[0]), .Y(ydec_b[0]));
inv_hvt I160_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I160_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I160_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I160_4_ ( .A(dec_trim_b[4]), .Y(dec_trim[4]));
inv_hvt I160_3_ ( .A(dec_trim_b[3]), .Y(dec_trim[3]));
inv_hvt I160_2_ ( .A(dec_trim_b[2]), .Y(dec_trim[2]));
inv_hvt I160_1_ ( .A(dec_trim_b[1]), .Y(dec_trim[1]));
inv_hvt I160_0_ ( .A(dec_trim_b[0]), .Y(dec_trim[0]));
inv_hvt I163 ( .A(net078), .Y(net080));
inv_hvt I162 ( .A(net076), .Y(net078));
inv_hvt I165 ( .A(net073), .Y(net071));
inv_hvt I166 ( .A(net075), .Y(net073));
inv_hvt I167 ( .A(fsm_tm_sdiode), .Y(net075));
inv_hvt I175 ( .A(net059), .Y(net061));
inv_hvt I176 ( .A(net037), .Y(net059));
inv_hvt I114 ( .A(net47), .Y(sa_high_res));
inv_hvt I161 ( .A(saen), .Y(net076));
inv_hvt I159_2_ ( .A(ydec_b[2]), .Y(ydec[2]));
inv_hvt I159_1_ ( .A(ydec_b[1]), .Y(ydec[1]));
inv_hvt I159_0_ ( .A(ydec_b[0]), .Y(ydec[0]));
inv_hvt I76_4_ ( .A(net48[0]), .Y(trim[4]));
inv_hvt I76_3_ ( .A(net48[1]), .Y(trim[3]));
inv_hvt I76_2_ ( .A(net48[2]), .Y(trim[2]));
inv_hvt I76_1_ ( .A(net48[3]), .Y(trim[1]));
inv_hvt I78_4_ ( .A(trim[4]), .Y(sa_ngate[4]));
inv_hvt I78_3_ ( .A(trim[3]), .Y(sa_ngate[3]));
inv_hvt I78_2_ ( .A(trim[2]), .Y(sa_ngate[2]));
inv_hvt I78_1_ ( .A(trim[1]), .Y(sa_ngate[1]));
ml_hv_invx3 I135 ( .sel_hv(net048), .sel_25(net048),
     .vddp_tieh(vddp_tieh), .out_b_hv(saen_b_vpxa), .in_hv(vpxa));
ml_hv_invx3 I168 ( .sel_hv(net0123), .sel_25(net0123),
     .vddp_tieh(vddp_tieh), .out_b_hv(sdiode_en_vpxa), .in_hv(vpxa));
ml_hv_invx3 I178 ( .sel_hv(net0109), .sel_25(net0109),
     .vddp_tieh(vddp_tieh), .out_b_hv(saprd_b_vpxa), .in_hv(vpxa));
ml_ls_vdd2vdd25 I136 ( .in(net053), .sup(vpxa), .out_vddio_b(net047),
     .out_vddio(net048), .in_b(net052));
ml_ls_vdd2vdd25 I137 ( .in(net078), .sup(vddp_), .out_vddio_b(net052),
     .out_vddio(net053), .in_b(net080));
ml_ls_vdd2vdd25 I172 ( .in(net0129), .sup(vpxa), .out_vddio_b(net0123),
     .out_vddio(net0124), .in_b(net0128));
ml_ls_vdd2vdd25 I173 ( .in(net073), .sup(vddp_), .out_vddio_b(net0128),
     .out_vddio(net0129), .in_b(net071));
ml_ls_vdd2vdd25 I180 ( .in(net0104), .sup(vpxa), .out_vddio_b(net0108),
     .out_vddio(net0109), .in_b(net0103));
ml_ls_vdd2vdd25 I181 ( .in(net059), .sup(vddp_), .out_vddio_b(net0103),
     .out_vddio(net0104), .in_b(net061));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl, View - schematic
// LAST TIME SAVED: Aug  3 19:29:02 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25, gred_25,
     gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25,
     gwlb_en_25, pgminhi_dmmy_b_25, s_25, s_rd_b_hv, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, bgr, bl_pgm_glb,
     gwl_b_sup_25, gwp_sup_hv, srdsup_hv, vddp_tieh, vpp_int, vpxa,
     wr_sup_25, fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rprd, fsm_tm_trow,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, s_rdin_hv, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25;

inout  bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv, srdsup_hv, vddp_tieh,
     vpp_int, vpxa, wr_sup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [5:0]  gnv_b_25;
output [3:0]  s_25;
output [5:0]  gnv_25;
output [1:0]  gred_b_25;
output [4:1]  sa_ngate;
output [1:0]  gred_25;
output [3:0]  s_rd_b_hv;

input [2:0]  fsm_trim_rrefpgm;
input [7:0]  fsm_rowadd;
input [0:0]  fsm_coladd;
input [3:0]  fsm_trim_ipp;
input [3:0]  s_rdin_hv;
input [2:0]  fsm_trim_rrefrd;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  gred;

wire  [2:0]  sa_trim;

wire  [3:0]  s;

wire  [5:0]  gnv;



P_25_LP  M9 ( .D(vddp_tieh), .B(vddp_), .G(net0159), .S(vddp_));
N_11_LPHVT  M2 ( .D(net0159), .B(GND_), .G(net0159), .S(gnd_));
vdd_tielow I204 ( .gnd_tiel(net0165));
ml_rdhv_inv Iml_rdhv_inv_3_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[3]), .s_rd_b_hv(s_rd_b_hv[3]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_2_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[2]), .s_rd_b_hv(s_rd_b_hv[2]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_1_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[1]), .s_rd_b_hv(s_rd_b_hv[1]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_0_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[0]), .s_rd_b_hv(s_rd_b_hv[0]),
     .vddp_tieh(vddp_tieh));
ml_hvmux_hotswitch_enhance Ihvmux_gwpsup_hv ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwphv_vppint_25), .sel_hv_a_25(gwphv_vddp_25),
     .out_hv(gwp_sup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_gwlwr_ctrl_logic Igwlwr_ctrl_logic ( .fsm_tm_rprd(fsm_tm_rprd),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_pgmdisc(fsm_pgmdisc), .gwlb_en(gwlb_en),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_rd(fsm_rd), .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[0]), .wrsup_2vdd(wrsup_2vdd),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .testdec_prec_b(testdec_prec_b),
     .testdec_odd_b(testdec_odd_b), .testdec_even_b(testdec_even_b),
     .testdec_en_b(testdec_en_b), .saen(saen), .sa_trim(sa_trim[2:0]),
     .s(s[3:0]), .pgminhi_dmmy_b(net179), .gwphv_vppint(gwphv_vppint),
     .gwphv_vddp(gwphv_vddp), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vddp(gwlbsup_vddp), .gwlb_dis(gwlb_dis),
     .gwl_misc(gwl_misc), .gred(gred[1:0]), .gnv(gnv[5:0]));
ml_hvmux_hotswitch Ihvmux_gwlbsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwlbsup_vpxa_25), .sel_hv_a_25(gwlbsup_vddp_25),
     .out_hv(gwl_b_sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_gwlwr_bldrv Igwlwr_bldrv ( .fsm_din(fsm_din), .tm_dma(tm_dma),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .bl_frc_gnd(gnd_), .bgr(bgr),
     .bl_pgm_glb(bl_pgm_glb));
ml_gwlwr_ctrl_wr_sup Igwlwr_ctrl_wr_sup ( .wrsup_2vdd(wrsup_2vdd),
     .wrsup_2vdd_25(wrsup_2vdd_25), .wr_sup_25(wr_sup_25));
ml_gwlwr_ctrl_ls25 Igwlwr_ctrl_ls25 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_en(gwlb_en), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwlb_dis(gwlb_dis), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vpxa_25(gwlbsup_vpxa_25), .wrsup_2vdd_25(wrsup_2vdd_25),
     .wrsup_2vdd(wrsup_2vdd), .testdec_odd_b(testdec_odd_b),
     .testdec_even_b(testdec_even_b),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .pgminhi_dmmy_b(net179),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwphv_vddp(gwphv_vddp),
     .gwlbsup_vddp(gwlbsup_vddp), .gwphv_vppint(gwphv_vppint),
     .gwlbsup_vddp_25(gwlbsup_vddp_25),
     .gwphv_vppint_25(gwphv_vppint_25), .gwphv_vddp_25(gwphv_vddp_25),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .s(s[3:0]), .gwl_red(fsm_nv_rrow),
     .gwl_nvcm(fsm_nv_bstream), .gwl_misc(gwl_misc), .gred(gred[1:0]),
     .gnv(gnv[5:0]), .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]));
ml_core_sa_npgate_gen Icore_sa_npgate_gen ( .fsm_tm_sdiode(net0165),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .sdiode_en_vpxa(sdiode_en_vpxa), .sa_ngate(sa_ngate[4:1]),
     .fsm_tm_testdec(tm_testdec), .satrim(sa_trim[2:0]),
     .vddp_tieh(vddp_tieh), .saen(saen), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .vpxa(vpxa));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_top_384, View - schematic
// LAST TIME SAVED: Jan 18 18:03:26 2012
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_gwlwr_top_384 ( fsm_gwlbdis_b_25, gwl_b_25, gwl_b_sup_25,
     gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b, wr, bgr,
     bl_pgm_glb, srdsup_hv, vpp_int, vpxa, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     s_rdin_hv, tm_dma, tm_testdec, tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_b_sup_25, pgminhi_dmmy_b_25, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b;

inout  bgr, bl_pgm_glb, srdsup_hv, vpp_int, vpxa;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [27:0]  wr;
output [6:0]  gwl_b_25;
output [3:0]  s_rd_b_hv;
output [6:0]  gwp_hv;
output [4:1]  sa_ngate;

input [0:0]  fsm_coladd;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  s_rdin_hv;
input [3:0]  fsm_trim_ipp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  gnv_b_25;

wire  [1:0]  gred_25;

wire  [1:0]  gred_b_25;

wire  [3:0]  s_25;

wire  [5:0]  gnv_25;



ml_gwlwr_384 Igwlwr ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .wr_sup_25(wr_sup_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));
ml_gwlwr_ctrl Igwlwr_ctrl ( .saprd_b_vpxa(saprd_b_vpxa),
     .sdiode_en_vpxa(sdiode_en_vpxa), .srdsup_hv(srdsup_hv),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rdin_hv(s_rdin_hv[3:0]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_en_b(testdec_en_b), .testdec_prec_b(testdec_prec_b),
     .fsm_pgmdisc(fsm_pgmdisc), .gwlb_en_25(gwlb_en_25),
     .fsm_din(fsm_din), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_allwl_l(fsm_tm_allwl_l), .fsm_tm_allwl_h(fsm_tm_allwl_h),
     .fsm_tm_allbl_l(fsm_tm_allbl_l), .fsm_tm_allbl_h(fsm_tm_allbl_h),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .s_25(s_25[3:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_red_25(gwl_red_25), .gwl_nvcm_25(gwl_nvcm_25),
     .gwl_misc_25(gwl_misc_25), .gred_b_25(gred_b_25[1:0]),
     .gred_25(gred_25[1:0]), .gnv_b_25(gnv_b_25[5:0]),
     .gnv_25(gnv_25[5:0]), .wr_sup_25(wr_sup_25), .vpxa(vpxa),
     .vpp_int(vpp_int), .vddp_tieh(vddp_tieh), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr));

endmodule
// Library - NVCM_40nm, Cell - ml_core_bank_1_384, View - schematic
// LAST TIME SAVED: Jan 18 18:03:45 2012
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_core_bank_1_384 ( fsm_gwlbdis_b_25, gwl_b_25, gwp_hv,
     nv_dataout, pgminhi_dmmy_b_25, s_rd, s_rd_b_hv, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b, wr, bgr,
     bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     srdsup_hv, vblinhi_rde, vblinhi_rdo, vpp_int, vpxa, ysup_25,
     fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din, fsm_gwlbdis,
     fsm_lshven, fsm_multibl_read, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b,
     fsm_sample, fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, s_rdin_hv, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr );
output  fsm_gwlbdis_b_25, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b;

inout  bgr, bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     srdsup_hv, vblinhi_rde, vblinhi_rdo, vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [6:0]  gwl_b_25;
output [3:0]  s_rd;
output [4:1]  sa_ngate;
output [3:0]  s_rd_b_hv;
output [27:0]  wr;
output [8:4]  nv_dataout;
output [6:0]  gwp_hv;

input [1:0]  fsm_tm_ref;
input [2:0]  fsm_trim_rrefpgm;
input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
input [3:0]  s_rdin_hv;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_blkadd_b;
input [9:0]  fsm_coladd;
input [3:0]  fsm_trim_ipp;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net590;

wire  [3:0]  net596;

wire  [3:0]  net597;

wire  [3:0]  net591;

wire  [3:0]  net598;

wire  [3:0]  net595;



ml_gwlwr_top_384 Igwlwr_top_384 ( .gwl_b_25(gwl_b_25[6:0]),
     .gwp_hv(gwp_hv[6:0]), .wr(wr[27:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wgnden(fsm_wgnden), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_tm_allbl_h(tm_allbl_h),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_lshven(fsm_lshven), .fsm_wren(fsm_wren),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .testdec_en_b(testdec_en_b), .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sdiode_en_vpxa(sdiode_en_vpxa), .srdsup_hv(srdsup_hv),
     .vpxa(vpxa), .vpp_int(vpp_int), .bl_pgm_glb(bl_pgm_glb),
     .bgr(bgr), .gwl_b_sup_25(gwl_b_sup_25), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rdin_hv(s_rdin_hv[3:0]), .tm_testdec(fsm_tm_testdec),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .sa_ngate(sa_ngate[4:1]), .testdec_prec_b(testdec_prec_b),
     .fsm_wpen(fsm_wpen), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_tm_allwl_l(tm_allwl_l), .fsm_tm_allbl_l(tm_allbl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .fsm_din(fsm_din), .tm_dma(tm_dma));
ml_core_328x24_top_384 Iblk_4 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net590[0], net590[1], net590[2], net590[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[4]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_328x24_top_384 Iblk_7 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net596[0], net596[1], net596[2], net596[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd[1], fsm_blkadd[0]}), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .ysup_25(ysup_25), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .testdec_odd_b_25(testdec_odd_b_25),
     .vpxa(vpxa), .testdec_even_b_25(testdec_even_b_25),
     .saen_b_vpxa(saen_b_vpxa), .vblinhi_rdo(vblinhi_rdo),
     .saen_25(saen_25), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[7]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_328x24_top_384 blk_6 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net597[0], net597[1], net597[2], net597[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[6]),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_tm_trow(fsm_tm_trow),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_rd(fsm_rd),
     .bl_pgm_glb(bl_pgm_glb), .fsm_rowadd(fsm_rowadd[1:0]),
     .gwl_b_sup_25(gwl_b_sup_25), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .ngate_25(ngate_25), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .saen_25(saen_25), .vblinhi_rdo(vblinhi_rdo),
     .saen_b_vpxa(saen_b_vpxa), .testdec_even_b_25(testdec_even_b_25),
     .vpxa(vpxa), .testdec_odd_b_25(testdec_odd_b_25),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ysup_25(ysup_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd[2], fsm_blkadd[1],
     fsm_blkadd_b[0]}), .tm_testdec_wr(tm_testdec_wr),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_328x24_top_384 Iblk_5 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net598[0], net598[1], net598[2], net598[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[5]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_328x24_top_384 Iblk_8 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rd({net595[0], net595[1], net595[2], net595[3]}),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .sa_ngate(sa_ngate[4:1]),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[8]),
     .fsm_coladd(fsm_coladd[9:0]));
inv_hvt I66_3_ ( .A(net590[0]), .Y(net591[0]));
inv_hvt I66_2_ ( .A(net590[1]), .Y(net591[1]));
inv_hvt I66_1_ ( .A(net590[2]), .Y(net591[2]));
inv_hvt I66_0_ ( .A(net590[3]), .Y(net591[3]));
inv_hvt I6_3_ ( .A(net591[0]), .Y(s_rd[3]));
inv_hvt I6_2_ ( .A(net591[1]), .Y(s_rd[2]));
inv_hvt I6_1_ ( .A(net591[2]), .Y(s_rd[1]));
inv_hvt I6_0_ ( .A(net591[3]), .Y(s_rd[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_core_384, View - schematic
// LAST TIME SAVED: Jan 18 17:22:34 2012
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_chip_nvcm_core_384 ( nv_dataout, s_rd, bgr, ngate_25,
     sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi, vpp_int, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_multibl_read, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_ref,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_trim_ipp,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, s_rdin_hv, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi,
     vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [3:0]  s_rd;
output [8:0]  nv_dataout;

input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_trim_ipp;
input [7:0]  fsm_rowadd;
input [3:0]  s_rdin_hv;
input [1:0]  fsm_tm_ref;
input [2:0]  fsm_trim_rrefrd;
input [9:0]  fsm_coladd;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefpgm;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [6:0]  gwp_hv;

wire  [27:0]  wr;

wire  [6:0]  gwl_b_25;

wire  [3:0]  s_rd_b_hv;

wire  [4:1]  sa_ngate;



ml_core_bank_0_384 Ibank_0 ( .gwl_b_25(gwl_b_25[6:0]),
     .gwp_hv(gwp_hv[6:0]), .wr(wr[27:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .saen_25(saen_25), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .saen_b_vpxa(saen_b_vpxa),
     .saprd_b_vpxa(saprd_b_vxpa), .gwl_b_sup_25(gwl_b_sup_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .fsm_nvcmen(fsm_nvcmen), .fsm_pgm(fsm_pgm),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd(fsm_blkadd[3:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_tm_trow(fsm_tm_trow), .ngate_25(ngate_25),
     .nv_dataout(nv_dataout[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .tm_allbank_sel(tm_allbank_sel));
ml_core_bank_1_384 Ibank_1 ( .wr(wr[27:0]), .gwp_hv(gwp_hv[6:0]),
     .gwl_b_25(gwl_b_25[6:0]), .s_rdin_hv(s_rdin_hv[3:0]),
     .srdsup_hv(srdsup_hv), .sdiode_en_vpxa(net230),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_din(fsm_din), .fsm_wren(fsm_wren), .fsm_pgmhv(fsm_pgmhv),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_wgnden(fsm_wgnden), .bgr(bgr), .vpp_int(vpp_int),
     .sa_ngate(sa_ngate[4:1]), .testdec_prec_b(testdec_prec_b),
     .testdec_en_b(testdec_en_b), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .tm_allbank_sel(tm_allbank_sel), .saprd_b_vpxa(saprd_b_vxpa),
     .gwl_b_sup_25(gwl_b_sup_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .ngate_25(ngate_25),
     .s_rd(s_rd[3:0]), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .bl_pgm_glb(bl_pgm_glb),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd(fsm_blkadd[3:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_rprd(fsm_tm_rprd), .nv_dataout(nv_dataout[8:4]));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_buf, View - schematic
// LAST TIME SAVED: Aug  3 19:28:53 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_bgr_buf ( sa_out, en_25, inn, inp, sa_bias_25 );
inout  sa_out;

input  en_25, inn, inp, sa_bias_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M95 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M94 ( .D(net0119), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
P_25_LP  M96 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M71 ( .D(sa_mirr_25), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
P_25_LP  M101 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M102 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
P_25_LP  M98 ( .D(net0239), .B(vddp_), .G(net0239), .S(vddp_));
P_25_LP  M10 ( .D(sa_mirr_25), .B(vddp_), .G(en_25), .S(vddp_));
P_25_LP  M91 ( .D(sa_out), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
P_25_LP  M25 ( .D(sa_out), .B(vddp_), .G(en_25), .S(vddp_));
P_25_LP  M93 ( .D(net0123), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
N_25_LP  M46 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
N_25_LP  M92 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
N_25_LP  M97 ( .D(tie_low), .B(GND_), .G(net0239), .S(GND_));
N_25_LP  M3 ( .D(net436), .B(GND_), .G(sa_bias_25), .S(GND_));
N_25_LPNVT  M0 ( .D(sa_mirr_25), .B(GND_), .G(inp), .S(net436));
N_25_LPNVT  M1 ( .D(sa_out), .B(GND_), .G(inn), .S(net436));
N_25_LPNVT  M2 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
N_25_LPNVT  M4 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
N_25_LPNVT  M8 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
N_25_LPNVT  M7 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));

endmodule
// Library - sbtlibn65lp, Cell - nand4_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:55 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module nand4_25 ( Y, A, B, C, D, G, Gb, P, Pb );
output  Y;

input  A, B, C, D, G, Gb, P, Pb;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
P_25_LP  M0 ( .D(Y), .B(Pb), .G(B), .S(P));
P_25_LP  M3 ( .D(Y), .B(Pb), .G(D), .S(P));
P_25_LP  M2 ( .D(Y), .B(Pb), .G(C), .S(P));
N_25_LP  M6 ( .D(net14), .B(Gb), .G(C), .S(net10));
N_25_LP  M7 ( .D(net10), .B(Gb), .G(D), .S(G));
N_25_LP  M4 ( .D(Y), .B(Gb), .G(A), .S(net18));
N_25_LP  M5 ( .D(net18), .B(Gb), .G(B), .S(net14));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ref_sw, View - schematic
// LAST TIME SAVED: Aug  3 19:29:13 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_vpp_ref_sw ( in, out, sel_b_25 );
inout  in, out;

input  sel_b_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M14 ( .D(in), .B(vddp_), .G(sel_b_25), .S(out));
N_25_LP  M12 ( .D(out), .B(GND_), .G(net122), .S(in));
inv_25 I281 ( .IN(sel_b_25), .OUT(net122), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_res_100_ohm, View - schematic
// LAST TIME SAVED: Oct 18 18:17:24 2011
// NETLIST TIME: Jan 18 18:48:17 2012
`timescale 1ns / 1ns 

module ml_bgr_res_100_ohm ( b, t );
inout  b, t;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



RNPPO_LP_pcell2460 R0 ( .B(gnd_), .MINUS(b), .PLUS(t));
RNPPO_LP_pcell2460 R1 ( .B(gnd_), .MINUS(b), .PLUS(t));
RNPPO_LP_pcell2460 R2 ( .B(gnd_), .MINUS(b), .PLUS(t));
RNPPO_LP_pcell2460 R3 ( .B(gnd_), .MINUS(b), .PLUS(t));
RNPPO_LP_pcell2460 R4 ( .B(gnd_), .MINUS(b), .PLUS(t));
RNPPO_LP_pcell2460 R5 ( .B(gnd_), .MINUS(b), .PLUS(t));
RNPPO_LP_pcell2460 R6 ( .B(gnd_), .MINUS(net7), .PLUS(net7));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_sup_25, View - schematic
// LAST TIME SAVED: Aug  3 19:21:56 2011
// NETLIST TIME: Jan 18 18:48:16 2012
`timescale 1ns / 1ns 

module oai21x2_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply1 vdd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 gnd_;
supply0 GND_;
supply1 VDD_;



P_25_LP  M0 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));
P_25_LP  M3 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));
P_25_LP  M2 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
N_25_LP  M1 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
N_25_LP  M4 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
N_25_LP  M7 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));

endmodule
