// Library - ice8chip, Cell - fabric_buf_ice8p, View - schematic
// LAST TIME SAVED: Aug 13 15:11:11 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module fabric_buf_ice8p ( f_out, f_in );
output  f_out;

input  f_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I_inv_lvt_2 ( .A(net6), .Y(f_out));
inv_lvt I_inv_lvt_1 ( .A(f_in), .Y(net6));

endmodule
// Library - io, Cell - cebdffrqn, View - schematic
// LAST TIME SAVED: Apr 27 16:16:03 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module cebdffrqn ( q, qn, ceb, clk, d, r );
output  q, qn;

input  ceb, clk, d, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I43 ( .A(so), .Y(low_s));
inv_lvt I50 ( .A(clkb), .Y(clkd));
inv_lvt Iinv_ckfb ( .A(clatb), .Y(net50));
inv_lvt I40 ( .A(r), .Y(rstb));
inv_lvt I_q_inv ( .A(qn), .Y(q));
inv_lvt I39 ( .A(net77), .Y(qn));
txgate_lvt I52 ( .in(so), .out(mi), .pp(clkb), .nn(clkd));
txgate_lvt I44 ( .in(d), .out(si), .pp(clkd), .nn(clkb));
txgate_lvt I51 ( .in(si), .out(low_s), .pp(clkb), .nn(clkd));
txgate_lvt I53 ( .in(mi), .out(qn), .pp(clkd), .nn(clkb));
nand2_lvt I290 ( .A(clk), .Y(clkb), .B(clatb));
nand2_lvt I42 ( .A(si), .Y(so), .B(rstb));
nor2_lvt INAND2_m ( .A(r), .B(mi), .Y(net77));
anor21_lvt I54 ( .A(net50), .B(clk), .Y(clatb), .C(ceb));

endmodule
// Library - io, Cell - dffrckb, View - schematic
// LAST TIME SAVED: Aug 12 13:15:42 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module dffrckb ( q, qn, clk, d, e, r );
output  q, qn;

input  clk, d, e, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



oai21x2_lvt I57 ( .A1(clk), .Y(clat), .A0(clatb), .B0(e));
nor2_lvt I48 ( .B(clat), .A(clk), .Y(clkb));
nand2_lvt I54 ( .A(rstb), .Y(qn), .B(q));
nand2_lvt I42 ( .A(si), .B(rstb), .Y(so));
txgate_lvt I59 ( .in(d), .out(si), .pp(clkb), .nn(clkd));
txgate_lvt I64 ( .in(low_s), .out(si), .pp(clkd), .nn(clkb));
txgate_lvt I62 ( .in(qn), .out(mi), .pp(clkb), .nn(clkd));
txgate_lvt I60 ( .in(so), .out(mi), .pp(clkd), .nn(clkb));
inv_lvt I55 ( .A(mi), .Y(q));
inv_lvt I50 ( .A(clkb), .Y(clkd));
inv_lvt I56 ( .A(clat), .Y(clatb));
inv_lvt I43 ( .A(so), .Y(low_s));
inv_lvt I40 ( .A(r), .Y(rstb));

endmodule
// Library - io, Cell - in_logic_v1_imp, View - schematic
// LAST TIME SAVED: Dec 22 12:28:01 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module in_logic_v1_imp ( dout0, dout1, sdo, bs_en, cbit, cbitb, ceb,
     clk, cntl, din, mode, rstio, sdi, shift, tclk, ud );
output  dout0, dout1, sdo;

input  bs_en, ceb, clk, cntl, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



insel1_lvt_imp I_insel1 ( .in1(dinb), .in0(regb), .out(reg_),
     .sb({cbit1b, cbitb[0]}), .sel({cbit1, cbit[0]}), .in2(net037),
     .in3(net037));
mux2x1_hvt I_mux_mode ( .sel(mode), .in1(udd), .in0(reg_),
     .out(doutb));
mux2x1_hvt I_mux_clk ( .in1(tclk), .in0(clk), .out(ck2r0),
     .sel(bs_en));
mux2x1_hvt I_mux_data ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
mux2x1_hvt I_mux2_btw ( .in1(sdo), .in0(din), .out(net056),
     .sel(bs_en));
nand2_lvt I188 ( .A(cntl), .Y(cbit1b), .B(cbit[1]));
inv_lvt I_inv_dout0 ( .A(doutb), .Y(dout0));
inv_lvt I_inv_dout1 ( .A(udd), .Y(dout1));
inv_lvt I185 ( .A(cbit1b), .Y(cbit1));
inv_lvt I186 ( .A(dout0), .Y(net037));
inv_lvt I172 ( .A(din), .Y(dinb));
cebdffrqn I_dff0 ( .ceb(ceb), .clk(ck2r0), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff1 ( .e(ud), .clk(ck2r0), .qn(udd), .r(rstio), .q(net060),
     .d(net056));

endmodule
// Library - io, Cell - in_logic_v3_imp, View - schematic
// LAST TIME SAVED: Aug  9 13:26:43 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module in_logic_v3_imp ( dout0, dout1, sdo, sp12, bl, bs_en, ceb, clk,
     cntl, din, mode, pgate, prog, reset, rstio, sdi, shift, slfop,
     tclk, ud, vdd_cntl, wl );
output  dout0, dout1, sdo, sp12;


input  bs_en, ceb, clk, cntl, din, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
in_logic_v1_imp I_in_logic ( .ceb(ceb), .rstio(rstio), .din(din),
     .cntl(cntl), .dout1(dout1), .dout0(dout0), .shift(shift), .ud(ud),
     .clk(clk), .sdo(sdo), .sdi(sdi), .cbit({cbit[0], cbit[1]}),
     .cbitb({cbitb[0], cbitb[1]}), .tclk(tclk), .bs_en(bs_en),
     .mode(mode));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[3]), .sp12(sp12),
     .prog(prog));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - outsel1_lvt, View - schematic
// LAST TIME SAVED: Nov 22 19:11:18 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module outsel1_lvt ( out, clk, in0, in1, in2, sb, sel );
output  out;

input  clk, in0, in1, in2;

input [1:0]  sel;
input [1:0]  sb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I41 ( .A(in1), .Y(net036));
inv_lvt I40 ( .A(clk), .Y(clkb));
txgate_lvt I33 ( .in(whatever), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_lvt I_txgate1 ( .in(net036), .out(whatever), .pp(sb[0]),
     .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(whatever), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(ddr), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_lvt I38 ( .in(in2), .out(ddr), .pp(clkb), .nn(clk));
txgate_lvt I39 ( .in(in1), .out(ddr), .pp(clk), .nn(clkb));

endmodule
// Library - io, Cell - out_logic_v1, View - schematic
// LAST TIME SAVED: Aug 13 11:02:21 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module out_logic_v1 ( dout, sdo, bs_en, cbit, cbitb, ceb, clk, ddr0,
     ddr1, mode, rstio, sdi, shift, tclk, ud );
output  dout, sdo;

input  bs_en, ceb, clk, ddr0, ddr1, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



outsel1_lvt I169 ( .clk(ddrclk), .in2(udb), .sb(cbitb[1:0]),
     .sel(cbit[1:0]), .in1(net094), .in0(dinb), .out(muxob));
mux2x1_hvt I170 ( .sel(mode), .in1(udb), .in0(muxob), .out(doutb));
mux2x1_hvt I177 ( .in1(tclk), .in0(clk), .out(mux4clk), .sel(bs_en));
mux2x1_hvt I173 ( .in1(sdi), .in0(ddr0), .out(dd), .sel(shift));
mux2x1_hvt I176 ( .in1(sdo), .in0(ddr1), .out(mux4d), .sel(bs_en));
nor2_lvt I179 ( .A(mux4clk), .B(cbit[0]), .Y(ddrclk));
inv_lvt I171 ( .A(doutb), .Y(dout));
inv_lvt I172 ( .A(ddr0), .Y(dinb));
cebdffrqn I_reg0 ( .ceb(ceb), .clk(mux4clk), .qn(net094), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_reg1 ( .e(ud), .clk(mux4clk), .qn(udb), .r(rstio), .q(net44),
     .d(mux4d));

endmodule
// Library - io, Cell - out_logic_v3, View - schematic
// LAST TIME SAVED: Aug  9 13:26:57 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module out_logic_v3 ( dout, sdo, sp12, bl, bs_en, ceb, clk, ddr0, ddr1,
     mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk, ud,
     vdd_cntl, wl );
output  dout, sdo, sp12;


input  bs_en, ceb, clk, ddr0, ddr1, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;

wire  [3:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
out_logic_v1 I_outlogic_v1 ( .shift(shift), .ud(ud), .clk(clk),
     .sdo(sdo), .sdi(sdi), .ceb(ceb), .cbit({cbit[2], cbit[3]}),
     .cbitb({cbitb[2], cbitb[3]}), .dout(dout), .ddr0(ddr0),
     .tclk(tclk), .bs_en(bs_en), .rstio(rstio), .ddr1(ddr1),
     .mode(mode));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
odrv12 I_odrv12 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp12(sp12));

endmodule
// Library - io, Cell - ioesel_lvt, View - schematic
// LAST TIME SAVED: Dec  1 14:31:52 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioesel_lvt ( out, in0, in1, sb, sel );
output  out;

input  in0, in1;

input [1:0]  sb;
input [1:0]  sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I38 ( .A(sel[0]), .Y(net017));
txgate_lvt I33 ( .in(mid), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_lvt I_txgate1 ( .in(in1), .out(mid), .pp(sb[0]), .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(mid), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(net017), .out(out), .pp(sel[1]), .nn(sb[1]));

endmodule
// Library - io, Cell - ioe_logic_v1, View - schematic
// LAST TIME SAVED: Aug 13 14:52:51 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioe_logic_v1 ( outb, sdo, bs_en, cbit, cbitb, ceb, clk, din,
     mode, rstio, sdi, shift, tclk, ud );
output  outb, sdo;

input  bs_en, ceb, clk, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ioesel_lvt I_ioe_mux2 ( .sb(cbitb[1:0]), .sel(cbit[1:0]), .in1(regb),
     .in0(dinb), .out(regmuxb));
mux2x1_hvt I175 ( .in1(tclk), .in0(clk), .out(net039), .sel(bs_en));
mux2x1_hvt I170 ( .sel(mode), .in1(udd), .in0(regmuxb), .out(outb));
mux2x1_hvt I173 ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
inv_lvt I172 ( .A(din), .Y(dinb));
cebdffrqn I_dff_1 ( .ceb(ceb), .clk(net039), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I_dff_2 ( .e(ud), .clk(net039), .qn(udd), .r(rstio), .q(net44),
     .d(sdo));

endmodule
// Library - io, Cell - ioe_logic_v3, View - schematic
// LAST TIME SAVED: Aug 12 13:29:42 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioe_logic_v3 ( padeb, sdo, sp12, bl, bs_en, ceb, clk, din,
     hiz_b, mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk,
     ud, vdd_cntl, wl );
output  padeb, sdo, sp12;


input  bs_en, ceb, clk, din, hiz_b, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbit;

wire  [3:0]  cbitb;



inv_lvt I_inv ( .A(oeb), .Y(oed));
nand2_lvt I_nand2 ( .A(oed), .Y(padeb), .B(hiz_b));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
ioe_logic_v1 I_ioe_logic ( .shift(shift), .ud(ud), .clk(clk),
     .sdo(sdo), .sdi(sdi), .cbit(cbit[3:2]), .din(din),
     .cbitb(cbitb[3:2]), .ceb(ceb), .rstio(rstio), .bs_en(bs_en),
     .tclk(tclk), .outb(oeb), .mode(mode));
odrv12 I_odrv12x2 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp12(sp12));

endmodule
// Library - leafcell, Cell - dffs, View - schematic
// LAST TIME SAVED: Dec  3 13:08:03 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module dffs ( Q, QN, CLK, D, S );
output  Q, QN;

input  CLK, D, S;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net45), .Y(net38));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net42));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net49), .Y(net42));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net49), .Y(net38));
nand2_hvt I5 ( .A(net38), .Y(net45), .B(net26));
nand2_hvt I125 ( .A(net42), .Y(net49), .B(net26));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));
inv_hvt I146 ( .A(net38), .Y(Q));
inv_hvt I147 ( .A(net45), .Y(QN));
inv_hvt I2 ( .A(S), .Y(net26));
inv_hvt I131 ( .A(CLK), .Y(clk_b));

endmodule
// Library - io, Cell - odrv12x3, View - schematic
// LAST TIME SAVED: Aug  9 13:26:19 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module odrv12x3 ( sp12, bl, pgate, prog, reset, slfop, vdd_cntl, wl );


input  prog;

output [2:0]  sp12;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  reset;
input [2:0]  slfop;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12_2_ ( .slfop(slfop[2]), .cbitb(cbitb[2]),
     .sp12(sp12[2]), .prog(prog));
odrv12 I_odrv12_1_ ( .slfop(slfop[1]), .cbitb(cbitb[1]),
     .sp12(sp12[1]), .prog(prog));
odrv12 I_odrv12_0_ ( .slfop(slfop[0]), .cbitb(cbitb[0]),
     .sp12(sp12[0]), .prog(prog));
cram2x2 I_cram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioe_col2_v3, View - schematic
// LAST TIME SAVED: May 12 17:42:20 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioe_col2_v3 ( dout, padeb, pado, sdo, sp12_h_l, bl, bs_en, ceb,
     hiz_b, hold, inclk, mode, outclk, padin, pgate, prog, reset,
     rstio, sdi, shift, tclk, ti, update, vdd_cntl, wl );
output  sdo;


input  bs_en, ceb, hiz_b, hold, inclk, mode, outclk, prog, rstio, sdi,
     shift, tclk, update;

output [1:0]  pado;
output [23:0]  sp12_h_l;
output [3:0]  dout;
output [1:0]  padeb;

inout [1:0]  bl;

input [1:0]  padin;
input [5:0]  ti;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



in_logic_v3_imp I_in1 ( .slfop(dout[3]), .shift(shift),
     .dout1(dout[3]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[2]), .sp12(sp12_h_l[14]), .wl(wl[13:12]),
     .ceb(ceb), .reset(reset[13:12]), .sdo(s4), .sdi(s3),
     .vdd_cntl(vdd_cntl[13:12]), .pgate(pgate[13:12]), .din(padin[1]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode),
     .rstio(rstio));
in_logic_v3_imp I_in0 ( .slfop(dout[0]), .shift(shift),
     .dout1(dout[1]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[0]), .sp12(sp12_h_l[8]), .wl(wl[3:2]),
     .ceb(ceb), .reset(reset[3:2]), .sdo(s1), .sdi(s0),
     .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]), .din(padin[0]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode),
     .rstio(rstio));
out_logic_v3 I_out1 ( .shift(shift), .slfop(dout[3]), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .sp12(sp12_h_l[6]),
     .wl(wl[11:10]), .ceb(ceb), .reset(reset[11:10]), .sdo(s3),
     .sdi(s2), .vdd_cntl(vdd_cntl[11:10]), .pgate(pgate[11:10]),
     .dout(pado[1]), .tclk(tclk), .bs_en(bs_en), .rstio(rstio),
     .ddr1(ti[5]), .mode(mode), .ddr0(ti[4]));
out_logic_v3 I_out0 ( .shift(shift), .slfop(dout[0]), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .sp12(sp12_h_l[0]),
     .wl(wl[1:0]), .ceb(ceb), .reset(reset[1:0]), .sdo(s0), .sdi(sdi),
     .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]), .dout(pado[0]),
     .tclk(tclk), .bs_en(bs_en), .rstio(rstio), .ddr1(ti[2]),
     .mode(mode), .ddr0(ti[1]));
ioe_logic_v3 I_ioe0 ( .shift(shift), .hiz_b(hiz_b), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .padeb(padeb[0]),
     .slfop(dout[0]), .sp12(sp12_h_l[16]), .wl(wl[5:4]), .ceb(ceb),
     .reset(reset[5:4]), .sdo(s2), .sdi(s1), .pgate(pgate[5:4]),
     .din(ti[0]), .tclk(tclk), .vdd_cntl(vdd_cntl[5:4]), .bs_en(bs_en),
     .mode(mode), .rstio(rstio));
ioe_logic_v3 I_ioe1 ( .shift(shift), .hiz_b(hiz_b), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .padeb(padeb[1]),
     .slfop(dout[3]), .sp12(sp12_h_l[22]), .wl(wl[15:14]), .ceb(ceb),
     .reset(reset[15:14]), .sdo(sdo), .sdi(s4), .pgate(pgate[15:14]),
     .din(ti[3]), .tclk(tclk), .vdd_cntl(vdd_cntl[15:14]),
     .bs_en(bs_en), .mode(mode), .rstio(rstio));
odrv12x3 I_odrv12x3_1 ( .bl(bl[1:0]), .wl(wl[7:6]), .reset(reset[7:6]),
     .pgate(pgate[7:6]), .slfop({dout[1], dout[1], dout[1]}),
     .sp12({sp12_h_l[18], sp12_h_l[10], sp12_h_l[2]}),
     .vdd_cntl(vdd_cntl[7:6]), .prog(prog));
odrv12x3 I_odrv12x3_2 ( .bl(bl[1:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]), .slfop({dout[2], dout[2], dout[2]}),
     .sp12({sp12_h_l[20], sp12_h_l[12], sp12_h_l[4]}),
     .vdd_cntl(vdd_cntl[9:8]), .prog(prog));

endmodule
// Library - io, Cell - io_odrv4x5, View - schematic
// LAST TIME SAVED: Aug  9 13:55:12 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_odrv4x5 ( cbit, sp4_out, bl, pgate, prog,
     reset, slfop, vdd_cntl, wl );


input  prog, slfop;

output [4:0]  sp4_out;
output [7:5]  cbit;

inout [3:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
/* //////wire vddp_ = test.cds_globalsInst.vddp_; */ supply1 vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  cbitb;

wire  [1:0]  r_vdd;

wire [7:0] cbit_int;
assign cbit[7:5] = cbit_int[7:5];



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv4 I_odrv_4_ ( .cbitb(cbitb[4]), .sp4(sp4_out[4]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_3_ ( .cbitb(cbitb[3]), .sp4(sp4_out[3]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_2_ ( .cbitb(cbitb[2]), .sp4(sp4_out[2]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_1_ ( .cbitb(cbitb[1]), .sp4(sp4_out[1]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_0_ ( .cbitb(cbitb[0]), .sp4(sp4_out[0]), .slfop(slfop),
     .prog(prog));
cram2x2 Icram2x2_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset[1:0]), .q(cbit_int[7:4]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));
cram2x2 Icram2x2_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset[1:0]), .q(cbit_int[3:0]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - io_col_odrv4_x40bare_v3, View - schematic
// LAST TIME SAVED: Jun  2 10:03:19 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_col_odrv4_x40bare_v3 ( cf, bl, sp4_h_l,
     sp4_v_b, dout0, dout1,
     pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [23:0]  cf;

inout [3:0]  bl;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_b;

input [0:1]  dout1;
input [0:1]  dout0;
input [15:0]  wl;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
/* //////wire vddp_ = test.cds_globalsInst.vddp_; */ supply1 vddp_;
supply0 GND_;
supply1 VDD_;



io_odrv4x5 I_io_odrv4x5_6 ( cf[20:18], {sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6]}, bl[3:0], pgate[13:12],
     prog, reset[13:12], dout1[1], vdd_cntl[13:12], wl[13:12]);
io_odrv4x5 I_io_odrv4x5_4 ( cf[14:12], {sp4_h_l[36], sp4_h_l[28],
     sp4_h_l[20], sp4_h_l[12], sp4_h_l[4]}, bl[3:0], pgate[9:8], prog,
     reset[9:8], dout0[1], vdd_cntl[9:8], wl[9:8]);
io_odrv4x5 I_io_odrv4x5_7 ( cf[23:21], {sp4_v_b[15], sp4_v_b[11],
     sp4_v_b[7], sp4_v_b[3], sp4_h_l[46]}, bl[3:0], pgate[15:14], prog,
     reset[15:14], dout1[1], vdd_cntl[15:14], wl[15:14]);
io_odrv4x5 I_io_odrv4x5_3 ( cf[11:9], {sp4_v_b[13], sp4_v_b[9],
     sp4_v_b[5], sp4_v_b[1], sp4_h_l[42]}, bl[3:0], pgate[7:6], prog,
     reset[7:6], dout1[0], vdd_cntl[7:6], wl[7:6]);
io_odrv4x5 I_io_odrv4x5_2 ( cf[8:6], {sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2]}, bl[3:0], pgate[5:4], prog,
     reset[5:4], dout1[0], vdd_cntl[5:4], wl[5:4]);
io_odrv4x5 I_io_odrv4x5_0 ( cf[2:0], {sp4_h_l[32], sp4_h_l[24],
     sp4_h_l[16], sp4_h_l[8], sp4_h_l[0]}, bl[3:0], pgate[1:0], prog,
     reset[1:0], dout0[0], vdd_cntl[1:0], wl[1:0]);
io_odrv4x5 I_io_odrv4x5_1 ( cf[5:3], {sp4_v_b[12], sp4_v_b[8],
     sp4_v_b[4], sp4_v_b[0], sp4_h_l[40]}, bl[3:0], pgate[3:2], prog,
     reset[3:2], dout0[0], vdd_cntl[3:2], wl[3:2]);
io_odrv4x5 I_io_odrv4x5_5 ( cf[17:15], {sp4_v_b[14], sp4_v_b[10],
     sp4_v_b[6], sp4_v_b[2], sp4_h_l[44]}, bl[3:0], pgate[11:10], prog,
     reset[11:10], dout0[1], vdd_cntl[11:10], wl[11:10]);

endmodule
// Library - ice8chip, Cell - io_col4_rgt_ice8p_v2, View - schematic
// LAST TIME SAVED: Jan 12 14:59:31 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_col4_rgt_ice8p_v2 ( cbit_colcntl, cf, fabric_out, padeb,
     pado, sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t,
     sp12_h_l, bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold,
     lft_op, mode, padin, pgate, prog, r, reset, sdi, shift, spioeb,
     spiout, tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [23:0]  cf;
output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;
output [7:0]  cbit_colcntl;

inout [15:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;
inout [15:0]  sp4_v_t;
inout [23:0]  sp12_h_l;

input [1:0]  spioeb;
input [1:0]  spiout;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [15:0]  wl;
input [15:0]  reset;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [7:0]  glb_netwk;
input [1:0]  padin;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



rm7w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
sbox1_colbdlc_v4 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_gmux_x16bare_v4 I_io_gmux_x16bare_v4 (
     .cbit_colcntl(cbit_colcntl[7:0]), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});

endmodule
// Library - ice8chip, Cell - tckbufx32_ice8p, View - schematic
// LAST TIME SAVED: Aug 13 15:04:42 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module tckbufx32_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I_inv_lvt_1 ( .A(in), .Y(net4));
inv_lvt Iinv_lvt_2 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - tielo4x, View - schematic
// LAST TIME SAVED: May 18 10:31:28 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module tielo4x ( tielo );
output  tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - tiehi4x, View - schematic
// LAST TIME SAVED: May 18 10:33:00 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module tiehi4x ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - ice1chip, Cell - io_rgt_top_1x8_ice1f, View - schematic
// LAST TIME SAVED: Mar  4 20:34:44 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_rgt_top_1x8_ice1f ( cf_r, fabric_out_09, fabric_out_10,
     padeb, pado, sdo, slf_op_01, slf_op_02, slf_op_03, slf_op_04,
     slf_op_05, slf_op_06, slf_op_07, slf_op_08, tclk_o, SP4_h_l_01,
     SP4_h_l_02, SP4_h_l_03, SP4_h_l_04, SP4_h_l_05, SP4_h_l_06,
     SP4_h_l_07, SP4_h_l_08, SP12_h_l_01, SP12_h_l_02, SP12_h_l_03,
     SP12_h_l_04, SP12_h_l_05, SP12_h_l_06, SP12_h_l_07, SP12_h_l_08,
     bl, pgate, reset_b, sp4_v_b_13_09, sp4_v_t_08, vdd_cntl, wl,
     bnl_op_13_09, bs_en, ceb, glb_netwk_col, hiz_b, hold, lft_op_01,
     lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06, lft_op_07,
     lft_op_08, mode, padin, prog, r, sdi, shift, tclk, tnl_op_08,
     update );
output  fabric_out_09, fabric_out_10, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_03;
output [3:0]  slf_op_08;
output [3:0]  slf_op_06;
output [3:0]  slf_op_02;
output [24:13]  padeb;
output [24:13]  pado;
output [3:0]  slf_op_05;
output [3:0]  slf_op_07;
output [3:0]  slf_op_04;
output [191:0]  cf_r;
output [3:0]  slf_op_01;

inout [23:0]  SP12_h_l_08;
inout [47:0]  SP4_h_l_07;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_01;
inout [23:0]  SP12_h_l_03;
inout [23:0]  SP12_h_l_02;
inout [47:0]  SP4_h_l_03;
inout [15:0]  sp4_v_t_08;
inout [47:0]  SP4_h_l_02;
inout [127:0]  vdd_cntl;
inout [127:0]  reset_b;
inout [127:0]  pgate;
inout [23:0]  SP12_h_l_06;
inout [23:0]  SP12_h_l_01;
inout [23:0]  SP12_h_l_07;
inout [47:0]  SP4_h_l_04;
inout [23:0]  SP12_h_l_04;
inout [127:0]  wl;
inout [47:0]  SP4_h_l_08;
inout [47:0]  SP4_h_l_06;
inout [23:0]  SP12_h_l_05;
inout [15:0]  sp4_v_b_13_09;
inout [47:0]  SP4_h_l_05;

input [7:0]  lft_op_07;
input [7:0]  lft_op_02;
input [7:0]  bnl_op_13_09;
input [7:0]  tnl_op_08;
input [24:13]  padin;
input [7:0]  lft_op_03;
input [7:0]  lft_op_01;
input [7:0]  lft_op_05;
input [7:0]  lft_op_08;
input [7:0]  lft_op_04;
input [7:0]  glb_netwk_col;
input [7:0]  lft_op_06;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net632;

wire  [15:0]  net478;

wire  [7:0]  colbuf_cntl_t;

wire  [7:0]  colbuf_cntl_b;

wire  [7:0]  glb_netwk_b;

wire  [7:0]  glb_netwk_t;

wire  [15:0]  net586;

wire  [1:0]  net618;

wire  [1:0]  net630;

wire  [15:0]  net442;

wire  [7:0]  net633;

wire  [7:0]  net317;

wire  [7:0]  net461;

wire  [1:0]  net590;

wire  [1:0]  net624;

wire  [7:0]  net497;

wire  [1:0]  net625;

wire  [1:0]  net620;

wire  [15:0]  net370;

wire  [1:0]  net628;

wire  [1:0]  net476;

wire  [7:0]  net623;

wire  [1:0]  net616;

wire  [15:0]  net514;

wire  [1:0]  net477;

wire  [1:0]  net332;

wire  [1:0]  net629;

wire  [15:0]  net550;

wire  [15:0]  net406;



io_col4_rgt_ice8p_v2 I_io_00_08 ( .cbit_colcntl({net317[0], net317[1],
     net317[2], net317[3], net317[4], net317[5], net317[6],
     net317[7]}), .ceb(ceb), .sdo(sdo), .sdi(net355), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin({net332[0], net332[1]}),
     .pado({net332[0], net332[1]}), .padeb({net616[0], net616[1]}),
     .sp4_v_t(sp4_v_t_08[15:0]), .sp4_h_l(SP4_h_l_08[47:0]),
     .sp12_h_l(SP12_h_l_08[23:0]), .prog(prog),
     .spi_ss_in_b({net628[0], net628[1]}), .tnl_op(tnl_op_08[7:0]),
     .lft_op(lft_op_08[7:0]), .bnl_op(lft_op_07[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b({net370[0], net370[1], net370[2], net370[3], net370[4],
     net370[5], net370[6], net370[7], net370[8], net370[9], net370[10],
     net370[11], net370[12], net370[13], net370[14], net370[15]}),
     .wl(wl[127:112]), .cf(cf_r[191:168]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[127:112]), .slf_op(slf_op_08[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold), .fabric_out(net352));
io_col4_rgt_ice8p_v2 I_io_00_07 ( .cbit_colcntl({net632[0], net632[1],
     net632[2], net632[3], net632[4], net632[5], net632[6],
     net632[7]}), .ceb(ceb), .sdo(net355), .sdi(net427),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[24:23]), .pado(pado[24:23]), .padeb(padeb[24:23]),
     .sp4_v_t({net370[0], net370[1], net370[2], net370[3], net370[4],
     net370[5], net370[6], net370[7], net370[8], net370[9], net370[10],
     net370[11], net370[12], net370[13], net370[14], net370[15]}),
     .sp4_h_l(SP4_h_l_07[47:0]), .sp12_h_l(SP12_h_l_07[23:0]),
     .prog(prog), .spi_ss_in_b({net629[0], net629[1]}),
     .tnl_op(lft_op_08[7:0]), .lft_op(lft_op_07[7:0]),
     .bnl_op(lft_op_06[7:0]), .pgate(pgate[111:96]),
     .reset(reset_b[111:96]), .sp4_v_b({net442[0], net442[1],
     net442[2], net442[3], net442[4], net442[5], net442[6], net442[7],
     net442[8], net442[9], net442[10], net442[11], net442[12],
     net442[13], net442[14], net442[15]}), .wl(wl[111:96]),
     .cf(cf_r[167:144]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_07[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net388));
io_col4_rgt_ice8p_v2 I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net391), .sdi(net571), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[20:19]), .pado(pado[20:19]),
     .padeb(padeb[20:19]), .sp4_v_t({net406[0], net406[1], net406[2],
     net406[3], net406[4], net406[5], net406[6], net406[7], net406[8],
     net406[9], net406[10], net406[11], net406[12], net406[13],
     net406[14], net406[15]}), .sp4_h_l(SP4_h_l_05[47:0]),
     .sp12_h_l(SP12_h_l_05[23:0]), .prog(prog),
     .spi_ss_in_b({net618[0], net618[1]}), .tnl_op(lft_op_06[7:0]),
     .lft_op(lft_op_05[7:0]), .bnl_op(lft_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]), .sp4_v_b({net586[0],
     net586[1], net586[2], net586[3], net586[4], net586[5], net586[6],
     net586[7], net586[8], net586[9], net586[10], net586[11],
     net586[12], net586[13], net586[14], net586[15]}), .wl(wl[79:64]),
     .cf(cf_r[119:96]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net424));
io_col4_rgt_ice8p_v2 I_io_00_06 ( .cbit_colcntl({net633[0], net633[1],
     net633[2], net633[3], net633[4], net633[5], net633[6],
     net633[7]}), .ceb(ceb), .sdo(net427), .sdi(net391),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[22:21]), .pado(pado[22:21]), .padeb(padeb[22:21]),
     .sp4_v_t({net442[0], net442[1], net442[2], net442[3], net442[4],
     net442[5], net442[6], net442[7], net442[8], net442[9], net442[10],
     net442[11], net442[12], net442[13], net442[14], net442[15]}),
     .sp4_h_l(SP4_h_l_06[47:0]), .sp12_h_l(SP12_h_l_06[23:0]),
     .prog(prog), .spi_ss_in_b({net625[0], net625[1]}),
     .tnl_op(lft_op_07[7:0]), .lft_op(lft_op_06[7:0]),
     .bnl_op(lft_op_05[7:0]), .pgate(pgate[95:80]),
     .reset(reset_b[95:80]), .sp4_v_b({net406[0], net406[1], net406[2],
     net406[3], net406[4], net406[5], net406[6], net406[7], net406[8],
     net406[9], net406[10], net406[11], net406[12], net406[13],
     net406[14], net406[15]}), .wl(wl[95:80]), .cf(cf_r[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(net460));
io_col4_rgt_ice8p_v2 I_io_00_02 ( .cbit_colcntl({net461[0], net461[1],
     net461[2], net461[3], net461[4], net461[5], net461[6],
     net461[7]}), .ceb(ceb), .sdo(net463), .sdi(net499),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin({net476[0],
     net476[1]}), .pado({net476[0], net476[1]}), .padeb({net477[0],
     net477[1]}), .sp4_v_t({net478[0], net478[1], net478[2], net478[3],
     net478[4], net478[5], net478[6], net478[7], net478[8], net478[9],
     net478[10], net478[11], net478[12], net478[13], net478[14],
     net478[15]}), .sp4_h_l(SP4_h_l_02[47:0]),
     .sp12_h_l(SP12_h_l_02[23:0]), .prog(prog),
     .spi_ss_in_b({net630[0], net630[1]}), .tnl_op(lft_op_03[7:0]),
     .lft_op(lft_op_02[7:0]), .bnl_op(lft_op_01[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]), .sp4_v_b({net514[0],
     net514[1], net514[2], net514[3], net514[4], net514[5], net514[6],
     net514[7], net514[8], net514[9], net514[10], net514[11],
     net514[12], net514[13], net514[14], net514[15]}), .wl(wl[31:16]),
     .cf(cf_r[47:24]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fabric_out_10));
io_col4_rgt_ice8p_v2 I_io_00_01 ( .cbit_colcntl({net497[0], net497[1],
     net497[2], net497[3], net497[4], net497[5], net497[6],
     net497[7]}), .ceb(ceb), .sdo(net499), .sdi(sdi), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin(padin[14:13]),
     .pado(pado[14:13]), .padeb(padeb[14:13]), .sp4_v_t({net514[0],
     net514[1], net514[2], net514[3], net514[4], net514[5], net514[6],
     net514[7], net514[8], net514[9], net514[10], net514[11],
     net514[12], net514[13], net514[14], net514[15]}),
     .sp4_h_l(SP4_h_l_01[47:0]), .sp12_h_l(SP12_h_l_01[23:0]),
     .prog(prog), .spi_ss_in_b({net620[0], net620[1]}),
     .tnl_op(lft_op_02[7:0]), .lft_op(lft_op_01[7:0]),
     .bnl_op(bnl_op_13_09[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_13_09[15:0]),
     .wl(wl[15:0]), .cf(cf_r[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_09));
io_col4_rgt_ice8p_v2 I_io_00_03 ( .cbit_colcntl({net623[0], net623[1],
     net623[2], net623[3], net623[4], net623[5], net623[6],
     net623[7]}), .ceb(ceb), .sdo(net535), .sdi(net463),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[16:15]), .pado(pado[16:15]), .padeb(padeb[16:15]),
     .sp4_v_t({net550[0], net550[1], net550[2], net550[3], net550[4],
     net550[5], net550[6], net550[7], net550[8], net550[9], net550[10],
     net550[11], net550[12], net550[13], net550[14], net550[15]}),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b({net624[0], net624[1]}),
     .tnl_op(lft_op_04[7:0]), .lft_op(lft_op_03[7:0]),
     .bnl_op(lft_op_02[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b({net478[0], net478[1], net478[2],
     net478[3], net478[4], net478[5], net478[6], net478[7], net478[8],
     net478[9], net478[10], net478[11], net478[12], net478[13],
     net478[14], net478[15]}), .wl(wl[47:32]), .cf(cf_r[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net568));
io_col4_rgt_ice8p_v2 I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net571), .sdi(net535), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[18:17]), .pado(pado[18:17]),
     .padeb(padeb[18:17]), .sp4_v_t({net586[0], net586[1], net586[2],
     net586[3], net586[4], net586[5], net586[6], net586[7], net586[8],
     net586[9], net586[10], net586[11], net586[12], net586[13],
     net586[14], net586[15]}), .sp4_h_l(SP4_h_l_04[47:0]),
     .sp12_h_l(SP12_h_l_04[23:0]), .prog(prog),
     .spi_ss_in_b({net590[0], net590[1]}), .tnl_op(lft_op_05[7:0]),
     .lft_op(lft_op_04[7:0]), .bnl_op(lft_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]), .sp4_v_b({net550[0],
     net550[1], net550[2], net550[3], net550[4], net550[5], net550[6],
     net550[7], net550[8], net550[9], net550[10], net550[11],
     net550[12], net550[13], net550[14], net550[15]}), .wl(wl[63:48]),
     .cf(cf_r[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net604));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - bram_bufferx4x6, View - schematic
// LAST TIME SAVED: Sep 15 13:53:57 2008
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_bufferx4x6 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I4 ( .in(d1), .out(d2));
bram_bufferx4 I5 ( .in(d2), .out(d3));
bram_bufferx4 I6 ( .in(d3), .out(d4));
bram_bufferx4 I7 ( .in(d4), .out(out));
bram_bufferx4 I3 ( .in(d0), .out(d1));
bram_bufferx4 I0 ( .in(in), .out(d0));

endmodule
// Library - leafcell, Cell - pllphase_sr_40lp, View - schematic
// LAST TIME SAVED: Apr 20 09:43:38 2011
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pllphase_sr_40lp ( f_dvd2, f_dvd4_p0, f_dvd4_p90, f_out, CLK,
     cbit, sr, tiehi, tielo );
output  f_dvd2, f_dvd4_p0, f_dvd4_p90, f_out;

input  CLK, cbit, sr, tiehi, tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  qn;



mux2_hvt I_MUX4DIV7 ( .in1(net077), .in0(net051), .out(net038),
     .sel(cbit));
inv_tri_2_hvt I21 ( .Tb(net0136), .T(net0136), .A(net0136),
     .Y(net0113));
nor2_hvt I22 ( .A(net0113), .B(tielo), .Y(net0116));
inv_hvt I26 ( .A(net089), .Y(net086));
inv_hvt I27 ( .A(CLK), .Y(net089));
inv_hvt I23 ( .A(net0116), .Y(net044));
inv_hvt I20 ( .A(net0138), .Y(net0136));
inv_hvt I19 ( .A(net080), .Y(net0138));
inv_hvt I28 ( .A(net086), .Y(net057));
inv_hvt I29 ( .A(net057), .Y(net080));
inv_hvt I8 ( .A(qn[1]), .Y(f_dvd4_p90));
inv_hvt I7 ( .A(net0100), .Y(f_dvd2));
inv_hvt I6 ( .A(net044), .Y(f_out));
inv_hvt I5 ( .A(qn[0]), .Y(f_dvd4_p0));
pll_ml_dff I2 ( .R(sr), .D(net056), .CLK(CLK), .QN(qn[1]), .Q(net051));
pll_ml_dff I0 ( .R(sr), .D(net054), .CLK(CLK), .QN(qn[0]), .Q(net056));
pll_ml_dff I3 ( .R(sr), .D(net051), .CLK(CLK), .QN(net061),
     .Q(net040));
pll_ml_dff I12 ( .R(sr), .D(net0100), .CLK(CLK), .QN(net0100),
     .Q(net067));
dffs I10 ( .D(net082), .QN(net071), .Q(net054), .CLK(CLK), .S(sr));
dffs I9 ( .D(net053), .QN(net076), .Q(net077), .CLK(CLK), .S(sr));
dffs I11 ( .D(net038), .QN(net081), .Q(net082), .CLK(CLK), .S(sr));
dffs I4 ( .D(net040), .CLK(CLK), .QN(net087), .Q(net053), .S(sr));

endmodule
// Library - leafcell, Cell - lowla_modified, View - schematic
// LAST TIME SAVED: Aug 12 09:10:07 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module lowla_modified ( lao, clk, min );
output  lao;

input  clk, min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I249 ( .in(lao), .out(st2), .pp(cbitb), .nn(clkd));
txgate_hvt I248 ( .in(min), .out(st2), .pp(clkd), .nn(cbitb));
inv_hvt I289 ( .A(net29), .Y(lao));
inv_hvt I290 ( .A(st2), .Y(net29));
inv_hvt I_inv ( .A(clk), .Y(cbitb));
inv_hvt I_inv3 ( .A(cbitb), .Y(clkd));

endmodule
// Library - ice8chip, Cell - scan_buf_ice8p, View - schematic
// LAST TIME SAVED: Jun 28 09:23:39 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module scan_buf_ice8p ( bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo,
     shift_o, tclk_o, update_o, bs_en_i, ceb_i, hiz_b_i, mode_i, r_i,
     sdi, shift_i, tclk_i, update_i );
output  bs_en_o, ceb_o, hiz_b_o, mode_o, r_o, sdo, shift_o, tclk_o,
     update_o;

input  bs_en_i, ceb_i, hiz_b_i, mode_i, r_i, sdi, shift_i, tclk_i,
     update_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



tckbufx32_ice8p I_tclkbuf ( .in(tclk_i), .out(tclk_o));
bram_bufferx4 I_bs_enbuf ( .in(bs_en_i), .out(bs_en_o));
bram_bufferx4 I_cebbuf ( .in(ceb_i), .out(ceb_o));
bram_bufferx4 I_modebuf ( .in(mode_i), .out(mode_o));
bram_bufferx4 I_hiz_bbuf ( .in(hiz_b_i), .out(hiz_b_o));
bram_bufferx4 I_updatebuf ( .in(update_i), .out(update_o));
bram_bufferx4 I_shiftbuf ( .in(shift_i), .out(shift_o));
bram_bufferx4 I_rbuf ( .in(r_i), .out(r_o));
bram_bufferx4x6 I_sdibuf ( .in(sdi), .out(sdi_2));
lowla_modified I_lowla ( .clk(tclk_i), .min(sdi_2), .lao(sdo));

endmodule
// Library - io, Cell - ioinmx1mux2_imp, View - schematic
// LAST TIME SAVED: Aug 13 14:11:56 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioinmx1mux2_imp ( clk, mo, ti, bl, cdone_in, ce, ceb, in, min,
     pgate, prog, reset, spi, vdd_cntl, wl );
output  clk, ti;


input  cdone_in, ceb, prog;

output [1:0]  mo;

inout [5:0]  bl;

input [1:0]  spi;
input [11:0]  ce;
input [1:0]  in;
input [7:0]  min;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  moo;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  mob;

wire  [1:0]  r_vdd;



mux2x1_hvt I_emux_1_ ( .in1(in[1]), .in0(spi[1]), .out(moo[1]),
     .sel(cdone_in));
mux2x1_hvt I_emux_0_ ( .in1(in[0]), .in0(spi[0]), .out(moo[0]),
     .sel(cdone_in));
inv_lvt inv_1_1_ ( .A(moo[1]), .Y(mob[1]));
inv_lvt inv_1_0_ ( .A(moo[0]), .Y(mob[0]));
inv_lvt I_inv_2_1_ ( .A(mob[1]), .Y(mo[1]));
inv_lvt I_inv_2_0_ ( .A(mob[0]), .Y(mo[0]));
ioin_mux_v2 I_ioin_mux ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clk_mux12to1 I_clk_mux12to1 ( .prog(prog), .min(ce[11:0]), .clk(clk),
     .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7], cbitb[10],
     cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7], cbit[10],
     cbit[6], cbit[4]}), .cenb(ceb));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc, View - schematic
// LAST TIME SAVED: Aug 12 13:51:42 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  spi;
output [1:0]  ti;

inout [5:0]  bl;

input [7:0]  min1;
input [7:0]  min0;
input [1:0]  padin;
input [1:0]  pgate;
input [7:0]  min2;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



inv_lvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_lvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
nor2_lvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_lvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
ioin_mux_v2 I_ioin_mux_bankcntl ( bankcntl, {cbit[11], cbit[8], cbit[9],
     cbit[10]}, {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0],
     prog);
ioin_mux_v2 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v2 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nand2inv, View - schematic
// LAST TIME SAVED: Oct  8 16:13:18 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioinmx2nand2inv ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [7:0]  min0;
input [7:0]  ce;
input [1:0]  reset;
input [1:0]  wl;
input [7:0]  min1;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



nand2_lvt I180 ( .A(update_b), .Y(updt), .B(bs_en));
inv_lvt I181 ( .A(update), .Y(update_b));
ioin_mux_v2 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v2 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc_v3, View - schematic
// LAST TIME SAVED: May 12 17:30:59 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module sbox1_colbdlc_v3 ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  spi_ss_in_b;
output [1:0]  padeb;
output [5:0]  ti;
output [1:0]  pado;

inout [5:0]  bl;
inout [3:0]  t_mid;
inout [3:0]  sp4_v_b;
inout [3:0]  l;
inout [3:0]  r;

input [1:0]  out;
input [1:0]  padin;
input [11:0]  clk_in;
input [7:0]  min5;
input [1:0]  spiout;
input [7:0]  ceb_in;
input [7:0]  min4;
input [11:0]  inclk_in;
input [7:0]  min2;
input [1:0]  oeb;
input [7:0]  min1;
input [1:0]  spioeb;
input [7:0]  min3;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  min0;
input [7:0]  min6;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ioinmx1mux2_imp I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .in(out[1:0]), .ti(ti[2]), .min(min2[7:0]), .spi(spiout[1:0]),
     .wl(wl[9:8]), .reset(reset[9:8]), .pgate(pgate[9:8]),
     .cdone_in(cdone_in), .mo(pado[1:0]));
ioinmx1mux2_imp I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .in(oeb[1:0]), .ti(ti[5]), .min(min5[7:0]), .spi(spioeb[1:0]),
     .wl(wl[15:14]), .reset(reset[15:14]), .pgate(pgate[15:14]),
     .cdone_in(cdone_in), .mo(padeb[1:0]));
ioinmx2nor2invx2bdlc I5 ( .vdd_cntl(vdd_cntl[5:4]), .min2(min6[7:0]),
     .bankcntl(fabric_out), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx2nand2inv I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - io, Cell - io_gmux_x2v2, View - schematic
// LAST TIME SAVED: Jun  1 11:08:17 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_gmux_x2v2 ( .cbitb_colcntl({cbitb[11], cbitb[9]}), gout, bl,
     min0, min1, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [1:0]  gout;
output [11:0]  cbitb;

inout [5:0]  bl;

input [15:0]  min0;
input [1:0]  vdd_cntl;
input [15:0]  min1;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux I_g_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux I_g_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare_v3, View - schematic
// LAST TIME SAVED: Jun  2 10:52:40 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_gmux_x16bare_v3 ( cbitb_colcntl, lc_trk_g0, lc_trk_g1, bl,
     min0, min1, min2, min3, min4, min5, min6, min7, min8, min9, min10,
     min11, min12, min13, min14, min15, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  cbitb_colcntl;

inout [5:0]  bl;

input [15:0]  min7;
input [15:0]  min0;
input [15:0]  min9;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min15;
input [15:0]  min3;
input [15:0]  min14;
input [15:0]  min12;
input [15:0]  min6;
input [15:0]  min8;
input [15:0]  min5;
input [15:0]  min4;
input [15:0]  min11;
input [15:0]  min10;
input [15:0]  vdd_cntl;
input [15:0]  min2;
input [15:0]  reset;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net114;

wire  [1:0]  net187;

wire  [1:0]  net188;

wire  [1:0]  net124;



io_gmux_x2v2 I_io_gmux_x2_7 ( .cbitb_colcntl({net114[0], net114[1]}),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[15:14]));
io_gmux_x2v2 I_io_gmux_x2_6 ( .cbitb_colcntl({net124[0], net124[1]}),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[13:12]));
io_gmux_x2v2 I_io_gmux_x2_2 ( .cbitb_colcntl(cbitb_colcntl[5:4]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[5:4]));
io_gmux_x2v2 I_io_gmux_x2_0 ( .cbitb_colcntl(cbitb_colcntl[1:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[1:0]));
io_gmux_x2v2 _io_gmux_x2_1 ( .cbitb_colcntl(cbitb_colcntl[3:2]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[3:2]));
io_gmux_x2v2 I_io_gmux_x2_4 ( .cbitb_colcntl({net187[0], net187[1]}),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[9:8]));
io_gmux_x2v2 I_io_gmux_x2_5 ( .cbitb_colcntl({net188[0], net188[1]}),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[11:10]));
io_gmux_x2v2 I_io_gmux_x2_3 ( .cbitb_colcntl(cbitb_colcntl[7:6]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[7:6]));

endmodule
// Library - ice8chip, Cell - io_col4_top_ice8p, View - schematic
// LAST TIME SAVED: Jan 12 15:49:45 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_col4_top_ice8p ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  padeb;
output [1:0]  pado;
output [23:0]  cf;
output [3:0]  slf_op;
output [1:0]  spi_ss_in_b;

inout [15:0]  sp4_v_t;
inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [15:0]  sp4_v_b;
inout [47:0]  sp4_h_l;

input [1:0]  spioeb;
input [15:0]  wl;
input [7:0]  lft_op;
input [15:0]  reset;
input [1:0]  spiout;
input [15:0]  vdd_cntl;
input [7:0]  bnl_op;
input [15:0]  pgate;
input [7:0]  tnl_op;
input [1:0]  padin;
input [7:0]  glb_netwk;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  ti;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  om;

wire  [1:0]  oenm;

wire  [7:0]  net0100;



rm6w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
sbox1_colbdlc_v3 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
io_gmux_x16bare_v3 I_io_gmux_x16bare_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .cbitb_colcntl({net0100[0], net0100[1], net0100[2], net0100[3],
     net0100[4], net0100[5], net0100[6], net0100[7]}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));

endmodule
// Library - ice1chip, Cell - io_top_rgt_1x6_ice1f, View - schematic
// LAST TIME SAVED: Mar  8 10:17:00 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_top_rgt_1x6_ice1f ( bs_en_o, ceb_o, cf_t, fabric_out_07_17,
     fabric_out_08_17, hiz_b_o, mode_o, padeb_t_r, pado_t_r, r_o, sdo,
     shift_o, slf_op_01_17, slf_op_02_17, slf_op_03_17, slf_op_04_17,
     slf_op_05_17, slf_op_06_17, tclk_o, update_o, bl_01, bl_02, bl_03,
     bl_04, bl_05, bl_06, sp4_h_l_07_17, sp4_h_r_12_17, sp4_v_b_01_17,
     sp4_v_b_02_17, sp4_v_b_03_17, sp4_v_b_04_17, sp4_v_b_05_17,
     sp4_v_b_06_17, sp12_v_b_01_17, sp12_v_b_02_17, sp12_v_b_03_17,
     sp12_v_b_04_17, sp12_v_b_05_17, sp12_v_b_06_17, bnl_op_07_17,
     bnr_op_12_17, bs_en_i, ceb_i, glb_net_01, glb_net_02, glb_net_03,
     glb_net_04, glb_net_05, glb_net_06, hiz_b_i, hold_t_r,
     lft_op_01_17, lft_op_02_17, lft_op_03_17, lft_op_04_17,
     lft_op_05_17, lft_op_06_17, mode_i, padin_t_r, pgate_l, prog, r_i,
     reset_l, sdi, shift_i, tclk_i, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_07_17, fabric_out_08_17, hiz_b_o,
     mode_o, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_r, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_02_17;
output [3:0]  slf_op_06_17;
output [3:0]  slf_op_03_17;
output [143:0]  cf_t;
output [23:12]  padeb_t_r;
output [23:12]  pado_t_r;
output [3:0]  slf_op_04_17;
output [3:0]  slf_op_01_17;
output [3:0]  slf_op_05_17;

inout [47:0]  sp4_v_b_06_17;
inout [23:0]  sp12_v_b_06_17;
inout [23:0]  sp12_v_b_05_17;
inout [47:0]  sp4_v_b_05_17;
inout [47:0]  sp4_v_b_03_17;
inout [47:0]  sp4_v_b_01_17;
inout [23:0]  sp12_v_b_03_17;
inout [47:0]  sp4_v_b_02_17;
inout [47:0]  sp4_v_b_04_17;
inout [15:0]  sp4_h_l_07_17;
inout [23:0]  sp12_v_b_04_17;
inout [53:0]  bl_05;
inout [53:0]  bl_06;
inout [23:0]  sp12_v_b_02_17;
inout [41:0]  bl_04;
inout [53:0]  bl_03;
inout [15:0]  sp4_h_r_12_17;
inout [53:0]  bl_02;
inout [53:0]  bl_01;
inout [23:0]  sp12_v_b_01_17;

input [7:0]  bnr_op_12_17;
input [7:0]  glb_net_03;
input [7:0]  glb_net_01;
input [7:0]  lft_op_05_17;
input [7:0]  bnl_op_07_17;
input [7:0]  lft_op_03_17;
input [7:0]  lft_op_04_17;
input [7:0]  glb_net_06;
input [7:0]  lft_op_06_17;
input [7:0]  glb_net_02;
input [7:0]  glb_net_04;
input [23:12]  padin_t_r;
input [7:0]  lft_op_01_17;
input [15:0]  reset_l;
input [15:0]  wl_l;
input [7:0]  lft_op_02_17;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_05;
input [15:0]  pgate_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  net433;

wire  [1:0]  net472;

wire  [15:0]  net363;

wire  [1:0]  net290;

wire  [15:0]  net503;

wire  [1:0]  net507;

wire  [15:0]  net328;

wire  [15:0]  net398;

wire  [1:0]  net402;

wire  [1:0]  net332;

wire  [1:0]  net289;



tckbufx32_ice8p I_tck_halfbankcenter ( .in(net273), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));
scan_buf_ice8p I345 ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net273), .shift_o(shift_o),
     .sdo(net453), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_top_ice8p I_IO_08_17 ( .sdo(net383), .sdi(net313),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net398[0], net398[1], net398[2], net398[3],
     net398[4], net398[5], net398[6], net398[7], net398[8], net398[9],
     net398[10], net398[11], net398[12], net398[13], net398[14],
     net398[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_r[15:14]), .pado(pado_t_r[15:14]),
     .padeb(padeb_t_r[15:14]), .sp4_v_b({net328[0], net328[1],
     net328[2], net328[3], net328[4], net328[5], net328[6], net328[7],
     net328[8], net328[9], net328[10], net328[11], net328[12],
     net328[13], net328[14], net328[15]}),
     .sp4_h_l(sp4_v_b_02_17[47:0]), .sp12_h_l(sp12_v_b_02_17[23:0]),
     .prog(prog), .spi_ss_in_b({net332[0], net332[1]}),
     .tnl_op(lft_op_01_17[7:0]), .lft_op(lft_op_02_17[7:0]),
     .bnl_op(lft_op_03_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_t[47:24]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_17[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_t_r), .fabric_out(fabric_out_08_17));
io_col4_top_ice8p I_IO_10_17_bram ( .sdo(net488), .sdi(net348),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net503[0], net503[1], net503[2], net503[3],
     net503[4], net503[5], net503[6], net503[7], net503[8], net503[9],
     net503[10], net503[11], net503[12], net503[13], net503[14],
     net503[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_r[19:18]), .pado(pado_t_r[19:18]),
     .padeb(padeb_t_r[19:18]), .sp4_v_b({net363[0], net363[1],
     net363[2], net363[3], net363[4], net363[5], net363[6], net363[7],
     net363[8], net363[9], net363[10], net363[11], net363[12],
     net363[13], net363[14], net363[15]}),
     .sp4_h_l(sp4_v_b_04_17[47:0]), .sp12_h_l(sp12_v_b_04_17[23:0]),
     .prog(prog), .spi_ss_in_b({net289[0], net289[1]}),
     .tnl_op(lft_op_03_17[7:0]), .lft_op(lft_op_04_17[7:0]),
     .bnl_op(lft_op_05_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf(cf_t[71:48]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_17[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_t_r), .fabric_out(net381));
io_col4_top_ice8p I_IO_07_17 ( .sdo(sdo), .sdi(net383),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_07_17[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_r[13:12]),
     .pado(pado_t_r[13:12]), .padeb(padeb_t_r[13:12]),
     .sp4_v_b({net398[0], net398[1], net398[2], net398[3], net398[4],
     net398[5], net398[6], net398[7], net398[8], net398[9], net398[10],
     net398[11], net398[12], net398[13], net398[14], net398[15]}),
     .sp4_h_l(sp4_v_b_01_17[47:0]), .sp12_h_l(sp12_v_b_01_17[23:0]),
     .prog(prog), .spi_ss_in_b({net402[0], net402[1]}),
     .tnl_op(bnl_op_07_17[7:0]), .lft_op(lft_op_01_17[7:0]),
     .bnl_op(lft_op_02_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_t[23:0]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_17[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_t_r), .fabric_out(fabric_out_07_17));
io_col4_top_ice8p I_IO_11_17 ( .sdo(net348), .sdi(net418),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net363[0], net363[1], net363[2], net363[3],
     net363[4], net363[5], net363[6], net363[7], net363[8], net363[9],
     net363[10], net363[11], net363[12], net363[13], net363[14],
     net363[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_r[21:20]), .pado(pado_t_r[21:20]),
     .padeb(padeb_t_r[21:20]), .sp4_v_b({net433[0], net433[1],
     net433[2], net433[3], net433[4], net433[5], net433[6], net433[7],
     net433[8], net433[9], net433[10], net433[11], net433[12],
     net433[13], net433[14], net433[15]}),
     .sp4_h_l(sp4_v_b_05_17[47:0]), .sp12_h_l(sp12_v_b_05_17[23:0]),
     .prog(prog), .spi_ss_in_b({net290[0], net290[1]}),
     .tnl_op(lft_op_04_17[7:0]), .lft_op(lft_op_05_17[7:0]),
     .bnl_op(lft_op_06_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf(cf_t[119:96]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_17[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_t_r), .fabric_out(net451));
io_col4_top_ice8p I_IO_12_17 ( .sdo(net418), .sdi(net453),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net433[0], net433[1], net433[2], net433[3],
     net433[4], net433[5], net433[6], net433[7], net433[8], net433[9],
     net433[10], net433[11], net433[12], net433[13], net433[14],
     net433[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_r[23:22]), .pado(pado_t_r[23:22]),
     .padeb(padeb_t_r[23:22]), .sp4_v_b(sp4_h_r_12_17[15:0]),
     .sp4_h_l(sp4_v_b_06_17[47:0]), .sp12_h_l(sp12_v_b_06_17[23:0]),
     .prog(prog), .spi_ss_in_b({net472[0], net472[1]}),
     .tnl_op(lft_op_05_17[7:0]), .lft_op(lft_op_06_17[7:0]),
     .bnl_op(bnr_op_12_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_06[5], bl_06[4], bl_06[37],
     bl_06[36], bl_06[35], bl_06[34], bl_06[33], bl_06[32], bl_06[14],
     bl_06[20], bl_06[19], bl_06[18], bl_06[17], bl_06[16], bl_06[27],
     bl_06[26], bl_06[25], bl_06[23]}), .wl(wl_l[15:0]),
     .cf(cf_t[143:120]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_17[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_t_r), .fabric_out(net486));
io_col4_top_ice8p I_IO_09_17 ( .sdo(net313), .sdi(net488),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net328[0], net328[1], net328[2], net328[3],
     net328[4], net328[5], net328[6], net328[7], net328[8], net328[9],
     net328[10], net328[11], net328[12], net328[13], net328[14],
     net328[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_r[17:16]), .pado(pado_t_r[17:16]),
     .padeb(padeb_t_r[17:16]), .sp4_v_b({net503[0], net503[1],
     net503[2], net503[3], net503[4], net503[5], net503[6], net503[7],
     net503[8], net503[9], net503[10], net503[11], net503[12],
     net503[13], net503[14], net503[15]}),
     .sp4_h_l(sp4_v_b_03_17[47:0]), .sp12_h_l(sp12_v_b_03_17[23:0]),
     .prog(prog), .spi_ss_in_b({net507[0], net507[1]}),
     .tnl_op(lft_op_02_17[7:0]), .lft_op(lft_op_03_17[7:0]),
     .bnl_op(lft_op_04_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_t[95:72]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_17[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_t_r), .fabric_out(net521));

endmodule
// Library - leafcell, Cell - clkmux2buffer, View - schematic
// LAST TIME SAVED: Jun 29 15:54:22 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module clkmux2buffer ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate Itg20 ( .in(in1), .out(net16), .pp(net10), .nn(sel));
txgate I31 ( .in(in0), .out(net16), .pp(sel), .nn(net10));
inv I_inv1 ( .A(net16), .Y(outb));
inv I_inv2 ( .A(outb), .Y(out));
inv I1 ( .A(sel), .Y(net10));

endmodule
// Library - ice8chip, Cell - clk_quad_buf_ice8p, View - schematic
// LAST TIME SAVED: Aug 12 09:03:48 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module clk_quad_buf_ice8p ( clko, clki );
output  clko;

input  clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I19 ( .A(clkb), .Y(clko));
inv_lvt I22 ( .A(clki), .Y(clkb));

endmodule
// Library - ice8chip, Cell - clk_quad_buf_x8_ice8p, View - schematic
// LAST TIME SAVED: Jun 24 14:46:09 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module clk_quad_buf_x8_ice8p ( clko, clki );


output [7:0]  clko;

input [7:0]  clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_quad_buf_ice8p I_clk_quad_buf_ice8p_7_ ( .clki(clki[7]),
     .clko(clko[7]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_6_ ( .clki(clki[6]),
     .clko(clko[6]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_5_ ( .clki(clki[5]),
     .clko(clko[5]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_4_ ( .clki(clki[4]),
     .clko(clko[4]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_3_ ( .clki(clki[3]),
     .clko(clko[3]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_2_ ( .clki(clki[2]),
     .clko(clko[2]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_1_ ( .clki(clki[1]),
     .clko(clko[1]));
clk_quad_buf_ice8p I_clk_quad_buf_ice8p_0_ ( .clki(clki[0]),
     .clko(clko[0]));

endmodule
// Library - xpmem, Cell - cram_2x28, View - schematic
// LAST TIME SAVED: Jun 24 18:02:26 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module cram_2x28 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [55:0]  q;
output [55:0]  q_b;

inout [27:0]  bl;

input [1:0]  r_vdd;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 I_mstake_13_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[27:26]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[1:0]));
cram2x2 I_mstake_12_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[25:24]), .q_b(q_b[51:48]),
     .q(q[51:48]), .wl(wl[1:0]));
cram2x2 I_mstake_11_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[23:22]), .q_b(q_b[47:44]),
     .q(q[47:44]), .wl(wl[1:0]));
cram2x2 I_mstake_10_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[21:20]), .q_b(q_b[43:40]),
     .q(q[43:40]), .wl(wl[1:0]));
cram2x2 I_mstake_9_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[19:18]), .q_b(q_b[39:36]),
     .q(q[39:36]), .wl(wl[1:0]));
cram2x2 I_mstake_8_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[17:16]), .q_b(q_b[35:32]),
     .q(q[35:32]), .wl(wl[1:0]));
cram2x2 I_mstake_7_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[15:14]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[1:0]));
cram2x2 I_mstake_6_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[13:12]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[1:0]));
cram2x2 I_mstake_5_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 I_mstake_4_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 I_mstake_3_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 I_mstake_2_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 I_mstake_1_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 I_mstake_0_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - logic_cell_rev, View - schematic
// LAST TIME SAVED: Sep  3 10:41:29 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module logic_cell_rev ( carry_out, out, out_vic, carry_in, cbit, clk,
     clkb, in0, in1, in2, in3, prog, purst, s_r );
output  carry_out, out, out_vic;

input  carry_in, clk, clkb, in0, in1, in2, in3, prog, purst, s_r;

input [20:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clut4vic I_clut4 ( .lut4vic(out_vic), .in3b(in3b), .in3(in3),
     .in2b(in2b), .in2(in2), .in1b(in1b), .in1(in1), .in0b(in0b),
     .in0(in0), .cbit(cbit[15:0]), .lut4(LUT4_outd));
o_mux I_o_mux ( .prog(prog), .in1(rego), .in0(LUT4_outd),
     .cbit(cbit[19]), .out(out));
inv_lvt I196 ( .A(in3), .Y(in3b));
inv_lvt I189 ( .A(in0), .Y(in0b));
inv_lvt I194 ( .A(in1), .Y(in1b));
inv_lvt I195 ( .A(in2), .Y(in2b));
carry_logic_nand I_carry_logic ( .vg_en(cbit[20]), .carry_in(carry_in),
     .b_bar(in1b), .b(in1), .a_bar(in2b), .a(in2), .cout(carry_out));
coredffr I_coredffr ( .purst(purst), .d(LUT4_outd), .clkb(clkb),
     .clk(clk), .cbit(cbit[17:16]), .S_R(s_r), .q(rego));

endmodule
// Library - leafcell, Cell - lcmuxod3_0_0, View - schematic
// LAST TIME SAVED: Oct 18 13:59:54 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module lcmuxod3_0_0 ( carry_out, cbit, cbitb, op, op_vic, sp4_h_r,
     sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb,
     min0, min1, min2, min3, op_bot, pgate, prog, purst, reset_b, s_r,
     vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_h_r;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [2:0]  sp4_r_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_h_r;
output [55:0]  cbit;
output [55:0]  cbitb;
output [2:0]  sp4_v_b;

input [1:0]  wl;
input [27:0]  bl;
input [15:0]  min0;
input [1:0]  pgate;
input [15:0]  min1;
input [1:0]  vdd_cntl;
input [15:0]  min3;
input [15:0]  min2;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



in_mux_nand I_in2mux_nand ( .cbitb({cbitb[50], cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50], cbit[12],
     cbit[13], cbit[16], cbit[19], cbit[17]}), .op_bot(op_bot),
     .prog(prog), .inmuxo(in2), .min(min2[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_30 I_odrv30 ( .slfop(op), .prog(prog),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53], cbitb[55],
     cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44], cbitb[46],
     cbitb[43], cbitb[41], cbitb[42], cbitb[40]}), .sp12_h_r(sp12_h_r),
     .sp12_v_b(sp12_v_b[1:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
in_mux I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));

endmodule
// Library - leafcell, Cell - lcmuxod3_0, View - schematic
// LAST TIME SAVED: Jun 24 18:04:48 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module lcmuxod3_0 ( carry_out, op, op_vic, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, op_bot, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_h_r;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;

input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [15:0]  min2;
input [27:0]  bl;
input [15:0]  min1;
input [1:0]  pgate;
input [15:0]  min3;
input [1:0]  wl;
input [15:0]  min0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [1:0]  r_vdd;

wire  [55:0]  cbitb;



in_mux_nand I_in2mux_nand ( .cbitb({cbitb[50], cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50], cbit[12],
     cbit[13], cbit[16], cbit[19], cbit[17]}), .op_bot(op_bot),
     .prog(prog), .inmuxo(in2), .min(min2[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_30 I_odrv30 ( .slfop(op), .prog(prog),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53], cbitb[55],
     cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44], cbitb[46],
     cbitb[43], cbitb[41], cbitb[42], cbitb[40]}), .sp12_h_r(sp12_h_r),
     .sp12_v_b(sp12_v_b[1:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
in_mux I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));

endmodule
// Library - leafcell, Cell - lcmuxod7_4, View - schematic
// LAST TIME SAVED: Jun 24 18:10:24 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module lcmuxod7_4 ( carry_out, op, op_vic, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, op_bot, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, op_vic, sp12_v_b;

input  carry_in, clk, clkb, op_bot, prog, purst, s_r;

output [2:0]  sp4_v_b;
output [2:0]  sp4_r_v_b;
output [1:0]  sp12_h_r;
output [2:0]  sp4_h_r;

input [15:0]  min0;
input [15:0]  min3;
input [1:0]  vdd_cntl;
input [15:0]  min2;
input [15:0]  min1;
input [1:0]  reset_b;
input [27:0]  bl;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



in_mux_nand I_in2mux ( .cbitb({cbitb[50], cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .cbit({cbit[50], cbit[12],
     cbit[13], cbit[16], cbit[19], cbit[17]}), .op_bot(op_bot),
     .prog(prog), .inmuxo(in2), .min(min2[15:0]));
cram_2x28 I_cram_2x28 ( .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]), .reset(reset_b[1:0]),
     .q_b(cbitb[55:0]));
odrv12_74 I_odrv74 ( .slfop(op), .prog(prog), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));
in_mux I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
in_mux I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
logic_cell_rev I_LC ( .out_vic(op_vic), .carry_in(carry_in), .in1(in1),
     .in3(in3), .clk(clk), .out(op), .carry_out(carry_out), .in2(in2),
     .clkb(clkb), .prog(prog), .purst(purst), .in0(in0), .s_r(s_r),
     .cbit({cbit[38], cbit[39], cbit[39], cbit[37], cbit[36], cbit[22],
     cbit[20], cbit[21], cbit[23], cbit[26], cbit[24], cbit[25],
     cbit[27], cbit[35], cbit[33], cbit[32], cbit[34], cbit[31],
     cbit[29], cbit[28], cbit[30]}));

endmodule
// Library - leafcell, Cell - lccol_rev0, View - schematic
// LAST TIME SAVED: Oct 18 13:49:45 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module lccol_rev0 ( carry_out, op_vic, slf_op, bl, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, cin2local, clk, clkb, lc_trk_g0,
     lc_trk_g1, lc_trk_g2, lc_trk_g3, op_bot, pgate, prog, purst,
     reset_b, s_r, vdd_cntl, wl );
output  carry_out, op_vic;


input  cin2local, clk, clkb, op_bot, prog, purst, s_r;

output [7:0]  slf_op;

inout [27:0]  bl;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;

input [15:0]  reset_b;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g2;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  wl;
input [7:0]  lc_trk_g3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbitb;

wire  [55:0]  cbit;



lcmuxod3_0_0 I_LC_00 ( .cbitb(cbitb[55:0]), .cbit(cbit[55:0]),
     .op_bot(op_bot), .op_vic(net0118), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .carry_out(c_01),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], cin}),
     .reset_b(reset_b[1:0]), .vdd_cntl(vdd_cntl[1:0]), .wl(wl[1:0]),
     .op(slf_op[0]), .s_r(s_r), .sp4_h_r({sp4_h_r[32], sp4_h_r[16],
     sp4_h_r[0]}), .sp12_v_b({sp12_v_b[16], sp12_v_b[0]}),
     .sp4_r_v_b({sp4_r_v_b[33], sp4_r_v_b[17], sp4_r_v_b[1]}),
     .sp4_v_b({sp4_v_b[32], sp4_v_b[16], sp4_v_b[0]}), .carry_in(cin),
     .sp12_h_r(sp12_h_r[8]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[1:0]), .prog(prog));
lcmuxod3_0 I_LC_02 ( .op_bot(net0166), .op_vic(net094),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .carry_out(c_23), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_12}),
     .reset_b(reset_b[5:4]), .vdd_cntl(vdd_cntl[5:4]), .wl(wl[5:4]),
     .op(slf_op[2]), .s_r(s_r), .sp4_h_r({sp4_h_r[36], sp4_h_r[20],
     sp4_h_r[4]}), .sp12_v_b({sp12_v_b[20], sp12_v_b[4]}),
     .sp4_r_v_b({sp4_r_v_b[37], sp4_r_v_b[21], sp4_r_v_b[5]}),
     .sp4_v_b({sp4_v_b[36], sp4_v_b[20], sp4_v_b[4]}), .carry_in(c_12),
     .sp12_h_r(sp12_h_r[12]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[5:4]), .prog(prog));
lcmuxod3_0 I_LC_03 ( .op_bot(net094), .op_vic(net0142),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .carry_out(c_34), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_23}),
     .reset_b(reset_b[7:6]), .vdd_cntl(vdd_cntl[7:6]), .wl(wl[7:6]),
     .op(slf_op[3]), .s_r(s_r), .sp4_h_r({sp4_h_r[38], sp4_h_r[22],
     sp4_h_r[6]}), .sp12_v_b({sp12_v_b[22], sp12_v_b[6]}),
     .sp4_r_v_b({sp4_r_v_b[39], sp4_r_v_b[23], sp4_r_v_b[7]}),
     .sp4_v_b({sp4_v_b[38], sp4_v_b[22], sp4_v_b[6]}), .carry_in(c_23),
     .sp12_h_r(sp12_h_r[14]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[7:6]), .prog(prog));
lcmuxod3_0 I_LC_01 ( .op_bot(net0118), .op_vic(net0166),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .carry_out(c_12), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_01}),
     .reset_b(reset_b[3:2]), .vdd_cntl(vdd_cntl[3:2]), .wl(wl[3:2]),
     .op(slf_op[1]), .s_r(s_r), .sp4_h_r({sp4_h_r[34], sp4_h_r[18],
     sp4_h_r[2]}), .sp12_v_b({sp12_v_b[18], sp12_v_b[2]}),
     .sp4_r_v_b({sp4_r_v_b[35], sp4_r_v_b[19], sp4_r_v_b[3]}),
     .sp4_v_b({sp4_v_b[34], sp4_v_b[18], sp4_v_b[2]}), .carry_in(c_01),
     .sp12_h_r(sp12_h_r[10]), .clkb(clkb), .clk(clk), .bl(bl[27:0]),
     .purst(purst), .pgate(pgate[3:2]), .prog(prog));
lcmuxod7_4 I_LC_07 ( .op_vic(op_vic), .op_bot(net0261), .bl(bl[27:0]),
     .reset_b(reset_b[15:14]), .purst(purst), .wl(wl[15:14]),
     .vdd_cntl(vdd_cntl[15:14]), .sp4_r_v_b({sp4_r_v_b[47],
     sp4_r_v_b[31], sp4_r_v_b[15]}), .sp4_h_r({sp4_h_r[46],
     sp4_h_r[30], sp4_h_r[14]}), .sp4_v_b({sp4_v_b[46], sp4_v_b[30],
     sp4_v_b[14]}), .pgate(pgate[15:14]), .sp12_h_r({sp12_h_r[22],
     sp12_h_r[6]}), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_67}),
     .carry_out(carry_out), .op(slf_op[7]), .s_r(s_r),
     .sp12_v_b(sp12_v_b[14]), .clk(clk), .carry_in(c_67),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clkb(clkb), .prog(prog));
lcmuxod7_4 I_LC_04 ( .op_vic(net0213), .op_bot(net0142), .prog(prog),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_34}), .clkb(clkb),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .purst(purst),
     .sp4_h_r({sp4_h_r[40], sp4_h_r[24], sp4_h_r[8]}),
     .sp4_r_v_b({sp4_r_v_b[41], sp4_r_v_b[25], sp4_r_v_b[9]}),
     .sp12_v_b(sp12_v_b[8]), .reset_b(reset_b[9:8]),
     .vdd_cntl(vdd_cntl[9:8]), .bl(bl[27:0]), .pgate(pgate[9:8]),
     .wl(wl[9:8]), .sp4_v_b({sp4_v_b[40], sp4_v_b[24], sp4_v_b[8]}),
     .sp12_h_r({sp12_h_r[16], sp12_h_r[0]}), .carry_out(c_45),
     .carry_in(c_34), .op(slf_op[4]));
lcmuxod7_4 I_LC_05 ( .op_vic(net0237), .op_bot(net0213), .prog(prog),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_45}), .clkb(clkb),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .purst(purst),
     .sp4_h_r({sp4_h_r[42], sp4_h_r[26], sp4_h_r[10]}),
     .sp4_r_v_b({sp4_r_v_b[43], sp4_r_v_b[27], sp4_r_v_b[11]}),
     .sp12_v_b(sp12_v_b[10]), .reset_b(reset_b[11:10]),
     .vdd_cntl(vdd_cntl[11:10]), .bl(bl[27:0]), .pgate(pgate[11:10]),
     .wl(wl[11:10]), .sp4_v_b({sp4_v_b[42], sp4_v_b[26], sp4_v_b[10]}),
     .sp12_h_r({sp12_h_r[18], sp12_h_r[2]}), .carry_out(c_56),
     .carry_in(c_45), .op(slf_op[5]));
lcmuxod7_4 I_LC_06 ( .op_vic(net0261), .op_bot(net0237), .prog(prog),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_56}), .clkb(clkb),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .clk(clk), .s_r(s_r), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .purst(purst),
     .sp4_h_r({sp4_h_r[44], sp4_h_r[28], sp4_h_r[12]}),
     .sp4_r_v_b({sp4_r_v_b[45], sp4_r_v_b[29], sp4_r_v_b[13]}),
     .sp12_v_b(sp12_v_b[12]), .reset_b(reset_b[13:12]),
     .vdd_cntl(vdd_cntl[13:12]), .bl(bl[27:0]), .pgate(pgate[13:12]),
     .wl(wl[13:12]), .sp4_v_b({sp4_v_b[44], sp4_v_b[28], sp4_v_b[12]}),
     .sp12_h_r({sp12_h_r[20], sp12_h_r[4]}), .carry_out(c_67),
     .carry_in(c_56), .op(slf_op[6]));
mux_4carry I_carry_cnt ( .cin(cin2local), .lcl_cin(cin),
     .cbitb({cbitb[45], cbitb[48]}), .prog(prog), .cbit({cbit[45],
     cbit[48]}));

endmodule
// Library - ice8chip, Cell - ltile4_ice8p_v1, View - schematic
// LAST TIME SAVED: Apr 27 16:22:34 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module ltile4_ice8p_v1 ( carry_out, cntl_cbit, op_vic, slf_op, bl,
     sp4_h_l, sp4_h_r, sp4_r_v_b, sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r,
     sp12_v_b, sp12_v_t, bnl_op, bnr_op, bot_op, carry_in, glb_netwk,
     lft_op, op_bot, pgate, prog, purst, reset_b, rgt_op, tnl_op,
     tnr_op, top_op, vdd_cntl, wl );
output  carry_out, op_vic;


input  carry_in, op_bot, prog, purst;

output [7:0]  cntl_cbit;
output [7:0]  slf_op;

inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_t;
inout [53:0]  bl;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_t;

input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  bot_op;
input [7:0]  tnr_op;
input [15:0]  vdd_cntl;
input [7:0]  top_op;
input [7:0]  lft_op;
input [15:0]  pgate;
input [7:0]  bnr_op;
input [7:0]  bnl_op;
input [15:0]  reset_b;
input [15:0]  wl;
input [7:0]  glb_netwk;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net138;

wire  [3:0]  net_glb2local;

wire  [63:0]  cbitb_c;

wire  [63:0]  cbit_c;

wire  [7:0]  lc_trk_g0;

wire  [1:0]  sp12_h_r_mid;

wire  [7:0]  lc_trk_g3;

wire  [1:0]  sp12_v_b_mid;

wire  [7:0]  lc_trk_g1;

wire  [7:0]  lc_trk_g2;

wire  [7:0]  net139;



lccol_rev0 I_lccol_rev0 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .prog(progd), .purst(purstd), .op_bot(op_bot), .s_r(s_r),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .wl({wl[14], wl[15], wl[12], wl[13],
     wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2],
     wl[3], wl[0], wl[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .clkb(clkb), .clk(clk),
     .cin2local(carry_in), .slf_op(slf_op[7:0]), .carry_out(carry_out),
     .sp12_v_b(sp12_v_b[23:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .bl(bl[53:26]), .op_vic(op_vic));
rm7y  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7y  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7y  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7y  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7y  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7y  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7y  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7y  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7y  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7y  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7y  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7y  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7y  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7y  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7y  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7y  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7y  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7y  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7y  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7y  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7y  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7y  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7y  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7y  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
gmux_sp12to4 I_gmux_sp12to4 ( .reset_b({reset_b[14], reset_b[15],
     reset_b[12], reset_b[13], reset_b[10], reset_b[11], reset_b[8],
     reset_b[9], reset_b[6], reset_b[7], reset_b[4], reset_b[5],
     reset_b[2], reset_b[3], reset_b[0], reset_b[1]}),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .lft_op(lft_op[7:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .glb2local(net_glb2local[3:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .bnr_op(bnr_op[7:0]), .lc_trk_g2(lc_trk_g2[7:0]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .bl(bl[25:14]), .lc_trk_g3(lc_trk_g3[7:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .prog(progd));
misc_module4_v3 I_misc ( .wl({wl[14], wl[15], wl[12], wl[13], wl[10],
     wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3],
     wl[0], wl[1]}), .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18],
     sp12_h_r[16], sp12_h_r[14], sp12_h_r[12], sp12_h_r[10],
     sp12_h_r[8]}), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .b(sp12_v_b[1:0]), .lc_trk_g2(lc_trk_g2[5:0]),
     .lc_trk_g3(lc_trk_g3[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .glb2local(net_glb2local[3:0]), .bl(bl[3:0]),
     .min3(glb_netwk[7:0]), .cbitb(cbitb_c[63:0]), .clk(clk),
     .min2(glb_netwk[7:0]), .reset_b({reset_b[14], reset_b[15],
     reset_b[12], reset_b[13], reset_b[10], reset_b[11], reset_b[8],
     reset_b[9], reset_b[6], reset_b[7], reset_b[4], reset_b[5],
     reset_b[2], reset_b[3], reset_b[0], reset_b[1]}), .prog(progd),
     .m(sp12_v_b_mid[1:0]), .r(sp12_h_r[1:0]), .S_R(s_r),
     .sp4(sp4_h_r[23:16]), .clkb(clkb), .cbit({cbit_c[63:61],
     cntl_cbit[7], cbit_c[59:57], cntl_cbit[6], cbit_c[55:53],
     cntl_cbit[5], cbit_c[51:49], cntl_cbit[4], cbit_c[47:45],
     cntl_cbit[3], cbit_c[43:41], cntl_cbit[2], cbit_c[39:33],
     cntl_cbit[1], cbit_c[31:4], cntl_cbit[0], cbit_c[2:0]}),
     .lc_trk_g0(lc_trk_g0[5:0]), .glb_netwk(glb_netwk[7:0]),
     .min1(glb_netwk[7:0]), .min0(glb_netwk[7:0]),
     .l(sp12_h_r_mid[1:0]), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}));
span4_ice8p I_sp4_sw ( .bl(bl[13:4]), .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .pgate({pgate[14], pgate[15], pgate[12], pgate[13],
     pgate[10], pgate[11], pgate[8], pgate[9], pgate[6], pgate[7],
     pgate[4], pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .sp4_h_l(sp4_h_l[47:0]), .prog(progd), .sp4_v_b(sp4_v_b[47:0]),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .sp4_v_t(sp4_v_t[47:0]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .sp4_h_r(sp4_h_r[47:0]), .ccntrl_cbit({net139[0], net139[1],
     net139[2], net139[3], net139[4], net139[5], net139[6],
     net139[7]}), .bram_cbit({net138[0], net138[1], net138[2],
     net138[3], net138[4], net138[5], net138[6], net138[7]}));
rm8y  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm8y  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm8y  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm8y  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm8y  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm8y  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm8y  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm8y  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm8y  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm8y  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm8y  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm8y  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm8y  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm8y  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm8y  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm8y  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm8y  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm8y  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm8y  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm8y  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm8y  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm8y  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm8y  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm8y  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
inv_hvt I89 ( .A(progb), .Y(progd));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I97 ( .A(purst), .Y(purstb));
inv_hvt I98 ( .A(purstb), .Y(purstd));

endmodule
// Library - ice1chip, Cell - lt_1x8_top_ice1f, View - schematic
// LAST TIME SAVED: Mar  4 20:35:57 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module lt_1x8_top_ice1f ( carry_out, glb_netwk_b, glb_netwk_t, op_vic,
     slf_op_01, slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06,
     slf_op_07, slf_op_08, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02,
     sp4_h_l_03, sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07,
     sp4_h_l_08, sp4_h_r_01, sp4_h_r_02, sp4_h_r_03, sp4_h_r_04,
     sp4_h_r_05, sp4_h_r_06, sp4_h_r_07, sp4_h_r_08, sp4_r_v_b_01,
     sp4_r_v_b_02, sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05,
     sp4_r_v_b_06, sp4_r_v_b_07, sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02,
     sp4_v_b_03, sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07,
     sp4_v_b_08, sp4_v_t_08, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03,
     sp12_h_l_04, sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08,
     sp12_h_r_01, sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_h_r_05,
     sp12_h_r_06, sp12_h_r_07, sp12_h_r_08, sp12_v_b_01, sp12_v_t_08,
     vdd_cntl, wl, bnl_op_01, bnr_op_01, bot_op_01, carry_in,
     glb_netwk_col, lc_bot, lft_op_01, lft_op_02, lft_op_03, lft_op_04,
     lft_op_05, lft_op_06, lft_op_07, lft_op_08, prog, purst,
     rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04, rgt_op_05, rgt_op_06,
     rgt_op_07, rgt_op_08, tnl_op_08, tnr_op_08, top_op_08 );
output  carry_out, op_vic;


input  carry_in, lc_bot, prog, purst;

output [7:0]  slf_op_02;
output [7:0]  slf_op_08;
output [7:0]  slf_op_06;
output [7:0]  slf_op_01;
output [7:0]  slf_op_05;
output [7:0]  slf_op_07;
output [7:0]  glb_netwk_t;
output [7:0]  slf_op_04;
output [7:0]  glb_netwk_b;
output [7:0]  slf_op_03;

inout [47:0]  sp4_h_l_02;
inout [47:0]  sp4_h_l_07;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_v_b_05;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_h_r_03;
inout [23:0]  sp12_h_r_07;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_h_r_04;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_r_v_b_04;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_v_b_06;
inout [53:0]  bl;
inout [47:0]  sp4_h_l_06;
inout [47:0]  sp4_h_r_08;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_v_t_08;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_h_l_04;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_v_b_03;
inout [23:0]  sp12_h_l_05;
inout [23:0]  sp12_h_r_06;
inout [23:0]  sp12_h_l_03;
inout [23:0]  sp12_h_l_02;
inout [23:0]  sp12_h_r_04;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_r_v_b_05;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_r_v_b_08;
inout [23:0]  sp12_v_t_08;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_h_l_08;
inout [23:0]  sp12_v_b_01;
inout [23:0]  sp12_h_l_07;
inout [23:0]  sp12_h_r_08;
inout [127:0]  vdd_cntl;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_r_v_b_02;
inout [23:0]  sp12_h_l_06;
inout [127:0]  wl;
inout [127:0]  pgate;
inout [47:0]  sp4_v_b_02;
inout [127:0]  reset_b;

input [7:0]  lft_op_03;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_01;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_04;
input [7:0]  rgt_op_05;
input [7:0]  bot_op_01;
input [7:0]  lft_op_04;
input [7:0]  rgt_op_01;
input [7:0]  bnr_op_01;
input [7:0]  lft_op_07;
input [7:0]  lft_op_02;
input [7:0]  lft_op_05;
input [7:0]  bnl_op_01;
input [7:0]  top_op_08;
input [7:0]  lft_op_06;
input [7:0]  lft_op_08;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_02;
input [7:0]  rgt_op_08;
input [7:0]  tnr_op_08;
input [7:0]  tnl_op_08;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  colbuf_cntl_b;

wire  [23:0]  net990;

wire  [23:0]  net1083;

wire  [23:0]  net742;

wire  [23:0]  net649;

wire  [7:0]  net947;

wire  [7:0]  net1071;

wire  [23:0]  net680;

wire  [7:0]  net637;

wire  [7:0]  net978;

wire  [7:0]  colbuf_cntl_t;

wire  [23:0]  net959;

wire  [23:0]  net711;

wire  [7:0]  net0754;

wire  [7:0]  net668;



ltile4_ice8p_v1 I_LT06 ( .cntl_cbit({net637[0], net637[1], net637[2],
     net637[3], net637[4], net637[5], net637[6], net637[7]}),
     .op_bot(net732), .op_vic(net639), .prog(prog), .carry_out(net641),
     .lft_op(lft_op_06[7:0]), .sp12_h_l(sp12_h_l_06[23:0]),
     .sp4_h_l(sp4_h_l_06[47:0]), .sp4_v_b(sp4_v_b_06[47:0]),
     .sp12_v_b({net742[0], net742[1], net742[2], net742[3], net742[4],
     net742[5], net742[6], net742[7], net742[8], net742[9], net742[10],
     net742[11], net742[12], net742[13], net742[14], net742[15],
     net742[16], net742[17], net742[18], net742[19], net742[20],
     net742[21], net742[22], net742[23]}),
     .sp12_h_r(sp12_h_r_06[23:0]), .sp4_h_r(sp4_h_r_06[47:0]),
     .sp12_v_t({net649[0], net649[1], net649[2], net649[3], net649[4],
     net649[5], net649[6], net649[7], net649[8], net649[9], net649[10],
     net649[11], net649[12], net649[13], net649[14], net649[15],
     net649[16], net649[17], net649[18], net649[19], net649[20],
     net649[21], net649[22], net649[23]}), .sp4_v_t(sp4_v_b_07[47:0]),
     .sp4_r_v_b(sp4_r_v_b_06[47:0]), .wl(wl[95:80]),
     .top_op(slf_op_07[7:0]), .rgt_op(rgt_op_06[7:0]),
     .bot_op(slf_op_05[7:0]), .bl(bl[53:0]), .reset_b(reset_b[95:80]),
     .vdd_cntl(vdd_cntl[95:80]), .glb_netwk(glb_netwk_t[7:0]),
     .carry_in(net734), .purst(purst), .slf_op(slf_op_06[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_05[7:0]),
     .bnl_op(lft_op_05[7:0]), .tnr_op(rgt_op_07[7:0]),
     .tnl_op(lft_op_07[7:0]));
ltile4_ice8p_v1 I_LT03 ( .cntl_cbit({net668[0], net668[1], net668[2],
     net668[3], net668[4], net668[5], net668[6], net668[7]}),
     .op_bot(net980), .op_vic(net670), .prog(prog), .carry_out(net672),
     .lft_op(lft_op_03[7:0]), .sp12_h_l(sp12_h_l_03[23:0]),
     .sp4_h_l(sp4_h_l_03[47:0]), .sp4_v_b(sp4_v_b_03[47:0]),
     .sp12_v_b({net990[0], net990[1], net990[2], net990[3], net990[4],
     net990[5], net990[6], net990[7], net990[8], net990[9], net990[10],
     net990[11], net990[12], net990[13], net990[14], net990[15],
     net990[16], net990[17], net990[18], net990[19], net990[20],
     net990[21], net990[22], net990[23]}),
     .sp12_h_r(sp12_h_r_03[23:0]), .sp4_h_r(sp4_h_r_03[47:0]),
     .sp12_v_t({net680[0], net680[1], net680[2], net680[3], net680[4],
     net680[5], net680[6], net680[7], net680[8], net680[9], net680[10],
     net680[11], net680[12], net680[13], net680[14], net680[15],
     net680[16], net680[17], net680[18], net680[19], net680[20],
     net680[21], net680[22], net680[23]}), .sp4_v_t(sp4_v_b_04[47:0]),
     .sp4_r_v_b(sp4_r_v_b_03[47:0]), .wl(wl[47:32]),
     .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(net982), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4_ice8p_v1 I_LT04 ( .cntl_cbit(colbuf_cntl_b[7:0]),
     .op_bot(net670), .op_vic(net701), .prog(prog), .carry_out(net703),
     .lft_op(lft_op_04[7:0]), .sp12_h_l(sp12_h_l_04[23:0]),
     .sp4_h_l(sp4_h_l_04[47:0]), .sp4_v_b(sp4_v_b_04[47:0]),
     .sp12_v_b({net680[0], net680[1], net680[2], net680[3], net680[4],
     net680[5], net680[6], net680[7], net680[8], net680[9], net680[10],
     net680[11], net680[12], net680[13], net680[14], net680[15],
     net680[16], net680[17], net680[18], net680[19], net680[20],
     net680[21], net680[22], net680[23]}),
     .sp12_h_r(sp12_h_r_04[23:0]), .sp4_h_r(sp4_h_r_04[47:0]),
     .sp12_v_t({net711[0], net711[1], net711[2], net711[3], net711[4],
     net711[5], net711[6], net711[7], net711[8], net711[9], net711[10],
     net711[11], net711[12], net711[13], net711[14], net711[15],
     net711[16], net711[17], net711[18], net711[19], net711[20],
     net711[21], net711[22], net711[23]}), .sp4_v_t(sp4_v_b_05[47:0]),
     .sp4_r_v_b(sp4_r_v_b_04[47:0]), .wl(wl[63:48]),
     .top_op(slf_op_05[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(net672), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(rgt_op_05[7:0]),
     .tnl_op(lft_op_05[7:0]));
ltile4_ice8p_v1 I_LT05 ( .cntl_cbit(colbuf_cntl_t[7:0]),
     .op_bot(net701), .op_vic(net732), .prog(prog), .carry_out(net734),
     .lft_op(lft_op_05[7:0]), .sp12_h_l(sp12_h_l_05[23:0]),
     .sp4_h_l(sp4_h_l_05[47:0]), .sp4_v_b(sp4_v_b_05[47:0]),
     .sp12_v_b({net711[0], net711[1], net711[2], net711[3], net711[4],
     net711[5], net711[6], net711[7], net711[8], net711[9], net711[10],
     net711[11], net711[12], net711[13], net711[14], net711[15],
     net711[16], net711[17], net711[18], net711[19], net711[20],
     net711[21], net711[22], net711[23]}),
     .sp12_h_r(sp12_h_r_05[23:0]), .sp4_h_r(sp4_h_r_05[47:0]),
     .sp12_v_t({net742[0], net742[1], net742[2], net742[3], net742[4],
     net742[5], net742[6], net742[7], net742[8], net742[9], net742[10],
     net742[11], net742[12], net742[13], net742[14], net742[15],
     net742[16], net742[17], net742[18], net742[19], net742[20],
     net742[21], net742[22], net742[23]}), .sp4_v_t(sp4_v_b_06[47:0]),
     .sp4_r_v_b(sp4_r_v_b_05[47:0]), .wl(wl[79:64]),
     .top_op(slf_op_06[7:0]), .rgt_op(rgt_op_05[7:0]),
     .bot_op(slf_op_04[7:0]), .bl(bl[53:0]), .reset_b(reset_b[79:64]),
     .vdd_cntl(vdd_cntl[79:64]), .glb_netwk(glb_netwk_t[7:0]),
     .carry_in(net703), .purst(purst), .slf_op(slf_op_05[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_04[7:0]),
     .bnl_op(lft_op_04[7:0]), .tnr_op(rgt_op_06[7:0]),
     .tnl_op(lft_op_06[7:0]));
ltile4_ice8p_v1 I_LT01 ( .cntl_cbit({net947[0], net947[1], net947[2],
     net947[3], net947[4], net947[5], net947[6], net947[7]}),
     .op_bot(lc_bot), .op_vic(net949), .prog(prog), .carry_out(net951),
     .lft_op(lft_op_01[7:0]), .sp12_h_l(sp12_h_l_01[23:0]),
     .sp4_h_l(sp4_h_l_01[47:0]), .sp4_v_b(sp4_v_b_01[47:0]),
     .sp12_v_b(sp12_v_b_01[23:0]), .sp12_h_r(sp12_h_r_01[23:0]),
     .sp4_h_r(sp4_h_r_01[47:0]), .sp12_v_t({net959[0], net959[1],
     net959[2], net959[3], net959[4], net959[5], net959[6], net959[7],
     net959[8], net959[9], net959[10], net959[11], net959[12],
     net959[13], net959[14], net959[15], net959[16], net959[17],
     net959[18], net959[19], net959[20], net959[21], net959[22],
     net959[23]}), .sp4_v_t(sp4_v_b_02[47:0]),
     .sp4_r_v_b(sp4_r_v_b_01[47:0]), .wl(wl[15:0]),
     .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4_ice8p_v1 I_LT02 ( .cntl_cbit({net978[0], net978[1], net978[2],
     net978[3], net978[4], net978[5], net978[6], net978[7]}),
     .op_bot(net949), .op_vic(net980), .prog(prog), .carry_out(net982),
     .lft_op(lft_op_02[7:0]), .sp12_h_l(sp12_h_l_02[23:0]),
     .sp4_h_l(sp4_h_l_02[47:0]), .sp4_v_b(sp4_v_b_02[47:0]),
     .sp12_v_b({net959[0], net959[1], net959[2], net959[3], net959[4],
     net959[5], net959[6], net959[7], net959[8], net959[9], net959[10],
     net959[11], net959[12], net959[13], net959[14], net959[15],
     net959[16], net959[17], net959[18], net959[19], net959[20],
     net959[21], net959[22], net959[23]}),
     .sp12_h_r(sp12_h_r_02[23:0]), .sp4_h_r(sp4_h_r_02[47:0]),
     .sp12_v_t({net990[0], net990[1], net990[2], net990[3], net990[4],
     net990[5], net990[6], net990[7], net990[8], net990[9], net990[10],
     net990[11], net990[12], net990[13], net990[14], net990[15],
     net990[16], net990[17], net990[18], net990[19], net990[20],
     net990[21], net990[22], net990[23]}), .sp4_v_t(sp4_v_b_03[47:0]),
     .sp4_r_v_b(sp4_r_v_b_02[47:0]), .wl(wl[31:16]),
     .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk_b[7:0]),
     .carry_in(net951), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));
ltile4_ice8p_v1 I_LT08 ( .cntl_cbit({net0754[0], net0754[1],
     net0754[2], net0754[3], net0754[4], net0754[5], net0754[6],
     net0754[7]}), .op_bot(net1073), .op_vic(op_vic), .prog(prog),
     .carry_out(carry_out), .lft_op(lft_op_08[7:0]),
     .sp12_h_l(sp12_h_l_08[23:0]), .sp4_h_l(sp4_h_l_08[47:0]),
     .sp4_v_b(sp4_v_b_08[47:0]), .sp12_v_b({net1083[0], net1083[1],
     net1083[2], net1083[3], net1083[4], net1083[5], net1083[6],
     net1083[7], net1083[8], net1083[9], net1083[10], net1083[11],
     net1083[12], net1083[13], net1083[14], net1083[15], net1083[16],
     net1083[17], net1083[18], net1083[19], net1083[20], net1083[21],
     net1083[22], net1083[23]}), .sp12_h_r(sp12_h_r_08[23:0]),
     .sp4_h_r(sp4_h_r_08[47:0]), .sp12_v_t(sp12_v_t_08[23:0]),
     .sp4_v_t(sp4_v_t_08[47:0]), .sp4_r_v_b(sp4_r_v_b_08[47:0]),
     .wl(wl[127:112]), .top_op(top_op_08[7:0]),
     .rgt_op(rgt_op_08[7:0]), .bot_op(slf_op_07[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[127:112]), .vdd_cntl(vdd_cntl[127:112]),
     .glb_netwk(glb_netwk_t[7:0]), .carry_in(net1075), .purst(purst),
     .slf_op(slf_op_08[7:0]), .pgate(pgate[127:112]),
     .bnr_op(rgt_op_07[7:0]), .bnl_op(lft_op_07[7:0]),
     .tnr_op(tnr_op_08[7:0]), .tnl_op(tnl_op_08[7:0]));
ltile4_ice8p_v1 I_LT07 ( .cntl_cbit({net1071[0], net1071[1],
     net1071[2], net1071[3], net1071[4], net1071[5], net1071[6],
     net1071[7]}), .op_bot(net639), .op_vic(net1073), .prog(prog),
     .carry_out(net1075), .lft_op(lft_op_07[7:0]),
     .sp12_h_l(sp12_h_l_07[23:0]), .sp4_h_l(sp4_h_l_07[47:0]),
     .sp4_v_b(sp4_v_b_07[47:0]), .sp12_v_b({net649[0], net649[1],
     net649[2], net649[3], net649[4], net649[5], net649[6], net649[7],
     net649[8], net649[9], net649[10], net649[11], net649[12],
     net649[13], net649[14], net649[15], net649[16], net649[17],
     net649[18], net649[19], net649[20], net649[21], net649[22],
     net649[23]}), .sp12_h_r(sp12_h_r_07[23:0]),
     .sp4_h_r(sp4_h_r_07[47:0]), .sp12_v_t({net1083[0], net1083[1],
     net1083[2], net1083[3], net1083[4], net1083[5], net1083[6],
     net1083[7], net1083[8], net1083[9], net1083[10], net1083[11],
     net1083[12], net1083[13], net1083[14], net1083[15], net1083[16],
     net1083[17], net1083[18], net1083[19], net1083[20], net1083[21],
     net1083[22], net1083[23]}), .sp4_v_t(sp4_v_b_08[47:0]),
     .sp4_r_v_b(sp4_r_v_b_07[47:0]), .wl(wl[111:96]),
     .top_op(slf_op_08[7:0]), .rgt_op(rgt_op_07[7:0]),
     .bot_op(slf_op_06[7:0]), .bl(bl[53:0]), .reset_b(reset_b[111:96]),
     .vdd_cntl(vdd_cntl[111:96]), .glb_netwk(glb_netwk_t[7:0]),
     .carry_in(net641), .purst(purst), .slf_op(slf_op_07[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_06[7:0]),
     .bnl_op(lft_op_06[7:0]), .tnr_op(rgt_op_08[7:0]),
     .tnl_op(lft_op_08[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - clkbuffer500um, View - schematic
// LAST TIME SAVED: May 13 10:52:41 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module clkbuffer500um ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I4 ( .A(net6), .Y(out));
inv I3 ( .A(in), .Y(net6));

endmodule
// Library - ice1chip, Cell - quad_tr_ice1, View - schematic
// LAST TIME SAVED: Apr 26 17:01:49 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module quad_tr_ice1 ( bm_aa_2bot, bm_ab_2bot, bm_sdo_o, bs_en_o, ceb_o,
     cf_r, cf_t, fabric_out_07_17, fabric_out_08_17, fabric_out_13_09,
     fabric_out_13_10, hiz_b_o, mode_o, padeb_r, padeb_t_r,
     padin_07_17a, padin_13_09a, pado_r, pado_t_r, r_o, sdo, shift_o,
     slf_op_07_09, slf_op_07_10, slf_op_07_11, slf_op_07_12,
     slf_op_07_13, slf_op_07_14, slf_op_07_15, slf_op_07_16,
     slf_op_07_17, slf_op_08_09, slf_op_09_09, slf_op_10_09,
     slf_op_11_09, slf_op_12_09, slf_op_13_09, tclk_o, update_o, bl,
     pgate_r, reset_b_r, sp4_h_l_07_09, sp4_h_l_07_10, sp4_h_l_07_11,
     sp4_h_l_07_12, sp4_h_l_07_13, sp4_h_l_07_14, sp4_h_l_07_15,
     sp4_h_l_07_16, sp4_h_l_07_17, sp4_h_r_13_09, sp4_v_b_07_09,
     sp4_v_b_07_10, sp4_v_b_07_11, sp4_v_b_07_12, sp4_v_b_07_13,
     sp4_v_b_07_14, sp4_v_b_07_15, sp4_v_b_07_16, sp4_v_b_08_09,
     sp4_v_b_09_09, sp4_v_b_10_09, sp4_v_b_11_09, sp4_v_b_12_09,
     sp12_h_l_07_09, sp12_h_l_07_10, sp12_h_l_07_11, sp12_h_l_07_12,
     sp12_h_l_07_13, sp12_h_l_07_14, sp12_h_l_07_15, sp12_h_l_07_16,
     sp12_v_b_07_09, sp12_v_b_08_09, sp12_v_b_09_09, sp12_v_b_10_09,
     sp12_v_b_11_09, sp12_v_b_12_09, vdd_cntl_r, wl_r, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_07_09,
     bnl_op_08_09, bnl_op_09_09, bnl_op_10_09, bnl_op_11_09,
     bnl_op_12_09, bnl_op_13_09, bnr_op_07_09, bnr_op_08_09,
     bnr_op_09_09, bnr_op_10_09, bnr_op_11_09, bnr_op_12_09,
     bot_op_07_09, bot_op_08_09, bot_op_09_09, bot_op_10_09,
     bot_op_11_09, bot_op_12_09, bs_en_i, carry_in_07_09,
     carry_in_08_09, carry_in_09_09, carry_in_11_09, carry_in_12_09,
     ceb_i, glb_in, hiz_b_i, hold_r_t, hold_t_r, lc_bot_07_09,
     lc_bot_08_09, lc_bot_09_09, lc_bot_11_09, lc_bot_12_09,
     lft_op_07_09, lft_op_07_10, lft_op_07_11, lft_op_07_12,
     lft_op_07_13, lft_op_07_14, lft_op_07_15, lft_op_07_16, mode_i,
     padin_r, padin_t_r, prog, purst, r_i, sdi, shift_i, tclk_i,
     tnl_op_07_16, update_i );
output  bs_en_o, ceb_o, fabric_out_07_17, fabric_out_08_17,
     fabric_out_13_09, fabric_out_13_10, hiz_b_o, mode_o, padin_07_17a,
     padin_13_09a, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, carry_in_07_09, carry_in_08_09,
     carry_in_09_09, carry_in_11_09, carry_in_12_09, ceb_i, hiz_b_i,
     hold_r_t, hold_t_r, lc_bot_07_09, lc_bot_08_09, lc_bot_09_09,
     lc_bot_11_09, lc_bot_12_09, mode_i, prog, purst, r_i, sdi,
     shift_i, tclk_i, update_i;

output [23:12]  pado_t_r;
output [7:0]  slf_op_07_15;
output [7:0]  slf_op_08_09;
output [143:0]  cf_t;
output [191:0]  cf_r;
output [3:0]  slf_op_07_17;
output [23:12]  padeb_t_r;
output [3:0]  slf_op_13_09;
output [7:0]  slf_op_07_10;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_12_09;
output [7:0]  slf_op_07_11;
output [7:0]  slf_op_07_09;
output [7:0]  slf_op_07_12;
output [24:13]  padeb_r;
output [10:0]  bm_ab_2bot;
output [24:13]  pado_r;
output [7:0]  slf_op_07_13;
output [7:0]  slf_op_10_09;
output [10:0]  bm_aa_2bot;
output [7:0]  slf_op_07_16;
output [7:0]  slf_op_11_09;
output [7:0]  slf_op_09_09;
output [7:0]  slf_op_07_14;

inout [23:0]  sp12_v_b_11_09;
inout [47:0]  sp4_v_b_11_09;
inout [23:0]  sp12_h_l_07_15;
inout [47:0]  sp4_v_b_07_16;
inout [47:0]  sp4_h_l_07_09;
inout [47:0]  sp4_h_l_07_12;
inout [47:0]  sp4_h_l_07_13;
inout [47:0]  sp4_h_l_07_14;
inout [23:0]  sp12_v_b_10_09;
inout [23:0]  sp12_h_l_07_16;
inout [23:0]  sp12_v_b_07_09;
inout [47:0]  sp4_v_b_09_09;
inout [47:0]  sp4_v_b_07_10;
inout [47:0]  sp4_v_b_10_09;
inout [23:0]  sp12_v_b_09_09;
inout [23:0]  sp12_h_l_07_14;
inout [143:0]  wl_r;
inout [143:0]  vdd_cntl_r;
inout [23:0]  sp12_v_b_12_09;
inout [47:0]  sp4_v_b_07_12;
inout [15:0]  sp4_h_l_07_17;
inout [47:0]  sp4_h_l_07_16;
inout [47:0]  sp4_v_b_07_14;
inout [23:0]  sp12_h_l_07_10;
inout [47:0]  sp4_v_b_07_11;
inout [47:0]  sp4_v_b_07_15;
inout [23:0]  sp12_h_l_07_11;
inout [47:0]  sp4_h_l_07_15;
inout [143:0]  pgate_r;
inout [143:0]  reset_b_r;
inout [23:0]  sp12_h_l_07_12;
inout [47:0]  sp4_v_b_12_09;
inout [23:0]  sp12_h_l_07_09;
inout [47:0]  sp4_h_l_07_10;
inout [15:0]  sp4_h_r_13_09;
inout [23:0]  sp12_v_b_08_09;
inout [47:0]  sp4_v_b_07_09;
inout [23:0]  sp12_h_l_07_13;
inout [47:0]  sp4_h_l_07_11;
inout [47:0]  sp4_v_b_07_13;
inout [47:0]  sp4_v_b_08_09;
inout [329:0]  bl;

input [7:0]  bnl_op_13_09;
input [1:0]  bm_sweb_i;
input [7:0]  bnl_op_12_09;
input [7:0]  bnr_op_08_09;
input [7:0]  bot_op_12_09;
input [1:0]  bm_sclkrw_i;
input [7:0]  bm_sa_i;
input [7:0]  bnr_op_07_09;
input [7:0]  bnr_op_12_09;
input [7:0]  lft_op_07_13;
input [1:0]  bm_sdi_i;
input [7:0]  bnl_op_11_09;
input [7:0]  bnl_op_07_09;
input [7:0]  bnr_op_10_09;
input [7:0]  bot_op_09_09;
input [24:13]  padin_r;
input [7:0]  bot_op_11_09;
input [7:0]  bot_op_10_09;
input [7:0]  lft_op_07_15;
input [7:0]  lft_op_07_11;
input [7:0]  lft_op_07_16;
input [7:0]  lft_op_07_14;
input [7:0]  bot_op_08_09;
input [7:0]  bnr_op_09_09;
input [7:0]  bnl_op_08_09;
input [7:0]  lft_op_07_09;
input [23:12]  padin_t_r;
input [7:0]  bnl_op_09_09;
input [7:0]  lft_op_07_10;
input [7:0]  bnr_op_11_09;
input [3:0]  tnl_op_07_16;
input [7:0]  lft_op_07_12;
input [7:0]  glb_in;
input [7:0]  bot_op_07_09;
input [7:0]  bnl_op_10_09;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  net1153;

wire  [3:0]  slf_op_13_16;

wire  [3:0]  slf_op_13_12;

wire  [3:0]  slf_op_13_14;

wire  [0:0]  padinlat_t_r;

wire  [23:0]  net1014;

wire  [3:0]  slf_op_13_15;

wire  [47:0]  net1114;

wire  [3:0]  slf_op_13_10;

wire  [3:0]  slf_op_10_17;

wire  [3:0]  slf_op_08_17;

wire  [7:0]  clk_center;

wire  [7:0]  clk_tree_drv_tr;

wire  [3:0]  slf_op_12_17;

wire  [3:0]  slf_op_09_17;

wire  [1:0]  bm_sdi_b1_o;

wire  [3:0]  slf_op_11_17;

wire  [3:0]  slf_op_13_11;

wire  [3:0]  slf_op_13_13;

wire  [7:0]  net1224;

wire  [47:0]  net1111;

wire  [47:0]  net1365;

wire  [47:0]  net1400;

wire  [23:0]  net870;

wire  [7:0]  net1004;

wire  [47:0]  net938;

wire  [47:0]  net1157;

wire  [47:0]  net1402;

wire  [7:0]  net1405;

wire  [7:0]  net1190;

wire  [23:0]  net921;

wire  [47:0]  net996;

wire  [47:0]  net1067;

wire  [47:0]  net1220;

wire  [47:0]  net1032;

wire  [7:0]  net943;

wire  [23:0]  net1056;

wire  [23:0]  net1200;

wire  [47:0]  net1183;

wire  [47:0]  net1369;

wire  [7:0]  net1141;

wire  [47:0]  net1184;

wire  [23:0]  net1341;

wire  [47:0]  net879;

wire  [23:0]  net1107;

wire  [47:0]  net1430;

wire  [7:0]  net1407;

wire  [23:0]  net1150;

wire  [23:0]  net1297;

wire  [23:0]  net1109;

wire  [47:0]  net1252;

wire  [7:0]  net1284;

wire  [23:0]  net1108;

wire  [7:0]  net1130;

wire  [47:0]  net1368;

wire  [47:0]  net1062;

wire  [7:0]  net1227;

wire  [47:0]  net1090;

wire  [47:0]  net994;

wire  [47:0]  net1088;

wire  [47:0]  net1257;

wire  [47:0]  net1158;

wire  [47:0]  net1314;

wire  [23:0]  net965;

wire  [47:0]  net1069;

wire  [47:0]  net899;

wire  [47:0]  net1301;

wire  [47:0]  net973;

wire  [7:0]  net1131;

wire  [47:0]  net1431;

wire  [23:0]  net1377;

wire  [7:0]  net1097;

wire  [47:0]  net1020;

wire  [7:0]  net1225;

wire  [7:0]  net1191;

wire  [7:0]  net1098;

wire  [47:0]  net822;

wire  [47:0]  net1063;

wire  [47:0]  net1255;

wire  [47:0]  net1156;

wire  [7:0]  net813;

wire  [7:0]  net1192;

wire  [1:0]  net1387;

wire  [47:0]  net1019;

wire  [23:0]  net1013;

wire  [7:0]  net1095;

wire  [47:0]  net975;

wire  [47:0]  net817;

wire  [23:0]  net963;

wire  [7:0]  net1003;

wire  [7:0]  net1133;

wire  [47:0]  net1383;

wire  [47:0]  net1163;

wire  [23:0]  net934;

wire  [47:0]  net1432;

wire  [47:0]  net900;

wire  [47:0]  net824;

wire  [47:0]  net974;

wire  [23:0]  net918;

wire  [47:0]  net1256;

wire  [7:0]  net1408;

wire  [7:0]  net01228;

wire  [7:0]  net1047;

wire  [23:0]  net1151;

wire  [47:0]  net968;

wire  [47:0]  net995;

wire  [23:0]  net1393;

wire  [7:0]  net0848;

wire  [47:0]  net1361;

wire  [47:0]  net1428;

wire  [23:0]  net1216;

wire  [47:0]  net1207;

wire  [47:0]  net1161;

wire  [47:0]  net993;

wire  [47:0]  net972;

wire  [47:0]  net1087;

wire  [23:0]  net1244;

wire  [47:0]  net881;

wire  [23:0]  net868;

wire  [47:0]  net902;

wire  [47:0]  net1113;

wire  [7:0]  net953;

wire  [23:0]  net1294;

wire  [23:0]  net1201;

wire  [47:0]  net1371;

wire  [23:0]  net1386;

wire  [7:0]  net1039;

wire  [23:0]  net1106;

wire  [23:0]  net1059;

wire  [23:0]  net1245;

wire  [47:0]  net1182;

wire  [7:0]  net1318;

wire  [47:0]  net970;

wire  [7:0]  net1189;

wire  [47:0]  net1278;

wire  [47:0]  net0885;

wire  [47:0]  net1300;

wire  [7:0]  net1410;

wire  [47:0]  net878;

wire  [47:0]  net1160;

wire  [47:0]  net1018;

wire  [23:0]  net1203;

wire  [7:0]  net1285;

wire  [47:0]  net1427;

wire  [47:0]  net0882;

wire  [23:0]  net1355;

wire  [47:0]  net1089;

wire  [1:0]  net1380;

wire  [7:0]  net1404;

wire  [23:0]  net964;

wire  [47:0]  net1162;

wire  [23:0]  net1246;

wire  [47:0]  net1068;

wire  [23:0]  net1353;

wire  [23:0]  net1015;

wire  [47:0]  net1299;

wire  [7:0]  net01133;

wire  [7:0]  net1096;

wire  [23:0]  net1122;

wire  [47:0]  net820;

wire  [7:0]  net1036;

wire  [23:0]  net869;

wire  [47:0]  net1302;

wire  [15:0]  net793;

wire  [47:0]  net1254;

wire  [7:0]  net942;

wire  [47:0]  net821;

wire  [7:0]  net1001;

wire  [7:0]  net1409;

wire  [47:0]  net1372;

wire  [47:0]  net1205;

wire  [47:0]  net1275;

wire  [23:0]  net1385;

wire  [23:0]  net1295;

wire  [47:0]  net880;

wire  [7:0]  net1283;

wire  [47:0]  net1401;

wire  [23:0]  net1058;

wire  [47:0]  net1276;

wire  [47:0]  net1206;

wire  [7:0]  net01038;

wire  [7:0]  net1037;

wire  [47:0]  net1181;

wire  [23:0]  net919;

wire  [23:0]  net1202;

wire  [47:0]  net1017;

wire  [7:0]  net1423;

wire  [23:0]  net1152;

wire  [47:0]  net1064;

wire  [47:0]  net901;

wire  [7:0]  net1286;

wire  [7:0]  net1406;

wire  [47:0]  net1429;

wire  [7:0]  net1002;

wire  [23:0]  net1310;

wire  [23:0]  net1358;

wire  [47:0]  net1208;

wire  [47:0]  net969;

wire  [47:0]  net1250;

wire  [23:0]  net871;

wire  [47:0]  net1251;

wire  [23:0]  net1296;

wire  [7:0]  net1235;

wire  [23:0]  net1012;

wire  [47:0]  net1126;

wire  [23:0]  net1057;

wire  [7:0]  net1422;

wire  [23:0]  net1357;

wire  [7:0]  net0943;

wire  [23:0]  net1247;

wire  [23:0]  net1028;

wire  [23:0]  net920;

wire  [47:0]  net1066;

wire  [23:0]  net962;

wire  [47:0]  net823;

wire  [7:0]  net945;

wire  [47:0]  net1112;

wire  [47:0]  net1277;



bram1x4_ice1f I_lt_col_t10 ( .glb_netwk_top({net1423[0], net1423[1],
     net1423[2], net1423[3], net1423[4], net1423[5], net1423[6],
     net1423[7]}), .prog(prog), .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .reset_b(reset_b_r[127:0]), .bm_wdummymux_en_o(net1328),
     .bm_sreb_o(net1329), .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(net809),
     .bm_sa_o({net813[0], net813[1], net813[2], net813[3], net813[4],
     net813[5], net813[6], net813[7]}), .bm_rcapmux_en_o(net1333),
     .bm_init_o(net814), .lft_op_05({net1192[0], net1192[1],
     net1192[2], net1192[3], net1192[4], net1192[5], net1192[6],
     net1192[7]}), .bl(bl[203:162]), .sp4_h_l_06({net995[0], net995[1],
     net995[2], net995[3], net995[4], net995[5], net995[6], net995[7],
     net995[8], net995[9], net995[10], net995[11], net995[12],
     net995[13], net995[14], net995[15], net995[16], net995[17],
     net995[18], net995[19], net995[20], net995[21], net995[22],
     net995[23], net995[24], net995[25], net995[26], net995[27],
     net995[28], net995[29], net995[30], net995[31], net995[32],
     net995[33], net995[34], net995[35], net995[36], net995[37],
     net995[38], net995[39], net995[40], net995[41], net995[42],
     net995[43], net995[44], net995[45], net995[46], net995[47]}),
     .sp12_h_l_02({net964[0], net964[1], net964[2], net964[3],
     net964[4], net964[5], net964[6], net964[7], net964[8], net964[9],
     net964[10], net964[11], net964[12], net964[13], net964[14],
     net964[15], net964[16], net964[17], net964[18], net964[19],
     net964[20], net964[21], net964[22], net964[23]}),
     .lft_op_06({net1191[0], net1191[1], net1191[2], net1191[3],
     net1191[4], net1191[5], net1191[6], net1191[7]}),
     .sp12_h_l_03({net963[0], net963[1], net963[2], net963[3],
     net963[4], net963[5], net963[6], net963[7], net963[8], net963[9],
     net963[10], net963[11], net963[12], net963[13], net963[14],
     net963[15], net963[16], net963[17], net963[18], net963[19],
     net963[20], net963[21], net963[22], net963[23]}),
     .sp12_h_r_03({net1341[0], net1341[1], net1341[2], net1341[3],
     net1341[4], net1341[5], net1341[6], net1341[7], net1341[8],
     net1341[9], net1341[10], net1341[11], net1341[12], net1341[13],
     net1341[14], net1341[15], net1341[16], net1341[17], net1341[18],
     net1341[19], net1341[20], net1341[21], net1341[22], net1341[23]}),
     .sp12_h_l_01({net965[0], net965[1], net965[2], net965[3],
     net965[4], net965[5], net965[6], net965[7], net965[8], net965[9],
     net965[10], net965[11], net965[12], net965[13], net965[14],
     net965[15], net965[16], net965[17], net965[18], net965[19],
     net965[20], net965[21], net965[22], net965[23]}),
     .sp4_v_b_04({net968[0], net968[1], net968[2], net968[3],
     net968[4], net968[5], net968[6], net968[7], net968[8], net968[9],
     net968[10], net968[11], net968[12], net968[13], net968[14],
     net968[15], net968[16], net968[17], net968[18], net968[19],
     net968[20], net968[21], net968[22], net968[23], net968[24],
     net968[25], net968[26], net968[27], net968[28], net968[29],
     net968[30], net968[31], net968[32], net968[33], net968[34],
     net968[35], net968[36], net968[37], net968[38], net968[39],
     net968[40], net968[41], net968[42], net968[43], net968[44],
     net968[45], net968[46], net968[47]}), .sp4_v_b_05({net1017[0],
     net1017[1], net1017[2], net1017[3], net1017[4], net1017[5],
     net1017[6], net1017[7], net1017[8], net1017[9], net1017[10],
     net1017[11], net1017[12], net1017[13], net1017[14], net1017[15],
     net1017[16], net1017[17], net1017[18], net1017[19], net1017[20],
     net1017[21], net1017[22], net1017[23], net1017[24], net1017[25],
     net1017[26], net1017[27], net1017[28], net1017[29], net1017[30],
     net1017[31], net1017[32], net1017[33], net1017[34], net1017[35],
     net1017[36], net1017[37], net1017[38], net1017[39], net1017[40],
     net1017[41], net1017[42], net1017[43], net1017[44], net1017[45],
     net1017[46], net1017[47]}), .lft_op_07({net1190[0], net1190[1],
     net1190[2], net1190[3], net1190[4], net1190[5], net1190[6],
     net1190[7]}), .sp4_v_b_06({net1018[0], net1018[1], net1018[2],
     net1018[3], net1018[4], net1018[5], net1018[6], net1018[7],
     net1018[8], net1018[9], net1018[10], net1018[11], net1018[12],
     net1018[13], net1018[14], net1018[15], net1018[16], net1018[17],
     net1018[18], net1018[19], net1018[20], net1018[21], net1018[22],
     net1018[23], net1018[24], net1018[25], net1018[26], net1018[27],
     net1018[28], net1018[29], net1018[30], net1018[31], net1018[32],
     net1018[33], net1018[34], net1018[35], net1018[36], net1018[37],
     net1018[38], net1018[39], net1018[40], net1018[41], net1018[42],
     net1018[43], net1018[44], net1018[45], net1018[46], net1018[47]}),
     .sp4_v_b_08({net1020[0], net1020[1], net1020[2], net1020[3],
     net1020[4], net1020[5], net1020[6], net1020[7], net1020[8],
     net1020[9], net1020[10], net1020[11], net1020[12], net1020[13],
     net1020[14], net1020[15], net1020[16], net1020[17], net1020[18],
     net1020[19], net1020[20], net1020[21], net1020[22], net1020[23],
     net1020[24], net1020[25], net1020[26], net1020[27], net1020[28],
     net1020[29], net1020[30], net1020[31], net1020[32], net1020[33],
     net1020[34], net1020[35], net1020[36], net1020[37], net1020[38],
     net1020[39], net1020[40], net1020[41], net1020[42], net1020[43],
     net1020[44], net1020[45], net1020[46], net1020[47]}),
     .sp4_v_b_07({net1019[0], net1019[1], net1019[2], net1019[3],
     net1019[4], net1019[5], net1019[6], net1019[7], net1019[8],
     net1019[9], net1019[10], net1019[11], net1019[12], net1019[13],
     net1019[14], net1019[15], net1019[16], net1019[17], net1019[18],
     net1019[19], net1019[20], net1019[21], net1019[22], net1019[23],
     net1019[24], net1019[25], net1019[26], net1019[27], net1019[28],
     net1019[29], net1019[30], net1019[31], net1019[32], net1019[33],
     net1019[34], net1019[35], net1019[36], net1019[37], net1019[38],
     net1019[39], net1019[40], net1019[41], net1019[42], net1019[43],
     net1019[44], net1019[45], net1019[46], net1019[47]}),
     .lft_op_03({net1131[0], net1131[1], net1131[2], net1131[3],
     net1131[4], net1131[5], net1131[6], net1131[7]}),
     .lft_op_01(slf_op_09_09[7:0]), .sp4_h_l_02({net974[0], net974[1],
     net974[2], net974[3], net974[4], net974[5], net974[6], net974[7],
     net974[8], net974[9], net974[10], net974[11], net974[12],
     net974[13], net974[14], net974[15], net974[16], net974[17],
     net974[18], net974[19], net974[20], net974[21], net974[22],
     net974[23], net974[24], net974[25], net974[26], net974[27],
     net974[28], net974[29], net974[30], net974[31], net974[32],
     net974[33], net974[34], net974[35], net974[36], net974[37],
     net974[38], net974[39], net974[40], net974[41], net974[42],
     net974[43], net974[44], net974[45], net974[46], net974[47]}),
     .sp12_h_l_06({net1013[0], net1013[1], net1013[2], net1013[3],
     net1013[4], net1013[5], net1013[6], net1013[7], net1013[8],
     net1013[9], net1013[10], net1013[11], net1013[12], net1013[13],
     net1013[14], net1013[15], net1013[16], net1013[17], net1013[18],
     net1013[19], net1013[20], net1013[21], net1013[22], net1013[23]}),
     .sp12_h_r_07({net1353[0], net1353[1], net1353[2], net1353[3],
     net1353[4], net1353[5], net1353[6], net1353[7], net1353[8],
     net1353[9], net1353[10], net1353[11], net1353[12], net1353[13],
     net1353[14], net1353[15], net1353[16], net1353[17], net1353[18],
     net1353[19], net1353[20], net1353[21], net1353[22], net1353[23]}),
     .sp12_h_l_05({net1012[0], net1012[1], net1012[2], net1012[3],
     net1012[4], net1012[5], net1012[6], net1012[7], net1012[8],
     net1012[9], net1012[10], net1012[11], net1012[12], net1012[13],
     net1012[14], net1012[15], net1012[16], net1012[17], net1012[18],
     net1012[19], net1012[20], net1012[21], net1012[22], net1012[23]}),
     .sp12_h_r_06({net1355[0], net1355[1], net1355[2], net1355[3],
     net1355[4], net1355[5], net1355[6], net1355[7], net1355[8],
     net1355[9], net1355[10], net1355[11], net1355[12], net1355[13],
     net1355[14], net1355[15], net1355[16], net1355[17], net1355[18],
     net1355[19], net1355[20], net1355[21], net1355[22], net1355[23]}),
     .sp12_h_l_04({net962[0], net962[1], net962[2], net962[3],
     net962[4], net962[5], net962[6], net962[7], net962[8], net962[9],
     net962[10], net962[11], net962[12], net962[13], net962[14],
     net962[15], net962[16], net962[17], net962[18], net962[19],
     net962[20], net962[21], net962[22], net962[23]}),
     .sp12_h_r_05({net1357[0], net1357[1], net1357[2], net1357[3],
     net1357[4], net1357[5], net1357[6], net1357[7], net1357[8],
     net1357[9], net1357[10], net1357[11], net1357[12], net1357[13],
     net1357[14], net1357[15], net1357[16], net1357[17], net1357[18],
     net1357[19], net1357[20], net1357[21], net1357[22], net1357[23]}),
     .sp12_h_r_08({net1358[0], net1358[1], net1358[2], net1358[3],
     net1358[4], net1358[5], net1358[6], net1358[7], net1358[8],
     net1358[9], net1358[10], net1358[11], net1358[12], net1358[13],
     net1358[14], net1358[15], net1358[16], net1358[17], net1358[18],
     net1358[19], net1358[20], net1358[21], net1358[22], net1358[23]}),
     .sp12_h_l_07({net1014[0], net1014[1], net1014[2], net1014[3],
     net1014[4], net1014[5], net1014[6], net1014[7], net1014[8],
     net1014[9], net1014[10], net1014[11], net1014[12], net1014[13],
     net1014[14], net1014[15], net1014[16], net1014[17], net1014[18],
     net1014[19], net1014[20], net1014[21], net1014[22], net1014[23]}),
     .sp12_h_l_08({net1015[0], net1015[1], net1015[2], net1015[3],
     net1015[4], net1015[5], net1015[6], net1015[7], net1015[8],
     net1015[9], net1015[10], net1015[11], net1015[12], net1015[13],
     net1015[14], net1015[15], net1015[16], net1015[17], net1015[18],
     net1015[19], net1015[20], net1015[21], net1015[22], net1015[23]}),
     .sp4_r_v_b_03({net1361[0], net1361[1], net1361[2], net1361[3],
     net1361[4], net1361[5], net1361[6], net1361[7], net1361[8],
     net1361[9], net1361[10], net1361[11], net1361[12], net1361[13],
     net1361[14], net1361[15], net1361[16], net1361[17], net1361[18],
     net1361[19], net1361[20], net1361[21], net1361[22], net1361[23],
     net1361[24], net1361[25], net1361[26], net1361[27], net1361[28],
     net1361[29], net1361[30], net1361[31], net1361[32], net1361[33],
     net1361[34], net1361[35], net1361[36], net1361[37], net1361[38],
     net1361[39], net1361[40], net1361[41], net1361[42], net1361[43],
     net1361[44], net1361[45], net1361[46], net1361[47]}),
     .vdd_cntl(vdd_cntl_r[127:0]), .pgate(pgate_r[127:0]),
     .bot_op_01(bot_op_10_09[7:0]), .sp4_r_v_b_04({net1365[0],
     net1365[1], net1365[2], net1365[3], net1365[4], net1365[5],
     net1365[6], net1365[7], net1365[8], net1365[9], net1365[10],
     net1365[11], net1365[12], net1365[13], net1365[14], net1365[15],
     net1365[16], net1365[17], net1365[18], net1365[19], net1365[20],
     net1365[21], net1365[22], net1365[23], net1365[24], net1365[25],
     net1365[26], net1365[27], net1365[28], net1365[29], net1365[30],
     net1365[31], net1365[32], net1365[33], net1365[34], net1365[35],
     net1365[36], net1365[37], net1365[38], net1365[39], net1365[40],
     net1365[41], net1365[42], net1365[43], net1365[44], net1365[45],
     net1365[46], net1365[47]}), .sp4_v_b_01(sp4_v_b_10_09[47:0]),
     .sp4_v_b_03({net969[0], net969[1], net969[2], net969[3],
     net969[4], net969[5], net969[6], net969[7], net969[8], net969[9],
     net969[10], net969[11], net969[12], net969[13], net969[14],
     net969[15], net969[16], net969[17], net969[18], net969[19],
     net969[20], net969[21], net969[22], net969[23], net969[24],
     net969[25], net969[26], net969[27], net969[28], net969[29],
     net969[30], net969[31], net969[32], net969[33], net969[34],
     net969[35], net969[36], net969[37], net969[38], net969[39],
     net969[40], net969[41], net969[42], net969[43], net969[44],
     net969[45], net969[46], net969[47]}), .sp4_h_r_08({net1368[0],
     net1368[1], net1368[2], net1368[3], net1368[4], net1368[5],
     net1368[6], net1368[7], net1368[8], net1368[9], net1368[10],
     net1368[11], net1368[12], net1368[13], net1368[14], net1368[15],
     net1368[16], net1368[17], net1368[18], net1368[19], net1368[20],
     net1368[21], net1368[22], net1368[23], net1368[24], net1368[25],
     net1368[26], net1368[27], net1368[28], net1368[29], net1368[30],
     net1368[31], net1368[32], net1368[33], net1368[34], net1368[35],
     net1368[36], net1368[37], net1368[38], net1368[39], net1368[40],
     net1368[41], net1368[42], net1368[43], net1368[44], net1368[45],
     net1368[46], net1368[47]}), .sp4_r_v_b_05({net1369[0], net1369[1],
     net1369[2], net1369[3], net1369[4], net1369[5], net1369[6],
     net1369[7], net1369[8], net1369[9], net1369[10], net1369[11],
     net1369[12], net1369[13], net1369[14], net1369[15], net1369[16],
     net1369[17], net1369[18], net1369[19], net1369[20], net1369[21],
     net1369[22], net1369[23], net1369[24], net1369[25], net1369[26],
     net1369[27], net1369[28], net1369[29], net1369[30], net1369[31],
     net1369[32], net1369[33], net1369[34], net1369[35], net1369[36],
     net1369[37], net1369[38], net1369[39], net1369[40], net1369[41],
     net1369[42], net1369[43], net1369[44], net1369[45], net1369[46],
     net1369[47]}), .sp4_v_b_02({net970[0], net970[1], net970[2],
     net970[3], net970[4], net970[5], net970[6], net970[7], net970[8],
     net970[9], net970[10], net970[11], net970[12], net970[13],
     net970[14], net970[15], net970[16], net970[17], net970[18],
     net970[19], net970[20], net970[21], net970[22], net970[23],
     net970[24], net970[25], net970[26], net970[27], net970[28],
     net970[29], net970[30], net970[31], net970[32], net970[33],
     net970[34], net970[35], net970[36], net970[37], net970[38],
     net970[39], net970[40], net970[41], net970[42], net970[43],
     net970[44], net970[45], net970[46], net970[47]}),
     .sp4_v_t_08({net1371[0], net1371[1], net1371[2], net1371[3],
     net1371[4], net1371[5], net1371[6], net1371[7], net1371[8],
     net1371[9], net1371[10], net1371[11], net1371[12], net1371[13],
     net1371[14], net1371[15], net1371[16], net1371[17], net1371[18],
     net1371[19], net1371[20], net1371[21], net1371[22], net1371[23],
     net1371[24], net1371[25], net1371[26], net1371[27], net1371[28],
     net1371[29], net1371[30], net1371[31], net1371[32], net1371[33],
     net1371[34], net1371[35], net1371[36], net1371[37], net1371[38],
     net1371[39], net1371[40], net1371[41], net1371[42], net1371[43],
     net1371[44], net1371[45], net1371[46], net1371[47]}),
     .sp4_r_v_b_02({net1372[0], net1372[1], net1372[2], net1372[3],
     net1372[4], net1372[5], net1372[6], net1372[7], net1372[8],
     net1372[9], net1372[10], net1372[11], net1372[12], net1372[13],
     net1372[14], net1372[15], net1372[16], net1372[17], net1372[18],
     net1372[19], net1372[20], net1372[21], net1372[22], net1372[23],
     net1372[24], net1372[25], net1372[26], net1372[27], net1372[28],
     net1372[29], net1372[30], net1372[31], net1372[32], net1372[33],
     net1372[34], net1372[35], net1372[36], net1372[37], net1372[38],
     net1372[39], net1372[40], net1372[41], net1372[42], net1372[43],
     net1372[44], net1372[45], net1372[46], net1372[47]}),
     .bnr_op_01(bnr_op_10_09[7:0]), .bm_sdi_o(bm_sdi_b1_o[1:0]),
     .sp4_h_l_04({net972[0], net972[1], net972[2], net972[3],
     net972[4], net972[5], net972[6], net972[7], net972[8], net972[9],
     net972[10], net972[11], net972[12], net972[13], net972[14],
     net972[15], net972[16], net972[17], net972[18], net972[19],
     net972[20], net972[21], net972[22], net972[23], net972[24],
     net972[25], net972[26], net972[27], net972[28], net972[29],
     net972[30], net972[31], net972[32], net972[33], net972[34],
     net972[35], net972[36], net972[37], net972[38], net972[39],
     net972[40], net972[41], net972[42], net972[43], net972[44],
     net972[45], net972[46], net972[47]}), .lft_op_08({net1189[0],
     net1189[1], net1189[2], net1189[3], net1189[4], net1189[5],
     net1189[6], net1189[7]}), .sp12_h_r_01({net1377[0], net1377[1],
     net1377[2], net1377[3], net1377[4], net1377[5], net1377[6],
     net1377[7], net1377[8], net1377[9], net1377[10], net1377[11],
     net1377[12], net1377[13], net1377[14], net1377[15], net1377[16],
     net1377[17], net1377[18], net1377[19], net1377[20], net1377[21],
     net1377[22], net1377[23]}), .bm_sdo_i({tiegnd_bram_t,
     bm_sdi_b1_o[0]}), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sweb_o({net1380[0], net1380[1]}), .sp4_h_l_03({net973[0],
     net973[1], net973[2], net973[3], net973[4], net973[5], net973[6],
     net973[7], net973[8], net973[9], net973[10], net973[11],
     net973[12], net973[13], net973[14], net973[15], net973[16],
     net973[17], net973[18], net973[19], net973[20], net973[21],
     net973[22], net973[23], net973[24], net973[25], net973[26],
     net973[27], net973[28], net973[29], net973[30], net973[31],
     net973[32], net973[33], net973[34], net973[35], net973[36],
     net973[37], net973[38], net973[39], net973[40], net973[41],
     net973[42], net973[43], net973[44], net973[45], net973[46],
     net973[47]}), .sp4_h_l_01({net975[0], net975[1], net975[2],
     net975[3], net975[4], net975[5], net975[6], net975[7], net975[8],
     net975[9], net975[10], net975[11], net975[12], net975[13],
     net975[14], net975[15], net975[16], net975[17], net975[18],
     net975[19], net975[20], net975[21], net975[22], net975[23],
     net975[24], net975[25], net975[26], net975[27], net975[28],
     net975[29], net975[30], net975[31], net975[32], net975[33],
     net975[34], net975[35], net975[36], net975[37], net975[38],
     net975[39], net975[40], net975[41], net975[42], net975[43],
     net975[44], net975[45], net975[46], net975[47]}),
     .sp4_h_r_01({net1383[0], net1383[1], net1383[2], net1383[3],
     net1383[4], net1383[5], net1383[6], net1383[7], net1383[8],
     net1383[9], net1383[10], net1383[11], net1383[12], net1383[13],
     net1383[14], net1383[15], net1383[16], net1383[17], net1383[18],
     net1383[19], net1383[20], net1383[21], net1383[22], net1383[23],
     net1383[24], net1383[25], net1383[26], net1383[27], net1383[28],
     net1383[29], net1383[30], net1383[31], net1383[32], net1383[33],
     net1383[34], net1383[35], net1383[36], net1383[37], net1383[38],
     net1383[39], net1383[40], net1383[41], net1383[42], net1383[43],
     net1383[44], net1383[45], net1383[46], net1383[47]}),
     .tnr_op_08({slf_op_11_17[3], slf_op_11_17[2], slf_op_11_17[1],
     slf_op_11_17[0], slf_op_11_17[3], slf_op_11_17[2],
     slf_op_11_17[1], slf_op_11_17[0]}), .sp12_h_r_02({net1385[0],
     net1385[1], net1385[2], net1385[3], net1385[4], net1385[5],
     net1385[6], net1385[7], net1385[8], net1385[9], net1385[10],
     net1385[11], net1385[12], net1385[13], net1385[14], net1385[15],
     net1385[16], net1385[17], net1385[18], net1385[19], net1385[20],
     net1385[21], net1385[22], net1385[23]}), .sp12_h_r_04({net1386[0],
     net1386[1], net1386[2], net1386[3], net1386[4], net1386[5],
     net1386[6], net1386[7], net1386[8], net1386[9], net1386[10],
     net1386[11], net1386[12], net1386[13], net1386[14], net1386[15],
     net1386[16], net1386[17], net1386[18], net1386[19], net1386[20],
     net1386[21], net1386[22], net1386[23]}), .bm_sclkrw_o({net1387[0],
     net1387[1]}), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .lft_op_02({net1133[0], net1133[1], net1133[2], net1133[3],
     net1133[4], net1133[5], net1133[6], net1133[7]}),
     .lft_op_04({net1141[0], net1141[1], net1141[2], net1141[3],
     net1141[4], net1141[5], net1141[6], net1141[7]}),
     .bm_sweb_i(bm_sweb_i[1:0]), .bnl_op_01(bnl_op_10_09[7:0]),
     .sp12_v_t_08({net1393[0], net1393[1], net1393[2], net1393[3],
     net1393[4], net1393[5], net1393[6], net1393[7], net1393[8],
     net1393[9], net1393[10], net1393[11], net1393[12], net1393[13],
     net1393[14], net1393[15], net1393[16], net1393[17], net1393[18],
     net1393[19], net1393[20], net1393[21], net1393[22], net1393[23]}),
     .wl(wl_r[127:0]), .tnl_op_08({slf_op_09_17[3], slf_op_09_17[2],
     slf_op_09_17[1], slf_op_09_17[0], slf_op_09_17[3],
     slf_op_09_17[2], slf_op_09_17[1], slf_op_09_17[0]}),
     .top_op_08({slf_op_10_17[3], slf_op_10_17[2], slf_op_10_17[1],
     slf_op_10_17[0], slf_op_10_17[3], slf_op_10_17[2],
     slf_op_10_17[1], slf_op_10_17[0]}), .bm_ab_2bot(bm_ab_2bot[10:0]),
     .bm_aa_2bot(bm_aa_2bot[10:0]), .sp12_v_b_01(sp12_v_b_10_09[23:0]),
     .sp4_r_v_b_08({net1400[0], net1400[1], net1400[2], net1400[3],
     net1400[4], net1400[5], net1400[6], net1400[7], net1400[8],
     net1400[9], net1400[10], net1400[11], net1400[12], net1400[13],
     net1400[14], net1400[15], net1400[16], net1400[17], net1400[18],
     net1400[19], net1400[20], net1400[21], net1400[22], net1400[23],
     net1400[24], net1400[25], net1400[26], net1400[27], net1400[28],
     net1400[29], net1400[30], net1400[31], net1400[32], net1400[33],
     net1400[34], net1400[35], net1400[36], net1400[37], net1400[38],
     net1400[39], net1400[40], net1400[41], net1400[42], net1400[43],
     net1400[44], net1400[45], net1400[46], net1400[47]}),
     .sp4_r_v_b_07({net1401[0], net1401[1], net1401[2], net1401[3],
     net1401[4], net1401[5], net1401[6], net1401[7], net1401[8],
     net1401[9], net1401[10], net1401[11], net1401[12], net1401[13],
     net1401[14], net1401[15], net1401[16], net1401[17], net1401[18],
     net1401[19], net1401[20], net1401[21], net1401[22], net1401[23],
     net1401[24], net1401[25], net1401[26], net1401[27], net1401[28],
     net1401[29], net1401[30], net1401[31], net1401[32], net1401[33],
     net1401[34], net1401[35], net1401[36], net1401[37], net1401[38],
     net1401[39], net1401[40], net1401[41], net1401[42], net1401[43],
     net1401[44], net1401[45], net1401[46], net1401[47]}),
     .sp4_r_v_b_06({net1402[0], net1402[1], net1402[2], net1402[3],
     net1402[4], net1402[5], net1402[6], net1402[7], net1402[8],
     net1402[9], net1402[10], net1402[11], net1402[12], net1402[13],
     net1402[14], net1402[15], net1402[16], net1402[17], net1402[18],
     net1402[19], net1402[20], net1402[21], net1402[22], net1402[23],
     net1402[24], net1402[25], net1402[26], net1402[27], net1402[28],
     net1402[29], net1402[30], net1402[31], net1402[32], net1402[33],
     net1402[34], net1402[35], net1402[36], net1402[37], net1402[38],
     net1402[39], net1402[40], net1402[41], net1402[42], net1402[43],
     net1402[44], net1402[45], net1402[46], net1402[47]}),
     .sp4_r_v_b_01(sp4_v_b_11_09[47:0]), .rgt_op_08({net1404[0],
     net1404[1], net1404[2], net1404[3], net1404[4], net1404[5],
     net1404[6], net1404[7]}), .rgt_op_07({net1405[0], net1405[1],
     net1405[2], net1405[3], net1405[4], net1405[5], net1405[6],
     net1405[7]}), .rgt_op_06({net1406[0], net1406[1], net1406[2],
     net1406[3], net1406[4], net1406[5], net1406[6], net1406[7]}),
     .rgt_op_05({net1407[0], net1407[1], net1407[2], net1407[3],
     net1407[4], net1407[5], net1407[6], net1407[7]}),
     .rgt_op_04({net1408[0], net1408[1], net1408[2], net1408[3],
     net1408[4], net1408[5], net1408[6], net1408[7]}),
     .rgt_op_03({net1409[0], net1409[1], net1409[2], net1409[3],
     net1409[4], net1409[5], net1409[6], net1409[7]}),
     .rgt_op_02({net1410[0], net1410[1], net1410[2], net1410[3],
     net1410[4], net1410[5], net1410[6], net1410[7]}),
     .rgt_op_01(slf_op_11_09[7:0]), .slf_op_02({net945[0], net945[1],
     net945[2], net945[3], net945[4], net945[5], net945[6],
     net945[7]}), .slf_op_01(slf_op_10_09[7:0]), .slf_op_03({net943[0],
     net943[1], net943[2], net943[3], net943[4], net943[5], net943[6],
     net943[7]}), .slf_op_04({net953[0], net953[1], net953[2],
     net953[3], net953[4], net953[5], net953[6], net953[7]}),
     .slf_op_05({net1004[0], net1004[1], net1004[2], net1004[3],
     net1004[4], net1004[5], net1004[6], net1004[7]}),
     .slf_op_06({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7]}),
     .slf_op_07({net1002[0], net1002[1], net1002[2], net1002[3],
     net1002[4], net1002[5], net1002[6], net1002[7]}),
     .slf_op_08({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7]}),
     .bm_ab_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .bm_aa_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .glb_netwk_bot({net1422[0], net1422[1], net1422[2], net1422[3],
     net1422[4], net1422[5], net1422[6], net1422[7]}),
     .sp4_h_l_08({net993[0], net993[1], net993[2], net993[3],
     net993[4], net993[5], net993[6], net993[7], net993[8], net993[9],
     net993[10], net993[11], net993[12], net993[13], net993[14],
     net993[15], net993[16], net993[17], net993[18], net993[19],
     net993[20], net993[21], net993[22], net993[23], net993[24],
     net993[25], net993[26], net993[27], net993[28], net993[29],
     net993[30], net993[31], net993[32], net993[33], net993[34],
     net993[35], net993[36], net993[37], net993[38], net993[39],
     net993[40], net993[41], net993[42], net993[43], net993[44],
     net993[45], net993[46], net993[47]}), .sp4_h_l_07({net994[0],
     net994[1], net994[2], net994[3], net994[4], net994[5], net994[6],
     net994[7], net994[8], net994[9], net994[10], net994[11],
     net994[12], net994[13], net994[14], net994[15], net994[16],
     net994[17], net994[18], net994[19], net994[20], net994[21],
     net994[22], net994[23], net994[24], net994[25], net994[26],
     net994[27], net994[28], net994[29], net994[30], net994[31],
     net994[32], net994[33], net994[34], net994[35], net994[36],
     net994[37], net994[38], net994[39], net994[40], net994[41],
     net994[42], net994[43], net994[44], net994[45], net994[46],
     net994[47]}), .sp4_h_l_05({net996[0], net996[1], net996[2],
     net996[3], net996[4], net996[5], net996[6], net996[7], net996[8],
     net996[9], net996[10], net996[11], net996[12], net996[13],
     net996[14], net996[15], net996[16], net996[17], net996[18],
     net996[19], net996[20], net996[21], net996[22], net996[23],
     net996[24], net996[25], net996[26], net996[27], net996[28],
     net996[29], net996[30], net996[31], net996[32], net996[33],
     net996[34], net996[35], net996[36], net996[37], net996[38],
     net996[39], net996[40], net996[41], net996[42], net996[43],
     net996[44], net996[45], net996[46], net996[47]}),
     .sp4_h_r_02({net1427[0], net1427[1], net1427[2], net1427[3],
     net1427[4], net1427[5], net1427[6], net1427[7], net1427[8],
     net1427[9], net1427[10], net1427[11], net1427[12], net1427[13],
     net1427[14], net1427[15], net1427[16], net1427[17], net1427[18],
     net1427[19], net1427[20], net1427[21], net1427[22], net1427[23],
     net1427[24], net1427[25], net1427[26], net1427[27], net1427[28],
     net1427[29], net1427[30], net1427[31], net1427[32], net1427[33],
     net1427[34], net1427[35], net1427[36], net1427[37], net1427[38],
     net1427[39], net1427[40], net1427[41], net1427[42], net1427[43],
     net1427[44], net1427[45], net1427[46], net1427[47]}),
     .sp4_h_r_03({net1428[0], net1428[1], net1428[2], net1428[3],
     net1428[4], net1428[5], net1428[6], net1428[7], net1428[8],
     net1428[9], net1428[10], net1428[11], net1428[12], net1428[13],
     net1428[14], net1428[15], net1428[16], net1428[17], net1428[18],
     net1428[19], net1428[20], net1428[21], net1428[22], net1428[23],
     net1428[24], net1428[25], net1428[26], net1428[27], net1428[28],
     net1428[29], net1428[30], net1428[31], net1428[32], net1428[33],
     net1428[34], net1428[35], net1428[36], net1428[37], net1428[38],
     net1428[39], net1428[40], net1428[41], net1428[42], net1428[43],
     net1428[44], net1428[45], net1428[46], net1428[47]}),
     .sp4_h_r_04({net1429[0], net1429[1], net1429[2], net1429[3],
     net1429[4], net1429[5], net1429[6], net1429[7], net1429[8],
     net1429[9], net1429[10], net1429[11], net1429[12], net1429[13],
     net1429[14], net1429[15], net1429[16], net1429[17], net1429[18],
     net1429[19], net1429[20], net1429[21], net1429[22], net1429[23],
     net1429[24], net1429[25], net1429[26], net1429[27], net1429[28],
     net1429[29], net1429[30], net1429[31], net1429[32], net1429[33],
     net1429[34], net1429[35], net1429[36], net1429[37], net1429[38],
     net1429[39], net1429[40], net1429[41], net1429[42], net1429[43],
     net1429[44], net1429[45], net1429[46], net1429[47]}),
     .sp4_h_r_05({net1430[0], net1430[1], net1430[2], net1430[3],
     net1430[4], net1430[5], net1430[6], net1430[7], net1430[8],
     net1430[9], net1430[10], net1430[11], net1430[12], net1430[13],
     net1430[14], net1430[15], net1430[16], net1430[17], net1430[18],
     net1430[19], net1430[20], net1430[21], net1430[22], net1430[23],
     net1430[24], net1430[25], net1430[26], net1430[27], net1430[28],
     net1430[29], net1430[30], net1430[31], net1430[32], net1430[33],
     net1430[34], net1430[35], net1430[36], net1430[37], net1430[38],
     net1430[39], net1430[40], net1430[41], net1430[42], net1430[43],
     net1430[44], net1430[45], net1430[46], net1430[47]}),
     .sp4_h_r_06({net1431[0], net1431[1], net1431[2], net1431[3],
     net1431[4], net1431[5], net1431[6], net1431[7], net1431[8],
     net1431[9], net1431[10], net1431[11], net1431[12], net1431[13],
     net1431[14], net1431[15], net1431[16], net1431[17], net1431[18],
     net1431[19], net1431[20], net1431[21], net1431[22], net1431[23],
     net1431[24], net1431[25], net1431[26], net1431[27], net1431[28],
     net1431[29], net1431[30], net1431[31], net1431[32], net1431[33],
     net1431[34], net1431[35], net1431[36], net1431[37], net1431[38],
     net1431[39], net1431[40], net1431[41], net1431[42], net1431[43],
     net1431[44], net1431[45], net1431[46], net1431[47]}),
     .sp4_h_r_07({net1432[0], net1432[1], net1432[2], net1432[3],
     net1432[4], net1432[5], net1432[6], net1432[7], net1432[8],
     net1432[9], net1432[10], net1432[11], net1432[12], net1432[13],
     net1432[14], net1432[15], net1432[16], net1432[17], net1432[18],
     net1432[19], net1432[20], net1432[21], net1432[22], net1432[23],
     net1432[24], net1432[25], net1432[26], net1432[27], net1432[28],
     net1432[29], net1432[30], net1432[31], net1432[32], net1432[33],
     net1432[34], net1432[35], net1432[36], net1432[37], net1432[38],
     net1432[39], net1432[40], net1432[41], net1432[42], net1432[43],
     net1432[44], net1432[45], net1432[46], net1432[47]}));
fabric_buf_ice8p I461 ( .f_in(net01448), .f_out(padin_13_09a));
fabric_buf_ice8p I_fabric_buf_8p_r_32 ( .f_in(net_fabric_out_13_09),
     .f_out(fabric_out_13_09));
fabric_buf_ice8p I451 ( .f_in(net_fabric_out_13_10),
     .f_out(fabric_out_13_10));
fabric_buf_ice8p I453 ( .f_in(net_fabric_out_07_17),
     .f_out(fabric_out_07_17));
fabric_buf_ice8p I454 ( .f_in(padinlat_t_r[0]), .f_out(padin_07_17a));
fabric_buf_ice8p I452 ( .f_in(net_fabric_out_08_17),
     .f_out(fabric_out_08_17));
io_rgt_top_1x8_ice1f I_lt_col_t13 ( .cf_r(cf_r[191:0]),
     .shift(shift_i), .bs_en(bs_en_i), .mode(mode_i), .sdi(sdi),
     .hiz_b(hiz_b_i), .prog(prog), .hold(hold_r_t), .update(update_i),
     .r(r_i), .SP4_h_l_05({net902[0], net902[1], net902[2], net902[3],
     net902[4], net902[5], net902[6], net902[7], net902[8], net902[9],
     net902[10], net902[11], net902[12], net902[13], net902[14],
     net902[15], net902[16], net902[17], net902[18], net902[19],
     net902[20], net902[21], net902[22], net902[23], net902[24],
     net902[25], net902[26], net902[27], net902[28], net902[29],
     net902[30], net902[31], net902[32], net902[33], net902[34],
     net902[35], net902[36], net902[37], net902[38], net902[39],
     net902[40], net902[41], net902[42], net902[43], net902[44],
     net902[45], net902[46], net902[47]}),
     .slf_op_05(slf_op_13_13[3:0]), .slf_op_01(slf_op_13_09[3:0]),
     .slf_op_06(slf_op_13_14[3:0]), .slf_op_02(slf_op_13_10[3:0]),
     .sdo(net680), .bl(bl[329:312]), .tclk(tclk_i),
     .reset_b(reset_b_r[127:0]), .lft_op_07({net1096[0], net1096[1],
     net1096[2], net1096[3], net1096[4], net1096[5], net1096[6],
     net1096[7]}), .SP4_h_l_06({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15], net901[16], net901[17], net901[18],
     net901[19], net901[20], net901[21], net901[22], net901[23],
     net901[24], net901[25], net901[26], net901[27], net901[28],
     net901[29], net901[30], net901[31], net901[32], net901[33],
     net901[34], net901[35], net901[36], net901[37], net901[38],
     net901[39], net901[40], net901[41], net901[42], net901[43],
     net901[44], net901[45], net901[46], net901[47]}),
     .sp4_v_t_08({net793[0], net793[1], net793[2], net793[3],
     net793[4], net793[5], net793[6], net793[7], net793[8], net793[9],
     net793[10], net793[11], net793[12], net793[13], net793[14],
     net793[15]}), .slf_op_04(slf_op_13_12[3:0]),
     .slf_op_03(slf_op_13_11[3:0]), .slf_op_07(slf_op_13_15[3:0]),
     .slf_op_08(slf_op_13_16[3:0]), .SP4_h_l_08({net899[0], net899[1],
     net899[2], net899[3], net899[4], net899[5], net899[6], net899[7],
     net899[8], net899[9], net899[10], net899[11], net899[12],
     net899[13], net899[14], net899[15], net899[16], net899[17],
     net899[18], net899[19], net899[20], net899[21], net899[22],
     net899[23], net899[24], net899[25], net899[26], net899[27],
     net899[28], net899[29], net899[30], net899[31], net899[32],
     net899[33], net899[34], net899[35], net899[36], net899[37],
     net899[38], net899[39], net899[40], net899[41], net899[42],
     net899[43], net899[44], net899[45], net899[46], net899[47]}),
     .SP4_h_l_07({net900[0], net900[1], net900[2], net900[3],
     net900[4], net900[5], net900[6], net900[7], net900[8], net900[9],
     net900[10], net900[11], net900[12], net900[13], net900[14],
     net900[15], net900[16], net900[17], net900[18], net900[19],
     net900[20], net900[21], net900[22], net900[23], net900[24],
     net900[25], net900[26], net900[27], net900[28], net900[29],
     net900[30], net900[31], net900[32], net900[33], net900[34],
     net900[35], net900[36], net900[37], net900[38], net900[39],
     net900[40], net900[41], net900[42], net900[43], net900[44],
     net900[45], net900[46], net900[47]}), .SP4_h_l_03({net879[0],
     net879[1], net879[2], net879[3], net879[4], net879[5], net879[6],
     net879[7], net879[8], net879[9], net879[10], net879[11],
     net879[12], net879[13], net879[14], net879[15], net879[16],
     net879[17], net879[18], net879[19], net879[20], net879[21],
     net879[22], net879[23], net879[24], net879[25], net879[26],
     net879[27], net879[28], net879[29], net879[30], net879[31],
     net879[32], net879[33], net879[34], net879[35], net879[36],
     net879[37], net879[38], net879[39], net879[40], net879[41],
     net879[42], net879[43], net879[44], net879[45], net879[46],
     net879[47]}), .SP4_h_l_04({net878[0], net878[1], net878[2],
     net878[3], net878[4], net878[5], net878[6], net878[7], net878[8],
     net878[9], net878[10], net878[11], net878[12], net878[13],
     net878[14], net878[15], net878[16], net878[17], net878[18],
     net878[19], net878[20], net878[21], net878[22], net878[23],
     net878[24], net878[25], net878[26], net878[27], net878[28],
     net878[29], net878[30], net878[31], net878[32], net878[33],
     net878[34], net878[35], net878[36], net878[37], net878[38],
     net878[39], net878[40], net878[41], net878[42], net878[43],
     net878[44], net878[45], net878[46], net878[47]}),
     .SP4_h_l_02({net880[0], net880[1], net880[2], net880[3],
     net880[4], net880[5], net880[6], net880[7], net880[8], net880[9],
     net880[10], net880[11], net880[12], net880[13], net880[14],
     net880[15], net880[16], net880[17], net880[18], net880[19],
     net880[20], net880[21], net880[22], net880[23], net880[24],
     net880[25], net880[26], net880[27], net880[28], net880[29],
     net880[30], net880[31], net880[32], net880[33], net880[34],
     net880[35], net880[36], net880[37], net880[38], net880[39],
     net880[40], net880[41], net880[42], net880[43], net880[44],
     net880[45], net880[46], net880[47]}), .SP4_h_l_01({net881[0],
     net881[1], net881[2], net881[3], net881[4], net881[5], net881[6],
     net881[7], net881[8], net881[9], net881[10], net881[11],
     net881[12], net881[13], net881[14], net881[15], net881[16],
     net881[17], net881[18], net881[19], net881[20], net881[21],
     net881[22], net881[23], net881[24], net881[25], net881[26],
     net881[27], net881[28], net881[29], net881[30], net881[31],
     net881[32], net881[33], net881[34], net881[35], net881[36],
     net881[37], net881[38], net881[39], net881[40], net881[41],
     net881[42], net881[43], net881[44], net881[45], net881[46],
     net881[47]}), .lft_op_04({net1047[0], net1047[1], net1047[2],
     net1047[3], net1047[4], net1047[5], net1047[6], net1047[7]}),
     .lft_op_06({net1097[0], net1097[1], net1097[2], net1097[3],
     net1097[4], net1097[5], net1097[6], net1097[7]}),
     .lft_op_01(slf_op_12_09[7:0]), .lft_op_08({net1095[0], net1095[1],
     net1095[2], net1095[3], net1095[4], net1095[5], net1095[6],
     net1095[7]}), .lft_op_02({net1039[0], net1039[1], net1039[2],
     net1039[3], net1039[4], net1039[5], net1039[6], net1039[7]}),
     .pgate(pgate_r[127:0]), .vdd_cntl(vdd_cntl_r[127:0]),
     .tnl_op_08({slf_op_12_17[3], slf_op_12_17[2], slf_op_12_17[1],
     slf_op_12_17[0], slf_op_12_17[3], slf_op_12_17[2],
     slf_op_12_17[1], slf_op_12_17[0]}), .wl(wl_r[127:0]),
     .tclk_o(net707), .ceb(ceb_i),
     .fabric_out_09(net_fabric_out_13_09), .SP12_h_l_02({net870[0],
     net870[1], net870[2], net870[3], net870[4], net870[5], net870[6],
     net870[7], net870[8], net870[9], net870[10], net870[11],
     net870[12], net870[13], net870[14], net870[15], net870[16],
     net870[17], net870[18], net870[19], net870[20], net870[21],
     net870[22], net870[23]}), .SP12_h_l_04({net868[0], net868[1],
     net868[2], net868[3], net868[4], net868[5], net868[6], net868[7],
     net868[8], net868[9], net868[10], net868[11], net868[12],
     net868[13], net868[14], net868[15], net868[16], net868[17],
     net868[18], net868[19], net868[20], net868[21], net868[22],
     net868[23]}), .SP12_h_l_08({net921[0], net921[1], net921[2],
     net921[3], net921[4], net921[5], net921[6], net921[7], net921[8],
     net921[9], net921[10], net921[11], net921[12], net921[13],
     net921[14], net921[15], net921[16], net921[17], net921[18],
     net921[19], net921[20], net921[21], net921[22], net921[23]}),
     .SP12_h_l_06({net919[0], net919[1], net919[2], net919[3],
     net919[4], net919[5], net919[6], net919[7], net919[8], net919[9],
     net919[10], net919[11], net919[12], net919[13], net919[14],
     net919[15], net919[16], net919[17], net919[18], net919[19],
     net919[20], net919[21], net919[22], net919[23]}),
     .glb_netwk_col(clk_tree_drv_tr[7:0]), .SP12_h_l_05({net918[0],
     net918[1], net918[2], net918[3], net918[4], net918[5], net918[6],
     net918[7], net918[8], net918[9], net918[10], net918[11],
     net918[12], net918[13], net918[14], net918[15], net918[16],
     net918[17], net918[18], net918[19], net918[20], net918[21],
     net918[22], net918[23]}), .SP12_h_l_01({net871[0], net871[1],
     net871[2], net871[3], net871[4], net871[5], net871[6], net871[7],
     net871[8], net871[9], net871[10], net871[11], net871[12],
     net871[13], net871[14], net871[15], net871[16], net871[17],
     net871[18], net871[19], net871[20], net871[21], net871[22],
     net871[23]}), .SP12_h_l_03({net869[0], net869[1], net869[2],
     net869[3], net869[4], net869[5], net869[6], net869[7], net869[8],
     net869[9], net869[10], net869[11], net869[12], net869[13],
     net869[14], net869[15], net869[16], net869[17], net869[18],
     net869[19], net869[20], net869[21], net869[22], net869[23]}),
     .SP12_h_l_07({net920[0], net920[1], net920[2], net920[3],
     net920[4], net920[5], net920[6], net920[7], net920[8], net920[9],
     net920[10], net920[11], net920[12], net920[13], net920[14],
     net920[15], net920[16], net920[17], net920[18], net920[19],
     net920[20], net920[21], net920[22], net920[23]}),
     .fabric_out_10(net_fabric_out_13_10), .padin(padin_r[24:13]),
     .pado(pado_r[24:13]), .padeb(padeb_r[24:13]),
     .lft_op_03({net1037[0], net1037[1], net1037[2], net1037[3],
     net1037[4], net1037[5], net1037[6], net1037[7]}),
     .bnl_op_13_09(bnl_op_13_09[7:0]), .lft_op_05({net1098[0],
     net1098[1], net1098[2], net1098[3], net1098[4], net1098[5],
     net1098[6], net1098[7]}), .sp4_v_b_13_09(sp4_h_r_13_09[15:0]));
io_top_rgt_1x6_ice1f I_preio_top_l ( .pado_t_r(pado_t_r[23:12]),
     .padeb_t_r(padeb_t_r[23:12]), .padin_t_r(padin_t_r[23:12]),
     .cf_t(cf_t[143:0]), .fabric_out_08_17(net_fabric_out_08_17),
     .hold_t_r(hold_t_r), .wl_l({wl_r[142], wl_r[143], wl_r[141],
     wl_r[140], wl_r[138], wl_r[139], wl_r[137], wl_r[136], wl_r[134],
     wl_r[135], wl_r[133], wl_r[132], wl_r[130], wl_r[131], wl_r[129],
     wl_r[128]}), .lft_op_01_17(slf_op_07_16[7:0]),
     .vdd_cntl_l({vdd_cntl_r[142], vdd_cntl_r[143], vdd_cntl_r[141],
     vdd_cntl_r[140], vdd_cntl_r[138], vdd_cntl_r[139],
     vdd_cntl_r[137], vdd_cntl_r[136], vdd_cntl_r[134],
     vdd_cntl_r[135], vdd_cntl_r[133], vdd_cntl_r[132],
     vdd_cntl_r[130], vdd_cntl_r[131], vdd_cntl_r[129],
     vdd_cntl_r[128]}), .update_i(net736), .tclk_i(net737),
     .shift_i(net738), .sdi(net739), .reset_l({reset_b_r[142],
     reset_b_r[143], reset_b_r[141], reset_b_r[140], reset_b_r[138],
     reset_b_r[139], reset_b_r[137], reset_b_r[136], reset_b_r[134],
     reset_b_r[135], reset_b_r[133], reset_b_r[132], reset_b_r[130],
     reset_b_r[131], reset_b_r[129], reset_b_r[128]}), .r_i(net741),
     .prog(prog), .pgate_l({pgate_r[142], pgate_r[143], pgate_r[141],
     pgate_r[140], pgate_r[138], pgate_r[139], pgate_r[137],
     pgate_r[136], pgate_r[134], pgate_r[135], pgate_r[133],
     pgate_r[132], pgate_r[130], pgate_r[131], pgate_r[129],
     pgate_r[128]}), .mode_i(net744), .hiz_b_i(net745),
     .bs_en_i(net746), .update_o(update_o), .tclk_o(tclk_o),
     .shift_o(shift_o), .sdo(sdo), .r_o(r_o), .mode_o(mode_o),
     .hiz_b_o(hiz_b_o), .glb_net_06({net942[0], net942[1], net942[2],
     net942[3], net942[4], net942[5], net942[6], net942[7]}),
     .glb_net_05({net1130[0], net1130[1], net1130[2], net1130[3],
     net1130[4], net1130[5], net1130[6], net1130[7]}),
     .glb_net_04({net1423[0], net1423[1], net1423[2], net1423[3],
     net1423[4], net1423[5], net1423[6], net1423[7]}),
     .glb_net_03({net1036[0], net1036[1], net1036[2], net1036[3],
     net1036[4], net1036[5], net1036[6], net1036[7]}),
     .glb_net_02({net1224[0], net1224[1], net1224[2], net1224[3],
     net1224[4], net1224[5], net1224[6], net1224[7]}),
     .glb_net_01({net1318[0], net1318[1], net1318[2], net1318[3],
     net1318[4], net1318[5], net1318[6], net1318[7]}),
     .bs_en_o(bs_en_o), .bl_06(bl[311:258]), .bl_05(bl[257:204]),
     .bl_02(bl[107:54]), .bl_01(bl[53:0]), .lft_op_03_17({net1189[0],
     net1189[1], net1189[2], net1189[3], net1189[4], net1189[5],
     net1189[6], net1189[7]}), .sp4_v_b_04_17({net1371[0], net1371[1],
     net1371[2], net1371[3], net1371[4], net1371[5], net1371[6],
     net1371[7], net1371[8], net1371[9], net1371[10], net1371[11],
     net1371[12], net1371[13], net1371[14], net1371[15], net1371[16],
     net1371[17], net1371[18], net1371[19], net1371[20], net1371[21],
     net1371[22], net1371[23], net1371[24], net1371[25], net1371[26],
     net1371[27], net1371[28], net1371[29], net1371[30], net1371[31],
     net1371[32], net1371[33], net1371[34], net1371[35], net1371[36],
     net1371[37], net1371[38], net1371[39], net1371[40], net1371[41],
     net1371[42], net1371[43], net1371[44], net1371[45], net1371[46],
     net1371[47]}), .lft_op_02_17({net1283[0], net1283[1], net1283[2],
     net1283[3], net1283[4], net1283[5], net1283[6], net1283[7]}),
     .lft_op_04_17({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7]}),
     .sp4_v_b_06_17({net938[0], net938[1], net938[2], net938[3],
     net938[4], net938[5], net938[6], net938[7], net938[8], net938[9],
     net938[10], net938[11], net938[12], net938[13], net938[14],
     net938[15], net938[16], net938[17], net938[18], net938[19],
     net938[20], net938[21], net938[22], net938[23], net938[24],
     net938[25], net938[26], net938[27], net938[28], net938[29],
     net938[30], net938[31], net938[32], net938[33], net938[34],
     net938[35], net938[36], net938[37], net938[38], net938[39],
     net938[40], net938[41], net938[42], net938[43], net938[44],
     net938[45], net938[46], net938[47]}), .sp12_v_b_04_17({net1393[0],
     net1393[1], net1393[2], net1393[3], net1393[4], net1393[5],
     net1393[6], net1393[7], net1393[8], net1393[9], net1393[10],
     net1393[11], net1393[12], net1393[13], net1393[14], net1393[15],
     net1393[16], net1393[17], net1393[18], net1393[19], net1393[20],
     net1393[21], net1393[22], net1393[23]}),
     .sp4_v_b_02_17({net1220[0], net1220[1], net1220[2], net1220[3],
     net1220[4], net1220[5], net1220[6], net1220[7], net1220[8],
     net1220[9], net1220[10], net1220[11], net1220[12], net1220[13],
     net1220[14], net1220[15], net1220[16], net1220[17], net1220[18],
     net1220[19], net1220[20], net1220[21], net1220[22], net1220[23],
     net1220[24], net1220[25], net1220[26], net1220[27], net1220[28],
     net1220[29], net1220[30], net1220[31], net1220[32], net1220[33],
     net1220[34], net1220[35], net1220[36], net1220[37], net1220[38],
     net1220[39], net1220[40], net1220[41], net1220[42], net1220[43],
     net1220[44], net1220[45], net1220[46], net1220[47]}),
     .sp12_v_b_05_17({net1122[0], net1122[1], net1122[2], net1122[3],
     net1122[4], net1122[5], net1122[6], net1122[7], net1122[8],
     net1122[9], net1122[10], net1122[11], net1122[12], net1122[13],
     net1122[14], net1122[15], net1122[16], net1122[17], net1122[18],
     net1122[19], net1122[20], net1122[21], net1122[22], net1122[23]}),
     .lft_op_06_17({net1095[0], net1095[1], net1095[2], net1095[3],
     net1095[4], net1095[5], net1095[6], net1095[7]}),
     .slf_op_04_17(slf_op_10_17[3:0]), .sp4_v_b_05_17({net1126[0],
     net1126[1], net1126[2], net1126[3], net1126[4], net1126[5],
     net1126[6], net1126[7], net1126[8], net1126[9], net1126[10],
     net1126[11], net1126[12], net1126[13], net1126[14], net1126[15],
     net1126[16], net1126[17], net1126[18], net1126[19], net1126[20],
     net1126[21], net1126[22], net1126[23], net1126[24], net1126[25],
     net1126[26], net1126[27], net1126[28], net1126[29], net1126[30],
     net1126[31], net1126[32], net1126[33], net1126[34], net1126[35],
     net1126[36], net1126[37], net1126[38], net1126[39], net1126[40],
     net1126[41], net1126[42], net1126[43], net1126[44], net1126[45],
     net1126[46], net1126[47]}), .sp12_v_b_03_17({net1028[0],
     net1028[1], net1028[2], net1028[3], net1028[4], net1028[5],
     net1028[6], net1028[7], net1028[8], net1028[9], net1028[10],
     net1028[11], net1028[12], net1028[13], net1028[14], net1028[15],
     net1028[16], net1028[17], net1028[18], net1028[19], net1028[20],
     net1028[21], net1028[22], net1028[23]}),
     .slf_op_01_17(slf_op_07_17[3:0]), .sp4_v_b_01_17({net1314[0],
     net1314[1], net1314[2], net1314[3], net1314[4], net1314[5],
     net1314[6], net1314[7], net1314[8], net1314[9], net1314[10],
     net1314[11], net1314[12], net1314[13], net1314[14], net1314[15],
     net1314[16], net1314[17], net1314[18], net1314[19], net1314[20],
     net1314[21], net1314[22], net1314[23], net1314[24], net1314[25],
     net1314[26], net1314[27], net1314[28], net1314[29], net1314[30],
     net1314[31], net1314[32], net1314[33], net1314[34], net1314[35],
     net1314[36], net1314[37], net1314[38], net1314[39], net1314[40],
     net1314[41], net1314[42], net1314[43], net1314[44], net1314[45],
     net1314[46], net1314[47]}), .sp4_v_b_03_17({net1032[0],
     net1032[1], net1032[2], net1032[3], net1032[4], net1032[5],
     net1032[6], net1032[7], net1032[8], net1032[9], net1032[10],
     net1032[11], net1032[12], net1032[13], net1032[14], net1032[15],
     net1032[16], net1032[17], net1032[18], net1032[19], net1032[20],
     net1032[21], net1032[22], net1032[23], net1032[24], net1032[25],
     net1032[26], net1032[27], net1032[28], net1032[29], net1032[30],
     net1032[31], net1032[32], net1032[33], net1032[34], net1032[35],
     net1032[36], net1032[37], net1032[38], net1032[39], net1032[40],
     net1032[41], net1032[42], net1032[43], net1032[44], net1032[45],
     net1032[46], net1032[47]}), .slf_op_03_17(slf_op_09_17[3:0]),
     .lft_op_05_17({net1404[0], net1404[1], net1404[2], net1404[3],
     net1404[4], net1404[5], net1404[6], net1404[7]}),
     .sp12_v_b_01_17({net1310[0], net1310[1], net1310[2], net1310[3],
     net1310[4], net1310[5], net1310[6], net1310[7], net1310[8],
     net1310[9], net1310[10], net1310[11], net1310[12], net1310[13],
     net1310[14], net1310[15], net1310[16], net1310[17], net1310[18],
     net1310[19], net1310[20], net1310[21], net1310[22], net1310[23]}),
     .slf_op_06_17(slf_op_12_17[3:0]), .sp12_v_b_06_17({net934[0],
     net934[1], net934[2], net934[3], net934[4], net934[5], net934[6],
     net934[7], net934[8], net934[9], net934[10], net934[11],
     net934[12], net934[13], net934[14], net934[15], net934[16],
     net934[17], net934[18], net934[19], net934[20], net934[21],
     net934[22], net934[23]}), .slf_op_02_17(slf_op_08_17[3:0]),
     .sp12_v_b_02_17({net1216[0], net1216[1], net1216[2], net1216[3],
     net1216[4], net1216[5], net1216[6], net1216[7], net1216[8],
     net1216[9], net1216[10], net1216[11], net1216[12], net1216[13],
     net1216[14], net1216[15], net1216[16], net1216[17], net1216[18],
     net1216[19], net1216[20], net1216[21], net1216[22], net1216[23]}),
     .bl_03(bl[161:108]), .bl_04(bl[203:162]), .ceb_o(ceb_o),
     .slf_op_05_17(slf_op_11_17[3:0]), .ceb_i(net791),
     .fabric_out_07_17(net_fabric_out_07_17),
     .sp4_h_r_12_17({net793[0], net793[1], net793[2], net793[3],
     net793[4], net793[5], net793[6], net793[7], net793[8], net793[9],
     net793[10], net793[11], net793[12], net793[13], net793[14],
     net793[15]}), .bnr_op_12_17({slf_op_13_16[3], slf_op_13_16[2],
     slf_op_13_16[1], slf_op_13_16[0], slf_op_13_16[3],
     slf_op_13_16[2], slf_op_13_16[1], slf_op_13_16[0]}),
     .sp4_h_l_07_17(sp4_h_l_07_17[15:0]),
     .bnl_op_07_17(lft_op_07_16[7:0]));
clk_quad_buf_x8_ice8p I428 ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));
clk_quad_buf_x8_ice8p I427 ( .clko(clk_tree_drv_tr[7:0]),
     .clki(clk_center[7:0]));
scan_buf_ice8p I446 ( .update_i(update_i), .tclk_i(net707),
     .shift_i(shift_i), .sdi(net680), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net736), .tclk_o(net737), .shift_o(net738),
     .sdo(net739), .r_o(net741), .mode_o(net744), .hiz_b_o(net745),
     .ceb_o(net791), .bs_en_o(net746));
tielo I430 ( .tielo(tiegnd_bram_t));
tielo I450 ( .tielo(net848));
lt_1x8_top_ice1f I_lt_col_t12 ( .glb_netwk_b({net0848[0], net0848[1],
     net0848[2], net0848[3], net0848[4], net0848[5], net0848[6],
     net0848[7]}), .rgt_op_03({slf_op_13_11[3], slf_op_13_11[2],
     slf_op_13_11[1], slf_op_13_11[0], slf_op_13_11[3],
     slf_op_13_11[2], slf_op_13_11[1], slf_op_13_11[0]}),
     .slf_op_02({net1039[0], net1039[1], net1039[2], net1039[3],
     net1039[4], net1039[5], net1039[6], net1039[7]}),
     .rgt_op_02({slf_op_13_10[3], slf_op_13_10[2], slf_op_13_10[1],
     slf_op_13_10[0], slf_op_13_10[3], slf_op_13_10[2],
     slf_op_13_10[1], slf_op_13_10[0]}), .rgt_op_01({slf_op_13_09[3],
     slf_op_13_09[2], slf_op_13_09[1], slf_op_13_09[0],
     slf_op_13_09[3], slf_op_13_09[2], slf_op_13_09[1],
     slf_op_13_09[0]}), .purst(purst), .prog(prog),
     .lft_op_04({net1408[0], net1408[1], net1408[2], net1408[3],
     net1408[4], net1408[5], net1408[6], net1408[7]}),
     .lft_op_03({net1409[0], net1409[1], net1409[2], net1409[3],
     net1409[4], net1409[5], net1409[6], net1409[7]}),
     .lft_op_02({net1410[0], net1410[1], net1410[2], net1410[3],
     net1410[4], net1410[5], net1410[6], net1410[7]}),
     .lft_op_01(slf_op_11_09[7:0]), .rgt_op_04({slf_op_13_12[3],
     slf_op_13_12[2], slf_op_13_12[1], slf_op_13_12[0],
     slf_op_13_12[3], slf_op_13_12[2], slf_op_13_12[1],
     slf_op_13_12[0]}), .carry_in(carry_in_12_09),
     .bnl_op_01(bnl_op_12_09[7:0]), .slf_op_04({net1047[0], net1047[1],
     net1047[2], net1047[3], net1047[4], net1047[5], net1047[6],
     net1047[7]}), .slf_op_03({net1037[0], net1037[1], net1037[2],
     net1037[3], net1037[4], net1037[5], net1037[6], net1037[7]}),
     .slf_op_01(slf_op_12_09[7:0]), .sp4_h_l_04({net1066[0],
     net1066[1], net1066[2], net1066[3], net1066[4], net1066[5],
     net1066[6], net1066[7], net1066[8], net1066[9], net1066[10],
     net1066[11], net1066[12], net1066[13], net1066[14], net1066[15],
     net1066[16], net1066[17], net1066[18], net1066[19], net1066[20],
     net1066[21], net1066[22], net1066[23], net1066[24], net1066[25],
     net1066[26], net1066[27], net1066[28], net1066[29], net1066[30],
     net1066[31], net1066[32], net1066[33], net1066[34], net1066[35],
     net1066[36], net1066[37], net1066[38], net1066[39], net1066[40],
     net1066[41], net1066[42], net1066[43], net1066[44], net1066[45],
     net1066[46], net1066[47]}), .carry_out(net866),
     .vdd_cntl(vdd_cntl_r[127:0]), .sp12_h_r_04({net868[0], net868[1],
     net868[2], net868[3], net868[4], net868[5], net868[6], net868[7],
     net868[8], net868[9], net868[10], net868[11], net868[12],
     net868[13], net868[14], net868[15], net868[16], net868[17],
     net868[18], net868[19], net868[20], net868[21], net868[22],
     net868[23]}), .sp12_h_r_03({net869[0], net869[1], net869[2],
     net869[3], net869[4], net869[5], net869[6], net869[7], net869[8],
     net869[9], net869[10], net869[11], net869[12], net869[13],
     net869[14], net869[15], net869[16], net869[17], net869[18],
     net869[19], net869[20], net869[21], net869[22], net869[23]}),
     .sp12_h_r_02({net870[0], net870[1], net870[2], net870[3],
     net870[4], net870[5], net870[6], net870[7], net870[8], net870[9],
     net870[10], net870[11], net870[12], net870[13], net870[14],
     net870[15], net870[16], net870[17], net870[18], net870[19],
     net870[20], net870[21], net870[22], net870[23]}),
     .sp12_h_r_01({net871[0], net871[1], net871[2], net871[3],
     net871[4], net871[5], net871[6], net871[7], net871[8], net871[9],
     net871[10], net871[11], net871[12], net871[13], net871[14],
     net871[15], net871[16], net871[17], net871[18], net871[19],
     net871[20], net871[21], net871[22], net871[23]}),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_12_09[47:0]), .sp4_r_v_b_04({net0882[0],
     net0882[1], net0882[2], net0882[3], net0882[4], net0882[5],
     net0882[6], net0882[7], net0882[8], net0882[9], net0882[10],
     net0882[11], net0882[12], net0882[13], net0882[14], net0882[15],
     net0882[16], net0882[17], net0882[18], net0882[19], net0882[20],
     net0882[21], net0882[22], net0882[23], net0882[24], net0882[25],
     net0882[26], net0882[27], net0882[28], net0882[29], net0882[30],
     net0882[31], net0882[32], net0882[33], net0882[34], net0882[35],
     net0882[36], net0882[37], net0882[38], net0882[39], net0882[40],
     net0882[41], net0882[42], net0882[43], net0882[44], net0882[45],
     net0882[46], net0882[47]}), .sp4_r_v_b_03({net820[0], net820[1],
     net820[2], net820[3], net820[4], net820[5], net820[6], net820[7],
     net820[8], net820[9], net820[10], net820[11], net820[12],
     net820[13], net820[14], net820[15], net820[16], net820[17],
     net820[18], net820[19], net820[20], net820[21], net820[22],
     net820[23], net820[24], net820[25], net820[26], net820[27],
     net820[28], net820[29], net820[30], net820[31], net820[32],
     net820[33], net820[34], net820[35], net820[36], net820[37],
     net820[38], net820[39], net820[40], net820[41], net820[42],
     net820[43], net820[44], net820[45], net820[46], net820[47]}),
     .sp4_r_v_b_02({net817[0], net817[1], net817[2], net817[3],
     net817[4], net817[5], net817[6], net817[7], net817[8], net817[9],
     net817[10], net817[11], net817[12], net817[13], net817[14],
     net817[15], net817[16], net817[17], net817[18], net817[19],
     net817[20], net817[21], net817[22], net817[23], net817[24],
     net817[25], net817[26], net817[27], net817[28], net817[29],
     net817[30], net817[31], net817[32], net817[33], net817[34],
     net817[35], net817[36], net817[37], net817[38], net817[39],
     net817[40], net817[41], net817[42], net817[43], net817[44],
     net817[45], net817[46], net817[47]}), .sp4_r_v_b_01({net0885[0],
     net0885[1], net0885[2], net0885[3], net0885[4], net0885[5],
     net0885[6], net0885[7], net0885[8], net0885[9], net0885[10],
     net0885[11], net0885[12], net0885[13], net0885[14], net0885[15],
     net0885[16], net0885[17], net0885[18], net0885[19], net0885[20],
     net0885[21], net0885[22], net0885[23], net0885[24], net0885[25],
     net0885[26], net0885[27], net0885[28], net0885[29], net0885[30],
     net0885[31], net0885[32], net0885[33], net0885[34], net0885[35],
     net0885[36], net0885[37], net0885[38], net0885[39], net0885[40],
     net0885[41], net0885[42], net0885[43], net0885[44], net0885[45],
     net0885[46], net0885[47]}), .sp4_h_r_04({net878[0], net878[1],
     net878[2], net878[3], net878[4], net878[5], net878[6], net878[7],
     net878[8], net878[9], net878[10], net878[11], net878[12],
     net878[13], net878[14], net878[15], net878[16], net878[17],
     net878[18], net878[19], net878[20], net878[21], net878[22],
     net878[23], net878[24], net878[25], net878[26], net878[27],
     net878[28], net878[29], net878[30], net878[31], net878[32],
     net878[33], net878[34], net878[35], net878[36], net878[37],
     net878[38], net878[39], net878[40], net878[41], net878[42],
     net878[43], net878[44], net878[45], net878[46], net878[47]}),
     .sp4_h_r_03({net879[0], net879[1], net879[2], net879[3],
     net879[4], net879[5], net879[6], net879[7], net879[8], net879[9],
     net879[10], net879[11], net879[12], net879[13], net879[14],
     net879[15], net879[16], net879[17], net879[18], net879[19],
     net879[20], net879[21], net879[22], net879[23], net879[24],
     net879[25], net879[26], net879[27], net879[28], net879[29],
     net879[30], net879[31], net879[32], net879[33], net879[34],
     net879[35], net879[36], net879[37], net879[38], net879[39],
     net879[40], net879[41], net879[42], net879[43], net879[44],
     net879[45], net879[46], net879[47]}), .sp4_h_r_02({net880[0],
     net880[1], net880[2], net880[3], net880[4], net880[5], net880[6],
     net880[7], net880[8], net880[9], net880[10], net880[11],
     net880[12], net880[13], net880[14], net880[15], net880[16],
     net880[17], net880[18], net880[19], net880[20], net880[21],
     net880[22], net880[23], net880[24], net880[25], net880[26],
     net880[27], net880[28], net880[29], net880[30], net880[31],
     net880[32], net880[33], net880[34], net880[35], net880[36],
     net880[37], net880[38], net880[39], net880[40], net880[41],
     net880[42], net880[43], net880[44], net880[45], net880[46],
     net880[47]}), .sp4_h_r_01({net881[0], net881[1], net881[2],
     net881[3], net881[4], net881[5], net881[6], net881[7], net881[8],
     net881[9], net881[10], net881[11], net881[12], net881[13],
     net881[14], net881[15], net881[16], net881[17], net881[18],
     net881[19], net881[20], net881[21], net881[22], net881[23],
     net881[24], net881[25], net881[26], net881[27], net881[28],
     net881[29], net881[30], net881[31], net881[32], net881[33],
     net881[34], net881[35], net881[36], net881[37], net881[38],
     net881[39], net881[40], net881[41], net881[42], net881[43],
     net881[44], net881[45], net881[46], net881[47]}),
     .sp4_h_l_03({net1067[0], net1067[1], net1067[2], net1067[3],
     net1067[4], net1067[5], net1067[6], net1067[7], net1067[8],
     net1067[9], net1067[10], net1067[11], net1067[12], net1067[13],
     net1067[14], net1067[15], net1067[16], net1067[17], net1067[18],
     net1067[19], net1067[20], net1067[21], net1067[22], net1067[23],
     net1067[24], net1067[25], net1067[26], net1067[27], net1067[28],
     net1067[29], net1067[30], net1067[31], net1067[32], net1067[33],
     net1067[34], net1067[35], net1067[36], net1067[37], net1067[38],
     net1067[39], net1067[40], net1067[41], net1067[42], net1067[43],
     net1067[44], net1067[45], net1067[46], net1067[47]}),
     .sp4_h_l_02({net1068[0], net1068[1], net1068[2], net1068[3],
     net1068[4], net1068[5], net1068[6], net1068[7], net1068[8],
     net1068[9], net1068[10], net1068[11], net1068[12], net1068[13],
     net1068[14], net1068[15], net1068[16], net1068[17], net1068[18],
     net1068[19], net1068[20], net1068[21], net1068[22], net1068[23],
     net1068[24], net1068[25], net1068[26], net1068[27], net1068[28],
     net1068[29], net1068[30], net1068[31], net1068[32], net1068[33],
     net1068[34], net1068[35], net1068[36], net1068[37], net1068[38],
     net1068[39], net1068[40], net1068[41], net1068[42], net1068[43],
     net1068[44], net1068[45], net1068[46], net1068[47]}),
     .sp4_h_l_01({net1069[0], net1069[1], net1069[2], net1069[3],
     net1069[4], net1069[5], net1069[6], net1069[7], net1069[8],
     net1069[9], net1069[10], net1069[11], net1069[12], net1069[13],
     net1069[14], net1069[15], net1069[16], net1069[17], net1069[18],
     net1069[19], net1069[20], net1069[21], net1069[22], net1069[23],
     net1069[24], net1069[25], net1069[26], net1069[27], net1069[28],
     net1069[29], net1069[30], net1069[31], net1069[32], net1069[33],
     net1069[34], net1069[35], net1069[36], net1069[37], net1069[38],
     net1069[39], net1069[40], net1069[41], net1069[42], net1069[43],
     net1069[44], net1069[45], net1069[46], net1069[47]}),
     .bl(bl[311:258]), .bot_op_01(bot_op_12_09[7:0]),
     .sp12_h_l_01({net1059[0], net1059[1], net1059[2], net1059[3],
     net1059[4], net1059[5], net1059[6], net1059[7], net1059[8],
     net1059[9], net1059[10], net1059[11], net1059[12], net1059[13],
     net1059[14], net1059[15], net1059[16], net1059[17], net1059[18],
     net1059[19], net1059[20], net1059[21], net1059[22], net1059[23]}),
     .sp12_h_l_02({net1058[0], net1058[1], net1058[2], net1058[3],
     net1058[4], net1058[5], net1058[6], net1058[7], net1058[8],
     net1058[9], net1058[10], net1058[11], net1058[12], net1058[13],
     net1058[14], net1058[15], net1058[16], net1058[17], net1058[18],
     net1058[19], net1058[20], net1058[21], net1058[22], net1058[23]}),
     .sp12_h_l_03({net1057[0], net1057[1], net1057[2], net1057[3],
     net1057[4], net1057[5], net1057[6], net1057[7], net1057[8],
     net1057[9], net1057[10], net1057[11], net1057[12], net1057[13],
     net1057[14], net1057[15], net1057[16], net1057[17], net1057[18],
     net1057[19], net1057[20], net1057[21], net1057[22], net1057[23]}),
     .sp12_h_l_04({net1056[0], net1056[1], net1056[2], net1056[3],
     net1056[4], net1056[5], net1056[6], net1056[7], net1056[8],
     net1056[9], net1056[10], net1056[11], net1056[12], net1056[13],
     net1056[14], net1056[15], net1056[16], net1056[17], net1056[18],
     net1056[19], net1056[20], net1056[21], net1056[22], net1056[23]}),
     .sp4_v_b_04({net1062[0], net1062[1], net1062[2], net1062[3],
     net1062[4], net1062[5], net1062[6], net1062[7], net1062[8],
     net1062[9], net1062[10], net1062[11], net1062[12], net1062[13],
     net1062[14], net1062[15], net1062[16], net1062[17], net1062[18],
     net1062[19], net1062[20], net1062[21], net1062[22], net1062[23],
     net1062[24], net1062[25], net1062[26], net1062[27], net1062[28],
     net1062[29], net1062[30], net1062[31], net1062[32], net1062[33],
     net1062[34], net1062[35], net1062[36], net1062[37], net1062[38],
     net1062[39], net1062[40], net1062[41], net1062[42], net1062[43],
     net1062[44], net1062[45], net1062[46], net1062[47]}),
     .sp4_v_b_03({net1063[0], net1063[1], net1063[2], net1063[3],
     net1063[4], net1063[5], net1063[6], net1063[7], net1063[8],
     net1063[9], net1063[10], net1063[11], net1063[12], net1063[13],
     net1063[14], net1063[15], net1063[16], net1063[17], net1063[18],
     net1063[19], net1063[20], net1063[21], net1063[22], net1063[23],
     net1063[24], net1063[25], net1063[26], net1063[27], net1063[28],
     net1063[29], net1063[30], net1063[31], net1063[32], net1063[33],
     net1063[34], net1063[35], net1063[36], net1063[37], net1063[38],
     net1063[39], net1063[40], net1063[41], net1063[42], net1063[43],
     net1063[44], net1063[45], net1063[46], net1063[47]}),
     .sp4_v_b_02({net1064[0], net1064[1], net1064[2], net1064[3],
     net1064[4], net1064[5], net1064[6], net1064[7], net1064[8],
     net1064[9], net1064[10], net1064[11], net1064[12], net1064[13],
     net1064[14], net1064[15], net1064[16], net1064[17], net1064[18],
     net1064[19], net1064[20], net1064[21], net1064[22], net1064[23],
     net1064[24], net1064[25], net1064[26], net1064[27], net1064[28],
     net1064[29], net1064[30], net1064[31], net1064[32], net1064[33],
     net1064[34], net1064[35], net1064[36], net1064[37], net1064[38],
     net1064[39], net1064[40], net1064[41], net1064[42], net1064[43],
     net1064[44], net1064[45], net1064[46], net1064[47]}),
     .bnr_op_01(bnr_op_12_09[7:0]), .sp4_h_l_05({net1090[0],
     net1090[1], net1090[2], net1090[3], net1090[4], net1090[5],
     net1090[6], net1090[7], net1090[8], net1090[9], net1090[10],
     net1090[11], net1090[12], net1090[13], net1090[14], net1090[15],
     net1090[16], net1090[17], net1090[18], net1090[19], net1090[20],
     net1090[21], net1090[22], net1090[23], net1090[24], net1090[25],
     net1090[26], net1090[27], net1090[28], net1090[29], net1090[30],
     net1090[31], net1090[32], net1090[33], net1090[34], net1090[35],
     net1090[36], net1090[37], net1090[38], net1090[39], net1090[40],
     net1090[41], net1090[42], net1090[43], net1090[44], net1090[45],
     net1090[46], net1090[47]}), .sp4_h_l_06({net1089[0], net1089[1],
     net1089[2], net1089[3], net1089[4], net1089[5], net1089[6],
     net1089[7], net1089[8], net1089[9], net1089[10], net1089[11],
     net1089[12], net1089[13], net1089[14], net1089[15], net1089[16],
     net1089[17], net1089[18], net1089[19], net1089[20], net1089[21],
     net1089[22], net1089[23], net1089[24], net1089[25], net1089[26],
     net1089[27], net1089[28], net1089[29], net1089[30], net1089[31],
     net1089[32], net1089[33], net1089[34], net1089[35], net1089[36],
     net1089[37], net1089[38], net1089[39], net1089[40], net1089[41],
     net1089[42], net1089[43], net1089[44], net1089[45], net1089[46],
     net1089[47]}), .sp4_h_l_07({net1088[0], net1088[1], net1088[2],
     net1088[3], net1088[4], net1088[5], net1088[6], net1088[7],
     net1088[8], net1088[9], net1088[10], net1088[11], net1088[12],
     net1088[13], net1088[14], net1088[15], net1088[16], net1088[17],
     net1088[18], net1088[19], net1088[20], net1088[21], net1088[22],
     net1088[23], net1088[24], net1088[25], net1088[26], net1088[27],
     net1088[28], net1088[29], net1088[30], net1088[31], net1088[32],
     net1088[33], net1088[34], net1088[35], net1088[36], net1088[37],
     net1088[38], net1088[39], net1088[40], net1088[41], net1088[42],
     net1088[43], net1088[44], net1088[45], net1088[46], net1088[47]}),
     .sp4_h_l_08({net1087[0], net1087[1], net1087[2], net1087[3],
     net1087[4], net1087[5], net1087[6], net1087[7], net1087[8],
     net1087[9], net1087[10], net1087[11], net1087[12], net1087[13],
     net1087[14], net1087[15], net1087[16], net1087[17], net1087[18],
     net1087[19], net1087[20], net1087[21], net1087[22], net1087[23],
     net1087[24], net1087[25], net1087[26], net1087[27], net1087[28],
     net1087[29], net1087[30], net1087[31], net1087[32], net1087[33],
     net1087[34], net1087[35], net1087[36], net1087[37], net1087[38],
     net1087[39], net1087[40], net1087[41], net1087[42], net1087[43],
     net1087[44], net1087[45], net1087[46], net1087[47]}),
     .sp4_h_r_08({net899[0], net899[1], net899[2], net899[3],
     net899[4], net899[5], net899[6], net899[7], net899[8], net899[9],
     net899[10], net899[11], net899[12], net899[13], net899[14],
     net899[15], net899[16], net899[17], net899[18], net899[19],
     net899[20], net899[21], net899[22], net899[23], net899[24],
     net899[25], net899[26], net899[27], net899[28], net899[29],
     net899[30], net899[31], net899[32], net899[33], net899[34],
     net899[35], net899[36], net899[37], net899[38], net899[39],
     net899[40], net899[41], net899[42], net899[43], net899[44],
     net899[45], net899[46], net899[47]}), .sp4_h_r_07({net900[0],
     net900[1], net900[2], net900[3], net900[4], net900[5], net900[6],
     net900[7], net900[8], net900[9], net900[10], net900[11],
     net900[12], net900[13], net900[14], net900[15], net900[16],
     net900[17], net900[18], net900[19], net900[20], net900[21],
     net900[22], net900[23], net900[24], net900[25], net900[26],
     net900[27], net900[28], net900[29], net900[30], net900[31],
     net900[32], net900[33], net900[34], net900[35], net900[36],
     net900[37], net900[38], net900[39], net900[40], net900[41],
     net900[42], net900[43], net900[44], net900[45], net900[46],
     net900[47]}), .sp4_h_r_06({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15], net901[16], net901[17], net901[18],
     net901[19], net901[20], net901[21], net901[22], net901[23],
     net901[24], net901[25], net901[26], net901[27], net901[28],
     net901[29], net901[30], net901[31], net901[32], net901[33],
     net901[34], net901[35], net901[36], net901[37], net901[38],
     net901[39], net901[40], net901[41], net901[42], net901[43],
     net901[44], net901[45], net901[46], net901[47]}),
     .sp4_h_r_05({net902[0], net902[1], net902[2], net902[3],
     net902[4], net902[5], net902[6], net902[7], net902[8], net902[9],
     net902[10], net902[11], net902[12], net902[13], net902[14],
     net902[15], net902[16], net902[17], net902[18], net902[19],
     net902[20], net902[21], net902[22], net902[23], net902[24],
     net902[25], net902[26], net902[27], net902[28], net902[29],
     net902[30], net902[31], net902[32], net902[33], net902[34],
     net902[35], net902[36], net902[37], net902[38], net902[39],
     net902[40], net902[41], net902[42], net902[43], net902[44],
     net902[45], net902[46], net902[47]}), .slf_op_05({net1098[0],
     net1098[1], net1098[2], net1098[3], net1098[4], net1098[5],
     net1098[6], net1098[7]}), .slf_op_06({net1097[0], net1097[1],
     net1097[2], net1097[3], net1097[4], net1097[5], net1097[6],
     net1097[7]}), .slf_op_07({net1096[0], net1096[1], net1096[2],
     net1096[3], net1096[4], net1096[5], net1096[6], net1096[7]}),
     .slf_op_08({net1095[0], net1095[1], net1095[2], net1095[3],
     net1095[4], net1095[5], net1095[6], net1095[7]}),
     .rgt_op_08({slf_op_13_16[3], slf_op_13_16[2], slf_op_13_16[1],
     slf_op_13_16[0], slf_op_13_16[3], slf_op_13_16[2],
     slf_op_13_16[1], slf_op_13_16[0]}), .rgt_op_07({slf_op_13_15[3],
     slf_op_13_15[2], slf_op_13_15[1], slf_op_13_15[0],
     slf_op_13_15[3], slf_op_13_15[2], slf_op_13_15[1],
     slf_op_13_15[0]}), .rgt_op_06({slf_op_13_14[3], slf_op_13_14[2],
     slf_op_13_14[1], slf_op_13_14[0], slf_op_13_14[3],
     slf_op_13_14[2], slf_op_13_14[1], slf_op_13_14[0]}),
     .rgt_op_05({slf_op_13_13[3], slf_op_13_13[2], slf_op_13_13[1],
     slf_op_13_13[0], slf_op_13_13[3], slf_op_13_13[2],
     slf_op_13_13[1], slf_op_13_13[0]}), .lft_op_08({net1404[0],
     net1404[1], net1404[2], net1404[3], net1404[4], net1404[5],
     net1404[6], net1404[7]}), .lft_op_07({net1405[0], net1405[1],
     net1405[2], net1405[3], net1405[4], net1405[5], net1405[6],
     net1405[7]}), .lft_op_06({net1406[0], net1406[1], net1406[2],
     net1406[3], net1406[4], net1406[5], net1406[6], net1406[7]}),
     .lft_op_05({net1407[0], net1407[1], net1407[2], net1407[3],
     net1407[4], net1407[5], net1407[6], net1407[7]}),
     .sp12_h_l_08({net1109[0], net1109[1], net1109[2], net1109[3],
     net1109[4], net1109[5], net1109[6], net1109[7], net1109[8],
     net1109[9], net1109[10], net1109[11], net1109[12], net1109[13],
     net1109[14], net1109[15], net1109[16], net1109[17], net1109[18],
     net1109[19], net1109[20], net1109[21], net1109[22], net1109[23]}),
     .sp12_h_l_07({net1108[0], net1108[1], net1108[2], net1108[3],
     net1108[4], net1108[5], net1108[6], net1108[7], net1108[8],
     net1108[9], net1108[10], net1108[11], net1108[12], net1108[13],
     net1108[14], net1108[15], net1108[16], net1108[17], net1108[18],
     net1108[19], net1108[20], net1108[21], net1108[22], net1108[23]}),
     .sp12_h_l_06({net1107[0], net1107[1], net1107[2], net1107[3],
     net1107[4], net1107[5], net1107[6], net1107[7], net1107[8],
     net1107[9], net1107[10], net1107[11], net1107[12], net1107[13],
     net1107[14], net1107[15], net1107[16], net1107[17], net1107[18],
     net1107[19], net1107[20], net1107[21], net1107[22], net1107[23]}),
     .sp12_h_r_05({net918[0], net918[1], net918[2], net918[3],
     net918[4], net918[5], net918[6], net918[7], net918[8], net918[9],
     net918[10], net918[11], net918[12], net918[13], net918[14],
     net918[15], net918[16], net918[17], net918[18], net918[19],
     net918[20], net918[21], net918[22], net918[23]}),
     .sp12_h_r_06({net919[0], net919[1], net919[2], net919[3],
     net919[4], net919[5], net919[6], net919[7], net919[8], net919[9],
     net919[10], net919[11], net919[12], net919[13], net919[14],
     net919[15], net919[16], net919[17], net919[18], net919[19],
     net919[20], net919[21], net919[22], net919[23]}),
     .sp12_h_r_07({net920[0], net920[1], net920[2], net920[3],
     net920[4], net920[5], net920[6], net920[7], net920[8], net920[9],
     net920[10], net920[11], net920[12], net920[13], net920[14],
     net920[15], net920[16], net920[17], net920[18], net920[19],
     net920[20], net920[21], net920[22], net920[23]}),
     .sp12_h_r_08({net921[0], net921[1], net921[2], net921[3],
     net921[4], net921[5], net921[6], net921[7], net921[8], net921[9],
     net921[10], net921[11], net921[12], net921[13], net921[14],
     net921[15], net921[16], net921[17], net921[18], net921[19],
     net921[20], net921[21], net921[22], net921[23]}),
     .sp12_h_l_05({net1106[0], net1106[1], net1106[2], net1106[3],
     net1106[4], net1106[5], net1106[6], net1106[7], net1106[8],
     net1106[9], net1106[10], net1106[11], net1106[12], net1106[13],
     net1106[14], net1106[15], net1106[16], net1106[17], net1106[18],
     net1106[19], net1106[20], net1106[21], net1106[22], net1106[23]}),
     .sp4_r_v_b_05({net824[0], net824[1], net824[2], net824[3],
     net824[4], net824[5], net824[6], net824[7], net824[8], net824[9],
     net824[10], net824[11], net824[12], net824[13], net824[14],
     net824[15], net824[16], net824[17], net824[18], net824[19],
     net824[20], net824[21], net824[22], net824[23], net824[24],
     net824[25], net824[26], net824[27], net824[28], net824[29],
     net824[30], net824[31], net824[32], net824[33], net824[34],
     net824[35], net824[36], net824[37], net824[38], net824[39],
     net824[40], net824[41], net824[42], net824[43], net824[44],
     net824[45], net824[46], net824[47]}), .sp4_r_v_b_06({net823[0],
     net823[1], net823[2], net823[3], net823[4], net823[5], net823[6],
     net823[7], net823[8], net823[9], net823[10], net823[11],
     net823[12], net823[13], net823[14], net823[15], net823[16],
     net823[17], net823[18], net823[19], net823[20], net823[21],
     net823[22], net823[23], net823[24], net823[25], net823[26],
     net823[27], net823[28], net823[29], net823[30], net823[31],
     net823[32], net823[33], net823[34], net823[35], net823[36],
     net823[37], net823[38], net823[39], net823[40], net823[41],
     net823[42], net823[43], net823[44], net823[45], net823[46],
     net823[47]}), .sp4_r_v_b_07({net821[0], net821[1], net821[2],
     net821[3], net821[4], net821[5], net821[6], net821[7], net821[8],
     net821[9], net821[10], net821[11], net821[12], net821[13],
     net821[14], net821[15], net821[16], net821[17], net821[18],
     net821[19], net821[20], net821[21], net821[22], net821[23],
     net821[24], net821[25], net821[26], net821[27], net821[28],
     net821[29], net821[30], net821[31], net821[32], net821[33],
     net821[34], net821[35], net821[36], net821[37], net821[38],
     net821[39], net821[40], net821[41], net821[42], net821[43],
     net821[44], net821[45], net821[46], net821[47]}),
     .sp4_r_v_b_08({net822[0], net822[1], net822[2], net822[3],
     net822[4], net822[5], net822[6], net822[7], net822[8], net822[9],
     net822[10], net822[11], net822[12], net822[13], net822[14],
     net822[15], net822[16], net822[17], net822[18], net822[19],
     net822[20], net822[21], net822[22], net822[23], net822[24],
     net822[25], net822[26], net822[27], net822[28], net822[29],
     net822[30], net822[31], net822[32], net822[33], net822[34],
     net822[35], net822[36], net822[37], net822[38], net822[39],
     net822[40], net822[41], net822[42], net822[43], net822[44],
     net822[45], net822[46], net822[47]}), .sp4_v_b_08({net1114[0],
     net1114[1], net1114[2], net1114[3], net1114[4], net1114[5],
     net1114[6], net1114[7], net1114[8], net1114[9], net1114[10],
     net1114[11], net1114[12], net1114[13], net1114[14], net1114[15],
     net1114[16], net1114[17], net1114[18], net1114[19], net1114[20],
     net1114[21], net1114[22], net1114[23], net1114[24], net1114[25],
     net1114[26], net1114[27], net1114[28], net1114[29], net1114[30],
     net1114[31], net1114[32], net1114[33], net1114[34], net1114[35],
     net1114[36], net1114[37], net1114[38], net1114[39], net1114[40],
     net1114[41], net1114[42], net1114[43], net1114[44], net1114[45],
     net1114[46], net1114[47]}), .sp4_v_b_07({net1113[0], net1113[1],
     net1113[2], net1113[3], net1113[4], net1113[5], net1113[6],
     net1113[7], net1113[8], net1113[9], net1113[10], net1113[11],
     net1113[12], net1113[13], net1113[14], net1113[15], net1113[16],
     net1113[17], net1113[18], net1113[19], net1113[20], net1113[21],
     net1113[22], net1113[23], net1113[24], net1113[25], net1113[26],
     net1113[27], net1113[28], net1113[29], net1113[30], net1113[31],
     net1113[32], net1113[33], net1113[34], net1113[35], net1113[36],
     net1113[37], net1113[38], net1113[39], net1113[40], net1113[41],
     net1113[42], net1113[43], net1113[44], net1113[45], net1113[46],
     net1113[47]}), .sp4_v_b_06({net1112[0], net1112[1], net1112[2],
     net1112[3], net1112[4], net1112[5], net1112[6], net1112[7],
     net1112[8], net1112[9], net1112[10], net1112[11], net1112[12],
     net1112[13], net1112[14], net1112[15], net1112[16], net1112[17],
     net1112[18], net1112[19], net1112[20], net1112[21], net1112[22],
     net1112[23], net1112[24], net1112[25], net1112[26], net1112[27],
     net1112[28], net1112[29], net1112[30], net1112[31], net1112[32],
     net1112[33], net1112[34], net1112[35], net1112[36], net1112[37],
     net1112[38], net1112[39], net1112[40], net1112[41], net1112[42],
     net1112[43], net1112[44], net1112[45], net1112[46], net1112[47]}),
     .sp4_v_b_05({net1111[0], net1111[1], net1111[2], net1111[3],
     net1111[4], net1111[5], net1111[6], net1111[7], net1111[8],
     net1111[9], net1111[10], net1111[11], net1111[12], net1111[13],
     net1111[14], net1111[15], net1111[16], net1111[17], net1111[18],
     net1111[19], net1111[20], net1111[21], net1111[22], net1111[23],
     net1111[24], net1111[25], net1111[26], net1111[27], net1111[28],
     net1111[29], net1111[30], net1111[31], net1111[32], net1111[33],
     net1111[34], net1111[35], net1111[36], net1111[37], net1111[38],
     net1111[39], net1111[40], net1111[41], net1111[42], net1111[43],
     net1111[44], net1111[45], net1111[46], net1111[47]}),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .wl(wl_r[127:0]), .sp12_v_t_08({net934[0], net934[1], net934[2],
     net934[3], net934[4], net934[5], net934[6], net934[7], net934[8],
     net934[9], net934[10], net934[11], net934[12], net934[13],
     net934[14], net934[15], net934[16], net934[17], net934[18],
     net934[19], net934[20], net934[21], net934[22], net934[23]}),
     .tnr_op_08({net848, net848, net848, net848, net848, net848,
     net848, net848}), .top_op_08({slf_op_12_17[3], slf_op_12_17[2],
     slf_op_12_17[1], slf_op_12_17[0], slf_op_12_17[3],
     slf_op_12_17[2], slf_op_12_17[1], slf_op_12_17[0]}),
     .tnl_op_08({slf_op_11_17[3], slf_op_11_17[2], slf_op_11_17[1],
     slf_op_11_17[0], slf_op_11_17[3], slf_op_11_17[2],
     slf_op_11_17[1], slf_op_11_17[0]}), .sp4_v_t_08({net938[0],
     net938[1], net938[2], net938[3], net938[4], net938[5], net938[6],
     net938[7], net938[8], net938[9], net938[10], net938[11],
     net938[12], net938[13], net938[14], net938[15], net938[16],
     net938[17], net938[18], net938[19], net938[20], net938[21],
     net938[22], net938[23], net938[24], net938[25], net938[26],
     net938[27], net938[28], net938[29], net938[30], net938[31],
     net938[32], net938[33], net938[34], net938[35], net938[36],
     net938[37], net938[38], net938[39], net938[40], net938[41],
     net938[42], net938[43], net938[44], net938[45], net938[46],
     net938[47]}), .lc_bot(lc_bot_12_09), .op_vic(net940),
     .sp12_v_b_01(sp12_v_b_12_09[23:0]), .glb_netwk_t({net942[0],
     net942[1], net942[2], net942[3], net942[4], net942[5], net942[6],
     net942[7]}));
lt_1x8_top_ice1f I_lt_col_t09 ( .glb_netwk_b({net0943[0], net0943[1],
     net0943[2], net0943[3], net0943[4], net0943[5], net0943[6],
     net0943[7]}), .rgt_op_03({net943[0], net943[1], net943[2],
     net943[3], net943[4], net943[5], net943[6], net943[7]}),
     .slf_op_02({net1133[0], net1133[1], net1133[2], net1133[3],
     net1133[4], net1133[5], net1133[6], net1133[7]}),
     .rgt_op_02({net945[0], net945[1], net945[2], net945[3], net945[4],
     net945[5], net945[6], net945[7]}), .rgt_op_01(slf_op_10_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04({net1235[0], net1235[1],
     net1235[2], net1235[3], net1235[4], net1235[5], net1235[6],
     net1235[7]}), .lft_op_03({net1225[0], net1225[1], net1225[2],
     net1225[3], net1225[4], net1225[5], net1225[6], net1225[7]}),
     .lft_op_02({net1227[0], net1227[1], net1227[2], net1227[3],
     net1227[4], net1227[5], net1227[6], net1227[7]}),
     .lft_op_01(slf_op_08_09[7:0]), .rgt_op_04({net953[0], net953[1],
     net953[2], net953[3], net953[4], net953[5], net953[6],
     net953[7]}), .carry_in(carry_in_09_09),
     .bnl_op_01(bnl_op_09_09[7:0]), .slf_op_04({net1141[0], net1141[1],
     net1141[2], net1141[3], net1141[4], net1141[5], net1141[6],
     net1141[7]}), .slf_op_03({net1131[0], net1131[1], net1131[2],
     net1131[3], net1131[4], net1131[5], net1131[6], net1131[7]}),
     .slf_op_01(slf_op_09_09[7:0]), .sp4_h_l_04({net1160[0],
     net1160[1], net1160[2], net1160[3], net1160[4], net1160[5],
     net1160[6], net1160[7], net1160[8], net1160[9], net1160[10],
     net1160[11], net1160[12], net1160[13], net1160[14], net1160[15],
     net1160[16], net1160[17], net1160[18], net1160[19], net1160[20],
     net1160[21], net1160[22], net1160[23], net1160[24], net1160[25],
     net1160[26], net1160[27], net1160[28], net1160[29], net1160[30],
     net1160[31], net1160[32], net1160[33], net1160[34], net1160[35],
     net1160[36], net1160[37], net1160[38], net1160[39], net1160[40],
     net1160[41], net1160[42], net1160[43], net1160[44], net1160[45],
     net1160[46], net1160[47]}), .carry_out(net960),
     .vdd_cntl(vdd_cntl_r[127:0]), .sp12_h_r_04({net962[0], net962[1],
     net962[2], net962[3], net962[4], net962[5], net962[6], net962[7],
     net962[8], net962[9], net962[10], net962[11], net962[12],
     net962[13], net962[14], net962[15], net962[16], net962[17],
     net962[18], net962[19], net962[20], net962[21], net962[22],
     net962[23]}), .sp12_h_r_03({net963[0], net963[1], net963[2],
     net963[3], net963[4], net963[5], net963[6], net963[7], net963[8],
     net963[9], net963[10], net963[11], net963[12], net963[13],
     net963[14], net963[15], net963[16], net963[17], net963[18],
     net963[19], net963[20], net963[21], net963[22], net963[23]}),
     .sp12_h_r_02({net964[0], net964[1], net964[2], net964[3],
     net964[4], net964[5], net964[6], net964[7], net964[8], net964[9],
     net964[10], net964[11], net964[12], net964[13], net964[14],
     net964[15], net964[16], net964[17], net964[18], net964[19],
     net964[20], net964[21], net964[22], net964[23]}),
     .sp12_h_r_01({net965[0], net965[1], net965[2], net965[3],
     net965[4], net965[5], net965[6], net965[7], net965[8], net965[9],
     net965[10], net965[11], net965[12], net965[13], net965[14],
     net965[15], net965[16], net965[17], net965[18], net965[19],
     net965[20], net965[21], net965[22], net965[23]}),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_09_09[47:0]), .sp4_r_v_b_04({net968[0],
     net968[1], net968[2], net968[3], net968[4], net968[5], net968[6],
     net968[7], net968[8], net968[9], net968[10], net968[11],
     net968[12], net968[13], net968[14], net968[15], net968[16],
     net968[17], net968[18], net968[19], net968[20], net968[21],
     net968[22], net968[23], net968[24], net968[25], net968[26],
     net968[27], net968[28], net968[29], net968[30], net968[31],
     net968[32], net968[33], net968[34], net968[35], net968[36],
     net968[37], net968[38], net968[39], net968[40], net968[41],
     net968[42], net968[43], net968[44], net968[45], net968[46],
     net968[47]}), .sp4_r_v_b_03({net969[0], net969[1], net969[2],
     net969[3], net969[4], net969[5], net969[6], net969[7], net969[8],
     net969[9], net969[10], net969[11], net969[12], net969[13],
     net969[14], net969[15], net969[16], net969[17], net969[18],
     net969[19], net969[20], net969[21], net969[22], net969[23],
     net969[24], net969[25], net969[26], net969[27], net969[28],
     net969[29], net969[30], net969[31], net969[32], net969[33],
     net969[34], net969[35], net969[36], net969[37], net969[38],
     net969[39], net969[40], net969[41], net969[42], net969[43],
     net969[44], net969[45], net969[46], net969[47]}),
     .sp4_r_v_b_02({net970[0], net970[1], net970[2], net970[3],
     net970[4], net970[5], net970[6], net970[7], net970[8], net970[9],
     net970[10], net970[11], net970[12], net970[13], net970[14],
     net970[15], net970[16], net970[17], net970[18], net970[19],
     net970[20], net970[21], net970[22], net970[23], net970[24],
     net970[25], net970[26], net970[27], net970[28], net970[29],
     net970[30], net970[31], net970[32], net970[33], net970[34],
     net970[35], net970[36], net970[37], net970[38], net970[39],
     net970[40], net970[41], net970[42], net970[43], net970[44],
     net970[45], net970[46], net970[47]}),
     .sp4_r_v_b_01(sp4_v_b_10_09[47:0]), .sp4_h_r_04({net972[0],
     net972[1], net972[2], net972[3], net972[4], net972[5], net972[6],
     net972[7], net972[8], net972[9], net972[10], net972[11],
     net972[12], net972[13], net972[14], net972[15], net972[16],
     net972[17], net972[18], net972[19], net972[20], net972[21],
     net972[22], net972[23], net972[24], net972[25], net972[26],
     net972[27], net972[28], net972[29], net972[30], net972[31],
     net972[32], net972[33], net972[34], net972[35], net972[36],
     net972[37], net972[38], net972[39], net972[40], net972[41],
     net972[42], net972[43], net972[44], net972[45], net972[46],
     net972[47]}), .sp4_h_r_03({net973[0], net973[1], net973[2],
     net973[3], net973[4], net973[5], net973[6], net973[7], net973[8],
     net973[9], net973[10], net973[11], net973[12], net973[13],
     net973[14], net973[15], net973[16], net973[17], net973[18],
     net973[19], net973[20], net973[21], net973[22], net973[23],
     net973[24], net973[25], net973[26], net973[27], net973[28],
     net973[29], net973[30], net973[31], net973[32], net973[33],
     net973[34], net973[35], net973[36], net973[37], net973[38],
     net973[39], net973[40], net973[41], net973[42], net973[43],
     net973[44], net973[45], net973[46], net973[47]}),
     .sp4_h_r_02({net974[0], net974[1], net974[2], net974[3],
     net974[4], net974[5], net974[6], net974[7], net974[8], net974[9],
     net974[10], net974[11], net974[12], net974[13], net974[14],
     net974[15], net974[16], net974[17], net974[18], net974[19],
     net974[20], net974[21], net974[22], net974[23], net974[24],
     net974[25], net974[26], net974[27], net974[28], net974[29],
     net974[30], net974[31], net974[32], net974[33], net974[34],
     net974[35], net974[36], net974[37], net974[38], net974[39],
     net974[40], net974[41], net974[42], net974[43], net974[44],
     net974[45], net974[46], net974[47]}), .sp4_h_r_01({net975[0],
     net975[1], net975[2], net975[3], net975[4], net975[5], net975[6],
     net975[7], net975[8], net975[9], net975[10], net975[11],
     net975[12], net975[13], net975[14], net975[15], net975[16],
     net975[17], net975[18], net975[19], net975[20], net975[21],
     net975[22], net975[23], net975[24], net975[25], net975[26],
     net975[27], net975[28], net975[29], net975[30], net975[31],
     net975[32], net975[33], net975[34], net975[35], net975[36],
     net975[37], net975[38], net975[39], net975[40], net975[41],
     net975[42], net975[43], net975[44], net975[45], net975[46],
     net975[47]}), .sp4_h_l_03({net1161[0], net1161[1], net1161[2],
     net1161[3], net1161[4], net1161[5], net1161[6], net1161[7],
     net1161[8], net1161[9], net1161[10], net1161[11], net1161[12],
     net1161[13], net1161[14], net1161[15], net1161[16], net1161[17],
     net1161[18], net1161[19], net1161[20], net1161[21], net1161[22],
     net1161[23], net1161[24], net1161[25], net1161[26], net1161[27],
     net1161[28], net1161[29], net1161[30], net1161[31], net1161[32],
     net1161[33], net1161[34], net1161[35], net1161[36], net1161[37],
     net1161[38], net1161[39], net1161[40], net1161[41], net1161[42],
     net1161[43], net1161[44], net1161[45], net1161[46], net1161[47]}),
     .sp4_h_l_02({net1162[0], net1162[1], net1162[2], net1162[3],
     net1162[4], net1162[5], net1162[6], net1162[7], net1162[8],
     net1162[9], net1162[10], net1162[11], net1162[12], net1162[13],
     net1162[14], net1162[15], net1162[16], net1162[17], net1162[18],
     net1162[19], net1162[20], net1162[21], net1162[22], net1162[23],
     net1162[24], net1162[25], net1162[26], net1162[27], net1162[28],
     net1162[29], net1162[30], net1162[31], net1162[32], net1162[33],
     net1162[34], net1162[35], net1162[36], net1162[37], net1162[38],
     net1162[39], net1162[40], net1162[41], net1162[42], net1162[43],
     net1162[44], net1162[45], net1162[46], net1162[47]}),
     .sp4_h_l_01({net1163[0], net1163[1], net1163[2], net1163[3],
     net1163[4], net1163[5], net1163[6], net1163[7], net1163[8],
     net1163[9], net1163[10], net1163[11], net1163[12], net1163[13],
     net1163[14], net1163[15], net1163[16], net1163[17], net1163[18],
     net1163[19], net1163[20], net1163[21], net1163[22], net1163[23],
     net1163[24], net1163[25], net1163[26], net1163[27], net1163[28],
     net1163[29], net1163[30], net1163[31], net1163[32], net1163[33],
     net1163[34], net1163[35], net1163[36], net1163[37], net1163[38],
     net1163[39], net1163[40], net1163[41], net1163[42], net1163[43],
     net1163[44], net1163[45], net1163[46], net1163[47]}),
     .bl(bl[161:108]), .bot_op_01(bot_op_09_09[7:0]),
     .sp12_h_l_01({net1153[0], net1153[1], net1153[2], net1153[3],
     net1153[4], net1153[5], net1153[6], net1153[7], net1153[8],
     net1153[9], net1153[10], net1153[11], net1153[12], net1153[13],
     net1153[14], net1153[15], net1153[16], net1153[17], net1153[18],
     net1153[19], net1153[20], net1153[21], net1153[22], net1153[23]}),
     .sp12_h_l_02({net1152[0], net1152[1], net1152[2], net1152[3],
     net1152[4], net1152[5], net1152[6], net1152[7], net1152[8],
     net1152[9], net1152[10], net1152[11], net1152[12], net1152[13],
     net1152[14], net1152[15], net1152[16], net1152[17], net1152[18],
     net1152[19], net1152[20], net1152[21], net1152[22], net1152[23]}),
     .sp12_h_l_03({net1151[0], net1151[1], net1151[2], net1151[3],
     net1151[4], net1151[5], net1151[6], net1151[7], net1151[8],
     net1151[9], net1151[10], net1151[11], net1151[12], net1151[13],
     net1151[14], net1151[15], net1151[16], net1151[17], net1151[18],
     net1151[19], net1151[20], net1151[21], net1151[22], net1151[23]}),
     .sp12_h_l_04({net1150[0], net1150[1], net1150[2], net1150[3],
     net1150[4], net1150[5], net1150[6], net1150[7], net1150[8],
     net1150[9], net1150[10], net1150[11], net1150[12], net1150[13],
     net1150[14], net1150[15], net1150[16], net1150[17], net1150[18],
     net1150[19], net1150[20], net1150[21], net1150[22], net1150[23]}),
     .sp4_v_b_04({net1156[0], net1156[1], net1156[2], net1156[3],
     net1156[4], net1156[5], net1156[6], net1156[7], net1156[8],
     net1156[9], net1156[10], net1156[11], net1156[12], net1156[13],
     net1156[14], net1156[15], net1156[16], net1156[17], net1156[18],
     net1156[19], net1156[20], net1156[21], net1156[22], net1156[23],
     net1156[24], net1156[25], net1156[26], net1156[27], net1156[28],
     net1156[29], net1156[30], net1156[31], net1156[32], net1156[33],
     net1156[34], net1156[35], net1156[36], net1156[37], net1156[38],
     net1156[39], net1156[40], net1156[41], net1156[42], net1156[43],
     net1156[44], net1156[45], net1156[46], net1156[47]}),
     .sp4_v_b_03({net1157[0], net1157[1], net1157[2], net1157[3],
     net1157[4], net1157[5], net1157[6], net1157[7], net1157[8],
     net1157[9], net1157[10], net1157[11], net1157[12], net1157[13],
     net1157[14], net1157[15], net1157[16], net1157[17], net1157[18],
     net1157[19], net1157[20], net1157[21], net1157[22], net1157[23],
     net1157[24], net1157[25], net1157[26], net1157[27], net1157[28],
     net1157[29], net1157[30], net1157[31], net1157[32], net1157[33],
     net1157[34], net1157[35], net1157[36], net1157[37], net1157[38],
     net1157[39], net1157[40], net1157[41], net1157[42], net1157[43],
     net1157[44], net1157[45], net1157[46], net1157[47]}),
     .sp4_v_b_02({net1158[0], net1158[1], net1158[2], net1158[3],
     net1158[4], net1158[5], net1158[6], net1158[7], net1158[8],
     net1158[9], net1158[10], net1158[11], net1158[12], net1158[13],
     net1158[14], net1158[15], net1158[16], net1158[17], net1158[18],
     net1158[19], net1158[20], net1158[21], net1158[22], net1158[23],
     net1158[24], net1158[25], net1158[26], net1158[27], net1158[28],
     net1158[29], net1158[30], net1158[31], net1158[32], net1158[33],
     net1158[34], net1158[35], net1158[36], net1158[37], net1158[38],
     net1158[39], net1158[40], net1158[41], net1158[42], net1158[43],
     net1158[44], net1158[45], net1158[46], net1158[47]}),
     .bnr_op_01(bnr_op_09_09[7:0]), .sp4_h_l_05({net1184[0],
     net1184[1], net1184[2], net1184[3], net1184[4], net1184[5],
     net1184[6], net1184[7], net1184[8], net1184[9], net1184[10],
     net1184[11], net1184[12], net1184[13], net1184[14], net1184[15],
     net1184[16], net1184[17], net1184[18], net1184[19], net1184[20],
     net1184[21], net1184[22], net1184[23], net1184[24], net1184[25],
     net1184[26], net1184[27], net1184[28], net1184[29], net1184[30],
     net1184[31], net1184[32], net1184[33], net1184[34], net1184[35],
     net1184[36], net1184[37], net1184[38], net1184[39], net1184[40],
     net1184[41], net1184[42], net1184[43], net1184[44], net1184[45],
     net1184[46], net1184[47]}), .sp4_h_l_06({net1183[0], net1183[1],
     net1183[2], net1183[3], net1183[4], net1183[5], net1183[6],
     net1183[7], net1183[8], net1183[9], net1183[10], net1183[11],
     net1183[12], net1183[13], net1183[14], net1183[15], net1183[16],
     net1183[17], net1183[18], net1183[19], net1183[20], net1183[21],
     net1183[22], net1183[23], net1183[24], net1183[25], net1183[26],
     net1183[27], net1183[28], net1183[29], net1183[30], net1183[31],
     net1183[32], net1183[33], net1183[34], net1183[35], net1183[36],
     net1183[37], net1183[38], net1183[39], net1183[40], net1183[41],
     net1183[42], net1183[43], net1183[44], net1183[45], net1183[46],
     net1183[47]}), .sp4_h_l_07({net1182[0], net1182[1], net1182[2],
     net1182[3], net1182[4], net1182[5], net1182[6], net1182[7],
     net1182[8], net1182[9], net1182[10], net1182[11], net1182[12],
     net1182[13], net1182[14], net1182[15], net1182[16], net1182[17],
     net1182[18], net1182[19], net1182[20], net1182[21], net1182[22],
     net1182[23], net1182[24], net1182[25], net1182[26], net1182[27],
     net1182[28], net1182[29], net1182[30], net1182[31], net1182[32],
     net1182[33], net1182[34], net1182[35], net1182[36], net1182[37],
     net1182[38], net1182[39], net1182[40], net1182[41], net1182[42],
     net1182[43], net1182[44], net1182[45], net1182[46], net1182[47]}),
     .sp4_h_l_08({net1181[0], net1181[1], net1181[2], net1181[3],
     net1181[4], net1181[5], net1181[6], net1181[7], net1181[8],
     net1181[9], net1181[10], net1181[11], net1181[12], net1181[13],
     net1181[14], net1181[15], net1181[16], net1181[17], net1181[18],
     net1181[19], net1181[20], net1181[21], net1181[22], net1181[23],
     net1181[24], net1181[25], net1181[26], net1181[27], net1181[28],
     net1181[29], net1181[30], net1181[31], net1181[32], net1181[33],
     net1181[34], net1181[35], net1181[36], net1181[37], net1181[38],
     net1181[39], net1181[40], net1181[41], net1181[42], net1181[43],
     net1181[44], net1181[45], net1181[46], net1181[47]}),
     .sp4_h_r_08({net993[0], net993[1], net993[2], net993[3],
     net993[4], net993[5], net993[6], net993[7], net993[8], net993[9],
     net993[10], net993[11], net993[12], net993[13], net993[14],
     net993[15], net993[16], net993[17], net993[18], net993[19],
     net993[20], net993[21], net993[22], net993[23], net993[24],
     net993[25], net993[26], net993[27], net993[28], net993[29],
     net993[30], net993[31], net993[32], net993[33], net993[34],
     net993[35], net993[36], net993[37], net993[38], net993[39],
     net993[40], net993[41], net993[42], net993[43], net993[44],
     net993[45], net993[46], net993[47]}), .sp4_h_r_07({net994[0],
     net994[1], net994[2], net994[3], net994[4], net994[5], net994[6],
     net994[7], net994[8], net994[9], net994[10], net994[11],
     net994[12], net994[13], net994[14], net994[15], net994[16],
     net994[17], net994[18], net994[19], net994[20], net994[21],
     net994[22], net994[23], net994[24], net994[25], net994[26],
     net994[27], net994[28], net994[29], net994[30], net994[31],
     net994[32], net994[33], net994[34], net994[35], net994[36],
     net994[37], net994[38], net994[39], net994[40], net994[41],
     net994[42], net994[43], net994[44], net994[45], net994[46],
     net994[47]}), .sp4_h_r_06({net995[0], net995[1], net995[2],
     net995[3], net995[4], net995[5], net995[6], net995[7], net995[8],
     net995[9], net995[10], net995[11], net995[12], net995[13],
     net995[14], net995[15], net995[16], net995[17], net995[18],
     net995[19], net995[20], net995[21], net995[22], net995[23],
     net995[24], net995[25], net995[26], net995[27], net995[28],
     net995[29], net995[30], net995[31], net995[32], net995[33],
     net995[34], net995[35], net995[36], net995[37], net995[38],
     net995[39], net995[40], net995[41], net995[42], net995[43],
     net995[44], net995[45], net995[46], net995[47]}),
     .sp4_h_r_05({net996[0], net996[1], net996[2], net996[3],
     net996[4], net996[5], net996[6], net996[7], net996[8], net996[9],
     net996[10], net996[11], net996[12], net996[13], net996[14],
     net996[15], net996[16], net996[17], net996[18], net996[19],
     net996[20], net996[21], net996[22], net996[23], net996[24],
     net996[25], net996[26], net996[27], net996[28], net996[29],
     net996[30], net996[31], net996[32], net996[33], net996[34],
     net996[35], net996[36], net996[37], net996[38], net996[39],
     net996[40], net996[41], net996[42], net996[43], net996[44],
     net996[45], net996[46], net996[47]}), .slf_op_05({net1192[0],
     net1192[1], net1192[2], net1192[3], net1192[4], net1192[5],
     net1192[6], net1192[7]}), .slf_op_06({net1191[0], net1191[1],
     net1191[2], net1191[3], net1191[4], net1191[5], net1191[6],
     net1191[7]}), .slf_op_07({net1190[0], net1190[1], net1190[2],
     net1190[3], net1190[4], net1190[5], net1190[6], net1190[7]}),
     .slf_op_08({net1189[0], net1189[1], net1189[2], net1189[3],
     net1189[4], net1189[5], net1189[6], net1189[7]}),
     .rgt_op_08({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7]}),
     .rgt_op_07({net1002[0], net1002[1], net1002[2], net1002[3],
     net1002[4], net1002[5], net1002[6], net1002[7]}),
     .rgt_op_06({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7]}),
     .rgt_op_05({net1004[0], net1004[1], net1004[2], net1004[3],
     net1004[4], net1004[5], net1004[6], net1004[7]}),
     .lft_op_08({net1283[0], net1283[1], net1283[2], net1283[3],
     net1283[4], net1283[5], net1283[6], net1283[7]}),
     .lft_op_07({net1284[0], net1284[1], net1284[2], net1284[3],
     net1284[4], net1284[5], net1284[6], net1284[7]}),
     .lft_op_06({net1285[0], net1285[1], net1285[2], net1285[3],
     net1285[4], net1285[5], net1285[6], net1285[7]}),
     .lft_op_05({net1286[0], net1286[1], net1286[2], net1286[3],
     net1286[4], net1286[5], net1286[6], net1286[7]}),
     .sp12_h_l_08({net1203[0], net1203[1], net1203[2], net1203[3],
     net1203[4], net1203[5], net1203[6], net1203[7], net1203[8],
     net1203[9], net1203[10], net1203[11], net1203[12], net1203[13],
     net1203[14], net1203[15], net1203[16], net1203[17], net1203[18],
     net1203[19], net1203[20], net1203[21], net1203[22], net1203[23]}),
     .sp12_h_l_07({net1202[0], net1202[1], net1202[2], net1202[3],
     net1202[4], net1202[5], net1202[6], net1202[7], net1202[8],
     net1202[9], net1202[10], net1202[11], net1202[12], net1202[13],
     net1202[14], net1202[15], net1202[16], net1202[17], net1202[18],
     net1202[19], net1202[20], net1202[21], net1202[22], net1202[23]}),
     .sp12_h_l_06({net1201[0], net1201[1], net1201[2], net1201[3],
     net1201[4], net1201[5], net1201[6], net1201[7], net1201[8],
     net1201[9], net1201[10], net1201[11], net1201[12], net1201[13],
     net1201[14], net1201[15], net1201[16], net1201[17], net1201[18],
     net1201[19], net1201[20], net1201[21], net1201[22], net1201[23]}),
     .sp12_h_r_05({net1012[0], net1012[1], net1012[2], net1012[3],
     net1012[4], net1012[5], net1012[6], net1012[7], net1012[8],
     net1012[9], net1012[10], net1012[11], net1012[12], net1012[13],
     net1012[14], net1012[15], net1012[16], net1012[17], net1012[18],
     net1012[19], net1012[20], net1012[21], net1012[22], net1012[23]}),
     .sp12_h_r_06({net1013[0], net1013[1], net1013[2], net1013[3],
     net1013[4], net1013[5], net1013[6], net1013[7], net1013[8],
     net1013[9], net1013[10], net1013[11], net1013[12], net1013[13],
     net1013[14], net1013[15], net1013[16], net1013[17], net1013[18],
     net1013[19], net1013[20], net1013[21], net1013[22], net1013[23]}),
     .sp12_h_r_07({net1014[0], net1014[1], net1014[2], net1014[3],
     net1014[4], net1014[5], net1014[6], net1014[7], net1014[8],
     net1014[9], net1014[10], net1014[11], net1014[12], net1014[13],
     net1014[14], net1014[15], net1014[16], net1014[17], net1014[18],
     net1014[19], net1014[20], net1014[21], net1014[22], net1014[23]}),
     .sp12_h_r_08({net1015[0], net1015[1], net1015[2], net1015[3],
     net1015[4], net1015[5], net1015[6], net1015[7], net1015[8],
     net1015[9], net1015[10], net1015[11], net1015[12], net1015[13],
     net1015[14], net1015[15], net1015[16], net1015[17], net1015[18],
     net1015[19], net1015[20], net1015[21], net1015[22], net1015[23]}),
     .sp12_h_l_05({net1200[0], net1200[1], net1200[2], net1200[3],
     net1200[4], net1200[5], net1200[6], net1200[7], net1200[8],
     net1200[9], net1200[10], net1200[11], net1200[12], net1200[13],
     net1200[14], net1200[15], net1200[16], net1200[17], net1200[18],
     net1200[19], net1200[20], net1200[21], net1200[22], net1200[23]}),
     .sp4_r_v_b_05({net1017[0], net1017[1], net1017[2], net1017[3],
     net1017[4], net1017[5], net1017[6], net1017[7], net1017[8],
     net1017[9], net1017[10], net1017[11], net1017[12], net1017[13],
     net1017[14], net1017[15], net1017[16], net1017[17], net1017[18],
     net1017[19], net1017[20], net1017[21], net1017[22], net1017[23],
     net1017[24], net1017[25], net1017[26], net1017[27], net1017[28],
     net1017[29], net1017[30], net1017[31], net1017[32], net1017[33],
     net1017[34], net1017[35], net1017[36], net1017[37], net1017[38],
     net1017[39], net1017[40], net1017[41], net1017[42], net1017[43],
     net1017[44], net1017[45], net1017[46], net1017[47]}),
     .sp4_r_v_b_06({net1018[0], net1018[1], net1018[2], net1018[3],
     net1018[4], net1018[5], net1018[6], net1018[7], net1018[8],
     net1018[9], net1018[10], net1018[11], net1018[12], net1018[13],
     net1018[14], net1018[15], net1018[16], net1018[17], net1018[18],
     net1018[19], net1018[20], net1018[21], net1018[22], net1018[23],
     net1018[24], net1018[25], net1018[26], net1018[27], net1018[28],
     net1018[29], net1018[30], net1018[31], net1018[32], net1018[33],
     net1018[34], net1018[35], net1018[36], net1018[37], net1018[38],
     net1018[39], net1018[40], net1018[41], net1018[42], net1018[43],
     net1018[44], net1018[45], net1018[46], net1018[47]}),
     .sp4_r_v_b_07({net1019[0], net1019[1], net1019[2], net1019[3],
     net1019[4], net1019[5], net1019[6], net1019[7], net1019[8],
     net1019[9], net1019[10], net1019[11], net1019[12], net1019[13],
     net1019[14], net1019[15], net1019[16], net1019[17], net1019[18],
     net1019[19], net1019[20], net1019[21], net1019[22], net1019[23],
     net1019[24], net1019[25], net1019[26], net1019[27], net1019[28],
     net1019[29], net1019[30], net1019[31], net1019[32], net1019[33],
     net1019[34], net1019[35], net1019[36], net1019[37], net1019[38],
     net1019[39], net1019[40], net1019[41], net1019[42], net1019[43],
     net1019[44], net1019[45], net1019[46], net1019[47]}),
     .sp4_r_v_b_08({net1020[0], net1020[1], net1020[2], net1020[3],
     net1020[4], net1020[5], net1020[6], net1020[7], net1020[8],
     net1020[9], net1020[10], net1020[11], net1020[12], net1020[13],
     net1020[14], net1020[15], net1020[16], net1020[17], net1020[18],
     net1020[19], net1020[20], net1020[21], net1020[22], net1020[23],
     net1020[24], net1020[25], net1020[26], net1020[27], net1020[28],
     net1020[29], net1020[30], net1020[31], net1020[32], net1020[33],
     net1020[34], net1020[35], net1020[36], net1020[37], net1020[38],
     net1020[39], net1020[40], net1020[41], net1020[42], net1020[43],
     net1020[44], net1020[45], net1020[46], net1020[47]}),
     .sp4_v_b_08({net1208[0], net1208[1], net1208[2], net1208[3],
     net1208[4], net1208[5], net1208[6], net1208[7], net1208[8],
     net1208[9], net1208[10], net1208[11], net1208[12], net1208[13],
     net1208[14], net1208[15], net1208[16], net1208[17], net1208[18],
     net1208[19], net1208[20], net1208[21], net1208[22], net1208[23],
     net1208[24], net1208[25], net1208[26], net1208[27], net1208[28],
     net1208[29], net1208[30], net1208[31], net1208[32], net1208[33],
     net1208[34], net1208[35], net1208[36], net1208[37], net1208[38],
     net1208[39], net1208[40], net1208[41], net1208[42], net1208[43],
     net1208[44], net1208[45], net1208[46], net1208[47]}),
     .sp4_v_b_07({net1207[0], net1207[1], net1207[2], net1207[3],
     net1207[4], net1207[5], net1207[6], net1207[7], net1207[8],
     net1207[9], net1207[10], net1207[11], net1207[12], net1207[13],
     net1207[14], net1207[15], net1207[16], net1207[17], net1207[18],
     net1207[19], net1207[20], net1207[21], net1207[22], net1207[23],
     net1207[24], net1207[25], net1207[26], net1207[27], net1207[28],
     net1207[29], net1207[30], net1207[31], net1207[32], net1207[33],
     net1207[34], net1207[35], net1207[36], net1207[37], net1207[38],
     net1207[39], net1207[40], net1207[41], net1207[42], net1207[43],
     net1207[44], net1207[45], net1207[46], net1207[47]}),
     .sp4_v_b_06({net1206[0], net1206[1], net1206[2], net1206[3],
     net1206[4], net1206[5], net1206[6], net1206[7], net1206[8],
     net1206[9], net1206[10], net1206[11], net1206[12], net1206[13],
     net1206[14], net1206[15], net1206[16], net1206[17], net1206[18],
     net1206[19], net1206[20], net1206[21], net1206[22], net1206[23],
     net1206[24], net1206[25], net1206[26], net1206[27], net1206[28],
     net1206[29], net1206[30], net1206[31], net1206[32], net1206[33],
     net1206[34], net1206[35], net1206[36], net1206[37], net1206[38],
     net1206[39], net1206[40], net1206[41], net1206[42], net1206[43],
     net1206[44], net1206[45], net1206[46], net1206[47]}),
     .sp4_v_b_05({net1205[0], net1205[1], net1205[2], net1205[3],
     net1205[4], net1205[5], net1205[6], net1205[7], net1205[8],
     net1205[9], net1205[10], net1205[11], net1205[12], net1205[13],
     net1205[14], net1205[15], net1205[16], net1205[17], net1205[18],
     net1205[19], net1205[20], net1205[21], net1205[22], net1205[23],
     net1205[24], net1205[25], net1205[26], net1205[27], net1205[28],
     net1205[29], net1205[30], net1205[31], net1205[32], net1205[33],
     net1205[34], net1205[35], net1205[36], net1205[37], net1205[38],
     net1205[39], net1205[40], net1205[41], net1205[42], net1205[43],
     net1205[44], net1205[45], net1205[46], net1205[47]}),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .wl(wl_r[127:0]), .sp12_v_t_08({net1028[0], net1028[1],
     net1028[2], net1028[3], net1028[4], net1028[5], net1028[6],
     net1028[7], net1028[8], net1028[9], net1028[10], net1028[11],
     net1028[12], net1028[13], net1028[14], net1028[15], net1028[16],
     net1028[17], net1028[18], net1028[19], net1028[20], net1028[21],
     net1028[22], net1028[23]}), .tnr_op_08({slf_op_10_17[3],
     slf_op_10_17[2], slf_op_10_17[1], slf_op_10_17[0],
     slf_op_10_17[3], slf_op_10_17[2], slf_op_10_17[1],
     slf_op_10_17[0]}), .top_op_08({slf_op_09_17[3], slf_op_09_17[2],
     slf_op_09_17[1], slf_op_09_17[0], slf_op_09_17[3],
     slf_op_09_17[2], slf_op_09_17[1], slf_op_09_17[0]}),
     .tnl_op_08({slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0], slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0]}), .sp4_v_t_08({net1032[0],
     net1032[1], net1032[2], net1032[3], net1032[4], net1032[5],
     net1032[6], net1032[7], net1032[8], net1032[9], net1032[10],
     net1032[11], net1032[12], net1032[13], net1032[14], net1032[15],
     net1032[16], net1032[17], net1032[18], net1032[19], net1032[20],
     net1032[21], net1032[22], net1032[23], net1032[24], net1032[25],
     net1032[26], net1032[27], net1032[28], net1032[29], net1032[30],
     net1032[31], net1032[32], net1032[33], net1032[34], net1032[35],
     net1032[36], net1032[37], net1032[38], net1032[39], net1032[40],
     net1032[41], net1032[42], net1032[43], net1032[44], net1032[45],
     net1032[46], net1032[47]}), .lc_bot(lc_bot_09_09),
     .op_vic(net1034), .sp12_v_b_01(sp12_v_b_09_09[23:0]),
     .glb_netwk_t({net1036[0], net1036[1], net1036[2], net1036[3],
     net1036[4], net1036[5], net1036[6], net1036[7]}));
lt_1x8_top_ice1f I_lt_col_t11 ( .glb_netwk_b({net01038[0], net01038[1],
     net01038[2], net01038[3], net01038[4], net01038[5], net01038[6],
     net01038[7]}), .rgt_op_03({net1037[0], net1037[1], net1037[2],
     net1037[3], net1037[4], net1037[5], net1037[6], net1037[7]}),
     .slf_op_02({net1410[0], net1410[1], net1410[2], net1410[3],
     net1410[4], net1410[5], net1410[6], net1410[7]}),
     .rgt_op_02({net1039[0], net1039[1], net1039[2], net1039[3],
     net1039[4], net1039[5], net1039[6], net1039[7]}),
     .rgt_op_01(slf_op_12_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04({net953[0], net953[1], net953[2], net953[3], net953[4],
     net953[5], net953[6], net953[7]}), .lft_op_03({net943[0],
     net943[1], net943[2], net943[3], net943[4], net943[5], net943[6],
     net943[7]}), .lft_op_02({net945[0], net945[1], net945[2],
     net945[3], net945[4], net945[5], net945[6], net945[7]}),
     .lft_op_01(slf_op_10_09[7:0]), .rgt_op_04({net1047[0], net1047[1],
     net1047[2], net1047[3], net1047[4], net1047[5], net1047[6],
     net1047[7]}), .carry_in(carry_in_11_09),
     .bnl_op_01(bnl_op_11_09[7:0]), .slf_op_04({net1408[0], net1408[1],
     net1408[2], net1408[3], net1408[4], net1408[5], net1408[6],
     net1408[7]}), .slf_op_03({net1409[0], net1409[1], net1409[2],
     net1409[3], net1409[4], net1409[5], net1409[6], net1409[7]}),
     .slf_op_01(slf_op_11_09[7:0]), .sp4_h_l_04({net1429[0],
     net1429[1], net1429[2], net1429[3], net1429[4], net1429[5],
     net1429[6], net1429[7], net1429[8], net1429[9], net1429[10],
     net1429[11], net1429[12], net1429[13], net1429[14], net1429[15],
     net1429[16], net1429[17], net1429[18], net1429[19], net1429[20],
     net1429[21], net1429[22], net1429[23], net1429[24], net1429[25],
     net1429[26], net1429[27], net1429[28], net1429[29], net1429[30],
     net1429[31], net1429[32], net1429[33], net1429[34], net1429[35],
     net1429[36], net1429[37], net1429[38], net1429[39], net1429[40],
     net1429[41], net1429[42], net1429[43], net1429[44], net1429[45],
     net1429[46], net1429[47]}), .carry_out(net1054),
     .vdd_cntl(vdd_cntl_r[127:0]), .sp12_h_r_04({net1056[0],
     net1056[1], net1056[2], net1056[3], net1056[4], net1056[5],
     net1056[6], net1056[7], net1056[8], net1056[9], net1056[10],
     net1056[11], net1056[12], net1056[13], net1056[14], net1056[15],
     net1056[16], net1056[17], net1056[18], net1056[19], net1056[20],
     net1056[21], net1056[22], net1056[23]}), .sp12_h_r_03({net1057[0],
     net1057[1], net1057[2], net1057[3], net1057[4], net1057[5],
     net1057[6], net1057[7], net1057[8], net1057[9], net1057[10],
     net1057[11], net1057[12], net1057[13], net1057[14], net1057[15],
     net1057[16], net1057[17], net1057[18], net1057[19], net1057[20],
     net1057[21], net1057[22], net1057[23]}), .sp12_h_r_02({net1058[0],
     net1058[1], net1058[2], net1058[3], net1058[4], net1058[5],
     net1058[6], net1058[7], net1058[8], net1058[9], net1058[10],
     net1058[11], net1058[12], net1058[13], net1058[14], net1058[15],
     net1058[16], net1058[17], net1058[18], net1058[19], net1058[20],
     net1058[21], net1058[22], net1058[23]}), .sp12_h_r_01({net1059[0],
     net1059[1], net1059[2], net1059[3], net1059[4], net1059[5],
     net1059[6], net1059[7], net1059[8], net1059[9], net1059[10],
     net1059[11], net1059[12], net1059[13], net1059[14], net1059[15],
     net1059[16], net1059[17], net1059[18], net1059[19], net1059[20],
     net1059[21], net1059[22], net1059[23]}),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_11_09[47:0]), .sp4_r_v_b_04({net1062[0],
     net1062[1], net1062[2], net1062[3], net1062[4], net1062[5],
     net1062[6], net1062[7], net1062[8], net1062[9], net1062[10],
     net1062[11], net1062[12], net1062[13], net1062[14], net1062[15],
     net1062[16], net1062[17], net1062[18], net1062[19], net1062[20],
     net1062[21], net1062[22], net1062[23], net1062[24], net1062[25],
     net1062[26], net1062[27], net1062[28], net1062[29], net1062[30],
     net1062[31], net1062[32], net1062[33], net1062[34], net1062[35],
     net1062[36], net1062[37], net1062[38], net1062[39], net1062[40],
     net1062[41], net1062[42], net1062[43], net1062[44], net1062[45],
     net1062[46], net1062[47]}), .sp4_r_v_b_03({net1063[0], net1063[1],
     net1063[2], net1063[3], net1063[4], net1063[5], net1063[6],
     net1063[7], net1063[8], net1063[9], net1063[10], net1063[11],
     net1063[12], net1063[13], net1063[14], net1063[15], net1063[16],
     net1063[17], net1063[18], net1063[19], net1063[20], net1063[21],
     net1063[22], net1063[23], net1063[24], net1063[25], net1063[26],
     net1063[27], net1063[28], net1063[29], net1063[30], net1063[31],
     net1063[32], net1063[33], net1063[34], net1063[35], net1063[36],
     net1063[37], net1063[38], net1063[39], net1063[40], net1063[41],
     net1063[42], net1063[43], net1063[44], net1063[45], net1063[46],
     net1063[47]}), .sp4_r_v_b_02({net1064[0], net1064[1], net1064[2],
     net1064[3], net1064[4], net1064[5], net1064[6], net1064[7],
     net1064[8], net1064[9], net1064[10], net1064[11], net1064[12],
     net1064[13], net1064[14], net1064[15], net1064[16], net1064[17],
     net1064[18], net1064[19], net1064[20], net1064[21], net1064[22],
     net1064[23], net1064[24], net1064[25], net1064[26], net1064[27],
     net1064[28], net1064[29], net1064[30], net1064[31], net1064[32],
     net1064[33], net1064[34], net1064[35], net1064[36], net1064[37],
     net1064[38], net1064[39], net1064[40], net1064[41], net1064[42],
     net1064[43], net1064[44], net1064[45], net1064[46], net1064[47]}),
     .sp4_r_v_b_01(sp4_v_b_12_09[47:0]), .sp4_h_r_04({net1066[0],
     net1066[1], net1066[2], net1066[3], net1066[4], net1066[5],
     net1066[6], net1066[7], net1066[8], net1066[9], net1066[10],
     net1066[11], net1066[12], net1066[13], net1066[14], net1066[15],
     net1066[16], net1066[17], net1066[18], net1066[19], net1066[20],
     net1066[21], net1066[22], net1066[23], net1066[24], net1066[25],
     net1066[26], net1066[27], net1066[28], net1066[29], net1066[30],
     net1066[31], net1066[32], net1066[33], net1066[34], net1066[35],
     net1066[36], net1066[37], net1066[38], net1066[39], net1066[40],
     net1066[41], net1066[42], net1066[43], net1066[44], net1066[45],
     net1066[46], net1066[47]}), .sp4_h_r_03({net1067[0], net1067[1],
     net1067[2], net1067[3], net1067[4], net1067[5], net1067[6],
     net1067[7], net1067[8], net1067[9], net1067[10], net1067[11],
     net1067[12], net1067[13], net1067[14], net1067[15], net1067[16],
     net1067[17], net1067[18], net1067[19], net1067[20], net1067[21],
     net1067[22], net1067[23], net1067[24], net1067[25], net1067[26],
     net1067[27], net1067[28], net1067[29], net1067[30], net1067[31],
     net1067[32], net1067[33], net1067[34], net1067[35], net1067[36],
     net1067[37], net1067[38], net1067[39], net1067[40], net1067[41],
     net1067[42], net1067[43], net1067[44], net1067[45], net1067[46],
     net1067[47]}), .sp4_h_r_02({net1068[0], net1068[1], net1068[2],
     net1068[3], net1068[4], net1068[5], net1068[6], net1068[7],
     net1068[8], net1068[9], net1068[10], net1068[11], net1068[12],
     net1068[13], net1068[14], net1068[15], net1068[16], net1068[17],
     net1068[18], net1068[19], net1068[20], net1068[21], net1068[22],
     net1068[23], net1068[24], net1068[25], net1068[26], net1068[27],
     net1068[28], net1068[29], net1068[30], net1068[31], net1068[32],
     net1068[33], net1068[34], net1068[35], net1068[36], net1068[37],
     net1068[38], net1068[39], net1068[40], net1068[41], net1068[42],
     net1068[43], net1068[44], net1068[45], net1068[46], net1068[47]}),
     .sp4_h_r_01({net1069[0], net1069[1], net1069[2], net1069[3],
     net1069[4], net1069[5], net1069[6], net1069[7], net1069[8],
     net1069[9], net1069[10], net1069[11], net1069[12], net1069[13],
     net1069[14], net1069[15], net1069[16], net1069[17], net1069[18],
     net1069[19], net1069[20], net1069[21], net1069[22], net1069[23],
     net1069[24], net1069[25], net1069[26], net1069[27], net1069[28],
     net1069[29], net1069[30], net1069[31], net1069[32], net1069[33],
     net1069[34], net1069[35], net1069[36], net1069[37], net1069[38],
     net1069[39], net1069[40], net1069[41], net1069[42], net1069[43],
     net1069[44], net1069[45], net1069[46], net1069[47]}),
     .sp4_h_l_03({net1428[0], net1428[1], net1428[2], net1428[3],
     net1428[4], net1428[5], net1428[6], net1428[7], net1428[8],
     net1428[9], net1428[10], net1428[11], net1428[12], net1428[13],
     net1428[14], net1428[15], net1428[16], net1428[17], net1428[18],
     net1428[19], net1428[20], net1428[21], net1428[22], net1428[23],
     net1428[24], net1428[25], net1428[26], net1428[27], net1428[28],
     net1428[29], net1428[30], net1428[31], net1428[32], net1428[33],
     net1428[34], net1428[35], net1428[36], net1428[37], net1428[38],
     net1428[39], net1428[40], net1428[41], net1428[42], net1428[43],
     net1428[44], net1428[45], net1428[46], net1428[47]}),
     .sp4_h_l_02({net1427[0], net1427[1], net1427[2], net1427[3],
     net1427[4], net1427[5], net1427[6], net1427[7], net1427[8],
     net1427[9], net1427[10], net1427[11], net1427[12], net1427[13],
     net1427[14], net1427[15], net1427[16], net1427[17], net1427[18],
     net1427[19], net1427[20], net1427[21], net1427[22], net1427[23],
     net1427[24], net1427[25], net1427[26], net1427[27], net1427[28],
     net1427[29], net1427[30], net1427[31], net1427[32], net1427[33],
     net1427[34], net1427[35], net1427[36], net1427[37], net1427[38],
     net1427[39], net1427[40], net1427[41], net1427[42], net1427[43],
     net1427[44], net1427[45], net1427[46], net1427[47]}),
     .sp4_h_l_01({net1383[0], net1383[1], net1383[2], net1383[3],
     net1383[4], net1383[5], net1383[6], net1383[7], net1383[8],
     net1383[9], net1383[10], net1383[11], net1383[12], net1383[13],
     net1383[14], net1383[15], net1383[16], net1383[17], net1383[18],
     net1383[19], net1383[20], net1383[21], net1383[22], net1383[23],
     net1383[24], net1383[25], net1383[26], net1383[27], net1383[28],
     net1383[29], net1383[30], net1383[31], net1383[32], net1383[33],
     net1383[34], net1383[35], net1383[36], net1383[37], net1383[38],
     net1383[39], net1383[40], net1383[41], net1383[42], net1383[43],
     net1383[44], net1383[45], net1383[46], net1383[47]}),
     .bl(bl[257:204]), .bot_op_01(bot_op_11_09[7:0]),
     .sp12_h_l_01({net1377[0], net1377[1], net1377[2], net1377[3],
     net1377[4], net1377[5], net1377[6], net1377[7], net1377[8],
     net1377[9], net1377[10], net1377[11], net1377[12], net1377[13],
     net1377[14], net1377[15], net1377[16], net1377[17], net1377[18],
     net1377[19], net1377[20], net1377[21], net1377[22], net1377[23]}),
     .sp12_h_l_02({net1385[0], net1385[1], net1385[2], net1385[3],
     net1385[4], net1385[5], net1385[6], net1385[7], net1385[8],
     net1385[9], net1385[10], net1385[11], net1385[12], net1385[13],
     net1385[14], net1385[15], net1385[16], net1385[17], net1385[18],
     net1385[19], net1385[20], net1385[21], net1385[22], net1385[23]}),
     .sp12_h_l_03({net1341[0], net1341[1], net1341[2], net1341[3],
     net1341[4], net1341[5], net1341[6], net1341[7], net1341[8],
     net1341[9], net1341[10], net1341[11], net1341[12], net1341[13],
     net1341[14], net1341[15], net1341[16], net1341[17], net1341[18],
     net1341[19], net1341[20], net1341[21], net1341[22], net1341[23]}),
     .sp12_h_l_04({net1386[0], net1386[1], net1386[2], net1386[3],
     net1386[4], net1386[5], net1386[6], net1386[7], net1386[8],
     net1386[9], net1386[10], net1386[11], net1386[12], net1386[13],
     net1386[14], net1386[15], net1386[16], net1386[17], net1386[18],
     net1386[19], net1386[20], net1386[21], net1386[22], net1386[23]}),
     .sp4_v_b_04({net1365[0], net1365[1], net1365[2], net1365[3],
     net1365[4], net1365[5], net1365[6], net1365[7], net1365[8],
     net1365[9], net1365[10], net1365[11], net1365[12], net1365[13],
     net1365[14], net1365[15], net1365[16], net1365[17], net1365[18],
     net1365[19], net1365[20], net1365[21], net1365[22], net1365[23],
     net1365[24], net1365[25], net1365[26], net1365[27], net1365[28],
     net1365[29], net1365[30], net1365[31], net1365[32], net1365[33],
     net1365[34], net1365[35], net1365[36], net1365[37], net1365[38],
     net1365[39], net1365[40], net1365[41], net1365[42], net1365[43],
     net1365[44], net1365[45], net1365[46], net1365[47]}),
     .sp4_v_b_03({net1361[0], net1361[1], net1361[2], net1361[3],
     net1361[4], net1361[5], net1361[6], net1361[7], net1361[8],
     net1361[9], net1361[10], net1361[11], net1361[12], net1361[13],
     net1361[14], net1361[15], net1361[16], net1361[17], net1361[18],
     net1361[19], net1361[20], net1361[21], net1361[22], net1361[23],
     net1361[24], net1361[25], net1361[26], net1361[27], net1361[28],
     net1361[29], net1361[30], net1361[31], net1361[32], net1361[33],
     net1361[34], net1361[35], net1361[36], net1361[37], net1361[38],
     net1361[39], net1361[40], net1361[41], net1361[42], net1361[43],
     net1361[44], net1361[45], net1361[46], net1361[47]}),
     .sp4_v_b_02({net1372[0], net1372[1], net1372[2], net1372[3],
     net1372[4], net1372[5], net1372[6], net1372[7], net1372[8],
     net1372[9], net1372[10], net1372[11], net1372[12], net1372[13],
     net1372[14], net1372[15], net1372[16], net1372[17], net1372[18],
     net1372[19], net1372[20], net1372[21], net1372[22], net1372[23],
     net1372[24], net1372[25], net1372[26], net1372[27], net1372[28],
     net1372[29], net1372[30], net1372[31], net1372[32], net1372[33],
     net1372[34], net1372[35], net1372[36], net1372[37], net1372[38],
     net1372[39], net1372[40], net1372[41], net1372[42], net1372[43],
     net1372[44], net1372[45], net1372[46], net1372[47]}),
     .bnr_op_01(bnr_op_11_09[7:0]), .sp4_h_l_05({net1430[0],
     net1430[1], net1430[2], net1430[3], net1430[4], net1430[5],
     net1430[6], net1430[7], net1430[8], net1430[9], net1430[10],
     net1430[11], net1430[12], net1430[13], net1430[14], net1430[15],
     net1430[16], net1430[17], net1430[18], net1430[19], net1430[20],
     net1430[21], net1430[22], net1430[23], net1430[24], net1430[25],
     net1430[26], net1430[27], net1430[28], net1430[29], net1430[30],
     net1430[31], net1430[32], net1430[33], net1430[34], net1430[35],
     net1430[36], net1430[37], net1430[38], net1430[39], net1430[40],
     net1430[41], net1430[42], net1430[43], net1430[44], net1430[45],
     net1430[46], net1430[47]}), .sp4_h_l_06({net1431[0], net1431[1],
     net1431[2], net1431[3], net1431[4], net1431[5], net1431[6],
     net1431[7], net1431[8], net1431[9], net1431[10], net1431[11],
     net1431[12], net1431[13], net1431[14], net1431[15], net1431[16],
     net1431[17], net1431[18], net1431[19], net1431[20], net1431[21],
     net1431[22], net1431[23], net1431[24], net1431[25], net1431[26],
     net1431[27], net1431[28], net1431[29], net1431[30], net1431[31],
     net1431[32], net1431[33], net1431[34], net1431[35], net1431[36],
     net1431[37], net1431[38], net1431[39], net1431[40], net1431[41],
     net1431[42], net1431[43], net1431[44], net1431[45], net1431[46],
     net1431[47]}), .sp4_h_l_07({net1432[0], net1432[1], net1432[2],
     net1432[3], net1432[4], net1432[5], net1432[6], net1432[7],
     net1432[8], net1432[9], net1432[10], net1432[11], net1432[12],
     net1432[13], net1432[14], net1432[15], net1432[16], net1432[17],
     net1432[18], net1432[19], net1432[20], net1432[21], net1432[22],
     net1432[23], net1432[24], net1432[25], net1432[26], net1432[27],
     net1432[28], net1432[29], net1432[30], net1432[31], net1432[32],
     net1432[33], net1432[34], net1432[35], net1432[36], net1432[37],
     net1432[38], net1432[39], net1432[40], net1432[41], net1432[42],
     net1432[43], net1432[44], net1432[45], net1432[46], net1432[47]}),
     .sp4_h_l_08({net1368[0], net1368[1], net1368[2], net1368[3],
     net1368[4], net1368[5], net1368[6], net1368[7], net1368[8],
     net1368[9], net1368[10], net1368[11], net1368[12], net1368[13],
     net1368[14], net1368[15], net1368[16], net1368[17], net1368[18],
     net1368[19], net1368[20], net1368[21], net1368[22], net1368[23],
     net1368[24], net1368[25], net1368[26], net1368[27], net1368[28],
     net1368[29], net1368[30], net1368[31], net1368[32], net1368[33],
     net1368[34], net1368[35], net1368[36], net1368[37], net1368[38],
     net1368[39], net1368[40], net1368[41], net1368[42], net1368[43],
     net1368[44], net1368[45], net1368[46], net1368[47]}),
     .sp4_h_r_08({net1087[0], net1087[1], net1087[2], net1087[3],
     net1087[4], net1087[5], net1087[6], net1087[7], net1087[8],
     net1087[9], net1087[10], net1087[11], net1087[12], net1087[13],
     net1087[14], net1087[15], net1087[16], net1087[17], net1087[18],
     net1087[19], net1087[20], net1087[21], net1087[22], net1087[23],
     net1087[24], net1087[25], net1087[26], net1087[27], net1087[28],
     net1087[29], net1087[30], net1087[31], net1087[32], net1087[33],
     net1087[34], net1087[35], net1087[36], net1087[37], net1087[38],
     net1087[39], net1087[40], net1087[41], net1087[42], net1087[43],
     net1087[44], net1087[45], net1087[46], net1087[47]}),
     .sp4_h_r_07({net1088[0], net1088[1], net1088[2], net1088[3],
     net1088[4], net1088[5], net1088[6], net1088[7], net1088[8],
     net1088[9], net1088[10], net1088[11], net1088[12], net1088[13],
     net1088[14], net1088[15], net1088[16], net1088[17], net1088[18],
     net1088[19], net1088[20], net1088[21], net1088[22], net1088[23],
     net1088[24], net1088[25], net1088[26], net1088[27], net1088[28],
     net1088[29], net1088[30], net1088[31], net1088[32], net1088[33],
     net1088[34], net1088[35], net1088[36], net1088[37], net1088[38],
     net1088[39], net1088[40], net1088[41], net1088[42], net1088[43],
     net1088[44], net1088[45], net1088[46], net1088[47]}),
     .sp4_h_r_06({net1089[0], net1089[1], net1089[2], net1089[3],
     net1089[4], net1089[5], net1089[6], net1089[7], net1089[8],
     net1089[9], net1089[10], net1089[11], net1089[12], net1089[13],
     net1089[14], net1089[15], net1089[16], net1089[17], net1089[18],
     net1089[19], net1089[20], net1089[21], net1089[22], net1089[23],
     net1089[24], net1089[25], net1089[26], net1089[27], net1089[28],
     net1089[29], net1089[30], net1089[31], net1089[32], net1089[33],
     net1089[34], net1089[35], net1089[36], net1089[37], net1089[38],
     net1089[39], net1089[40], net1089[41], net1089[42], net1089[43],
     net1089[44], net1089[45], net1089[46], net1089[47]}),
     .sp4_h_r_05({net1090[0], net1090[1], net1090[2], net1090[3],
     net1090[4], net1090[5], net1090[6], net1090[7], net1090[8],
     net1090[9], net1090[10], net1090[11], net1090[12], net1090[13],
     net1090[14], net1090[15], net1090[16], net1090[17], net1090[18],
     net1090[19], net1090[20], net1090[21], net1090[22], net1090[23],
     net1090[24], net1090[25], net1090[26], net1090[27], net1090[28],
     net1090[29], net1090[30], net1090[31], net1090[32], net1090[33],
     net1090[34], net1090[35], net1090[36], net1090[37], net1090[38],
     net1090[39], net1090[40], net1090[41], net1090[42], net1090[43],
     net1090[44], net1090[45], net1090[46], net1090[47]}),
     .slf_op_05({net1407[0], net1407[1], net1407[2], net1407[3],
     net1407[4], net1407[5], net1407[6], net1407[7]}),
     .slf_op_06({net1406[0], net1406[1], net1406[2], net1406[3],
     net1406[4], net1406[5], net1406[6], net1406[7]}),
     .slf_op_07({net1405[0], net1405[1], net1405[2], net1405[3],
     net1405[4], net1405[5], net1405[6], net1405[7]}),
     .slf_op_08({net1404[0], net1404[1], net1404[2], net1404[3],
     net1404[4], net1404[5], net1404[6], net1404[7]}),
     .rgt_op_08({net1095[0], net1095[1], net1095[2], net1095[3],
     net1095[4], net1095[5], net1095[6], net1095[7]}),
     .rgt_op_07({net1096[0], net1096[1], net1096[2], net1096[3],
     net1096[4], net1096[5], net1096[6], net1096[7]}),
     .rgt_op_06({net1097[0], net1097[1], net1097[2], net1097[3],
     net1097[4], net1097[5], net1097[6], net1097[7]}),
     .rgt_op_05({net1098[0], net1098[1], net1098[2], net1098[3],
     net1098[4], net1098[5], net1098[6], net1098[7]}),
     .lft_op_08({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7]}),
     .lft_op_07({net1002[0], net1002[1], net1002[2], net1002[3],
     net1002[4], net1002[5], net1002[6], net1002[7]}),
     .lft_op_06({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7]}),
     .lft_op_05({net1004[0], net1004[1], net1004[2], net1004[3],
     net1004[4], net1004[5], net1004[6], net1004[7]}),
     .sp12_h_l_08({net1358[0], net1358[1], net1358[2], net1358[3],
     net1358[4], net1358[5], net1358[6], net1358[7], net1358[8],
     net1358[9], net1358[10], net1358[11], net1358[12], net1358[13],
     net1358[14], net1358[15], net1358[16], net1358[17], net1358[18],
     net1358[19], net1358[20], net1358[21], net1358[22], net1358[23]}),
     .sp12_h_l_07({net1353[0], net1353[1], net1353[2], net1353[3],
     net1353[4], net1353[5], net1353[6], net1353[7], net1353[8],
     net1353[9], net1353[10], net1353[11], net1353[12], net1353[13],
     net1353[14], net1353[15], net1353[16], net1353[17], net1353[18],
     net1353[19], net1353[20], net1353[21], net1353[22], net1353[23]}),
     .sp12_h_l_06({net1355[0], net1355[1], net1355[2], net1355[3],
     net1355[4], net1355[5], net1355[6], net1355[7], net1355[8],
     net1355[9], net1355[10], net1355[11], net1355[12], net1355[13],
     net1355[14], net1355[15], net1355[16], net1355[17], net1355[18],
     net1355[19], net1355[20], net1355[21], net1355[22], net1355[23]}),
     .sp12_h_r_05({net1106[0], net1106[1], net1106[2], net1106[3],
     net1106[4], net1106[5], net1106[6], net1106[7], net1106[8],
     net1106[9], net1106[10], net1106[11], net1106[12], net1106[13],
     net1106[14], net1106[15], net1106[16], net1106[17], net1106[18],
     net1106[19], net1106[20], net1106[21], net1106[22], net1106[23]}),
     .sp12_h_r_06({net1107[0], net1107[1], net1107[2], net1107[3],
     net1107[4], net1107[5], net1107[6], net1107[7], net1107[8],
     net1107[9], net1107[10], net1107[11], net1107[12], net1107[13],
     net1107[14], net1107[15], net1107[16], net1107[17], net1107[18],
     net1107[19], net1107[20], net1107[21], net1107[22], net1107[23]}),
     .sp12_h_r_07({net1108[0], net1108[1], net1108[2], net1108[3],
     net1108[4], net1108[5], net1108[6], net1108[7], net1108[8],
     net1108[9], net1108[10], net1108[11], net1108[12], net1108[13],
     net1108[14], net1108[15], net1108[16], net1108[17], net1108[18],
     net1108[19], net1108[20], net1108[21], net1108[22], net1108[23]}),
     .sp12_h_r_08({net1109[0], net1109[1], net1109[2], net1109[3],
     net1109[4], net1109[5], net1109[6], net1109[7], net1109[8],
     net1109[9], net1109[10], net1109[11], net1109[12], net1109[13],
     net1109[14], net1109[15], net1109[16], net1109[17], net1109[18],
     net1109[19], net1109[20], net1109[21], net1109[22], net1109[23]}),
     .sp12_h_l_05({net1357[0], net1357[1], net1357[2], net1357[3],
     net1357[4], net1357[5], net1357[6], net1357[7], net1357[8],
     net1357[9], net1357[10], net1357[11], net1357[12], net1357[13],
     net1357[14], net1357[15], net1357[16], net1357[17], net1357[18],
     net1357[19], net1357[20], net1357[21], net1357[22], net1357[23]}),
     .sp4_r_v_b_05({net1111[0], net1111[1], net1111[2], net1111[3],
     net1111[4], net1111[5], net1111[6], net1111[7], net1111[8],
     net1111[9], net1111[10], net1111[11], net1111[12], net1111[13],
     net1111[14], net1111[15], net1111[16], net1111[17], net1111[18],
     net1111[19], net1111[20], net1111[21], net1111[22], net1111[23],
     net1111[24], net1111[25], net1111[26], net1111[27], net1111[28],
     net1111[29], net1111[30], net1111[31], net1111[32], net1111[33],
     net1111[34], net1111[35], net1111[36], net1111[37], net1111[38],
     net1111[39], net1111[40], net1111[41], net1111[42], net1111[43],
     net1111[44], net1111[45], net1111[46], net1111[47]}),
     .sp4_r_v_b_06({net1112[0], net1112[1], net1112[2], net1112[3],
     net1112[4], net1112[5], net1112[6], net1112[7], net1112[8],
     net1112[9], net1112[10], net1112[11], net1112[12], net1112[13],
     net1112[14], net1112[15], net1112[16], net1112[17], net1112[18],
     net1112[19], net1112[20], net1112[21], net1112[22], net1112[23],
     net1112[24], net1112[25], net1112[26], net1112[27], net1112[28],
     net1112[29], net1112[30], net1112[31], net1112[32], net1112[33],
     net1112[34], net1112[35], net1112[36], net1112[37], net1112[38],
     net1112[39], net1112[40], net1112[41], net1112[42], net1112[43],
     net1112[44], net1112[45], net1112[46], net1112[47]}),
     .sp4_r_v_b_07({net1113[0], net1113[1], net1113[2], net1113[3],
     net1113[4], net1113[5], net1113[6], net1113[7], net1113[8],
     net1113[9], net1113[10], net1113[11], net1113[12], net1113[13],
     net1113[14], net1113[15], net1113[16], net1113[17], net1113[18],
     net1113[19], net1113[20], net1113[21], net1113[22], net1113[23],
     net1113[24], net1113[25], net1113[26], net1113[27], net1113[28],
     net1113[29], net1113[30], net1113[31], net1113[32], net1113[33],
     net1113[34], net1113[35], net1113[36], net1113[37], net1113[38],
     net1113[39], net1113[40], net1113[41], net1113[42], net1113[43],
     net1113[44], net1113[45], net1113[46], net1113[47]}),
     .sp4_r_v_b_08({net1114[0], net1114[1], net1114[2], net1114[3],
     net1114[4], net1114[5], net1114[6], net1114[7], net1114[8],
     net1114[9], net1114[10], net1114[11], net1114[12], net1114[13],
     net1114[14], net1114[15], net1114[16], net1114[17], net1114[18],
     net1114[19], net1114[20], net1114[21], net1114[22], net1114[23],
     net1114[24], net1114[25], net1114[26], net1114[27], net1114[28],
     net1114[29], net1114[30], net1114[31], net1114[32], net1114[33],
     net1114[34], net1114[35], net1114[36], net1114[37], net1114[38],
     net1114[39], net1114[40], net1114[41], net1114[42], net1114[43],
     net1114[44], net1114[45], net1114[46], net1114[47]}),
     .sp4_v_b_08({net1400[0], net1400[1], net1400[2], net1400[3],
     net1400[4], net1400[5], net1400[6], net1400[7], net1400[8],
     net1400[9], net1400[10], net1400[11], net1400[12], net1400[13],
     net1400[14], net1400[15], net1400[16], net1400[17], net1400[18],
     net1400[19], net1400[20], net1400[21], net1400[22], net1400[23],
     net1400[24], net1400[25], net1400[26], net1400[27], net1400[28],
     net1400[29], net1400[30], net1400[31], net1400[32], net1400[33],
     net1400[34], net1400[35], net1400[36], net1400[37], net1400[38],
     net1400[39], net1400[40], net1400[41], net1400[42], net1400[43],
     net1400[44], net1400[45], net1400[46], net1400[47]}),
     .sp4_v_b_07({net1401[0], net1401[1], net1401[2], net1401[3],
     net1401[4], net1401[5], net1401[6], net1401[7], net1401[8],
     net1401[9], net1401[10], net1401[11], net1401[12], net1401[13],
     net1401[14], net1401[15], net1401[16], net1401[17], net1401[18],
     net1401[19], net1401[20], net1401[21], net1401[22], net1401[23],
     net1401[24], net1401[25], net1401[26], net1401[27], net1401[28],
     net1401[29], net1401[30], net1401[31], net1401[32], net1401[33],
     net1401[34], net1401[35], net1401[36], net1401[37], net1401[38],
     net1401[39], net1401[40], net1401[41], net1401[42], net1401[43],
     net1401[44], net1401[45], net1401[46], net1401[47]}),
     .sp4_v_b_06({net1402[0], net1402[1], net1402[2], net1402[3],
     net1402[4], net1402[5], net1402[6], net1402[7], net1402[8],
     net1402[9], net1402[10], net1402[11], net1402[12], net1402[13],
     net1402[14], net1402[15], net1402[16], net1402[17], net1402[18],
     net1402[19], net1402[20], net1402[21], net1402[22], net1402[23],
     net1402[24], net1402[25], net1402[26], net1402[27], net1402[28],
     net1402[29], net1402[30], net1402[31], net1402[32], net1402[33],
     net1402[34], net1402[35], net1402[36], net1402[37], net1402[38],
     net1402[39], net1402[40], net1402[41], net1402[42], net1402[43],
     net1402[44], net1402[45], net1402[46], net1402[47]}),
     .sp4_v_b_05({net1369[0], net1369[1], net1369[2], net1369[3],
     net1369[4], net1369[5], net1369[6], net1369[7], net1369[8],
     net1369[9], net1369[10], net1369[11], net1369[12], net1369[13],
     net1369[14], net1369[15], net1369[16], net1369[17], net1369[18],
     net1369[19], net1369[20], net1369[21], net1369[22], net1369[23],
     net1369[24], net1369[25], net1369[26], net1369[27], net1369[28],
     net1369[29], net1369[30], net1369[31], net1369[32], net1369[33],
     net1369[34], net1369[35], net1369[36], net1369[37], net1369[38],
     net1369[39], net1369[40], net1369[41], net1369[42], net1369[43],
     net1369[44], net1369[45], net1369[46], net1369[47]}),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .wl(wl_r[127:0]), .sp12_v_t_08({net1122[0], net1122[1],
     net1122[2], net1122[3], net1122[4], net1122[5], net1122[6],
     net1122[7], net1122[8], net1122[9], net1122[10], net1122[11],
     net1122[12], net1122[13], net1122[14], net1122[15], net1122[16],
     net1122[17], net1122[18], net1122[19], net1122[20], net1122[21],
     net1122[22], net1122[23]}), .tnr_op_08({slf_op_12_17[3],
     slf_op_12_17[2], slf_op_12_17[1], slf_op_12_17[0],
     slf_op_12_17[3], slf_op_12_17[2], slf_op_12_17[1],
     slf_op_12_17[0]}), .top_op_08({slf_op_11_17[3], slf_op_11_17[2],
     slf_op_11_17[1], slf_op_11_17[0], slf_op_11_17[3],
     slf_op_11_17[2], slf_op_11_17[1], slf_op_11_17[0]}),
     .tnl_op_08({slf_op_10_17[3], slf_op_10_17[2], slf_op_10_17[1],
     slf_op_10_17[0], slf_op_10_17[3], slf_op_10_17[2],
     slf_op_10_17[1], slf_op_10_17[0]}), .sp4_v_t_08({net1126[0],
     net1126[1], net1126[2], net1126[3], net1126[4], net1126[5],
     net1126[6], net1126[7], net1126[8], net1126[9], net1126[10],
     net1126[11], net1126[12], net1126[13], net1126[14], net1126[15],
     net1126[16], net1126[17], net1126[18], net1126[19], net1126[20],
     net1126[21], net1126[22], net1126[23], net1126[24], net1126[25],
     net1126[26], net1126[27], net1126[28], net1126[29], net1126[30],
     net1126[31], net1126[32], net1126[33], net1126[34], net1126[35],
     net1126[36], net1126[37], net1126[38], net1126[39], net1126[40],
     net1126[41], net1126[42], net1126[43], net1126[44], net1126[45],
     net1126[46], net1126[47]}), .lc_bot(lc_bot_11_09),
     .op_vic(net1128), .sp12_v_b_01(sp12_v_b_11_09[23:0]),
     .glb_netwk_t({net1130[0], net1130[1], net1130[2], net1130[3],
     net1130[4], net1130[5], net1130[6], net1130[7]}));
lt_1x8_top_ice1f I_lt_col_t08 ( .glb_netwk_b({net01133[0], net01133[1],
     net01133[2], net01133[3], net01133[4], net01133[5], net01133[6],
     net01133[7]}), .rgt_op_03({net1131[0], net1131[1], net1131[2],
     net1131[3], net1131[4], net1131[5], net1131[6], net1131[7]}),
     .slf_op_02({net1227[0], net1227[1], net1227[2], net1227[3],
     net1227[4], net1227[5], net1227[6], net1227[7]}),
     .rgt_op_02({net1133[0], net1133[1], net1133[2], net1133[3],
     net1133[4], net1133[5], net1133[6], net1133[7]}),
     .rgt_op_01(slf_op_09_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(slf_op_07_12[7:0]), .lft_op_03(slf_op_07_11[7:0]),
     .lft_op_02(slf_op_07_10[7:0]), .lft_op_01(slf_op_07_09[7:0]),
     .rgt_op_04({net1141[0], net1141[1], net1141[2], net1141[3],
     net1141[4], net1141[5], net1141[6], net1141[7]}),
     .carry_in(carry_in_08_09), .bnl_op_01(bnl_op_08_09[7:0]),
     .slf_op_04({net1235[0], net1235[1], net1235[2], net1235[3],
     net1235[4], net1235[5], net1235[6], net1235[7]}),
     .slf_op_03({net1225[0], net1225[1], net1225[2], net1225[3],
     net1225[4], net1225[5], net1225[6], net1225[7]}),
     .slf_op_01(slf_op_08_09[7:0]), .sp4_h_l_04({net1254[0],
     net1254[1], net1254[2], net1254[3], net1254[4], net1254[5],
     net1254[6], net1254[7], net1254[8], net1254[9], net1254[10],
     net1254[11], net1254[12], net1254[13], net1254[14], net1254[15],
     net1254[16], net1254[17], net1254[18], net1254[19], net1254[20],
     net1254[21], net1254[22], net1254[23], net1254[24], net1254[25],
     net1254[26], net1254[27], net1254[28], net1254[29], net1254[30],
     net1254[31], net1254[32], net1254[33], net1254[34], net1254[35],
     net1254[36], net1254[37], net1254[38], net1254[39], net1254[40],
     net1254[41], net1254[42], net1254[43], net1254[44], net1254[45],
     net1254[46], net1254[47]}), .carry_out(net1148),
     .vdd_cntl(vdd_cntl_r[127:0]), .sp12_h_r_04({net1150[0],
     net1150[1], net1150[2], net1150[3], net1150[4], net1150[5],
     net1150[6], net1150[7], net1150[8], net1150[9], net1150[10],
     net1150[11], net1150[12], net1150[13], net1150[14], net1150[15],
     net1150[16], net1150[17], net1150[18], net1150[19], net1150[20],
     net1150[21], net1150[22], net1150[23]}), .sp12_h_r_03({net1151[0],
     net1151[1], net1151[2], net1151[3], net1151[4], net1151[5],
     net1151[6], net1151[7], net1151[8], net1151[9], net1151[10],
     net1151[11], net1151[12], net1151[13], net1151[14], net1151[15],
     net1151[16], net1151[17], net1151[18], net1151[19], net1151[20],
     net1151[21], net1151[22], net1151[23]}), .sp12_h_r_02({net1152[0],
     net1152[1], net1152[2], net1152[3], net1152[4], net1152[5],
     net1152[6], net1152[7], net1152[8], net1152[9], net1152[10],
     net1152[11], net1152[12], net1152[13], net1152[14], net1152[15],
     net1152[16], net1152[17], net1152[18], net1152[19], net1152[20],
     net1152[21], net1152[22], net1152[23]}), .sp12_h_r_01({net1153[0],
     net1153[1], net1153[2], net1153[3], net1153[4], net1153[5],
     net1153[6], net1153[7], net1153[8], net1153[9], net1153[10],
     net1153[11], net1153[12], net1153[13], net1153[14], net1153[15],
     net1153[16], net1153[17], net1153[18], net1153[19], net1153[20],
     net1153[21], net1153[22], net1153[23]}),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_08_09[47:0]), .sp4_r_v_b_04({net1156[0],
     net1156[1], net1156[2], net1156[3], net1156[4], net1156[5],
     net1156[6], net1156[7], net1156[8], net1156[9], net1156[10],
     net1156[11], net1156[12], net1156[13], net1156[14], net1156[15],
     net1156[16], net1156[17], net1156[18], net1156[19], net1156[20],
     net1156[21], net1156[22], net1156[23], net1156[24], net1156[25],
     net1156[26], net1156[27], net1156[28], net1156[29], net1156[30],
     net1156[31], net1156[32], net1156[33], net1156[34], net1156[35],
     net1156[36], net1156[37], net1156[38], net1156[39], net1156[40],
     net1156[41], net1156[42], net1156[43], net1156[44], net1156[45],
     net1156[46], net1156[47]}), .sp4_r_v_b_03({net1157[0], net1157[1],
     net1157[2], net1157[3], net1157[4], net1157[5], net1157[6],
     net1157[7], net1157[8], net1157[9], net1157[10], net1157[11],
     net1157[12], net1157[13], net1157[14], net1157[15], net1157[16],
     net1157[17], net1157[18], net1157[19], net1157[20], net1157[21],
     net1157[22], net1157[23], net1157[24], net1157[25], net1157[26],
     net1157[27], net1157[28], net1157[29], net1157[30], net1157[31],
     net1157[32], net1157[33], net1157[34], net1157[35], net1157[36],
     net1157[37], net1157[38], net1157[39], net1157[40], net1157[41],
     net1157[42], net1157[43], net1157[44], net1157[45], net1157[46],
     net1157[47]}), .sp4_r_v_b_02({net1158[0], net1158[1], net1158[2],
     net1158[3], net1158[4], net1158[5], net1158[6], net1158[7],
     net1158[8], net1158[9], net1158[10], net1158[11], net1158[12],
     net1158[13], net1158[14], net1158[15], net1158[16], net1158[17],
     net1158[18], net1158[19], net1158[20], net1158[21], net1158[22],
     net1158[23], net1158[24], net1158[25], net1158[26], net1158[27],
     net1158[28], net1158[29], net1158[30], net1158[31], net1158[32],
     net1158[33], net1158[34], net1158[35], net1158[36], net1158[37],
     net1158[38], net1158[39], net1158[40], net1158[41], net1158[42],
     net1158[43], net1158[44], net1158[45], net1158[46], net1158[47]}),
     .sp4_r_v_b_01(sp4_v_b_09_09[47:0]), .sp4_h_r_04({net1160[0],
     net1160[1], net1160[2], net1160[3], net1160[4], net1160[5],
     net1160[6], net1160[7], net1160[8], net1160[9], net1160[10],
     net1160[11], net1160[12], net1160[13], net1160[14], net1160[15],
     net1160[16], net1160[17], net1160[18], net1160[19], net1160[20],
     net1160[21], net1160[22], net1160[23], net1160[24], net1160[25],
     net1160[26], net1160[27], net1160[28], net1160[29], net1160[30],
     net1160[31], net1160[32], net1160[33], net1160[34], net1160[35],
     net1160[36], net1160[37], net1160[38], net1160[39], net1160[40],
     net1160[41], net1160[42], net1160[43], net1160[44], net1160[45],
     net1160[46], net1160[47]}), .sp4_h_r_03({net1161[0], net1161[1],
     net1161[2], net1161[3], net1161[4], net1161[5], net1161[6],
     net1161[7], net1161[8], net1161[9], net1161[10], net1161[11],
     net1161[12], net1161[13], net1161[14], net1161[15], net1161[16],
     net1161[17], net1161[18], net1161[19], net1161[20], net1161[21],
     net1161[22], net1161[23], net1161[24], net1161[25], net1161[26],
     net1161[27], net1161[28], net1161[29], net1161[30], net1161[31],
     net1161[32], net1161[33], net1161[34], net1161[35], net1161[36],
     net1161[37], net1161[38], net1161[39], net1161[40], net1161[41],
     net1161[42], net1161[43], net1161[44], net1161[45], net1161[46],
     net1161[47]}), .sp4_h_r_02({net1162[0], net1162[1], net1162[2],
     net1162[3], net1162[4], net1162[5], net1162[6], net1162[7],
     net1162[8], net1162[9], net1162[10], net1162[11], net1162[12],
     net1162[13], net1162[14], net1162[15], net1162[16], net1162[17],
     net1162[18], net1162[19], net1162[20], net1162[21], net1162[22],
     net1162[23], net1162[24], net1162[25], net1162[26], net1162[27],
     net1162[28], net1162[29], net1162[30], net1162[31], net1162[32],
     net1162[33], net1162[34], net1162[35], net1162[36], net1162[37],
     net1162[38], net1162[39], net1162[40], net1162[41], net1162[42],
     net1162[43], net1162[44], net1162[45], net1162[46], net1162[47]}),
     .sp4_h_r_01({net1163[0], net1163[1], net1163[2], net1163[3],
     net1163[4], net1163[5], net1163[6], net1163[7], net1163[8],
     net1163[9], net1163[10], net1163[11], net1163[12], net1163[13],
     net1163[14], net1163[15], net1163[16], net1163[17], net1163[18],
     net1163[19], net1163[20], net1163[21], net1163[22], net1163[23],
     net1163[24], net1163[25], net1163[26], net1163[27], net1163[28],
     net1163[29], net1163[30], net1163[31], net1163[32], net1163[33],
     net1163[34], net1163[35], net1163[36], net1163[37], net1163[38],
     net1163[39], net1163[40], net1163[41], net1163[42], net1163[43],
     net1163[44], net1163[45], net1163[46], net1163[47]}),
     .sp4_h_l_03({net1255[0], net1255[1], net1255[2], net1255[3],
     net1255[4], net1255[5], net1255[6], net1255[7], net1255[8],
     net1255[9], net1255[10], net1255[11], net1255[12], net1255[13],
     net1255[14], net1255[15], net1255[16], net1255[17], net1255[18],
     net1255[19], net1255[20], net1255[21], net1255[22], net1255[23],
     net1255[24], net1255[25], net1255[26], net1255[27], net1255[28],
     net1255[29], net1255[30], net1255[31], net1255[32], net1255[33],
     net1255[34], net1255[35], net1255[36], net1255[37], net1255[38],
     net1255[39], net1255[40], net1255[41], net1255[42], net1255[43],
     net1255[44], net1255[45], net1255[46], net1255[47]}),
     .sp4_h_l_02({net1256[0], net1256[1], net1256[2], net1256[3],
     net1256[4], net1256[5], net1256[6], net1256[7], net1256[8],
     net1256[9], net1256[10], net1256[11], net1256[12], net1256[13],
     net1256[14], net1256[15], net1256[16], net1256[17], net1256[18],
     net1256[19], net1256[20], net1256[21], net1256[22], net1256[23],
     net1256[24], net1256[25], net1256[26], net1256[27], net1256[28],
     net1256[29], net1256[30], net1256[31], net1256[32], net1256[33],
     net1256[34], net1256[35], net1256[36], net1256[37], net1256[38],
     net1256[39], net1256[40], net1256[41], net1256[42], net1256[43],
     net1256[44], net1256[45], net1256[46], net1256[47]}),
     .sp4_h_l_01({net1257[0], net1257[1], net1257[2], net1257[3],
     net1257[4], net1257[5], net1257[6], net1257[7], net1257[8],
     net1257[9], net1257[10], net1257[11], net1257[12], net1257[13],
     net1257[14], net1257[15], net1257[16], net1257[17], net1257[18],
     net1257[19], net1257[20], net1257[21], net1257[22], net1257[23],
     net1257[24], net1257[25], net1257[26], net1257[27], net1257[28],
     net1257[29], net1257[30], net1257[31], net1257[32], net1257[33],
     net1257[34], net1257[35], net1257[36], net1257[37], net1257[38],
     net1257[39], net1257[40], net1257[41], net1257[42], net1257[43],
     net1257[44], net1257[45], net1257[46], net1257[47]}),
     .bl(bl[107:54]), .bot_op_01(bot_op_08_09[7:0]),
     .sp12_h_l_01({net1247[0], net1247[1], net1247[2], net1247[3],
     net1247[4], net1247[5], net1247[6], net1247[7], net1247[8],
     net1247[9], net1247[10], net1247[11], net1247[12], net1247[13],
     net1247[14], net1247[15], net1247[16], net1247[17], net1247[18],
     net1247[19], net1247[20], net1247[21], net1247[22], net1247[23]}),
     .sp12_h_l_02({net1246[0], net1246[1], net1246[2], net1246[3],
     net1246[4], net1246[5], net1246[6], net1246[7], net1246[8],
     net1246[9], net1246[10], net1246[11], net1246[12], net1246[13],
     net1246[14], net1246[15], net1246[16], net1246[17], net1246[18],
     net1246[19], net1246[20], net1246[21], net1246[22], net1246[23]}),
     .sp12_h_l_03({net1245[0], net1245[1], net1245[2], net1245[3],
     net1245[4], net1245[5], net1245[6], net1245[7], net1245[8],
     net1245[9], net1245[10], net1245[11], net1245[12], net1245[13],
     net1245[14], net1245[15], net1245[16], net1245[17], net1245[18],
     net1245[19], net1245[20], net1245[21], net1245[22], net1245[23]}),
     .sp12_h_l_04({net1244[0], net1244[1], net1244[2], net1244[3],
     net1244[4], net1244[5], net1244[6], net1244[7], net1244[8],
     net1244[9], net1244[10], net1244[11], net1244[12], net1244[13],
     net1244[14], net1244[15], net1244[16], net1244[17], net1244[18],
     net1244[19], net1244[20], net1244[21], net1244[22], net1244[23]}),
     .sp4_v_b_04({net1250[0], net1250[1], net1250[2], net1250[3],
     net1250[4], net1250[5], net1250[6], net1250[7], net1250[8],
     net1250[9], net1250[10], net1250[11], net1250[12], net1250[13],
     net1250[14], net1250[15], net1250[16], net1250[17], net1250[18],
     net1250[19], net1250[20], net1250[21], net1250[22], net1250[23],
     net1250[24], net1250[25], net1250[26], net1250[27], net1250[28],
     net1250[29], net1250[30], net1250[31], net1250[32], net1250[33],
     net1250[34], net1250[35], net1250[36], net1250[37], net1250[38],
     net1250[39], net1250[40], net1250[41], net1250[42], net1250[43],
     net1250[44], net1250[45], net1250[46], net1250[47]}),
     .sp4_v_b_03({net1251[0], net1251[1], net1251[2], net1251[3],
     net1251[4], net1251[5], net1251[6], net1251[7], net1251[8],
     net1251[9], net1251[10], net1251[11], net1251[12], net1251[13],
     net1251[14], net1251[15], net1251[16], net1251[17], net1251[18],
     net1251[19], net1251[20], net1251[21], net1251[22], net1251[23],
     net1251[24], net1251[25], net1251[26], net1251[27], net1251[28],
     net1251[29], net1251[30], net1251[31], net1251[32], net1251[33],
     net1251[34], net1251[35], net1251[36], net1251[37], net1251[38],
     net1251[39], net1251[40], net1251[41], net1251[42], net1251[43],
     net1251[44], net1251[45], net1251[46], net1251[47]}),
     .sp4_v_b_02({net1252[0], net1252[1], net1252[2], net1252[3],
     net1252[4], net1252[5], net1252[6], net1252[7], net1252[8],
     net1252[9], net1252[10], net1252[11], net1252[12], net1252[13],
     net1252[14], net1252[15], net1252[16], net1252[17], net1252[18],
     net1252[19], net1252[20], net1252[21], net1252[22], net1252[23],
     net1252[24], net1252[25], net1252[26], net1252[27], net1252[28],
     net1252[29], net1252[30], net1252[31], net1252[32], net1252[33],
     net1252[34], net1252[35], net1252[36], net1252[37], net1252[38],
     net1252[39], net1252[40], net1252[41], net1252[42], net1252[43],
     net1252[44], net1252[45], net1252[46], net1252[47]}),
     .bnr_op_01(bnr_op_08_09[7:0]), .sp4_h_l_05({net1278[0],
     net1278[1], net1278[2], net1278[3], net1278[4], net1278[5],
     net1278[6], net1278[7], net1278[8], net1278[9], net1278[10],
     net1278[11], net1278[12], net1278[13], net1278[14], net1278[15],
     net1278[16], net1278[17], net1278[18], net1278[19], net1278[20],
     net1278[21], net1278[22], net1278[23], net1278[24], net1278[25],
     net1278[26], net1278[27], net1278[28], net1278[29], net1278[30],
     net1278[31], net1278[32], net1278[33], net1278[34], net1278[35],
     net1278[36], net1278[37], net1278[38], net1278[39], net1278[40],
     net1278[41], net1278[42], net1278[43], net1278[44], net1278[45],
     net1278[46], net1278[47]}), .sp4_h_l_06({net1277[0], net1277[1],
     net1277[2], net1277[3], net1277[4], net1277[5], net1277[6],
     net1277[7], net1277[8], net1277[9], net1277[10], net1277[11],
     net1277[12], net1277[13], net1277[14], net1277[15], net1277[16],
     net1277[17], net1277[18], net1277[19], net1277[20], net1277[21],
     net1277[22], net1277[23], net1277[24], net1277[25], net1277[26],
     net1277[27], net1277[28], net1277[29], net1277[30], net1277[31],
     net1277[32], net1277[33], net1277[34], net1277[35], net1277[36],
     net1277[37], net1277[38], net1277[39], net1277[40], net1277[41],
     net1277[42], net1277[43], net1277[44], net1277[45], net1277[46],
     net1277[47]}), .sp4_h_l_07({net1276[0], net1276[1], net1276[2],
     net1276[3], net1276[4], net1276[5], net1276[6], net1276[7],
     net1276[8], net1276[9], net1276[10], net1276[11], net1276[12],
     net1276[13], net1276[14], net1276[15], net1276[16], net1276[17],
     net1276[18], net1276[19], net1276[20], net1276[21], net1276[22],
     net1276[23], net1276[24], net1276[25], net1276[26], net1276[27],
     net1276[28], net1276[29], net1276[30], net1276[31], net1276[32],
     net1276[33], net1276[34], net1276[35], net1276[36], net1276[37],
     net1276[38], net1276[39], net1276[40], net1276[41], net1276[42],
     net1276[43], net1276[44], net1276[45], net1276[46], net1276[47]}),
     .sp4_h_l_08({net1275[0], net1275[1], net1275[2], net1275[3],
     net1275[4], net1275[5], net1275[6], net1275[7], net1275[8],
     net1275[9], net1275[10], net1275[11], net1275[12], net1275[13],
     net1275[14], net1275[15], net1275[16], net1275[17], net1275[18],
     net1275[19], net1275[20], net1275[21], net1275[22], net1275[23],
     net1275[24], net1275[25], net1275[26], net1275[27], net1275[28],
     net1275[29], net1275[30], net1275[31], net1275[32], net1275[33],
     net1275[34], net1275[35], net1275[36], net1275[37], net1275[38],
     net1275[39], net1275[40], net1275[41], net1275[42], net1275[43],
     net1275[44], net1275[45], net1275[46], net1275[47]}),
     .sp4_h_r_08({net1181[0], net1181[1], net1181[2], net1181[3],
     net1181[4], net1181[5], net1181[6], net1181[7], net1181[8],
     net1181[9], net1181[10], net1181[11], net1181[12], net1181[13],
     net1181[14], net1181[15], net1181[16], net1181[17], net1181[18],
     net1181[19], net1181[20], net1181[21], net1181[22], net1181[23],
     net1181[24], net1181[25], net1181[26], net1181[27], net1181[28],
     net1181[29], net1181[30], net1181[31], net1181[32], net1181[33],
     net1181[34], net1181[35], net1181[36], net1181[37], net1181[38],
     net1181[39], net1181[40], net1181[41], net1181[42], net1181[43],
     net1181[44], net1181[45], net1181[46], net1181[47]}),
     .sp4_h_r_07({net1182[0], net1182[1], net1182[2], net1182[3],
     net1182[4], net1182[5], net1182[6], net1182[7], net1182[8],
     net1182[9], net1182[10], net1182[11], net1182[12], net1182[13],
     net1182[14], net1182[15], net1182[16], net1182[17], net1182[18],
     net1182[19], net1182[20], net1182[21], net1182[22], net1182[23],
     net1182[24], net1182[25], net1182[26], net1182[27], net1182[28],
     net1182[29], net1182[30], net1182[31], net1182[32], net1182[33],
     net1182[34], net1182[35], net1182[36], net1182[37], net1182[38],
     net1182[39], net1182[40], net1182[41], net1182[42], net1182[43],
     net1182[44], net1182[45], net1182[46], net1182[47]}),
     .sp4_h_r_06({net1183[0], net1183[1], net1183[2], net1183[3],
     net1183[4], net1183[5], net1183[6], net1183[7], net1183[8],
     net1183[9], net1183[10], net1183[11], net1183[12], net1183[13],
     net1183[14], net1183[15], net1183[16], net1183[17], net1183[18],
     net1183[19], net1183[20], net1183[21], net1183[22], net1183[23],
     net1183[24], net1183[25], net1183[26], net1183[27], net1183[28],
     net1183[29], net1183[30], net1183[31], net1183[32], net1183[33],
     net1183[34], net1183[35], net1183[36], net1183[37], net1183[38],
     net1183[39], net1183[40], net1183[41], net1183[42], net1183[43],
     net1183[44], net1183[45], net1183[46], net1183[47]}),
     .sp4_h_r_05({net1184[0], net1184[1], net1184[2], net1184[3],
     net1184[4], net1184[5], net1184[6], net1184[7], net1184[8],
     net1184[9], net1184[10], net1184[11], net1184[12], net1184[13],
     net1184[14], net1184[15], net1184[16], net1184[17], net1184[18],
     net1184[19], net1184[20], net1184[21], net1184[22], net1184[23],
     net1184[24], net1184[25], net1184[26], net1184[27], net1184[28],
     net1184[29], net1184[30], net1184[31], net1184[32], net1184[33],
     net1184[34], net1184[35], net1184[36], net1184[37], net1184[38],
     net1184[39], net1184[40], net1184[41], net1184[42], net1184[43],
     net1184[44], net1184[45], net1184[46], net1184[47]}),
     .slf_op_05({net1286[0], net1286[1], net1286[2], net1286[3],
     net1286[4], net1286[5], net1286[6], net1286[7]}),
     .slf_op_06({net1285[0], net1285[1], net1285[2], net1285[3],
     net1285[4], net1285[5], net1285[6], net1285[7]}),
     .slf_op_07({net1284[0], net1284[1], net1284[2], net1284[3],
     net1284[4], net1284[5], net1284[6], net1284[7]}),
     .slf_op_08({net1283[0], net1283[1], net1283[2], net1283[3],
     net1283[4], net1283[5], net1283[6], net1283[7]}),
     .rgt_op_08({net1189[0], net1189[1], net1189[2], net1189[3],
     net1189[4], net1189[5], net1189[6], net1189[7]}),
     .rgt_op_07({net1190[0], net1190[1], net1190[2], net1190[3],
     net1190[4], net1190[5], net1190[6], net1190[7]}),
     .rgt_op_06({net1191[0], net1191[1], net1191[2], net1191[3],
     net1191[4], net1191[5], net1191[6], net1191[7]}),
     .rgt_op_05({net1192[0], net1192[1], net1192[2], net1192[3],
     net1192[4], net1192[5], net1192[6], net1192[7]}),
     .lft_op_08(slf_op_07_16[7:0]), .lft_op_07(slf_op_07_15[7:0]),
     .lft_op_06(slf_op_07_14[7:0]), .lft_op_05(slf_op_07_13[7:0]),
     .sp12_h_l_08({net1297[0], net1297[1], net1297[2], net1297[3],
     net1297[4], net1297[5], net1297[6], net1297[7], net1297[8],
     net1297[9], net1297[10], net1297[11], net1297[12], net1297[13],
     net1297[14], net1297[15], net1297[16], net1297[17], net1297[18],
     net1297[19], net1297[20], net1297[21], net1297[22], net1297[23]}),
     .sp12_h_l_07({net1296[0], net1296[1], net1296[2], net1296[3],
     net1296[4], net1296[5], net1296[6], net1296[7], net1296[8],
     net1296[9], net1296[10], net1296[11], net1296[12], net1296[13],
     net1296[14], net1296[15], net1296[16], net1296[17], net1296[18],
     net1296[19], net1296[20], net1296[21], net1296[22], net1296[23]}),
     .sp12_h_l_06({net1295[0], net1295[1], net1295[2], net1295[3],
     net1295[4], net1295[5], net1295[6], net1295[7], net1295[8],
     net1295[9], net1295[10], net1295[11], net1295[12], net1295[13],
     net1295[14], net1295[15], net1295[16], net1295[17], net1295[18],
     net1295[19], net1295[20], net1295[21], net1295[22], net1295[23]}),
     .sp12_h_r_05({net1200[0], net1200[1], net1200[2], net1200[3],
     net1200[4], net1200[5], net1200[6], net1200[7], net1200[8],
     net1200[9], net1200[10], net1200[11], net1200[12], net1200[13],
     net1200[14], net1200[15], net1200[16], net1200[17], net1200[18],
     net1200[19], net1200[20], net1200[21], net1200[22], net1200[23]}),
     .sp12_h_r_06({net1201[0], net1201[1], net1201[2], net1201[3],
     net1201[4], net1201[5], net1201[6], net1201[7], net1201[8],
     net1201[9], net1201[10], net1201[11], net1201[12], net1201[13],
     net1201[14], net1201[15], net1201[16], net1201[17], net1201[18],
     net1201[19], net1201[20], net1201[21], net1201[22], net1201[23]}),
     .sp12_h_r_07({net1202[0], net1202[1], net1202[2], net1202[3],
     net1202[4], net1202[5], net1202[6], net1202[7], net1202[8],
     net1202[9], net1202[10], net1202[11], net1202[12], net1202[13],
     net1202[14], net1202[15], net1202[16], net1202[17], net1202[18],
     net1202[19], net1202[20], net1202[21], net1202[22], net1202[23]}),
     .sp12_h_r_08({net1203[0], net1203[1], net1203[2], net1203[3],
     net1203[4], net1203[5], net1203[6], net1203[7], net1203[8],
     net1203[9], net1203[10], net1203[11], net1203[12], net1203[13],
     net1203[14], net1203[15], net1203[16], net1203[17], net1203[18],
     net1203[19], net1203[20], net1203[21], net1203[22], net1203[23]}),
     .sp12_h_l_05({net1294[0], net1294[1], net1294[2], net1294[3],
     net1294[4], net1294[5], net1294[6], net1294[7], net1294[8],
     net1294[9], net1294[10], net1294[11], net1294[12], net1294[13],
     net1294[14], net1294[15], net1294[16], net1294[17], net1294[18],
     net1294[19], net1294[20], net1294[21], net1294[22], net1294[23]}),
     .sp4_r_v_b_05({net1205[0], net1205[1], net1205[2], net1205[3],
     net1205[4], net1205[5], net1205[6], net1205[7], net1205[8],
     net1205[9], net1205[10], net1205[11], net1205[12], net1205[13],
     net1205[14], net1205[15], net1205[16], net1205[17], net1205[18],
     net1205[19], net1205[20], net1205[21], net1205[22], net1205[23],
     net1205[24], net1205[25], net1205[26], net1205[27], net1205[28],
     net1205[29], net1205[30], net1205[31], net1205[32], net1205[33],
     net1205[34], net1205[35], net1205[36], net1205[37], net1205[38],
     net1205[39], net1205[40], net1205[41], net1205[42], net1205[43],
     net1205[44], net1205[45], net1205[46], net1205[47]}),
     .sp4_r_v_b_06({net1206[0], net1206[1], net1206[2], net1206[3],
     net1206[4], net1206[5], net1206[6], net1206[7], net1206[8],
     net1206[9], net1206[10], net1206[11], net1206[12], net1206[13],
     net1206[14], net1206[15], net1206[16], net1206[17], net1206[18],
     net1206[19], net1206[20], net1206[21], net1206[22], net1206[23],
     net1206[24], net1206[25], net1206[26], net1206[27], net1206[28],
     net1206[29], net1206[30], net1206[31], net1206[32], net1206[33],
     net1206[34], net1206[35], net1206[36], net1206[37], net1206[38],
     net1206[39], net1206[40], net1206[41], net1206[42], net1206[43],
     net1206[44], net1206[45], net1206[46], net1206[47]}),
     .sp4_r_v_b_07({net1207[0], net1207[1], net1207[2], net1207[3],
     net1207[4], net1207[5], net1207[6], net1207[7], net1207[8],
     net1207[9], net1207[10], net1207[11], net1207[12], net1207[13],
     net1207[14], net1207[15], net1207[16], net1207[17], net1207[18],
     net1207[19], net1207[20], net1207[21], net1207[22], net1207[23],
     net1207[24], net1207[25], net1207[26], net1207[27], net1207[28],
     net1207[29], net1207[30], net1207[31], net1207[32], net1207[33],
     net1207[34], net1207[35], net1207[36], net1207[37], net1207[38],
     net1207[39], net1207[40], net1207[41], net1207[42], net1207[43],
     net1207[44], net1207[45], net1207[46], net1207[47]}),
     .sp4_r_v_b_08({net1208[0], net1208[1], net1208[2], net1208[3],
     net1208[4], net1208[5], net1208[6], net1208[7], net1208[8],
     net1208[9], net1208[10], net1208[11], net1208[12], net1208[13],
     net1208[14], net1208[15], net1208[16], net1208[17], net1208[18],
     net1208[19], net1208[20], net1208[21], net1208[22], net1208[23],
     net1208[24], net1208[25], net1208[26], net1208[27], net1208[28],
     net1208[29], net1208[30], net1208[31], net1208[32], net1208[33],
     net1208[34], net1208[35], net1208[36], net1208[37], net1208[38],
     net1208[39], net1208[40], net1208[41], net1208[42], net1208[43],
     net1208[44], net1208[45], net1208[46], net1208[47]}),
     .sp4_v_b_08({net1302[0], net1302[1], net1302[2], net1302[3],
     net1302[4], net1302[5], net1302[6], net1302[7], net1302[8],
     net1302[9], net1302[10], net1302[11], net1302[12], net1302[13],
     net1302[14], net1302[15], net1302[16], net1302[17], net1302[18],
     net1302[19], net1302[20], net1302[21], net1302[22], net1302[23],
     net1302[24], net1302[25], net1302[26], net1302[27], net1302[28],
     net1302[29], net1302[30], net1302[31], net1302[32], net1302[33],
     net1302[34], net1302[35], net1302[36], net1302[37], net1302[38],
     net1302[39], net1302[40], net1302[41], net1302[42], net1302[43],
     net1302[44], net1302[45], net1302[46], net1302[47]}),
     .sp4_v_b_07({net1301[0], net1301[1], net1301[2], net1301[3],
     net1301[4], net1301[5], net1301[6], net1301[7], net1301[8],
     net1301[9], net1301[10], net1301[11], net1301[12], net1301[13],
     net1301[14], net1301[15], net1301[16], net1301[17], net1301[18],
     net1301[19], net1301[20], net1301[21], net1301[22], net1301[23],
     net1301[24], net1301[25], net1301[26], net1301[27], net1301[28],
     net1301[29], net1301[30], net1301[31], net1301[32], net1301[33],
     net1301[34], net1301[35], net1301[36], net1301[37], net1301[38],
     net1301[39], net1301[40], net1301[41], net1301[42], net1301[43],
     net1301[44], net1301[45], net1301[46], net1301[47]}),
     .sp4_v_b_06({net1300[0], net1300[1], net1300[2], net1300[3],
     net1300[4], net1300[5], net1300[6], net1300[7], net1300[8],
     net1300[9], net1300[10], net1300[11], net1300[12], net1300[13],
     net1300[14], net1300[15], net1300[16], net1300[17], net1300[18],
     net1300[19], net1300[20], net1300[21], net1300[22], net1300[23],
     net1300[24], net1300[25], net1300[26], net1300[27], net1300[28],
     net1300[29], net1300[30], net1300[31], net1300[32], net1300[33],
     net1300[34], net1300[35], net1300[36], net1300[37], net1300[38],
     net1300[39], net1300[40], net1300[41], net1300[42], net1300[43],
     net1300[44], net1300[45], net1300[46], net1300[47]}),
     .sp4_v_b_05({net1299[0], net1299[1], net1299[2], net1299[3],
     net1299[4], net1299[5], net1299[6], net1299[7], net1299[8],
     net1299[9], net1299[10], net1299[11], net1299[12], net1299[13],
     net1299[14], net1299[15], net1299[16], net1299[17], net1299[18],
     net1299[19], net1299[20], net1299[21], net1299[22], net1299[23],
     net1299[24], net1299[25], net1299[26], net1299[27], net1299[28],
     net1299[29], net1299[30], net1299[31], net1299[32], net1299[33],
     net1299[34], net1299[35], net1299[36], net1299[37], net1299[38],
     net1299[39], net1299[40], net1299[41], net1299[42], net1299[43],
     net1299[44], net1299[45], net1299[46], net1299[47]}),
     .pgate(pgate_r[127:0]), .reset_b(reset_b_r[127:0]),
     .wl(wl_r[127:0]), .sp12_v_t_08({net1216[0], net1216[1],
     net1216[2], net1216[3], net1216[4], net1216[5], net1216[6],
     net1216[7], net1216[8], net1216[9], net1216[10], net1216[11],
     net1216[12], net1216[13], net1216[14], net1216[15], net1216[16],
     net1216[17], net1216[18], net1216[19], net1216[20], net1216[21],
     net1216[22], net1216[23]}), .tnr_op_08({slf_op_09_17[3],
     slf_op_09_17[2], slf_op_09_17[1], slf_op_09_17[0],
     slf_op_09_17[3], slf_op_09_17[2], slf_op_09_17[1],
     slf_op_09_17[0]}), .top_op_08({slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0], slf_op_08_17[3],
     slf_op_08_17[2], slf_op_08_17[1], slf_op_08_17[0]}),
     .tnl_op_08({slf_op_07_17[3], slf_op_07_17[2], slf_op_07_17[1],
     slf_op_07_17[0], slf_op_07_17[3], slf_op_07_17[2],
     slf_op_07_17[1], slf_op_07_17[0]}), .sp4_v_t_08({net1220[0],
     net1220[1], net1220[2], net1220[3], net1220[4], net1220[5],
     net1220[6], net1220[7], net1220[8], net1220[9], net1220[10],
     net1220[11], net1220[12], net1220[13], net1220[14], net1220[15],
     net1220[16], net1220[17], net1220[18], net1220[19], net1220[20],
     net1220[21], net1220[22], net1220[23], net1220[24], net1220[25],
     net1220[26], net1220[27], net1220[28], net1220[29], net1220[30],
     net1220[31], net1220[32], net1220[33], net1220[34], net1220[35],
     net1220[36], net1220[37], net1220[38], net1220[39], net1220[40],
     net1220[41], net1220[42], net1220[43], net1220[44], net1220[45],
     net1220[46], net1220[47]}), .lc_bot(lc_bot_08_09),
     .op_vic(net1222), .sp12_v_b_01(sp12_v_b_08_09[23:0]),
     .glb_netwk_t({net1224[0], net1224[1], net1224[2], net1224[3],
     net1224[4], net1224[5], net1224[6], net1224[7]}));
lt_1x8_top_ice1f I_lt_col_t07 ( .glb_netwk_b({net01228[0], net01228[1],
     net01228[2], net01228[3], net01228[4], net01228[5], net01228[6],
     net01228[7]}), .rgt_op_03({net1225[0], net1225[1], net1225[2],
     net1225[3], net1225[4], net1225[5], net1225[6], net1225[7]}),
     .slf_op_02(slf_op_07_10[7:0]), .rgt_op_02({net1227[0], net1227[1],
     net1227[2], net1227[3], net1227[4], net1227[5], net1227[6],
     net1227[7]}), .rgt_op_01(slf_op_08_09[7:0]), .purst(purst),
     .prog(prog), .lft_op_04(lft_op_07_12[7:0]),
     .lft_op_03(lft_op_07_11[7:0]), .lft_op_02(lft_op_07_10[7:0]),
     .lft_op_01(lft_op_07_09[7:0]), .rgt_op_04({net1235[0], net1235[1],
     net1235[2], net1235[3], net1235[4], net1235[5], net1235[6],
     net1235[7]}), .carry_in(carry_in_07_09),
     .bnl_op_01(bnl_op_07_09[7:0]), .slf_op_04(slf_op_07_12[7:0]),
     .slf_op_03(slf_op_07_11[7:0]), .slf_op_01(slf_op_07_09[7:0]),
     .sp4_h_l_04(sp4_h_l_07_12[47:0]), .carry_out(net1242),
     .vdd_cntl(vdd_cntl_r[127:0]), .sp12_h_r_04({net1244[0],
     net1244[1], net1244[2], net1244[3], net1244[4], net1244[5],
     net1244[6], net1244[7], net1244[8], net1244[9], net1244[10],
     net1244[11], net1244[12], net1244[13], net1244[14], net1244[15],
     net1244[16], net1244[17], net1244[18], net1244[19], net1244[20],
     net1244[21], net1244[22], net1244[23]}), .sp12_h_r_03({net1245[0],
     net1245[1], net1245[2], net1245[3], net1245[4], net1245[5],
     net1245[6], net1245[7], net1245[8], net1245[9], net1245[10],
     net1245[11], net1245[12], net1245[13], net1245[14], net1245[15],
     net1245[16], net1245[17], net1245[18], net1245[19], net1245[20],
     net1245[21], net1245[22], net1245[23]}), .sp12_h_r_02({net1246[0],
     net1246[1], net1246[2], net1246[3], net1246[4], net1246[5],
     net1246[6], net1246[7], net1246[8], net1246[9], net1246[10],
     net1246[11], net1246[12], net1246[13], net1246[14], net1246[15],
     net1246[16], net1246[17], net1246[18], net1246[19], net1246[20],
     net1246[21], net1246[22], net1246[23]}), .sp12_h_r_01({net1247[0],
     net1247[1], net1247[2], net1247[3], net1247[4], net1247[5],
     net1247[6], net1247[7], net1247[8], net1247[9], net1247[10],
     net1247[11], net1247[12], net1247[13], net1247[14], net1247[15],
     net1247[16], net1247[17], net1247[18], net1247[19], net1247[20],
     net1247[21], net1247[22], net1247[23]}),
     .glb_netwk_col(clk_tree_drv_tr[7:0]),
     .sp4_v_b_01(sp4_v_b_07_09[47:0]), .sp4_r_v_b_04({net1250[0],
     net1250[1], net1250[2], net1250[3], net1250[4], net1250[5],
     net1250[6], net1250[7], net1250[8], net1250[9], net1250[10],
     net1250[11], net1250[12], net1250[13], net1250[14], net1250[15],
     net1250[16], net1250[17], net1250[18], net1250[19], net1250[20],
     net1250[21], net1250[22], net1250[23], net1250[24], net1250[25],
     net1250[26], net1250[27], net1250[28], net1250[29], net1250[30],
     net1250[31], net1250[32], net1250[33], net1250[34], net1250[35],
     net1250[36], net1250[37], net1250[38], net1250[39], net1250[40],
     net1250[41], net1250[42], net1250[43], net1250[44], net1250[45],
     net1250[46], net1250[47]}), .sp4_r_v_b_03({net1251[0], net1251[1],
     net1251[2], net1251[3], net1251[4], net1251[5], net1251[6],
     net1251[7], net1251[8], net1251[9], net1251[10], net1251[11],
     net1251[12], net1251[13], net1251[14], net1251[15], net1251[16],
     net1251[17], net1251[18], net1251[19], net1251[20], net1251[21],
     net1251[22], net1251[23], net1251[24], net1251[25], net1251[26],
     net1251[27], net1251[28], net1251[29], net1251[30], net1251[31],
     net1251[32], net1251[33], net1251[34], net1251[35], net1251[36],
     net1251[37], net1251[38], net1251[39], net1251[40], net1251[41],
     net1251[42], net1251[43], net1251[44], net1251[45], net1251[46],
     net1251[47]}), .sp4_r_v_b_02({net1252[0], net1252[1], net1252[2],
     net1252[3], net1252[4], net1252[5], net1252[6], net1252[7],
     net1252[8], net1252[9], net1252[10], net1252[11], net1252[12],
     net1252[13], net1252[14], net1252[15], net1252[16], net1252[17],
     net1252[18], net1252[19], net1252[20], net1252[21], net1252[22],
     net1252[23], net1252[24], net1252[25], net1252[26], net1252[27],
     net1252[28], net1252[29], net1252[30], net1252[31], net1252[32],
     net1252[33], net1252[34], net1252[35], net1252[36], net1252[37],
     net1252[38], net1252[39], net1252[40], net1252[41], net1252[42],
     net1252[43], net1252[44], net1252[45], net1252[46], net1252[47]}),
     .sp4_r_v_b_01(sp4_v_b_08_09[47:0]), .sp4_h_r_04({net1254[0],
     net1254[1], net1254[2], net1254[3], net1254[4], net1254[5],
     net1254[6], net1254[7], net1254[8], net1254[9], net1254[10],
     net1254[11], net1254[12], net1254[13], net1254[14], net1254[15],
     net1254[16], net1254[17], net1254[18], net1254[19], net1254[20],
     net1254[21], net1254[22], net1254[23], net1254[24], net1254[25],
     net1254[26], net1254[27], net1254[28], net1254[29], net1254[30],
     net1254[31], net1254[32], net1254[33], net1254[34], net1254[35],
     net1254[36], net1254[37], net1254[38], net1254[39], net1254[40],
     net1254[41], net1254[42], net1254[43], net1254[44], net1254[45],
     net1254[46], net1254[47]}), .sp4_h_r_03({net1255[0], net1255[1],
     net1255[2], net1255[3], net1255[4], net1255[5], net1255[6],
     net1255[7], net1255[8], net1255[9], net1255[10], net1255[11],
     net1255[12], net1255[13], net1255[14], net1255[15], net1255[16],
     net1255[17], net1255[18], net1255[19], net1255[20], net1255[21],
     net1255[22], net1255[23], net1255[24], net1255[25], net1255[26],
     net1255[27], net1255[28], net1255[29], net1255[30], net1255[31],
     net1255[32], net1255[33], net1255[34], net1255[35], net1255[36],
     net1255[37], net1255[38], net1255[39], net1255[40], net1255[41],
     net1255[42], net1255[43], net1255[44], net1255[45], net1255[46],
     net1255[47]}), .sp4_h_r_02({net1256[0], net1256[1], net1256[2],
     net1256[3], net1256[4], net1256[5], net1256[6], net1256[7],
     net1256[8], net1256[9], net1256[10], net1256[11], net1256[12],
     net1256[13], net1256[14], net1256[15], net1256[16], net1256[17],
     net1256[18], net1256[19], net1256[20], net1256[21], net1256[22],
     net1256[23], net1256[24], net1256[25], net1256[26], net1256[27],
     net1256[28], net1256[29], net1256[30], net1256[31], net1256[32],
     net1256[33], net1256[34], net1256[35], net1256[36], net1256[37],
     net1256[38], net1256[39], net1256[40], net1256[41], net1256[42],
     net1256[43], net1256[44], net1256[45], net1256[46], net1256[47]}),
     .sp4_h_r_01({net1257[0], net1257[1], net1257[2], net1257[3],
     net1257[4], net1257[5], net1257[6], net1257[7], net1257[8],
     net1257[9], net1257[10], net1257[11], net1257[12], net1257[13],
     net1257[14], net1257[15], net1257[16], net1257[17], net1257[18],
     net1257[19], net1257[20], net1257[21], net1257[22], net1257[23],
     net1257[24], net1257[25], net1257[26], net1257[27], net1257[28],
     net1257[29], net1257[30], net1257[31], net1257[32], net1257[33],
     net1257[34], net1257[35], net1257[36], net1257[37], net1257[38],
     net1257[39], net1257[40], net1257[41], net1257[42], net1257[43],
     net1257[44], net1257[45], net1257[46], net1257[47]}),
     .sp4_h_l_03(sp4_h_l_07_11[47:0]),
     .sp4_h_l_02(sp4_h_l_07_10[47:0]),
     .sp4_h_l_01(sp4_h_l_07_09[47:0]), .bl(bl[53:0]),
     .bot_op_01(bot_op_07_09[7:0]), .sp12_h_l_01(sp12_h_l_07_09[23:0]),
     .sp12_h_l_02(sp12_h_l_07_10[23:0]),
     .sp12_h_l_03(sp12_h_l_07_11[23:0]),
     .sp12_h_l_04(sp12_h_l_07_12[23:0]),
     .sp4_v_b_04(sp4_v_b_07_12[47:0]),
     .sp4_v_b_03(sp4_v_b_07_11[47:0]),
     .sp4_v_b_02(sp4_v_b_07_10[47:0]), .bnr_op_01(bnr_op_07_09[7:0]),
     .sp4_h_l_05(sp4_h_l_07_13[47:0]),
     .sp4_h_l_06(sp4_h_l_07_14[47:0]),
     .sp4_h_l_07(sp4_h_l_07_15[47:0]),
     .sp4_h_l_08(sp4_h_l_07_16[47:0]), .sp4_h_r_08({net1275[0],
     net1275[1], net1275[2], net1275[3], net1275[4], net1275[5],
     net1275[6], net1275[7], net1275[8], net1275[9], net1275[10],
     net1275[11], net1275[12], net1275[13], net1275[14], net1275[15],
     net1275[16], net1275[17], net1275[18], net1275[19], net1275[20],
     net1275[21], net1275[22], net1275[23], net1275[24], net1275[25],
     net1275[26], net1275[27], net1275[28], net1275[29], net1275[30],
     net1275[31], net1275[32], net1275[33], net1275[34], net1275[35],
     net1275[36], net1275[37], net1275[38], net1275[39], net1275[40],
     net1275[41], net1275[42], net1275[43], net1275[44], net1275[45],
     net1275[46], net1275[47]}), .sp4_h_r_07({net1276[0], net1276[1],
     net1276[2], net1276[3], net1276[4], net1276[5], net1276[6],
     net1276[7], net1276[8], net1276[9], net1276[10], net1276[11],
     net1276[12], net1276[13], net1276[14], net1276[15], net1276[16],
     net1276[17], net1276[18], net1276[19], net1276[20], net1276[21],
     net1276[22], net1276[23], net1276[24], net1276[25], net1276[26],
     net1276[27], net1276[28], net1276[29], net1276[30], net1276[31],
     net1276[32], net1276[33], net1276[34], net1276[35], net1276[36],
     net1276[37], net1276[38], net1276[39], net1276[40], net1276[41],
     net1276[42], net1276[43], net1276[44], net1276[45], net1276[46],
     net1276[47]}), .sp4_h_r_06({net1277[0], net1277[1], net1277[2],
     net1277[3], net1277[4], net1277[5], net1277[6], net1277[7],
     net1277[8], net1277[9], net1277[10], net1277[11], net1277[12],
     net1277[13], net1277[14], net1277[15], net1277[16], net1277[17],
     net1277[18], net1277[19], net1277[20], net1277[21], net1277[22],
     net1277[23], net1277[24], net1277[25], net1277[26], net1277[27],
     net1277[28], net1277[29], net1277[30], net1277[31], net1277[32],
     net1277[33], net1277[34], net1277[35], net1277[36], net1277[37],
     net1277[38], net1277[39], net1277[40], net1277[41], net1277[42],
     net1277[43], net1277[44], net1277[45], net1277[46], net1277[47]}),
     .sp4_h_r_05({net1278[0], net1278[1], net1278[2], net1278[3],
     net1278[4], net1278[5], net1278[6], net1278[7], net1278[8],
     net1278[9], net1278[10], net1278[11], net1278[12], net1278[13],
     net1278[14], net1278[15], net1278[16], net1278[17], net1278[18],
     net1278[19], net1278[20], net1278[21], net1278[22], net1278[23],
     net1278[24], net1278[25], net1278[26], net1278[27], net1278[28],
     net1278[29], net1278[30], net1278[31], net1278[32], net1278[33],
     net1278[34], net1278[35], net1278[36], net1278[37], net1278[38],
     net1278[39], net1278[40], net1278[41], net1278[42], net1278[43],
     net1278[44], net1278[45], net1278[46], net1278[47]}),
     .slf_op_05(slf_op_07_13[7:0]), .slf_op_06(slf_op_07_14[7:0]),
     .slf_op_07(slf_op_07_15[7:0]), .slf_op_08(slf_op_07_16[7:0]),
     .rgt_op_08({net1283[0], net1283[1], net1283[2], net1283[3],
     net1283[4], net1283[5], net1283[6], net1283[7]}),
     .rgt_op_07({net1284[0], net1284[1], net1284[2], net1284[3],
     net1284[4], net1284[5], net1284[6], net1284[7]}),
     .rgt_op_06({net1285[0], net1285[1], net1285[2], net1285[3],
     net1285[4], net1285[5], net1285[6], net1285[7]}),
     .rgt_op_05({net1286[0], net1286[1], net1286[2], net1286[3],
     net1286[4], net1286[5], net1286[6], net1286[7]}),
     .lft_op_08(lft_op_07_16[7:0]), .lft_op_07(lft_op_07_15[7:0]),
     .lft_op_06(lft_op_07_14[7:0]), .lft_op_05(lft_op_07_13[7:0]),
     .sp12_h_l_08(sp12_h_l_07_16[23:0]),
     .sp12_h_l_07(sp12_h_l_07_15[23:0]),
     .sp12_h_l_06(sp12_h_l_07_14[23:0]), .sp12_h_r_05({net1294[0],
     net1294[1], net1294[2], net1294[3], net1294[4], net1294[5],
     net1294[6], net1294[7], net1294[8], net1294[9], net1294[10],
     net1294[11], net1294[12], net1294[13], net1294[14], net1294[15],
     net1294[16], net1294[17], net1294[18], net1294[19], net1294[20],
     net1294[21], net1294[22], net1294[23]}), .sp12_h_r_06({net1295[0],
     net1295[1], net1295[2], net1295[3], net1295[4], net1295[5],
     net1295[6], net1295[7], net1295[8], net1295[9], net1295[10],
     net1295[11], net1295[12], net1295[13], net1295[14], net1295[15],
     net1295[16], net1295[17], net1295[18], net1295[19], net1295[20],
     net1295[21], net1295[22], net1295[23]}), .sp12_h_r_07({net1296[0],
     net1296[1], net1296[2], net1296[3], net1296[4], net1296[5],
     net1296[6], net1296[7], net1296[8], net1296[9], net1296[10],
     net1296[11], net1296[12], net1296[13], net1296[14], net1296[15],
     net1296[16], net1296[17], net1296[18], net1296[19], net1296[20],
     net1296[21], net1296[22], net1296[23]}), .sp12_h_r_08({net1297[0],
     net1297[1], net1297[2], net1297[3], net1297[4], net1297[5],
     net1297[6], net1297[7], net1297[8], net1297[9], net1297[10],
     net1297[11], net1297[12], net1297[13], net1297[14], net1297[15],
     net1297[16], net1297[17], net1297[18], net1297[19], net1297[20],
     net1297[21], net1297[22], net1297[23]}),
     .sp12_h_l_05(sp12_h_l_07_13[23:0]), .sp4_r_v_b_05({net1299[0],
     net1299[1], net1299[2], net1299[3], net1299[4], net1299[5],
     net1299[6], net1299[7], net1299[8], net1299[9], net1299[10],
     net1299[11], net1299[12], net1299[13], net1299[14], net1299[15],
     net1299[16], net1299[17], net1299[18], net1299[19], net1299[20],
     net1299[21], net1299[22], net1299[23], net1299[24], net1299[25],
     net1299[26], net1299[27], net1299[28], net1299[29], net1299[30],
     net1299[31], net1299[32], net1299[33], net1299[34], net1299[35],
     net1299[36], net1299[37], net1299[38], net1299[39], net1299[40],
     net1299[41], net1299[42], net1299[43], net1299[44], net1299[45],
     net1299[46], net1299[47]}), .sp4_r_v_b_06({net1300[0], net1300[1],
     net1300[2], net1300[3], net1300[4], net1300[5], net1300[6],
     net1300[7], net1300[8], net1300[9], net1300[10], net1300[11],
     net1300[12], net1300[13], net1300[14], net1300[15], net1300[16],
     net1300[17], net1300[18], net1300[19], net1300[20], net1300[21],
     net1300[22], net1300[23], net1300[24], net1300[25], net1300[26],
     net1300[27], net1300[28], net1300[29], net1300[30], net1300[31],
     net1300[32], net1300[33], net1300[34], net1300[35], net1300[36],
     net1300[37], net1300[38], net1300[39], net1300[40], net1300[41],
     net1300[42], net1300[43], net1300[44], net1300[45], net1300[46],
     net1300[47]}), .sp4_r_v_b_07({net1301[0], net1301[1], net1301[2],
     net1301[3], net1301[4], net1301[5], net1301[6], net1301[7],
     net1301[8], net1301[9], net1301[10], net1301[11], net1301[12],
     net1301[13], net1301[14], net1301[15], net1301[16], net1301[17],
     net1301[18], net1301[19], net1301[20], net1301[21], net1301[22],
     net1301[23], net1301[24], net1301[25], net1301[26], net1301[27],
     net1301[28], net1301[29], net1301[30], net1301[31], net1301[32],
     net1301[33], net1301[34], net1301[35], net1301[36], net1301[37],
     net1301[38], net1301[39], net1301[40], net1301[41], net1301[42],
     net1301[43], net1301[44], net1301[45], net1301[46], net1301[47]}),
     .sp4_r_v_b_08({net1302[0], net1302[1], net1302[2], net1302[3],
     net1302[4], net1302[5], net1302[6], net1302[7], net1302[8],
     net1302[9], net1302[10], net1302[11], net1302[12], net1302[13],
     net1302[14], net1302[15], net1302[16], net1302[17], net1302[18],
     net1302[19], net1302[20], net1302[21], net1302[22], net1302[23],
     net1302[24], net1302[25], net1302[26], net1302[27], net1302[28],
     net1302[29], net1302[30], net1302[31], net1302[32], net1302[33],
     net1302[34], net1302[35], net1302[36], net1302[37], net1302[38],
     net1302[39], net1302[40], net1302[41], net1302[42], net1302[43],
     net1302[44], net1302[45], net1302[46], net1302[47]}),
     .sp4_v_b_08(sp4_v_b_07_16[47:0]),
     .sp4_v_b_07(sp4_v_b_07_15[47:0]),
     .sp4_v_b_06(sp4_v_b_07_14[47:0]),
     .sp4_v_b_05(sp4_v_b_07_13[47:0]), .pgate(pgate_r[127:0]),
     .reset_b(reset_b_r[127:0]), .wl(wl_r[127:0]),
     .sp12_v_t_08({net1310[0], net1310[1], net1310[2], net1310[3],
     net1310[4], net1310[5], net1310[6], net1310[7], net1310[8],
     net1310[9], net1310[10], net1310[11], net1310[12], net1310[13],
     net1310[14], net1310[15], net1310[16], net1310[17], net1310[18],
     net1310[19], net1310[20], net1310[21], net1310[22], net1310[23]}),
     .tnr_op_08({slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0], slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0]}), .top_op_08({slf_op_07_17[3],
     slf_op_07_17[2], slf_op_07_17[1], slf_op_07_17[0],
     slf_op_07_17[3], slf_op_07_17[2], slf_op_07_17[1],
     slf_op_07_17[0]}), .tnl_op_08({tnl_op_07_16[3], tnl_op_07_16[2],
     tnl_op_07_16[1], tnl_op_07_16[0], tnl_op_07_16[3],
     tnl_op_07_16[2], tnl_op_07_16[1], tnl_op_07_16[0]}),
     .sp4_v_t_08({net1314[0], net1314[1], net1314[2], net1314[3],
     net1314[4], net1314[5], net1314[6], net1314[7], net1314[8],
     net1314[9], net1314[10], net1314[11], net1314[12], net1314[13],
     net1314[14], net1314[15], net1314[16], net1314[17], net1314[18],
     net1314[19], net1314[20], net1314[21], net1314[22], net1314[23],
     net1314[24], net1314[25], net1314[26], net1314[27], net1314[28],
     net1314[29], net1314[30], net1314[31], net1314[32], net1314[33],
     net1314[34], net1314[35], net1314[36], net1314[37], net1314[38],
     net1314[39], net1314[40], net1314[41], net1314[42], net1314[43],
     net1314[44], net1314[45], net1314[46], net1314[47]}),
     .lc_bot(lc_bot_07_09), .op_vic(net1316),
     .sp12_v_b_01(sp12_v_b_07_09[23:0]), .glb_netwk_t({net1318[0],
     net1318[1], net1318[2], net1318[3], net1318[4], net1318[5],
     net1318[6], net1318[7]}));
pinlatbuf12p I_pinlatbuf12p_r ( .pad_in(padin_r[13]),
     .icegate(hold_r_t), .cbit(cf_r[15]), .cout(net01448),
     .prog(prog));
pinlatbuf12p I_pinlatbuf12p ( .pad_in(padin_t_r[12]),
     .icegate(hold_t_r), .cbit(cf_t[15]), .cout(padinlat_t_r[0]),
     .prog(prog));

endmodule
// Library - ice8chip, Cell - io_col4_lft_ice8p_v2, View - schematic
// LAST TIME SAVED: Jan 12 15:05:42 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module io_col4_lft_ice8p_v2 ( cbit_colcntl, cf, fabric_out, padeb,
     pado, sdo, slf_op, spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t,
     sp12_h_l, bnl_op, bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold,
     lft_op, mode, padin, pgate, prog, r, reset, sdi, shift, spioeb,
     spiout, tclk, tnl_op, update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [7:0]  cbit_colcntl;
output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;
output [23:0]  cf;

inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;

input [7:0]  glb_netwk;
input [1:0]  padin;
input [15:0]  wl;
input [15:0]  reset;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [1:0]  spiout;
input [1:0]  spioeb;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  tnl_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [1:0]  om;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [3:0]  t_mid;



rm7w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
sbox1_colbdlc_v4 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
io_gmux_x16bare_v4 I_io_gmux_x16bare_v4 (
     .cbit_colcntl(cbit_colcntl[7:0]), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));

endmodule
// Library - ice1chip, Cell - io_lft_top_1x8_ice1f, View - schematic
// LAST TIME SAVED: Apr 11 16:00:35 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module io_lft_top_1x8_ice1f ( cf_l, fabric_out_09, fo_dlyadj, padeb,
     pado, sdo, slf_op_01, slf_op_02, slf_op_03, slf_op_04, slf_op_05,
     slf_op_06, slf_op_07, slf_op_08, tclk_o, SP4_h_l_01, SP4_h_l_02,
     SP4_h_l_03, SP4_h_l_04, SP4_h_l_05, SP4_h_l_06, SP4_h_l_07,
     SP4_h_l_08, SP12_h_l_01, SP12_h_l_02, SP12_h_l_03, SP12_h_l_04,
     SP12_h_l_05, SP12_h_l_06, SP12_h_l_07, SP12_h_l_08, bl, pgate,
     reset_b, sp4_v_b_00_09, sp4_v_t_08, vdd_cntl, wl, bnr_op_00_09,
     bs_en, ceb, glb_netwk_col, hiz_b, hold, jtag_rowtest_mode_rowu1_b,
     last_rsr, mode, padin, prog, r, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, sdi, shift,
     tclk, tnr_op_08, update );
output  fabric_out_09, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu1_b, mode, prog,
     r, sdi, shift, tclk, update;

output [3:0]  slf_op_03;
output [3:0]  slf_op_01;
output [3:0]  slf_op_02;
output [3:0]  slf_op_06;
output [3:0]  slf_op_07;
output [3:0]  slf_op_08;
output [3:0]  slf_op_05;
output [191:0]  cf_l;
output [3:0]  slf_op_04;
output [7:3]  fo_dlyadj;
output [23:12]  padeb;
output [23:12]  pado;

inout [47:0]  SP4_h_l_02;
inout [47:0]  SP4_h_l_08;
inout [23:0]  SP12_h_l_02;
inout [23:0]  SP12_h_l_08;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_06;
inout [23:0]  SP12_h_l_03;
inout [23:0]  SP12_h_l_07;
inout [47:0]  SP4_h_l_04;
inout [47:0]  SP4_h_l_05;
inout [47:0]  SP4_h_l_03;
inout [23:0]  SP12_h_l_05;
inout [23:0]  SP12_h_l_06;
inout [47:0]  SP4_h_l_01;
inout [47:0]  SP4_h_l_07;
inout [15:0]  sp4_v_t_08;
inout [23:0]  SP12_h_l_01;
inout [15:0]  sp4_v_b_00_09;
inout [127:0]  vdd_cntl;
inout [127:0]  pgate;
inout [127:0]  wl;
inout [127:0]  reset_b;
inout [23:0]  SP12_h_l_04;

input [7:0]  bnr_op_00_09;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_04;
input [1:1]  last_rsr;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_08;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_02;
input [23:12]  padin;
input [7:0]  rgt_op_07;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net1002;

wire  [1:0]  net1014;

wire  [1:0]  net1013;

wire  [7:0]  glb_netwk_b;

wire  [7:0]  net1016;

wire  [15:0]  net865;

wire  [7:0]  glb_netwk_t;

wire  [7:0]  net1017;

wire  [7:0]  net884;

wire  [7:0]  net1008;

wire  [1:0]  net1000;

wire  [7:0]  colbuf_cntl_b;

wire  [15:0]  net793;

wire  [1:0]  net1005;

wire  [15:0]  net757;

wire  [15:0]  net829;

wire  [7:0]  net1007;

wire  [1:0]  net1012;

wire  [1:0]  net719;

wire  [15:0]  net901;

wire  [7:0]  net704;

wire  [15:0]  net973;

wire  [1:0]  net1009;

wire  [15:0]  net937;

wire  [1:0]  net1010;

wire  [1:0]  net755;

wire  [1:0]  net1001;

wire  [1:0]  net1003;

wire  [7:0]  colbuf_cntl_t;



tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
io_col4_lft_ice8p_v2 I_io_00_08 ( .cbit_colcntl({net704[0], net704[1],
     net704[2], net704[3], net704[4], net704[5], net704[6],
     net704[7]}), .ceb(ceb), .sdo(net743), .sdi(sdi), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin({net719[0], net719[1]}),
     .pado({net719[0], net719[1]}), .padeb({net1000[0], net1000[1]}),
     .sp4_v_t(sp4_v_t_08[15:0]), .sp4_h_l(SP4_h_l_08[47:0]),
     .sp12_h_l(SP12_h_l_08[23:0]), .prog(prog),
     .spi_ss_in_b({net1012[0], net1012[1]}), .tnl_op(tnr_op_08[7:0]),
     .lft_op(rgt_op_08[7:0]), .bnl_op(rgt_op_07[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b({net757[0], net757[1], net757[2], net757[3], net757[4],
     net757[5], net757[6], net757[7], net757[8], net757[9], net757[10],
     net757[11], net757[12], net757[13], net757[14], net757[15]}),
     .wl(wl[127:112]), .cf(cf_l[191:168]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[127:112]), .slf_op(slf_op_08[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold), .fabric_out(net739));
io_col4_lft_ice8p_v2 I_io_00_07 ( .cbit_colcntl({net1016[0],
     net1016[1], net1016[2], net1016[3], net1016[4], net1016[5],
     net1016[6], net1016[7]}), .ceb(ceb), .sdo(net815), .sdi(net743),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin({net755[0],
     net755[1]}), .pado({net755[0], net755[1]}), .padeb({net1001[0],
     net1001[1]}), .sp4_v_t({net757[0], net757[1], net757[2],
     net757[3], net757[4], net757[5], net757[6], net757[7], net757[8],
     net757[9], net757[10], net757[11], net757[12], net757[13],
     net757[14], net757[15]}), .sp4_h_l(SP4_h_l_07[47:0]),
     .sp12_h_l(SP12_h_l_07[23:0]), .prog(prog),
     .spi_ss_in_b({net1013[0], net1013[1]}), .tnl_op(rgt_op_08[7:0]),
     .lft_op(rgt_op_07[7:0]), .bnl_op(rgt_op_06[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b({net829[0], net829[1], net829[2], net829[3], net829[4],
     net829[5], net829[6], net829[7], net829[8], net829[9], net829[10],
     net829[11], net829[12], net829[13], net829[14], net829[15]}),
     .wl(wl[111:96]), .cf(cf_l[167:144]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[111:96]), .slf_op(slf_op_07[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold), .fabric_out(net775));
io_col4_lft_ice8p_v2 I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net959), .sdi(net779), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[21:20]), .pado(pado[21:20]),
     .padeb(padeb[21:20]), .sp4_v_t({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7], net793[8],
     net793[9], net793[10], net793[11], net793[12], net793[13],
     net793[14], net793[15]}), .sp4_h_l(SP4_h_l_05[47:0]),
     .sp12_h_l(SP12_h_l_05[23:0]), .prog(prog),
     .spi_ss_in_b({net1003[0], net1003[1]}), .tnl_op(rgt_op_06[7:0]),
     .lft_op(rgt_op_05[7:0]), .bnl_op(rgt_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]), .sp4_v_b({net973[0],
     net973[1], net973[2], net973[3], net973[4], net973[5], net973[6],
     net973[7], net973[8], net973[9], net973[10], net973[11],
     net973[12], net973[13], net973[14], net973[15]}), .wl(wl[79:64]),
     .cf(cf_l[119:96]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[6]));
io_col4_lft_ice8p_v2 I_io_00_06 ( .cbit_colcntl({net1017[0],
     net1017[1], net1017[2], net1017[3], net1017[4], net1017[5],
     net1017[6], net1017[7]}), .ceb(ceb), .sdo(net779), .sdi(net815),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[23:22]), .pado(pado[23:22]), .padeb(padeb[23:22]),
     .sp4_v_t({net829[0], net829[1], net829[2], net829[3], net829[4],
     net829[5], net829[6], net829[7], net829[8], net829[9], net829[10],
     net829[11], net829[12], net829[13], net829[14], net829[15]}),
     .sp4_h_l(SP4_h_l_06[47:0]), .sp12_h_l(SP12_h_l_06[23:0]),
     .prog(prog), .spi_ss_in_b({net1010[0], net1010[1]}),
     .tnl_op(rgt_op_07[7:0]), .lft_op(rgt_op_06[7:0]),
     .bnl_op(rgt_op_05[7:0]), .pgate(pgate[95:80]),
     .reset(reset_b[95:80]), .sp4_v_b({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7], net793[8],
     net793[9], net793[10], net793[11], net793[12], net793[13],
     net793[14], net793[15]}), .wl(wl[95:80]), .cf(cf_l[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[7]));
io_col4_lft_ice8p_v2 I_io_00_02 ( .cbit_colcntl({net1007[0],
     net1007[1], net1007[2], net1007[3], net1007[4], net1007[5],
     net1007[6], net1007[7]}), .ceb(ceb), .sdo(net887), .sdi(net851),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[15:14]), .pado(pado[15:14]), .padeb(padeb[15:14]),
     .sp4_v_t({net865[0], net865[1], net865[2], net865[3], net865[4],
     net865[5], net865[6], net865[7], net865[8], net865[9], net865[10],
     net865[11], net865[12], net865[13], net865[14], net865[15]}),
     .sp4_h_l(SP4_h_l_02[47:0]), .sp12_h_l(SP12_h_l_02[23:0]),
     .prog(prog), .spi_ss_in_b({net1014[0], net1014[1]}),
     .tnl_op(rgt_op_03[7:0]), .lft_op(rgt_op_02[7:0]),
     .bnl_op(rgt_op_01[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15]}), .wl(wl[31:16]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[3]));
io_col4_lft_ice8p_v2 I_io_00_01 ( .cbit_colcntl({net884[0], net884[1],
     net884[2], net884[3], net884[4], net884[5], net884[6],
     net884[7]}), .ceb(ceb), .sdo(sdo), .sdi(net887), .spiout({tiegnd,
     last_rsr[1]}), .cdone_in(jtag_rowtest_mode_rowu1_b),
     .spioeb({tievdd, tiegnd}), .mode(mode), .shift(shift),
     .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[13:12]), .pado(pado[13:12]),
     .padeb(padeb[13:12]), .sp4_v_t({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15]}), .sp4_h_l(SP4_h_l_01[47:0]),
     .sp12_h_l(SP12_h_l_01[23:0]), .prog(prog),
     .spi_ss_in_b({net1005[0], net1005[1]}), .tnl_op(rgt_op_02[7:0]),
     .lft_op(rgt_op_01[7:0]), .bnl_op(bnr_op_00_09[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_v_b_00_09[15:0]), .wl(wl[15:0]), .cf(cf_l[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold),
     .fabric_out(fabric_out_09));
io_col4_lft_ice8p_v2 I_io_00_03 ( .cbit_colcntl({net1008[0],
     net1008[1], net1008[2], net1008[3], net1008[4], net1008[5],
     net1008[6], net1008[7]}), .ceb(ceb), .sdo(net851), .sdi(net923),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update),
     .padin(padin[17:16]), .pado(pado[17:16]), .padeb(padeb[17:16]),
     .sp4_v_t({net937[0], net937[1], net937[2], net937[3], net937[4],
     net937[5], net937[6], net937[7], net937[8], net937[9], net937[10],
     net937[11], net937[12], net937[13], net937[14], net937[15]}),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b({net1009[0], net1009[1]}),
     .tnl_op(rgt_op_04[7:0]), .lft_op(rgt_op_03[7:0]),
     .bnl_op(rgt_op_02[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b({net865[0], net865[1], net865[2],
     net865[3], net865[4], net865[5], net865[6], net865[7], net865[8],
     net865[9], net865[10], net865[11], net865[12], net865[13],
     net865[14], net865[15]}), .wl(wl[47:32]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[4]));
io_col4_lft_ice8p_v2 I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net923), .sdi(net959), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[19:18]), .pado(pado[19:18]),
     .padeb(padeb[19:18]), .sp4_v_t({net973[0], net973[1], net973[2],
     net973[3], net973[4], net973[5], net973[6], net973[7], net973[8],
     net973[9], net973[10], net973[11], net973[12], net973[13],
     net973[14], net973[15]}), .sp4_h_l(SP4_h_l_04[47:0]),
     .sp12_h_l(SP12_h_l_04[23:0]), .prog(prog),
     .spi_ss_in_b({net1002[0], net1002[1]}), .tnl_op(rgt_op_05[7:0]),
     .lft_op(rgt_op_04[7:0]), .bnl_op(rgt_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]), .sp4_v_b({net937[0],
     net937[1], net937[2], net937[3], net937[4], net937[5], net937[6],
     net937[7], net937[8], net937[9], net937[10], net937[11],
     net937[12], net937[13], net937[14], net937[15]}), .wl(wl[63:48]),
     .cf(cf_l[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[5]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - ice1chip, Cell - io_top_lft_1x6_ice1f, View - schematic
// LAST TIME SAVED: Mar  5 17:03:41 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module io_top_lft_1x6_ice1f ( bs_en_o, ceb_o, cf_top_l,
     fabric_out_06_17, hiz_b_o, mode_o, padeb_t_l, pado_t_l, r_o, sdo,
     shift_o, slf_op_01_17, slf_op_02_17, slf_op_03_17, slf_op_04_17,
     slf_op_05_17, slf_op_06_17, tclk_o, update_o, bl_01, bl_02, bl_03,
     bl_04, bl_05, bl_06, sp4_h_l_01_17, sp4_h_r_06_17, sp4_v_b_01_17,
     sp4_v_b_02_17, sp4_v_b_03_17, sp4_v_b_04_17, sp4_v_b_05_17,
     sp4_v_b_06_17, sp12_v_b_01_17, sp12_v_b_02_17, sp12_v_b_03_17,
     sp12_v_b_04_17, sp12_v_b_05_17, sp12_v_b_06_17, bnl_op_01_17,
     bnr_op_06_17, bs_en_i, ceb_i, glb_net_01, glb_net_02, glb_net_03,
     glb_net_04, glb_net_05, glb_net_06, hiz_b_i, hold_t_l,
     lft_op_01_17, lft_op_02_17, lft_op_03_17, lft_op_04_17,
     lft_op_05_17, lft_op_06_17, mode_i, padin_t_l, pgate_l, prog, r_i,
     reset_l, sdi, shift_i, tclk_i, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_06_17, hiz_b_o, mode_o, r_o, sdo,
     shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_01_17;
output [3:0]  slf_op_03_17;
output [3:0]  slf_op_04_17;
output [3:0]  slf_op_05_17;
output [11:0]  pado_t_l;
output [11:0]  padeb_t_l;
output [3:0]  slf_op_06_17;
output [3:0]  slf_op_02_17;
output [143:0]  cf_top_l;

inout [23:0]  sp12_v_b_04_17;
inout [23:0]  sp12_v_b_03_17;
inout [47:0]  sp4_v_b_01_17;
inout [23:0]  sp12_v_b_01_17;
inout [23:0]  sp12_v_b_05_17;
inout [15:0]  sp4_h_r_06_17;
inout [53:0]  bl_01;
inout [53:0]  bl_04;
inout [41:0]  bl_03;
inout [15:0]  sp4_h_l_01_17;
inout [53:0]  bl_05;
inout [53:0]  bl_06;
inout [23:0]  sp12_v_b_06_17;
inout [23:0]  sp12_v_b_02_17;
inout [47:0]  sp4_v_b_03_17;
inout [47:0]  sp4_v_b_06_17;
inout [47:0]  sp4_v_b_04_17;
inout [47:0]  sp4_v_b_02_17;
inout [47:0]  sp4_v_b_05_17;
inout [53:0]  bl_02;

input [7:0]  lft_op_03_17;
input [7:0]  glb_net_01;
input [7:0]  glb_net_03;
input [7:0]  bnl_op_01_17;
input [15:0]  wl_l;
input [7:0]  lft_op_01_17;
input [7:0]  glb_net_06;
input [7:0]  lft_op_05_17;
input [7:0]  lft_op_02_17;
input [11:0]  padin_t_l;
input [7:0]  glb_net_02;
input [15:0]  pgate_l;
input [7:0]  bnr_op_06_17;
input [7:0]  lft_op_04_17;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_04;
input [7:0]  lft_op_06_17;
input [7:0]  glb_net_05;
input [15:0]  reset_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  net1532;

wire  [1:0]  net1319;

wire  [15:0]  net1427;

wire  [1:0]  net1312;

wire  [1:0]  net1318;

wire  [1:0]  net1361;

wire  [15:0]  net1392;

wire  [15:0]  net1357;

wire  [1:0]  net1501;

wire  [1:0]  net1431;

wire  [15:0]  net1462;



tckbufx32_ice8p I_tck_halfbankcenter ( .in(net0262), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));
scan_buf_ice8p I345 ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net0262), .shift_o(shift_o),
     .sdo(net1482), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_top_ice8p I_IO_02_17 ( .sdo(net1412), .sdi(net1342),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1427[0], net1427[1], net1427[2],
     net1427[3], net1427[4], net1427[5], net1427[6], net1427[7],
     net1427[8], net1427[9], net1427[10], net1427[11], net1427[12],
     net1427[13], net1427[14], net1427[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[3:2]),
     .pado(pado_t_l[3:2]), .padeb(padeb_t_l[3:2]),
     .sp4_v_b({net1357[0], net1357[1], net1357[2], net1357[3],
     net1357[4], net1357[5], net1357[6], net1357[7], net1357[8],
     net1357[9], net1357[10], net1357[11], net1357[12], net1357[13],
     net1357[14], net1357[15]}), .sp4_h_l(sp4_v_b_02_17[47:0]),
     .sp12_h_l(sp12_v_b_02_17[23:0]), .prog(prog),
     .spi_ss_in_b({net1361[0], net1361[1]}),
     .tnl_op(lft_op_01_17[7:0]), .lft_op(lft_op_02_17[7:0]),
     .bnl_op(lft_op_03_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[47:24]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_17[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_t_l), .fabric_out(net1320));
io_col4_top_ice8p I_IO_03_17_bram ( .sdo(net1342), .sdi(net1377),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1357[0], net1357[1], net1357[2],
     net1357[3], net1357[4], net1357[5], net1357[6], net1357[7],
     net1357[8], net1357[9], net1357[10], net1357[11], net1357[12],
     net1357[13], net1357[14], net1357[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[5:4]),
     .pado(pado_t_l[5:4]), .padeb(padeb_t_l[5:4]),
     .sp4_v_b({net1392[0], net1392[1], net1392[2], net1392[3],
     net1392[4], net1392[5], net1392[6], net1392[7], net1392[8],
     net1392[9], net1392[10], net1392[11], net1392[12], net1392[13],
     net1392[14], net1392[15]}), .sp4_h_l(sp4_v_b_03_17[47:0]),
     .sp12_h_l(sp12_v_b_03_17[23:0]), .prog(prog),
     .spi_ss_in_b({net1318[0], net1318[1]}),
     .tnl_op(lft_op_02_17[7:0]), .lft_op(lft_op_03_17[7:0]),
     .bnl_op(lft_op_04_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[71:48]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_17[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_t_l), .fabric_out(net1410));
io_col4_top_ice8p I_IO_01_17 ( .sdo(sdo), .sdi(net1412),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_01_17[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[1:0]),
     .pado(pado_t_l[1:0]), .padeb(padeb_t_l[1:0]),
     .sp4_v_b({net1427[0], net1427[1], net1427[2], net1427[3],
     net1427[4], net1427[5], net1427[6], net1427[7], net1427[8],
     net1427[9], net1427[10], net1427[11], net1427[12], net1427[13],
     net1427[14], net1427[15]}), .sp4_h_l(sp4_v_b_01_17[47:0]),
     .sp12_h_l(sp12_v_b_01_17[23:0]), .prog(prog),
     .spi_ss_in_b({net1431[0], net1431[1]}),
     .tnl_op(bnl_op_01_17[7:0]), .lft_op(lft_op_01_17[7:0]),
     .bnl_op(lft_op_02_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[23:0]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_17[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_t_l), .fabric_out(net1445));
io_col4_top_ice8p I_IO_05_17 ( .sdo(net1517), .sdi(net1447),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1532[0], net1532[1], net1532[2],
     net1532[3], net1532[4], net1532[5], net1532[6], net1532[7],
     net1532[8], net1532[9], net1532[10], net1532[11], net1532[12],
     net1532[13], net1532[14], net1532[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[9:8]),
     .pado(pado_t_l[9:8]), .padeb(padeb_t_l[9:8]),
     .sp4_v_b({net1462[0], net1462[1], net1462[2], net1462[3],
     net1462[4], net1462[5], net1462[6], net1462[7], net1462[8],
     net1462[9], net1462[10], net1462[11], net1462[12], net1462[13],
     net1462[14], net1462[15]}), .sp4_h_l(sp4_v_b_05_17[47:0]),
     .sp12_h_l(sp12_v_b_05_17[23:0]), .prog(prog),
     .spi_ss_in_b({net1319[0], net1319[1]}),
     .tnl_op(lft_op_04_17[7:0]), .lft_op(lft_op_05_17[7:0]),
     .bnl_op(lft_op_06_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[119:96]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_17[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_t_l), .fabric_out(net1480));
io_col4_top_ice8p I_IO_06_17 ( .sdo(net1447), .sdi(net1482),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1462[0], net1462[1], net1462[2],
     net1462[3], net1462[4], net1462[5], net1462[6], net1462[7],
     net1462[8], net1462[9], net1462[10], net1462[11], net1462[12],
     net1462[13], net1462[14], net1462[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[11:10]),
     .pado(pado_t_l[11:10]), .padeb(padeb_t_l[11:10]),
     .sp4_v_b(sp4_h_r_06_17[15:0]), .sp4_h_l(sp4_v_b_06_17[47:0]),
     .sp12_h_l(sp12_v_b_06_17[23:0]), .prog(prog),
     .spi_ss_in_b({net1501[0], net1501[1]}),
     .tnl_op(lft_op_05_17[7:0]), .lft_op(lft_op_06_17[7:0]),
     .bnl_op(bnr_op_06_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_06[5], bl_06[4], bl_06[37],
     bl_06[36], bl_06[35], bl_06[34], bl_06[33], bl_06[32], bl_06[14],
     bl_06[20], bl_06[19], bl_06[18], bl_06[17], bl_06[16], bl_06[27],
     bl_06[26], bl_06[25], bl_06[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[143:120]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_17[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_t_l), .fabric_out(fabric_out_06_17));
io_col4_top_ice8p I_IO_04_17 ( .sdo(net1377), .sdi(net1517),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net1392[0], net1392[1], net1392[2],
     net1392[3], net1392[4], net1392[5], net1392[6], net1392[7],
     net1392[8], net1392[9], net1392[10], net1392[11], net1392[12],
     net1392[13], net1392[14], net1392[15]}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_t_l[7:6]),
     .pado(pado_t_l[7:6]), .padeb(padeb_t_l[7:6]),
     .sp4_v_b({net1532[0], net1532[1], net1532[2], net1532[3],
     net1532[4], net1532[5], net1532[6], net1532[7], net1532[8],
     net1532[9], net1532[10], net1532[11], net1532[12], net1532[13],
     net1532[14], net1532[15]}), .sp4_h_l(sp4_v_b_04_17[47:0]),
     .sp12_h_l(sp12_v_b_04_17[23:0]), .prog(prog),
     .spi_ss_in_b({net1312[0], net1312[1]}),
     .tnl_op(lft_op_03_17[7:0]), .lft_op(lft_op_04_17[7:0]),
     .bnl_op(lft_op_05_17[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf(cf_top_l[95:72]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_17[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_t_l), .fabric_out(net1313));

endmodule
// Library - ice1chip, Cell - quad_tl_ice1, View - schematic
// LAST TIME SAVED: Apr 26 17:02:35 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module quad_tl_ice1 ( bm_aa_2bot, bm_ab_2bot, bm_sdo_o, bs_en_o, ceb_o,
     cf_l, cf_t, fabric_out_00_09, fabric_out_06_17, fo_dlyadj,
     hiz_b_o, mode_o, padeb_l_t, padeb_t_l, padin_00_09a, padin_06_17b,
     pado_l_t, pado_t_l, r_o, sdo, shift_o, slf_op_00_09, slf_op_01_09,
     slf_op_02_09, slf_op_03_09, slf_op_04_09, slf_op_05_09,
     slf_op_06_09, slf_op_06_10, slf_op_06_11, slf_op_06_12,
     slf_op_06_13, slf_op_06_14, slf_op_06_15, slf_op_06_16,
     slf_op_06_17, tclk_o, update_o, bl, pgate_l, reset_b_l,
     sp4_h_r_06_09, sp4_h_r_06_10, sp4_h_r_06_11, sp4_h_r_06_12,
     sp4_h_r_06_13, sp4_h_r_06_14, sp4_h_r_06_15, sp4_h_r_06_16,
     sp4_h_r_06_17, sp4_r_v_b_06_09, sp4_r_v_b_06_10, sp4_r_v_b_06_11,
     sp4_r_v_b_06_12, sp4_r_v_b_06_13, sp4_r_v_b_06_14,
     sp4_r_v_b_06_15, sp4_r_v_b_06_16, sp4_v_b_00_09, sp4_v_b_01_09,
     sp4_v_b_02_09, sp4_v_b_03_09, sp4_v_b_04_09, sp4_v_b_05_09,
     sp4_v_b_06_09, sp12_h_r_06_09, sp12_h_r_06_10, sp12_h_r_06_11,
     sp12_h_r_06_12, sp12_h_r_06_13, sp12_h_r_06_14, sp12_h_r_06_15,
     sp12_h_r_06_16, sp12_v_b_01_09, sp12_v_b_02_09, sp12_v_b_03_09,
     sp12_v_b_04_09, sp12_v_b_05_09, sp12_v_b_06_09, vdd_cntl_l, wl_l,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_01_09,
     bnl_op_02_09, bnl_op_03_09, bnl_op_04_09, bnl_op_05_09,
     bnl_op_06_09, bnr_op_00_09, bnr_op_01_09, bnr_op_02_09,
     bnr_op_03_09, bnr_op_04_09, bnr_op_05_09, bnr_op_06_09,
     bot_op_01_09, bot_op_02_09, bot_op_03_09, bot_op_04_09,
     bot_op_05_09, bot_op_06_09, bs_en_i, carry_in_01_09,
     carry_in_02_09, carry_in_04_09, carry_in_05_09, carry_in_06_09,
     ceb_i, glb_in, hiz_b_i, hold_l_t, hold_t_l,
     jtag_rowtest_mode_rowu1_b, last_rsr, lc_bot_01_09, lc_bot_02_09,
     lc_bot_04_09, lc_bot_05_09, lc_bot_06_09, mode_i, padin_l_t,
     padin_t_l, prog, purst, r_i, rgt_op_06_09, rgt_op_06_10,
     rgt_op_06_11, rgt_op_06_12, rgt_op_06_13, rgt_op_06_14,
     rgt_op_06_15, rgt_op_06_16, sdi, shift_i, tclk_i, tnr_op_06_16,
     update_i );
output  bs_en_o, ceb_o, fabric_out_00_09, fabric_out_06_17, hiz_b_o,
     mode_o, padin_00_09a, padin_06_17b, r_o, sdo, shift_o, tclk_o,
     update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, carry_in_01_09, carry_in_02_09,
     carry_in_04_09, carry_in_05_09, carry_in_06_09, ceb_i, hiz_b_i,
     hold_l_t, hold_t_l, jtag_rowtest_mode_rowu1_b, lc_bot_01_09,
     lc_bot_02_09, lc_bot_04_09, lc_bot_05_09, lc_bot_06_09, mode_i,
     prog, purst, r_i, sdi, shift_i, tclk_i, update_i;

output [7:0]  slf_op_03_09;
output [23:12]  pado_l_t;
output [7:0]  slf_op_06_13;
output [7:0]  slf_op_02_09;
output [10:0]  bm_ab_2bot;
output [7:0]  slf_op_06_16;
output [7:0]  slf_op_06_12;
output [7:0]  slf_op_01_09;
output [7:0]  slf_op_05_09;
output [7:0]  slf_op_06_10;
output [3:0]  slf_op_06_17;
output [7:0]  slf_op_06_11;
output [7:3]  fo_dlyadj;
output [3:0]  slf_op_00_09;
output [10:0]  bm_aa_2bot;
output [7:0]  slf_op_06_09;
output [7:0]  slf_op_06_14;
output [23:12]  padeb_l_t;
output [11:0]  pado_t_l;
output [143:0]  cf_t;
output [191:0]  cf_l;
output [11:0]  padeb_t_l;
output [7:0]  slf_op_04_09;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_06_15;

inout [47:0]  sp4_r_v_b_06_10;
inout [47:0]  sp4_r_v_b_06_16;
inout [47:0]  sp4_v_b_01_09;
inout [47:0]  sp4_v_b_06_09;
inout [47:0]  sp4_h_r_06_13;
inout [47:0]  sp4_h_r_06_14;
inout [23:0]  sp12_h_r_06_15;
inout [15:0]  sp4_v_b_00_09;
inout [47:0]  sp4_r_v_b_06_09;
inout [47:0]  sp4_h_r_06_09;
inout [15:0]  sp4_h_r_06_17;
inout [23:0]  sp12_v_b_05_09;
inout [47:0]  sp4_r_v_b_06_13;
inout [143:0]  pgate_l;
inout [23:0]  sp12_h_r_06_12;
inout [23:0]  sp12_v_b_03_09;
inout [143:0]  vdd_cntl_l;
inout [23:0]  sp12_v_b_04_09;
inout [329:0]  bl;
inout [23:0]  sp12_h_r_06_13;
inout [23:0]  sp12_v_b_01_09;
inout [143:0]  reset_b_l;
inout [47:0]  sp4_r_v_b_06_11;
inout [23:0]  sp12_v_b_02_09;
inout [47:0]  sp4_h_r_06_11;
inout [47:0]  sp4_h_r_06_10;
inout [47:0]  sp4_h_r_06_16;
inout [23:0]  sp12_h_r_06_09;
inout [47:0]  sp4_r_v_b_06_14;
inout [23:0]  sp12_v_b_06_09;
inout [47:0]  sp4_v_b_02_09;
inout [47:0]  sp4_v_b_05_09;
inout [47:0]  sp4_v_b_03_09;
inout [47:0]  sp4_r_v_b_06_15;
inout [23:0]  sp12_h_r_06_10;
inout [23:0]  sp12_h_r_06_14;
inout [47:0]  sp4_h_r_06_15;
inout [47:0]  sp4_r_v_b_06_12;
inout [23:0]  sp12_h_r_06_11;
inout [23:0]  sp12_h_r_06_16;
inout [143:0]  wl_l;
inout [47:0]  sp4_h_r_06_12;
inout [47:0]  sp4_v_b_04_09;

input [7:0]  rgt_op_06_15;
input [1:0]  bm_sdi_i;
input [7:0]  rgt_op_06_14;
input [7:0]  rgt_op_06_11;
input [7:0]  bnl_op_05_09;
input [7:0]  bot_op_02_09;
input [7:0]  bm_sa_i;
input [7:0]  bnr_op_05_09;
input [1:0]  bm_sweb_i;
input [7:0]  bot_op_04_09;
input [7:0]  bot_op_05_09;
input [7:0]  bot_op_03_09;
input [1:0]  bm_sclkrw_i;
input [3:0]  tnr_op_06_16;
input [7:0]  bnr_op_02_09;
input [7:0]  bot_op_01_09;
input [11:0]  padin_t_l;
input [7:0]  glb_in;
input [7:0]  bnl_op_01_09;
input [7:0]  bnr_op_01_09;
input [7:0]  rgt_op_06_13;
input [7:0]  rgt_op_06_12;
input [7:0]  bnl_op_04_09;
input [7:0]  bnr_op_00_09;
input [7:0]  bnl_op_02_09;
input [1:1]  last_rsr;
input [7:0]  rgt_op_06_10;
input [7:0]  bnl_op_03_09;
input [7:0]  rgt_op_06_09;
input [23:12]  padin_l_t;
input [7:0]  rgt_op_06_16;
input [7:0]  bnr_op_03_09;
input [7:0]  bnl_op_06_09;
input [7:0]  bnr_op_04_09;
input [7:0]  bnr_op_06_09;
input [7:0]  bot_op_06_09;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [47:0]  net961;

wire  [1:0]  net1439;

wire  [7:0]  clk_tree_drv_tl;

wire  [3:0]  slf_op_02_17;

wire  [3:0]  slf_op_01_17;

wire  [3:0]  slf_op_05_17;

wire  [3:0]  slf_op_04_17;

wire  [7:0]  clk_center;

wire  [3:0]  slf_op_08_17;

wire  [3:0]  slf_op_00_15;

wire  [7:0]  net1274;

wire  [47:0]  net765;

wire  [7:0]  net1273;

wire  [3:0]  slf_op_00_11;

wire  [1:0]  bm_sdi_b1_o;

wire  [3:0]  slf_op_00_10;

wire  [3:0]  slf_op_00_12;

wire  [3:0]  slf_op_00_13;

wire  [3:0]  slf_op_00_14;

wire  [3:0]  slf_op_00_16;

wire  [7:0]  net1085;

wire  [7:0]  net1224;

wire  [47:0]  net1151;

wire  [23:0]  net1140;

wire  [47:0]  net956;

wire  [23:0]  net1000;

wire  [47:0]  net827;

wire  [47:0]  net819;

wire  [47:0]  net1196;

wire  [7:0]  net831;

wire  [47:0]  net1445;

wire  [47:0]  net795;

wire  [47:0]  net1049;

wire  [23:0]  net1191;

wire  [23:0]  net1190;

wire  [23:0]  net950;

wire  [47:0]  net763;

wire  [23:0]  net749;

wire  [47:0]  net1246;

wire  [23:0]  net1284;

wire  [47:0]  net1169;

wire  [23:0]  net855;

wire  [47:0]  net1450;

wire  [47:0]  net1172;

wire  [7:0]  net836;

wire  [7:0]  net1214;

wire  [23:0]  net1109;

wire  [7:0]  net832;

wire  [7:0]  net770;

wire  [47:0]  net746;

wire  [23:0]  net856;

wire  [7:0]  net834;

wire  [23:0]  net1233;

wire  [47:0]  net1050;

wire  [7:0]  net931;

wire  [7:0]  net1026;

wire  [7:0]  net833;

wire  [23:0]  net1188;

wire  [47:0]  net1144;

wire  [23:0]  net716;

wire  [7:0]  net769;

wire  [7:0]  net1460;

wire  [23:0]  net1014;

wire  [47:0]  net1303;

wire  [7:0]  net1034;

wire  [23:0]  net948;

wire  [47:0]  net1446;

wire  [47:0]  net1267;

wire  [23:0]  net1286;

wire  [23:0]  net1096;

wire  [23:0]  net851;

wire  [23:0]  net1234;

wire  [23:0]  net1043;

wire  [23:0]  net721;

wire  [47:0]  net979;

wire  [47:0]  net954;

wire  [23:0]  net1236;

wire  [47:0]  net1113;

wire  [47:0]  net1006;

wire  [47:0]  net828;

wire  [23:0]  net1394;

wire  [23:0]  net1283;

wire  [7:0]  net1024;

wire  [23:0]  net1046;

wire  [47:0]  net790;

wire  [23:0]  net1094;

wire  [47:0]  net1148;

wire  [23:0]  net949;

wire  [47:0]  net794;

wire  [23:0]  net748;

wire  [23:0]  net850;

wire  [47:0]  net1099;

wire  [47:0]  net735;

wire  [47:0]  net1193;

wire  [23:0]  net857;

wire  [23:0]  net1285;

wire  [47:0]  net1145;

wire  [47:0]  net1075;

wire  [47:0]  net959;

wire  [23:0]  net1001;

wire  [47:0]  net982;

wire  [47:0]  net1170;

wire  [47:0]  net791;

wire  [7:0]  net695;

wire  [7:0]  net786;

wire  [7:0]  net987;

wire  [7:0]  net989;

wire  [23:0]  net1044;

wire  [47:0]  net1003;

wire  [47:0]  net732;

wire  [23:0]  net740;

wire  [47:0]  net1208;

wire  [47:0]  net1076;

wire  [47:0]  net728;

wire  [7:0]  net1275;

wire  [23:0]  net1093;

wire  [23:0]  net1299;

wire  [7:0]  net773;

wire  [7:0]  net1117;

wire  [7:0]  net772;

wire  [47:0]  net1101;

wire  [7:0]  net1118;

wire  [47:0]  net1146;

wire  [7:0]  net1082;

wire  [47:0]  net1243;

wire  [47:0]  net1051;

wire  [47:0]  net1100;

wire  [7:0]  net1212;

wire  [23:0]  net1138;

wire  [47:0]  net793;

wire  [47:0]  net1194;

wire  [47:0]  net1240;

wire  [47:0]  net764;

wire  [23:0]  net852;

wire  [7:0]  net1307;

wire  [7:0]  net939;

wire  [47:0]  net1055;

wire  [47:0]  net1150;

wire  [23:0]  net1141;

wire  [47:0]  net1005;

wire  [47:0]  net960;

wire  [1:0]  net1441;

wire  [23:0]  net1189;

wire  [23:0]  net951;

wire  [47:0]  net1074;

wire  [47:0]  net1264;

wire  [23:0]  net1045;

wire  [47:0]  net731;

wire  [23:0]  net718;

wire  [7:0]  net990;

wire  [23:0]  net704;

wire  [7:0]  net988;

wire  [23:0]  net756;

wire  [47:0]  net830;

wire  [47:0]  net1288;

wire  [47:0]  net1265;

wire  [47:0]  net1195;

wire  [47:0]  net826;

wire  [23:0]  net1204;

wire  [47:0]  net724;

wire  [47:0]  net1018;

wire  [7:0]  net1451;

wire  [23:0]  net1139;

wire  [47:0]  net1245;

wire  [47:0]  net958;

wire  [47:0]  net825;

wire  [7:0]  net858;

wire  [47:0]  net734;

wire  [15:0]  net820;

wire  [47:0]  net955;

wire  [23:0]  net999;

wire  [7:0]  net1452;

wire  [7:0]  net1083;

wire  [47:0]  net1244;

wire  [47:0]  net1077;

wire  [47:0]  net1098;

wire  [47:0]  net1290;

wire  [47:0]  net980;

wire  [23:0]  net998;

wire  [7:0]  net1402;

wire  [47:0]  net981;

wire  [7:0]  net1332;

wire  [47:0]  net1398;

wire  [47:0]  net1289;

wire  [47:0]  net809;

wire  [47:0]  net1241;

wire  [7:0]  net1453;

wire  [7:0]  net767;

wire  [23:0]  net720;

wire  [47:0]  net1239;

wire  [7:0]  net929;

wire  [7:0]  net1022;

wire  [7:0]  net771;

wire  [47:0]  net792;

wire  [23:0]  net854;

wire  [47:0]  net1291;

wire  [7:0]  net1272;

wire  [7:0]  net768;

wire  [47:0]  net1171;

wire  [47:0]  net1053;

wire  [47:0]  net1149;

wire  [47:0]  net1449;

wire  [47:0]  net1004;

wire  [47:0]  net1056;

wire  [7:0]  net818;

wire  [23:0]  net849;

wire  [47:0]  net1443;

wire  [23:0]  net1095;

wire  [47:0]  net1448;

wire  [47:0]  net1054;

wire  [7:0]  net1216;

wire  [23:0]  net1235;

wire  [47:0]  net1266;

wire  [47:0]  net829;

wire  [7:0]  net1213;

wire  [47:0]  net1444;

wire  [7:0]  net1084;



bram1x4_ice1f I_bram_col_t03 ( .prog(prog),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .reset_b(reset_b_l[127:0]), .bm_wdummymux_en_o(net1440),
     .bm_sreb_o(net1436), .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(net694),
     .bm_sa_o({net695[0], net695[1], net695[2], net695[3], net695[4],
     net695[5], net695[6], net695[7]}), .bm_rcapmux_en_o(net1435),
     .bm_init_o(net697), .lft_op_05({net990[0], net990[1], net990[2],
     net990[3], net990[4], net990[5], net990[6], net990[7]}),
     .bl(bl[167:126]), .sp4_h_l_06({net1076[0], net1076[1], net1076[2],
     net1076[3], net1076[4], net1076[5], net1076[6], net1076[7],
     net1076[8], net1076[9], net1076[10], net1076[11], net1076[12],
     net1076[13], net1076[14], net1076[15], net1076[16], net1076[17],
     net1076[18], net1076[19], net1076[20], net1076[21], net1076[22],
     net1076[23], net1076[24], net1076[25], net1076[26], net1076[27],
     net1076[28], net1076[29], net1076[30], net1076[31], net1076[32],
     net1076[33], net1076[34], net1076[35], net1076[36], net1076[37],
     net1076[38], net1076[39], net1076[40], net1076[41], net1076[42],
     net1076[43], net1076[44], net1076[45], net1076[46], net1076[47]}),
     .sp12_h_l_02({net1045[0], net1045[1], net1045[2], net1045[3],
     net1045[4], net1045[5], net1045[6], net1045[7], net1045[8],
     net1045[9], net1045[10], net1045[11], net1045[12], net1045[13],
     net1045[14], net1045[15], net1045[16], net1045[17], net1045[18],
     net1045[19], net1045[20], net1045[21], net1045[22], net1045[23]}),
     .lft_op_06({net989[0], net989[1], net989[2], net989[3], net989[4],
     net989[5], net989[6], net989[7]}), .sp12_h_l_03({net1044[0],
     net1044[1], net1044[2], net1044[3], net1044[4], net1044[5],
     net1044[6], net1044[7], net1044[8], net1044[9], net1044[10],
     net1044[11], net1044[12], net1044[13], net1044[14], net1044[15],
     net1044[16], net1044[17], net1044[18], net1044[19], net1044[20],
     net1044[21], net1044[22], net1044[23]}), .sp12_h_r_03({net704[0],
     net704[1], net704[2], net704[3], net704[4], net704[5], net704[6],
     net704[7], net704[8], net704[9], net704[10], net704[11],
     net704[12], net704[13], net704[14], net704[15], net704[16],
     net704[17], net704[18], net704[19], net704[20], net704[21],
     net704[22], net704[23]}), .sp12_h_l_01({net1046[0], net1046[1],
     net1046[2], net1046[3], net1046[4], net1046[5], net1046[6],
     net1046[7], net1046[8], net1046[9], net1046[10], net1046[11],
     net1046[12], net1046[13], net1046[14], net1046[15], net1046[16],
     net1046[17], net1046[18], net1046[19], net1046[20], net1046[21],
     net1046[22], net1046[23]}), .sp4_v_b_04({net1049[0], net1049[1],
     net1049[2], net1049[3], net1049[4], net1049[5], net1049[6],
     net1049[7], net1049[8], net1049[9], net1049[10], net1049[11],
     net1049[12], net1049[13], net1049[14], net1049[15], net1049[16],
     net1049[17], net1049[18], net1049[19], net1049[20], net1049[21],
     net1049[22], net1049[23], net1049[24], net1049[25], net1049[26],
     net1049[27], net1049[28], net1049[29], net1049[30], net1049[31],
     net1049[32], net1049[33], net1049[34], net1049[35], net1049[36],
     net1049[37], net1049[38], net1049[39], net1049[40], net1049[41],
     net1049[42], net1049[43], net1049[44], net1049[45], net1049[46],
     net1049[47]}), .sp4_v_b_05({net1098[0], net1098[1], net1098[2],
     net1098[3], net1098[4], net1098[5], net1098[6], net1098[7],
     net1098[8], net1098[9], net1098[10], net1098[11], net1098[12],
     net1098[13], net1098[14], net1098[15], net1098[16], net1098[17],
     net1098[18], net1098[19], net1098[20], net1098[21], net1098[22],
     net1098[23], net1098[24], net1098[25], net1098[26], net1098[27],
     net1098[28], net1098[29], net1098[30], net1098[31], net1098[32],
     net1098[33], net1098[34], net1098[35], net1098[36], net1098[37],
     net1098[38], net1098[39], net1098[40], net1098[41], net1098[42],
     net1098[43], net1098[44], net1098[45], net1098[46], net1098[47]}),
     .lft_op_07({net988[0], net988[1], net988[2], net988[3], net988[4],
     net988[5], net988[6], net988[7]}), .sp4_v_b_06({net1099[0],
     net1099[1], net1099[2], net1099[3], net1099[4], net1099[5],
     net1099[6], net1099[7], net1099[8], net1099[9], net1099[10],
     net1099[11], net1099[12], net1099[13], net1099[14], net1099[15],
     net1099[16], net1099[17], net1099[18], net1099[19], net1099[20],
     net1099[21], net1099[22], net1099[23], net1099[24], net1099[25],
     net1099[26], net1099[27], net1099[28], net1099[29], net1099[30],
     net1099[31], net1099[32], net1099[33], net1099[34], net1099[35],
     net1099[36], net1099[37], net1099[38], net1099[39], net1099[40],
     net1099[41], net1099[42], net1099[43], net1099[44], net1099[45],
     net1099[46], net1099[47]}), .sp4_v_b_08({net1101[0], net1101[1],
     net1101[2], net1101[3], net1101[4], net1101[5], net1101[6],
     net1101[7], net1101[8], net1101[9], net1101[10], net1101[11],
     net1101[12], net1101[13], net1101[14], net1101[15], net1101[16],
     net1101[17], net1101[18], net1101[19], net1101[20], net1101[21],
     net1101[22], net1101[23], net1101[24], net1101[25], net1101[26],
     net1101[27], net1101[28], net1101[29], net1101[30], net1101[31],
     net1101[32], net1101[33], net1101[34], net1101[35], net1101[36],
     net1101[37], net1101[38], net1101[39], net1101[40], net1101[41],
     net1101[42], net1101[43], net1101[44], net1101[45], net1101[46],
     net1101[47]}), .sp4_v_b_07({net1100[0], net1100[1], net1100[2],
     net1100[3], net1100[4], net1100[5], net1100[6], net1100[7],
     net1100[8], net1100[9], net1100[10], net1100[11], net1100[12],
     net1100[13], net1100[14], net1100[15], net1100[16], net1100[17],
     net1100[18], net1100[19], net1100[20], net1100[21], net1100[22],
     net1100[23], net1100[24], net1100[25], net1100[26], net1100[27],
     net1100[28], net1100[29], net1100[30], net1100[31], net1100[32],
     net1100[33], net1100[34], net1100[35], net1100[36], net1100[37],
     net1100[38], net1100[39], net1100[40], net1100[41], net1100[42],
     net1100[43], net1100[44], net1100[45], net1100[46], net1100[47]}),
     .lft_op_03({net929[0], net929[1], net929[2], net929[3], net929[4],
     net929[5], net929[6], net929[7]}), .lft_op_01(slf_op_02_09[7:0]),
     .sp4_h_l_02({net1055[0], net1055[1], net1055[2], net1055[3],
     net1055[4], net1055[5], net1055[6], net1055[7], net1055[8],
     net1055[9], net1055[10], net1055[11], net1055[12], net1055[13],
     net1055[14], net1055[15], net1055[16], net1055[17], net1055[18],
     net1055[19], net1055[20], net1055[21], net1055[22], net1055[23],
     net1055[24], net1055[25], net1055[26], net1055[27], net1055[28],
     net1055[29], net1055[30], net1055[31], net1055[32], net1055[33],
     net1055[34], net1055[35], net1055[36], net1055[37], net1055[38],
     net1055[39], net1055[40], net1055[41], net1055[42], net1055[43],
     net1055[44], net1055[45], net1055[46], net1055[47]}),
     .sp12_h_l_06({net1094[0], net1094[1], net1094[2], net1094[3],
     net1094[4], net1094[5], net1094[6], net1094[7], net1094[8],
     net1094[9], net1094[10], net1094[11], net1094[12], net1094[13],
     net1094[14], net1094[15], net1094[16], net1094[17], net1094[18],
     net1094[19], net1094[20], net1094[21], net1094[22], net1094[23]}),
     .sp12_h_r_07({net716[0], net716[1], net716[2], net716[3],
     net716[4], net716[5], net716[6], net716[7], net716[8], net716[9],
     net716[10], net716[11], net716[12], net716[13], net716[14],
     net716[15], net716[16], net716[17], net716[18], net716[19],
     net716[20], net716[21], net716[22], net716[23]}),
     .sp12_h_l_05({net1093[0], net1093[1], net1093[2], net1093[3],
     net1093[4], net1093[5], net1093[6], net1093[7], net1093[8],
     net1093[9], net1093[10], net1093[11], net1093[12], net1093[13],
     net1093[14], net1093[15], net1093[16], net1093[17], net1093[18],
     net1093[19], net1093[20], net1093[21], net1093[22], net1093[23]}),
     .sp12_h_r_06({net718[0], net718[1], net718[2], net718[3],
     net718[4], net718[5], net718[6], net718[7], net718[8], net718[9],
     net718[10], net718[11], net718[12], net718[13], net718[14],
     net718[15], net718[16], net718[17], net718[18], net718[19],
     net718[20], net718[21], net718[22], net718[23]}),
     .sp12_h_l_04({net1043[0], net1043[1], net1043[2], net1043[3],
     net1043[4], net1043[5], net1043[6], net1043[7], net1043[8],
     net1043[9], net1043[10], net1043[11], net1043[12], net1043[13],
     net1043[14], net1043[15], net1043[16], net1043[17], net1043[18],
     net1043[19], net1043[20], net1043[21], net1043[22], net1043[23]}),
     .sp12_h_r_05({net720[0], net720[1], net720[2], net720[3],
     net720[4], net720[5], net720[6], net720[7], net720[8], net720[9],
     net720[10], net720[11], net720[12], net720[13], net720[14],
     net720[15], net720[16], net720[17], net720[18], net720[19],
     net720[20], net720[21], net720[22], net720[23]}),
     .sp12_h_r_08({net721[0], net721[1], net721[2], net721[3],
     net721[4], net721[5], net721[6], net721[7], net721[8], net721[9],
     net721[10], net721[11], net721[12], net721[13], net721[14],
     net721[15], net721[16], net721[17], net721[18], net721[19],
     net721[20], net721[21], net721[22], net721[23]}),
     .sp12_h_l_07({net1095[0], net1095[1], net1095[2], net1095[3],
     net1095[4], net1095[5], net1095[6], net1095[7], net1095[8],
     net1095[9], net1095[10], net1095[11], net1095[12], net1095[13],
     net1095[14], net1095[15], net1095[16], net1095[17], net1095[18],
     net1095[19], net1095[20], net1095[21], net1095[22], net1095[23]}),
     .sp12_h_l_08({net1096[0], net1096[1], net1096[2], net1096[3],
     net1096[4], net1096[5], net1096[6], net1096[7], net1096[8],
     net1096[9], net1096[10], net1096[11], net1096[12], net1096[13],
     net1096[14], net1096[15], net1096[16], net1096[17], net1096[18],
     net1096[19], net1096[20], net1096[21], net1096[22], net1096[23]}),
     .sp4_r_v_b_03({net724[0], net724[1], net724[2], net724[3],
     net724[4], net724[5], net724[6], net724[7], net724[8], net724[9],
     net724[10], net724[11], net724[12], net724[13], net724[14],
     net724[15], net724[16], net724[17], net724[18], net724[19],
     net724[20], net724[21], net724[22], net724[23], net724[24],
     net724[25], net724[26], net724[27], net724[28], net724[29],
     net724[30], net724[31], net724[32], net724[33], net724[34],
     net724[35], net724[36], net724[37], net724[38], net724[39],
     net724[40], net724[41], net724[42], net724[43], net724[44],
     net724[45], net724[46], net724[47]}),
     .vdd_cntl(vdd_cntl_l[127:0]), .pgate(pgate_l[127:0]),
     .bot_op_01(bot_op_03_09[7:0]), .sp4_r_v_b_04({net728[0],
     net728[1], net728[2], net728[3], net728[4], net728[5], net728[6],
     net728[7], net728[8], net728[9], net728[10], net728[11],
     net728[12], net728[13], net728[14], net728[15], net728[16],
     net728[17], net728[18], net728[19], net728[20], net728[21],
     net728[22], net728[23], net728[24], net728[25], net728[26],
     net728[27], net728[28], net728[29], net728[30], net728[31],
     net728[32], net728[33], net728[34], net728[35], net728[36],
     net728[37], net728[38], net728[39], net728[40], net728[41],
     net728[42], net728[43], net728[44], net728[45], net728[46],
     net728[47]}), .sp4_v_b_01(sp4_v_b_03_09[47:0]),
     .sp4_v_b_03({net1050[0], net1050[1], net1050[2], net1050[3],
     net1050[4], net1050[5], net1050[6], net1050[7], net1050[8],
     net1050[9], net1050[10], net1050[11], net1050[12], net1050[13],
     net1050[14], net1050[15], net1050[16], net1050[17], net1050[18],
     net1050[19], net1050[20], net1050[21], net1050[22], net1050[23],
     net1050[24], net1050[25], net1050[26], net1050[27], net1050[28],
     net1050[29], net1050[30], net1050[31], net1050[32], net1050[33],
     net1050[34], net1050[35], net1050[36], net1050[37], net1050[38],
     net1050[39], net1050[40], net1050[41], net1050[42], net1050[43],
     net1050[44], net1050[45], net1050[46], net1050[47]}),
     .sp4_h_r_08({net731[0], net731[1], net731[2], net731[3],
     net731[4], net731[5], net731[6], net731[7], net731[8], net731[9],
     net731[10], net731[11], net731[12], net731[13], net731[14],
     net731[15], net731[16], net731[17], net731[18], net731[19],
     net731[20], net731[21], net731[22], net731[23], net731[24],
     net731[25], net731[26], net731[27], net731[28], net731[29],
     net731[30], net731[31], net731[32], net731[33], net731[34],
     net731[35], net731[36], net731[37], net731[38], net731[39],
     net731[40], net731[41], net731[42], net731[43], net731[44],
     net731[45], net731[46], net731[47]}), .sp4_r_v_b_05({net732[0],
     net732[1], net732[2], net732[3], net732[4], net732[5], net732[6],
     net732[7], net732[8], net732[9], net732[10], net732[11],
     net732[12], net732[13], net732[14], net732[15], net732[16],
     net732[17], net732[18], net732[19], net732[20], net732[21],
     net732[22], net732[23], net732[24], net732[25], net732[26],
     net732[27], net732[28], net732[29], net732[30], net732[31],
     net732[32], net732[33], net732[34], net732[35], net732[36],
     net732[37], net732[38], net732[39], net732[40], net732[41],
     net732[42], net732[43], net732[44], net732[45], net732[46],
     net732[47]}), .sp4_v_b_02({net1051[0], net1051[1], net1051[2],
     net1051[3], net1051[4], net1051[5], net1051[6], net1051[7],
     net1051[8], net1051[9], net1051[10], net1051[11], net1051[12],
     net1051[13], net1051[14], net1051[15], net1051[16], net1051[17],
     net1051[18], net1051[19], net1051[20], net1051[21], net1051[22],
     net1051[23], net1051[24], net1051[25], net1051[26], net1051[27],
     net1051[28], net1051[29], net1051[30], net1051[31], net1051[32],
     net1051[33], net1051[34], net1051[35], net1051[36], net1051[37],
     net1051[38], net1051[39], net1051[40], net1051[41], net1051[42],
     net1051[43], net1051[44], net1051[45], net1051[46], net1051[47]}),
     .sp4_v_t_08({net734[0], net734[1], net734[2], net734[3],
     net734[4], net734[5], net734[6], net734[7], net734[8], net734[9],
     net734[10], net734[11], net734[12], net734[13], net734[14],
     net734[15], net734[16], net734[17], net734[18], net734[19],
     net734[20], net734[21], net734[22], net734[23], net734[24],
     net734[25], net734[26], net734[27], net734[28], net734[29],
     net734[30], net734[31], net734[32], net734[33], net734[34],
     net734[35], net734[36], net734[37], net734[38], net734[39],
     net734[40], net734[41], net734[42], net734[43], net734[44],
     net734[45], net734[46], net734[47]}), .sp4_r_v_b_02({net735[0],
     net735[1], net735[2], net735[3], net735[4], net735[5], net735[6],
     net735[7], net735[8], net735[9], net735[10], net735[11],
     net735[12], net735[13], net735[14], net735[15], net735[16],
     net735[17], net735[18], net735[19], net735[20], net735[21],
     net735[22], net735[23], net735[24], net735[25], net735[26],
     net735[27], net735[28], net735[29], net735[30], net735[31],
     net735[32], net735[33], net735[34], net735[35], net735[36],
     net735[37], net735[38], net735[39], net735[40], net735[41],
     net735[42], net735[43], net735[44], net735[45], net735[46],
     net735[47]}), .bnr_op_01(bnr_op_03_09[7:0]),
     .bm_sdi_o(bm_sdi_b1_o[1:0]), .sp4_h_l_04({net1053[0], net1053[1],
     net1053[2], net1053[3], net1053[4], net1053[5], net1053[6],
     net1053[7], net1053[8], net1053[9], net1053[10], net1053[11],
     net1053[12], net1053[13], net1053[14], net1053[15], net1053[16],
     net1053[17], net1053[18], net1053[19], net1053[20], net1053[21],
     net1053[22], net1053[23], net1053[24], net1053[25], net1053[26],
     net1053[27], net1053[28], net1053[29], net1053[30], net1053[31],
     net1053[32], net1053[33], net1053[34], net1053[35], net1053[36],
     net1053[37], net1053[38], net1053[39], net1053[40], net1053[41],
     net1053[42], net1053[43], net1053[44], net1053[45], net1053[46],
     net1053[47]}), .lft_op_08({net987[0], net987[1], net987[2],
     net987[3], net987[4], net987[5], net987[6], net987[7]}),
     .sp12_h_r_01({net740[0], net740[1], net740[2], net740[3],
     net740[4], net740[5], net740[6], net740[7], net740[8], net740[9],
     net740[10], net740[11], net740[12], net740[13], net740[14],
     net740[15], net740[16], net740[17], net740[18], net740[19],
     net740[20], net740[21], net740[22], net740[23]}),
     .bm_sdo_i({tiegnd_bram_t, bm_sdi_b1_o[0]}),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sweb_o({net1441[0], net1441[1]}),
     .sp4_h_l_03({net1054[0], net1054[1], net1054[2], net1054[3],
     net1054[4], net1054[5], net1054[6], net1054[7], net1054[8],
     net1054[9], net1054[10], net1054[11], net1054[12], net1054[13],
     net1054[14], net1054[15], net1054[16], net1054[17], net1054[18],
     net1054[19], net1054[20], net1054[21], net1054[22], net1054[23],
     net1054[24], net1054[25], net1054[26], net1054[27], net1054[28],
     net1054[29], net1054[30], net1054[31], net1054[32], net1054[33],
     net1054[34], net1054[35], net1054[36], net1054[37], net1054[38],
     net1054[39], net1054[40], net1054[41], net1054[42], net1054[43],
     net1054[44], net1054[45], net1054[46], net1054[47]}),
     .sp4_h_l_01({net1056[0], net1056[1], net1056[2], net1056[3],
     net1056[4], net1056[5], net1056[6], net1056[7], net1056[8],
     net1056[9], net1056[10], net1056[11], net1056[12], net1056[13],
     net1056[14], net1056[15], net1056[16], net1056[17], net1056[18],
     net1056[19], net1056[20], net1056[21], net1056[22], net1056[23],
     net1056[24], net1056[25], net1056[26], net1056[27], net1056[28],
     net1056[29], net1056[30], net1056[31], net1056[32], net1056[33],
     net1056[34], net1056[35], net1056[36], net1056[37], net1056[38],
     net1056[39], net1056[40], net1056[41], net1056[42], net1056[43],
     net1056[44], net1056[45], net1056[46], net1056[47]}),
     .sp4_h_r_01({net746[0], net746[1], net746[2], net746[3],
     net746[4], net746[5], net746[6], net746[7], net746[8], net746[9],
     net746[10], net746[11], net746[12], net746[13], net746[14],
     net746[15], net746[16], net746[17], net746[18], net746[19],
     net746[20], net746[21], net746[22], net746[23], net746[24],
     net746[25], net746[26], net746[27], net746[28], net746[29],
     net746[30], net746[31], net746[32], net746[33], net746[34],
     net746[35], net746[36], net746[37], net746[38], net746[39],
     net746[40], net746[41], net746[42], net746[43], net746[44],
     net746[45], net746[46], net746[47]}), .tnr_op_08({slf_op_04_17[3],
     slf_op_04_17[2], slf_op_04_17[1], slf_op_04_17[0],
     slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0]}), .sp12_h_r_02({net748[0], net748[1], net748[2],
     net748[3], net748[4], net748[5], net748[6], net748[7], net748[8],
     net748[9], net748[10], net748[11], net748[12], net748[13],
     net748[14], net748[15], net748[16], net748[17], net748[18],
     net748[19], net748[20], net748[21], net748[22], net748[23]}),
     .sp12_h_r_04({net749[0], net749[1], net749[2], net749[3],
     net749[4], net749[5], net749[6], net749[7], net749[8], net749[9],
     net749[10], net749[11], net749[12], net749[13], net749[14],
     net749[15], net749[16], net749[17], net749[18], net749[19],
     net749[20], net749[21], net749[22], net749[23]}),
     .bm_sclkrw_o({net1439[0], net1439[1]}),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .lft_op_02({net931[0], net931[1],
     net931[2], net931[3], net931[4], net931[5], net931[6],
     net931[7]}), .lft_op_04({net939[0], net939[1], net939[2],
     net939[3], net939[4], net939[5], net939[6], net939[7]}),
     .bm_sweb_i(bm_sweb_i[1:0]), .bnl_op_01(bnl_op_03_09[7:0]),
     .sp12_v_t_08({net756[0], net756[1], net756[2], net756[3],
     net756[4], net756[5], net756[6], net756[7], net756[8], net756[9],
     net756[10], net756[11], net756[12], net756[13], net756[14],
     net756[15], net756[16], net756[17], net756[18], net756[19],
     net756[20], net756[21], net756[22], net756[23]}),
     .wl(wl_l[127:0]), .tnl_op_08({slf_op_02_17[3], slf_op_02_17[2],
     slf_op_02_17[1], slf_op_02_17[0], slf_op_02_17[3],
     slf_op_02_17[2], slf_op_02_17[1], slf_op_02_17[0]}),
     .top_op_08({slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0], slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0]}), .bm_ab_2bot(bm_ab_2bot[10:0]),
     .bm_aa_2bot(bm_aa_2bot[10:0]), .sp12_v_b_01(sp12_v_b_03_09[23:0]),
     .sp4_r_v_b_08({net763[0], net763[1], net763[2], net763[3],
     net763[4], net763[5], net763[6], net763[7], net763[8], net763[9],
     net763[10], net763[11], net763[12], net763[13], net763[14],
     net763[15], net763[16], net763[17], net763[18], net763[19],
     net763[20], net763[21], net763[22], net763[23], net763[24],
     net763[25], net763[26], net763[27], net763[28], net763[29],
     net763[30], net763[31], net763[32], net763[33], net763[34],
     net763[35], net763[36], net763[37], net763[38], net763[39],
     net763[40], net763[41], net763[42], net763[43], net763[44],
     net763[45], net763[46], net763[47]}), .sp4_r_v_b_07({net764[0],
     net764[1], net764[2], net764[3], net764[4], net764[5], net764[6],
     net764[7], net764[8], net764[9], net764[10], net764[11],
     net764[12], net764[13], net764[14], net764[15], net764[16],
     net764[17], net764[18], net764[19], net764[20], net764[21],
     net764[22], net764[23], net764[24], net764[25], net764[26],
     net764[27], net764[28], net764[29], net764[30], net764[31],
     net764[32], net764[33], net764[34], net764[35], net764[36],
     net764[37], net764[38], net764[39], net764[40], net764[41],
     net764[42], net764[43], net764[44], net764[45], net764[46],
     net764[47]}), .sp4_r_v_b_06({net765[0], net765[1], net765[2],
     net765[3], net765[4], net765[5], net765[6], net765[7], net765[8],
     net765[9], net765[10], net765[11], net765[12], net765[13],
     net765[14], net765[15], net765[16], net765[17], net765[18],
     net765[19], net765[20], net765[21], net765[22], net765[23],
     net765[24], net765[25], net765[26], net765[27], net765[28],
     net765[29], net765[30], net765[31], net765[32], net765[33],
     net765[34], net765[35], net765[36], net765[37], net765[38],
     net765[39], net765[40], net765[41], net765[42], net765[43],
     net765[44], net765[45], net765[46], net765[47]}),
     .sp4_r_v_b_01(sp4_v_b_04_09[47:0]), .rgt_op_08({net767[0],
     net767[1], net767[2], net767[3], net767[4], net767[5], net767[6],
     net767[7]}), .rgt_op_07({net768[0], net768[1], net768[2],
     net768[3], net768[4], net768[5], net768[6], net768[7]}),
     .rgt_op_06({net769[0], net769[1], net769[2], net769[3], net769[4],
     net769[5], net769[6], net769[7]}), .rgt_op_05({net770[0],
     net770[1], net770[2], net770[3], net770[4], net770[5], net770[6],
     net770[7]}), .rgt_op_04({net771[0], net771[1], net771[2],
     net771[3], net771[4], net771[5], net771[6], net771[7]}),
     .rgt_op_03({net772[0], net772[1], net772[2], net772[3], net772[4],
     net772[5], net772[6], net772[7]}), .rgt_op_02({net773[0],
     net773[1], net773[2], net773[3], net773[4], net773[5], net773[6],
     net773[7]}), .rgt_op_01(slf_op_04_09[7:0]),
     .slf_op_02({net1026[0], net1026[1], net1026[2], net1026[3],
     net1026[4], net1026[5], net1026[6], net1026[7]}),
     .slf_op_01(slf_op_03_09[7:0]), .slf_op_03({net1024[0], net1024[1],
     net1024[2], net1024[3], net1024[4], net1024[5], net1024[6],
     net1024[7]}), .slf_op_04({net1034[0], net1034[1], net1034[2],
     net1034[3], net1034[4], net1034[5], net1034[6], net1034[7]}),
     .slf_op_05({net1085[0], net1085[1], net1085[2], net1085[3],
     net1085[4], net1085[5], net1085[6], net1085[7]}),
     .slf_op_06({net1084[0], net1084[1], net1084[2], net1084[3],
     net1084[4], net1084[5], net1084[6], net1084[7]}),
     .slf_op_07({net1083[0], net1083[1], net1083[2], net1083[3],
     net1083[4], net1083[5], net1083[6], net1083[7]}),
     .slf_op_08({net1082[0], net1082[1], net1082[2], net1082[3],
     net1082[4], net1082[5], net1082[6], net1082[7]}),
     .bm_ab_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .bm_aa_top({tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t,
     tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t, tiegnd_bram_t}),
     .glb_netwk_bot({net1453[0], net1453[1], net1453[2], net1453[3],
     net1453[4], net1453[5], net1453[6], net1453[7]}),
     .glb_netwk_top({net786[0], net786[1], net786[2], net786[3],
     net786[4], net786[5], net786[6], net786[7]}),
     .sp4_h_l_08({net1074[0], net1074[1], net1074[2], net1074[3],
     net1074[4], net1074[5], net1074[6], net1074[7], net1074[8],
     net1074[9], net1074[10], net1074[11], net1074[12], net1074[13],
     net1074[14], net1074[15], net1074[16], net1074[17], net1074[18],
     net1074[19], net1074[20], net1074[21], net1074[22], net1074[23],
     net1074[24], net1074[25], net1074[26], net1074[27], net1074[28],
     net1074[29], net1074[30], net1074[31], net1074[32], net1074[33],
     net1074[34], net1074[35], net1074[36], net1074[37], net1074[38],
     net1074[39], net1074[40], net1074[41], net1074[42], net1074[43],
     net1074[44], net1074[45], net1074[46], net1074[47]}),
     .sp4_h_l_07({net1075[0], net1075[1], net1075[2], net1075[3],
     net1075[4], net1075[5], net1075[6], net1075[7], net1075[8],
     net1075[9], net1075[10], net1075[11], net1075[12], net1075[13],
     net1075[14], net1075[15], net1075[16], net1075[17], net1075[18],
     net1075[19], net1075[20], net1075[21], net1075[22], net1075[23],
     net1075[24], net1075[25], net1075[26], net1075[27], net1075[28],
     net1075[29], net1075[30], net1075[31], net1075[32], net1075[33],
     net1075[34], net1075[35], net1075[36], net1075[37], net1075[38],
     net1075[39], net1075[40], net1075[41], net1075[42], net1075[43],
     net1075[44], net1075[45], net1075[46], net1075[47]}),
     .sp4_h_l_05({net1077[0], net1077[1], net1077[2], net1077[3],
     net1077[4], net1077[5], net1077[6], net1077[7], net1077[8],
     net1077[9], net1077[10], net1077[11], net1077[12], net1077[13],
     net1077[14], net1077[15], net1077[16], net1077[17], net1077[18],
     net1077[19], net1077[20], net1077[21], net1077[22], net1077[23],
     net1077[24], net1077[25], net1077[26], net1077[27], net1077[28],
     net1077[29], net1077[30], net1077[31], net1077[32], net1077[33],
     net1077[34], net1077[35], net1077[36], net1077[37], net1077[38],
     net1077[39], net1077[40], net1077[41], net1077[42], net1077[43],
     net1077[44], net1077[45], net1077[46], net1077[47]}),
     .sp4_h_r_02({net790[0], net790[1], net790[2], net790[3],
     net790[4], net790[5], net790[6], net790[7], net790[8], net790[9],
     net790[10], net790[11], net790[12], net790[13], net790[14],
     net790[15], net790[16], net790[17], net790[18], net790[19],
     net790[20], net790[21], net790[22], net790[23], net790[24],
     net790[25], net790[26], net790[27], net790[28], net790[29],
     net790[30], net790[31], net790[32], net790[33], net790[34],
     net790[35], net790[36], net790[37], net790[38], net790[39],
     net790[40], net790[41], net790[42], net790[43], net790[44],
     net790[45], net790[46], net790[47]}), .sp4_h_r_03({net791[0],
     net791[1], net791[2], net791[3], net791[4], net791[5], net791[6],
     net791[7], net791[8], net791[9], net791[10], net791[11],
     net791[12], net791[13], net791[14], net791[15], net791[16],
     net791[17], net791[18], net791[19], net791[20], net791[21],
     net791[22], net791[23], net791[24], net791[25], net791[26],
     net791[27], net791[28], net791[29], net791[30], net791[31],
     net791[32], net791[33], net791[34], net791[35], net791[36],
     net791[37], net791[38], net791[39], net791[40], net791[41],
     net791[42], net791[43], net791[44], net791[45], net791[46],
     net791[47]}), .sp4_h_r_04({net792[0], net792[1], net792[2],
     net792[3], net792[4], net792[5], net792[6], net792[7], net792[8],
     net792[9], net792[10], net792[11], net792[12], net792[13],
     net792[14], net792[15], net792[16], net792[17], net792[18],
     net792[19], net792[20], net792[21], net792[22], net792[23],
     net792[24], net792[25], net792[26], net792[27], net792[28],
     net792[29], net792[30], net792[31], net792[32], net792[33],
     net792[34], net792[35], net792[36], net792[37], net792[38],
     net792[39], net792[40], net792[41], net792[42], net792[43],
     net792[44], net792[45], net792[46], net792[47]}),
     .sp4_h_r_05({net793[0], net793[1], net793[2], net793[3],
     net793[4], net793[5], net793[6], net793[7], net793[8], net793[9],
     net793[10], net793[11], net793[12], net793[13], net793[14],
     net793[15], net793[16], net793[17], net793[18], net793[19],
     net793[20], net793[21], net793[22], net793[23], net793[24],
     net793[25], net793[26], net793[27], net793[28], net793[29],
     net793[30], net793[31], net793[32], net793[33], net793[34],
     net793[35], net793[36], net793[37], net793[38], net793[39],
     net793[40], net793[41], net793[42], net793[43], net793[44],
     net793[45], net793[46], net793[47]}), .sp4_h_r_06({net794[0],
     net794[1], net794[2], net794[3], net794[4], net794[5], net794[6],
     net794[7], net794[8], net794[9], net794[10], net794[11],
     net794[12], net794[13], net794[14], net794[15], net794[16],
     net794[17], net794[18], net794[19], net794[20], net794[21],
     net794[22], net794[23], net794[24], net794[25], net794[26],
     net794[27], net794[28], net794[29], net794[30], net794[31],
     net794[32], net794[33], net794[34], net794[35], net794[36],
     net794[37], net794[38], net794[39], net794[40], net794[41],
     net794[42], net794[43], net794[44], net794[45], net794[46],
     net794[47]}), .sp4_h_r_07({net795[0], net795[1], net795[2],
     net795[3], net795[4], net795[5], net795[6], net795[7], net795[8],
     net795[9], net795[10], net795[11], net795[12], net795[13],
     net795[14], net795[15], net795[16], net795[17], net795[18],
     net795[19], net795[20], net795[21], net795[22], net795[23],
     net795[24], net795[25], net795[26], net795[27], net795[28],
     net795[29], net795[30], net795[31], net795[32], net795[33],
     net795[34], net795[35], net795[36], net795[37], net795[38],
     net795[39], net795[40], net795[41], net795[42], net795[43],
     net795[44], net795[45], net795[46], net795[47]}));
pinlatbuf12p I389 ( .pad_in(padin_t_l[11]), .icegate(hold_t_l),
     .cbit(cf_t[135]), .cout(net675), .prog(prog));
pinlatbuf12p I_pinlatbuf12p_l ( .pad_in(padin_l_t[12]),
     .icegate(hold_l_t), .cbit(cf_l[15]), .cout(net1427), .prog(prog));
io_lft_top_1x8_ice1f I_preio_lt_t00 ( .padin(padin_l_t[23:12]),
     .pado(pado_l_t[23:12]), .padeb(padeb_l_t[23:12]),
     .fo_dlyadj(fo_dlyadj[7:3]), .sp4_v_b_00_09(sp4_v_b_00_09[15:0]),
     .bnr_op_00_09(bnr_op_00_09[7:0]), .tnr_op_08({slf_op_01_17[3],
     slf_op_01_17[2], slf_op_01_17[1], slf_op_01_17[0],
     slf_op_01_17[3], slf_op_01_17[2], slf_op_01_17[1],
     slf_op_01_17[0]}), .shift(shift_o), .bs_en(bs_en_o),
     .mode(mode_o), .sdi(net803), .hiz_b(hiz_b_o), .prog(prog),
     .hold(hold_l_t), .update(update_o), .r(r_o),
     .SP4_h_l_05({net809[0], net809[1], net809[2], net809[3],
     net809[4], net809[5], net809[6], net809[7], net809[8], net809[9],
     net809[10], net809[11], net809[12], net809[13], net809[14],
     net809[15], net809[16], net809[17], net809[18], net809[19],
     net809[20], net809[21], net809[22], net809[23], net809[24],
     net809[25], net809[26], net809[27], net809[28], net809[29],
     net809[30], net809[31], net809[32], net809[33], net809[34],
     net809[35], net809[36], net809[37], net809[38], net809[39],
     net809[40], net809[41], net809[42], net809[43], net809[44],
     net809[45], net809[46], net809[47]}),
     .slf_op_05(slf_op_00_13[3:0]), .slf_op_01(slf_op_00_09[3:0]),
     .slf_op_06(slf_op_00_14[3:0]), .slf_op_02(slf_op_00_10[3:0]),
     .sdo(sdo), .bl({bl[0], bl[1], bl[2], bl[3], bl[4], bl[5], bl[6],
     bl[7], bl[8], bl[9], bl[10], bl[11], bl[12], bl[13], bl[14],
     bl[15], bl[16], bl[17]}), .tclk(net816),
     .reset_b(reset_b_l[127:0]), .rgt_op_02({net818[0], net818[1],
     net818[2], net818[3], net818[4], net818[5], net818[6],
     net818[7]}), .SP4_h_l_06({net819[0], net819[1], net819[2],
     net819[3], net819[4], net819[5], net819[6], net819[7], net819[8],
     net819[9], net819[10], net819[11], net819[12], net819[13],
     net819[14], net819[15], net819[16], net819[17], net819[18],
     net819[19], net819[20], net819[21], net819[22], net819[23],
     net819[24], net819[25], net819[26], net819[27], net819[28],
     net819[29], net819[30], net819[31], net819[32], net819[33],
     net819[34], net819[35], net819[36], net819[37], net819[38],
     net819[39], net819[40], net819[41], net819[42], net819[43],
     net819[44], net819[45], net819[46], net819[47]}),
     .sp4_v_t_08({net820[0], net820[1], net820[2], net820[3],
     net820[4], net820[5], net820[6], net820[7], net820[8], net820[9],
     net820[10], net820[11], net820[12], net820[13], net820[14],
     net820[15]}), .slf_op_04(slf_op_00_12[3:0]),
     .slf_op_03(slf_op_00_11[3:0]), .slf_op_07(slf_op_00_15[3:0]),
     .slf_op_08(slf_op_00_16[3:0]), .SP4_h_l_08({net825[0], net825[1],
     net825[2], net825[3], net825[4], net825[5], net825[6], net825[7],
     net825[8], net825[9], net825[10], net825[11], net825[12],
     net825[13], net825[14], net825[15], net825[16], net825[17],
     net825[18], net825[19], net825[20], net825[21], net825[22],
     net825[23], net825[24], net825[25], net825[26], net825[27],
     net825[28], net825[29], net825[30], net825[31], net825[32],
     net825[33], net825[34], net825[35], net825[36], net825[37],
     net825[38], net825[39], net825[40], net825[41], net825[42],
     net825[43], net825[44], net825[45], net825[46], net825[47]}),
     .SP4_h_l_07({net826[0], net826[1], net826[2], net826[3],
     net826[4], net826[5], net826[6], net826[7], net826[8], net826[9],
     net826[10], net826[11], net826[12], net826[13], net826[14],
     net826[15], net826[16], net826[17], net826[18], net826[19],
     net826[20], net826[21], net826[22], net826[23], net826[24],
     net826[25], net826[26], net826[27], net826[28], net826[29],
     net826[30], net826[31], net826[32], net826[33], net826[34],
     net826[35], net826[36], net826[37], net826[38], net826[39],
     net826[40], net826[41], net826[42], net826[43], net826[44],
     net826[45], net826[46], net826[47]}), .SP4_h_l_03({net827[0],
     net827[1], net827[2], net827[3], net827[4], net827[5], net827[6],
     net827[7], net827[8], net827[9], net827[10], net827[11],
     net827[12], net827[13], net827[14], net827[15], net827[16],
     net827[17], net827[18], net827[19], net827[20], net827[21],
     net827[22], net827[23], net827[24], net827[25], net827[26],
     net827[27], net827[28], net827[29], net827[30], net827[31],
     net827[32], net827[33], net827[34], net827[35], net827[36],
     net827[37], net827[38], net827[39], net827[40], net827[41],
     net827[42], net827[43], net827[44], net827[45], net827[46],
     net827[47]}), .SP4_h_l_04({net828[0], net828[1], net828[2],
     net828[3], net828[4], net828[5], net828[6], net828[7], net828[8],
     net828[9], net828[10], net828[11], net828[12], net828[13],
     net828[14], net828[15], net828[16], net828[17], net828[18],
     net828[19], net828[20], net828[21], net828[22], net828[23],
     net828[24], net828[25], net828[26], net828[27], net828[28],
     net828[29], net828[30], net828[31], net828[32], net828[33],
     net828[34], net828[35], net828[36], net828[37], net828[38],
     net828[39], net828[40], net828[41], net828[42], net828[43],
     net828[44], net828[45], net828[46], net828[47]}),
     .SP4_h_l_02({net829[0], net829[1], net829[2], net829[3],
     net829[4], net829[5], net829[6], net829[7], net829[8], net829[9],
     net829[10], net829[11], net829[12], net829[13], net829[14],
     net829[15], net829[16], net829[17], net829[18], net829[19],
     net829[20], net829[21], net829[22], net829[23], net829[24],
     net829[25], net829[26], net829[27], net829[28], net829[29],
     net829[30], net829[31], net829[32], net829[33], net829[34],
     net829[35], net829[36], net829[37], net829[38], net829[39],
     net829[40], net829[41], net829[42], net829[43], net829[44],
     net829[45], net829[46], net829[47]}), .SP4_h_l_01({net830[0],
     net830[1], net830[2], net830[3], net830[4], net830[5], net830[6],
     net830[7], net830[8], net830[9], net830[10], net830[11],
     net830[12], net830[13], net830[14], net830[15], net830[16],
     net830[17], net830[18], net830[19], net830[20], net830[21],
     net830[22], net830[23], net830[24], net830[25], net830[26],
     net830[27], net830[28], net830[29], net830[30], net830[31],
     net830[32], net830[33], net830[34], net830[35], net830[36],
     net830[37], net830[38], net830[39], net830[40], net830[41],
     net830[42], net830[43], net830[44], net830[45], net830[46],
     net830[47]}), .rgt_op_07({net831[0], net831[1], net831[2],
     net831[3], net831[4], net831[5], net831[6], net831[7]}),
     .rgt_op_06({net832[0], net832[1], net832[2], net832[3], net832[4],
     net832[5], net832[6], net832[7]}), .rgt_op_05({net833[0],
     net833[1], net833[2], net833[3], net833[4], net833[5], net833[6],
     net833[7]}), .rgt_op_03({net834[0], net834[1], net834[2],
     net834[3], net834[4], net834[5], net834[6], net834[7]}),
     .rgt_op_01(slf_op_01_09[7:0]), .rgt_op_08({net836[0], net836[1],
     net836[2], net836[3], net836[4], net836[5], net836[6],
     net836[7]}), .pgate(pgate_l[127:0]), .vdd_cntl(vdd_cntl_l[127:0]),
     .last_rsr(last_rsr[1]),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .cf_l(cf_l[191:0]), .wl(wl_l[127:0]), .tclk_o(tclk_o),
     .ceb(ceb_o), .fabric_out_09(net1423), .SP12_h_l_02({net849[0],
     net849[1], net849[2], net849[3], net849[4], net849[5], net849[6],
     net849[7], net849[8], net849[9], net849[10], net849[11],
     net849[12], net849[13], net849[14], net849[15], net849[16],
     net849[17], net849[18], net849[19], net849[20], net849[21],
     net849[22], net849[23]}), .SP12_h_l_04({net850[0], net850[1],
     net850[2], net850[3], net850[4], net850[5], net850[6], net850[7],
     net850[8], net850[9], net850[10], net850[11], net850[12],
     net850[13], net850[14], net850[15], net850[16], net850[17],
     net850[18], net850[19], net850[20], net850[21], net850[22],
     net850[23]}), .SP12_h_l_08({net851[0], net851[1], net851[2],
     net851[3], net851[4], net851[5], net851[6], net851[7], net851[8],
     net851[9], net851[10], net851[11], net851[12], net851[13],
     net851[14], net851[15], net851[16], net851[17], net851[18],
     net851[19], net851[20], net851[21], net851[22], net851[23]}),
     .SP12_h_l_06({net852[0], net852[1], net852[2], net852[3],
     net852[4], net852[5], net852[6], net852[7], net852[8], net852[9],
     net852[10], net852[11], net852[12], net852[13], net852[14],
     net852[15], net852[16], net852[17], net852[18], net852[19],
     net852[20], net852[21], net852[22], net852[23]}),
     .glb_netwk_col(clk_tree_drv_tl[7:0]), .SP12_h_l_05({net854[0],
     net854[1], net854[2], net854[3], net854[4], net854[5], net854[6],
     net854[7], net854[8], net854[9], net854[10], net854[11],
     net854[12], net854[13], net854[14], net854[15], net854[16],
     net854[17], net854[18], net854[19], net854[20], net854[21],
     net854[22], net854[23]}), .SP12_h_l_01({net855[0], net855[1],
     net855[2], net855[3], net855[4], net855[5], net855[6], net855[7],
     net855[8], net855[9], net855[10], net855[11], net855[12],
     net855[13], net855[14], net855[15], net855[16], net855[17],
     net855[18], net855[19], net855[20], net855[21], net855[22],
     net855[23]}), .SP12_h_l_03({net856[0], net856[1], net856[2],
     net856[3], net856[4], net856[5], net856[6], net856[7], net856[8],
     net856[9], net856[10], net856[11], net856[12], net856[13],
     net856[14], net856[15], net856[16], net856[17], net856[18],
     net856[19], net856[20], net856[21], net856[22], net856[23]}),
     .SP12_h_l_07({net857[0], net857[1], net857[2], net857[3],
     net857[4], net857[5], net857[6], net857[7], net857[8], net857[9],
     net857[10], net857[11], net857[12], net857[13], net857[14],
     net857[15], net857[16], net857[17], net857[18], net857[19],
     net857[20], net857[21], net857[22], net857[23]}),
     .rgt_op_04({net858[0], net858[1], net858[2], net858[3], net858[4],
     net858[5], net858[6], net858[7]}));
io_top_lft_1x6_ice1f I_preio_top_l ( .fabric_out_06_17(net859),
     .cf_top_l(cf_t[143:0]), .wl_l({wl_l[142], wl_l[143], wl_l[141],
     wl_l[140], wl_l[138], wl_l[139], wl_l[137], wl_l[136], wl_l[134],
     wl_l[135], wl_l[133], wl_l[132], wl_l[130], wl_l[131], wl_l[129],
     wl_l[128]}), .lft_op_01_17({net836[0], net836[1], net836[2],
     net836[3], net836[4], net836[5], net836[6], net836[7]}),
     .vdd_cntl_l({vdd_cntl_l[142], vdd_cntl_l[143], vdd_cntl_l[141],
     vdd_cntl_l[140], vdd_cntl_l[138], vdd_cntl_l[139],
     vdd_cntl_l[137], vdd_cntl_l[136], vdd_cntl_l[134],
     vdd_cntl_l[135], vdd_cntl_l[133], vdd_cntl_l[132],
     vdd_cntl_l[130], vdd_cntl_l[131], vdd_cntl_l[129],
     vdd_cntl_l[128]}), .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .reset_l({reset_b_l[142],
     reset_b_l[143], reset_b_l[141], reset_b_l[140], reset_b_l[138],
     reset_b_l[139], reset_b_l[137], reset_b_l[136], reset_b_l[134],
     reset_b_l[135], reset_b_l[133], reset_b_l[132], reset_b_l[130],
     reset_b_l[131], reset_b_l[129], reset_b_l[128]}), .r_i(r_i),
     .prog(prog), .pgate_l({pgate_l[142], pgate_l[143], pgate_l[141],
     pgate_l[140], pgate_l[138], pgate_l[139], pgate_l[137],
     pgate_l[136], pgate_l[134], pgate_l[135], pgate_l[133],
     pgate_l[132], pgate_l[130], pgate_l[131], pgate_l[129],
     pgate_l[128]}), .mode_i(mode_i), .hiz_b_i(hiz_b_i),
     .bs_en_i(bs_en_i), .update_o(net1405), .tclk_o(net1406),
     .shift_o(net1407), .sdo(net1408), .r_o(net1409), .mode_o(net1410),
     .hiz_b_o(net1411), .glb_net_06({net1402[0], net1402[1],
     net1402[2], net1402[3], net1402[4], net1402[5], net1402[6],
     net1402[7]}), .glb_net_05({net1212[0], net1212[1], net1212[2],
     net1212[3], net1212[4], net1212[5], net1212[6], net1212[7]}),
     .glb_net_04({net1307[0], net1307[1], net1307[2], net1307[3],
     net1307[4], net1307[5], net1307[6], net1307[7]}),
     .glb_net_03({net786[0], net786[1], net786[2], net786[3],
     net786[4], net786[5], net786[6], net786[7]}),
     .glb_net_02({net1117[0], net1117[1], net1117[2], net1117[3],
     net1117[4], net1117[5], net1117[6], net1117[7]}),
     .glb_net_01({net1022[0], net1022[1], net1022[2], net1022[3],
     net1022[4], net1022[5], net1022[6], net1022[7]}),
     .bs_en_o(net1413), .sp4_h_r_06_17(sp4_h_r_06_17[15:0]),
     .bl_06(bl[329:276]), .bl_05(bl[275:222]), .bl_04(bl[221:168]),
     .bl_02(bl[125:72]), .bl_01(bl[71:18]), .sp4_h_l_01_17({net820[0],
     net820[1], net820[2], net820[3], net820[4], net820[5], net820[6],
     net820[7], net820[8], net820[9], net820[10], net820[11],
     net820[12], net820[13], net820[14], net820[15]}),
     .bnl_op_01_17({slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0], slf_op_00_16[3], slf_op_00_16[2],
     slf_op_00_16[1], slf_op_00_16[0]}), .padin_t_l(padin_t_l[11:0]),
     .lft_op_03_17({net1082[0], net1082[1], net1082[2], net1082[3],
     net1082[4], net1082[5], net1082[6], net1082[7]}),
     .sp4_v_b_04_17({net1303[0], net1303[1], net1303[2], net1303[3],
     net1303[4], net1303[5], net1303[6], net1303[7], net1303[8],
     net1303[9], net1303[10], net1303[11], net1303[12], net1303[13],
     net1303[14], net1303[15], net1303[16], net1303[17], net1303[18],
     net1303[19], net1303[20], net1303[21], net1303[22], net1303[23],
     net1303[24], net1303[25], net1303[26], net1303[27], net1303[28],
     net1303[29], net1303[30], net1303[31], net1303[32], net1303[33],
     net1303[34], net1303[35], net1303[36], net1303[37], net1303[38],
     net1303[39], net1303[40], net1303[41], net1303[42], net1303[43],
     net1303[44], net1303[45], net1303[46], net1303[47]}),
     .lft_op_02_17({net987[0], net987[1], net987[2], net987[3],
     net987[4], net987[5], net987[6], net987[7]}),
     .lft_op_04_17({net767[0], net767[1], net767[2], net767[3],
     net767[4], net767[5], net767[6], net767[7]}),
     .sp4_v_b_06_17({net1398[0], net1398[1], net1398[2], net1398[3],
     net1398[4], net1398[5], net1398[6], net1398[7], net1398[8],
     net1398[9], net1398[10], net1398[11], net1398[12], net1398[13],
     net1398[14], net1398[15], net1398[16], net1398[17], net1398[18],
     net1398[19], net1398[20], net1398[21], net1398[22], net1398[23],
     net1398[24], net1398[25], net1398[26], net1398[27], net1398[28],
     net1398[29], net1398[30], net1398[31], net1398[32], net1398[33],
     net1398[34], net1398[35], net1398[36], net1398[37], net1398[38],
     net1398[39], net1398[40], net1398[41], net1398[42], net1398[43],
     net1398[44], net1398[45], net1398[46], net1398[47]}),
     .sp12_v_b_04_17({net1299[0], net1299[1], net1299[2], net1299[3],
     net1299[4], net1299[5], net1299[6], net1299[7], net1299[8],
     net1299[9], net1299[10], net1299[11], net1299[12], net1299[13],
     net1299[14], net1299[15], net1299[16], net1299[17], net1299[18],
     net1299[19], net1299[20], net1299[21], net1299[22], net1299[23]}),
     .sp4_v_b_02_17({net1113[0], net1113[1], net1113[2], net1113[3],
     net1113[4], net1113[5], net1113[6], net1113[7], net1113[8],
     net1113[9], net1113[10], net1113[11], net1113[12], net1113[13],
     net1113[14], net1113[15], net1113[16], net1113[17], net1113[18],
     net1113[19], net1113[20], net1113[21], net1113[22], net1113[23],
     net1113[24], net1113[25], net1113[26], net1113[27], net1113[28],
     net1113[29], net1113[30], net1113[31], net1113[32], net1113[33],
     net1113[34], net1113[35], net1113[36], net1113[37], net1113[38],
     net1113[39], net1113[40], net1113[41], net1113[42], net1113[43],
     net1113[44], net1113[45], net1113[46], net1113[47]}),
     .sp12_v_b_05_17({net1204[0], net1204[1], net1204[2], net1204[3],
     net1204[4], net1204[5], net1204[6], net1204[7], net1204[8],
     net1204[9], net1204[10], net1204[11], net1204[12], net1204[13],
     net1204[14], net1204[15], net1204[16], net1204[17], net1204[18],
     net1204[19], net1204[20], net1204[21], net1204[22], net1204[23]}),
     .lft_op_06_17(slf_op_06_16[7:0]),
     .slf_op_04_17(slf_op_04_17[3:0]), .sp4_v_b_05_17({net1208[0],
     net1208[1], net1208[2], net1208[3], net1208[4], net1208[5],
     net1208[6], net1208[7], net1208[8], net1208[9], net1208[10],
     net1208[11], net1208[12], net1208[13], net1208[14], net1208[15],
     net1208[16], net1208[17], net1208[18], net1208[19], net1208[20],
     net1208[21], net1208[22], net1208[23], net1208[24], net1208[25],
     net1208[26], net1208[27], net1208[28], net1208[29], net1208[30],
     net1208[31], net1208[32], net1208[33], net1208[34], net1208[35],
     net1208[36], net1208[37], net1208[38], net1208[39], net1208[40],
     net1208[41], net1208[42], net1208[43], net1208[44], net1208[45],
     net1208[46], net1208[47]}), .sp12_v_b_03_17({net756[0], net756[1],
     net756[2], net756[3], net756[4], net756[5], net756[6], net756[7],
     net756[8], net756[9], net756[10], net756[11], net756[12],
     net756[13], net756[14], net756[15], net756[16], net756[17],
     net756[18], net756[19], net756[20], net756[21], net756[22],
     net756[23]}), .slf_op_01_17(slf_op_01_17[3:0]),
     .sp4_v_b_01_17({net1018[0], net1018[1], net1018[2], net1018[3],
     net1018[4], net1018[5], net1018[6], net1018[7], net1018[8],
     net1018[9], net1018[10], net1018[11], net1018[12], net1018[13],
     net1018[14], net1018[15], net1018[16], net1018[17], net1018[18],
     net1018[19], net1018[20], net1018[21], net1018[22], net1018[23],
     net1018[24], net1018[25], net1018[26], net1018[27], net1018[28],
     net1018[29], net1018[30], net1018[31], net1018[32], net1018[33],
     net1018[34], net1018[35], net1018[36], net1018[37], net1018[38],
     net1018[39], net1018[40], net1018[41], net1018[42], net1018[43],
     net1018[44], net1018[45], net1018[46], net1018[47]}),
     .sp4_v_b_03_17({net734[0], net734[1], net734[2], net734[3],
     net734[4], net734[5], net734[6], net734[7], net734[8], net734[9],
     net734[10], net734[11], net734[12], net734[13], net734[14],
     net734[15], net734[16], net734[17], net734[18], net734[19],
     net734[20], net734[21], net734[22], net734[23], net734[24],
     net734[25], net734[26], net734[27], net734[28], net734[29],
     net734[30], net734[31], net734[32], net734[33], net734[34],
     net734[35], net734[36], net734[37], net734[38], net734[39],
     net734[40], net734[41], net734[42], net734[43], net734[44],
     net734[45], net734[46], net734[47]}),
     .slf_op_03_17(slf_op_08_17[3:0]), .lft_op_05_17({net1272[0],
     net1272[1], net1272[2], net1272[3], net1272[4], net1272[5],
     net1272[6], net1272[7]}), .bnr_op_06_17(rgt_op_06_16[7:0]),
     .sp12_v_b_01_17({net1014[0], net1014[1], net1014[2], net1014[3],
     net1014[4], net1014[5], net1014[6], net1014[7], net1014[8],
     net1014[9], net1014[10], net1014[11], net1014[12], net1014[13],
     net1014[14], net1014[15], net1014[16], net1014[17], net1014[18],
     net1014[19], net1014[20], net1014[21], net1014[22], net1014[23]}),
     .slf_op_06_17(slf_op_06_17[3:0]), .sp12_v_b_06_17({net1394[0],
     net1394[1], net1394[2], net1394[3], net1394[4], net1394[5],
     net1394[6], net1394[7], net1394[8], net1394[9], net1394[10],
     net1394[11], net1394[12], net1394[13], net1394[14], net1394[15],
     net1394[16], net1394[17], net1394[18], net1394[19], net1394[20],
     net1394[21], net1394[22], net1394[23]}),
     .slf_op_02_17(slf_op_02_17[3:0]), .sp12_v_b_02_17({net1109[0],
     net1109[1], net1109[2], net1109[3], net1109[4], net1109[5],
     net1109[6], net1109[7], net1109[8], net1109[9], net1109[10],
     net1109[11], net1109[12], net1109[13], net1109[14], net1109[15],
     net1109[16], net1109[17], net1109[18], net1109[19], net1109[20],
     net1109[21], net1109[22], net1109[23]}),
     .padeb_t_l(padeb_t_l[11:0]), .bl_03(bl[167:126]), .ceb_o(net1412),
     .pado_t_l(pado_t_l[11:0]), .hold_t_l(hold_t_l),
     .slf_op_05_17(slf_op_05_17[3:0]), .ceb_i(ceb_i));
lt_1x8_top_ice1f I_lt_col_t01 ( .glb_netwk_b({net1451[0], net1451[1],
     net1451[2], net1451[3], net1451[4], net1451[5], net1451[6],
     net1451[7]}), .rgt_op_03({net929[0], net929[1], net929[2],
     net929[3], net929[4], net929[5], net929[6], net929[7]}),
     .slf_op_02({net818[0], net818[1], net818[2], net818[3], net818[4],
     net818[5], net818[6], net818[7]}), .rgt_op_02({net931[0],
     net931[1], net931[2], net931[3], net931[4], net931[5], net931[6],
     net931[7]}), .rgt_op_01(slf_op_02_09[7:0]), .purst(purst),
     .prog(prog), .lft_op_04({slf_op_00_12[3], slf_op_00_12[2],
     slf_op_00_12[1], slf_op_00_12[0], slf_op_00_12[3],
     slf_op_00_12[2], slf_op_00_12[1], slf_op_00_12[0]}),
     .lft_op_03({slf_op_00_11[3], slf_op_00_11[2], slf_op_00_11[1],
     slf_op_00_11[0], slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0]}), .lft_op_02({slf_op_00_10[3],
     slf_op_00_10[2], slf_op_00_10[1], slf_op_00_10[0],
     slf_op_00_10[3], slf_op_00_10[2], slf_op_00_10[1],
     slf_op_00_10[0]}), .lft_op_01({slf_op_00_09[3], slf_op_00_09[2],
     slf_op_00_09[1], slf_op_00_09[0], slf_op_00_09[3],
     slf_op_00_09[2], slf_op_00_09[1], slf_op_00_09[0]}),
     .rgt_op_04({net939[0], net939[1], net939[2], net939[3], net939[4],
     net939[5], net939[6], net939[7]}), .carry_in(carry_in_01_09),
     .bnl_op_01(bnl_op_01_09[7:0]), .slf_op_04({net858[0], net858[1],
     net858[2], net858[3], net858[4], net858[5], net858[6],
     net858[7]}), .slf_op_03({net834[0], net834[1], net834[2],
     net834[3], net834[4], net834[5], net834[6], net834[7]}),
     .slf_op_01(slf_op_01_09[7:0]), .sp4_h_l_04({net828[0], net828[1],
     net828[2], net828[3], net828[4], net828[5], net828[6], net828[7],
     net828[8], net828[9], net828[10], net828[11], net828[12],
     net828[13], net828[14], net828[15], net828[16], net828[17],
     net828[18], net828[19], net828[20], net828[21], net828[22],
     net828[23], net828[24], net828[25], net828[26], net828[27],
     net828[28], net828[29], net828[30], net828[31], net828[32],
     net828[33], net828[34], net828[35], net828[36], net828[37],
     net828[38], net828[39], net828[40], net828[41], net828[42],
     net828[43], net828[44], net828[45], net828[46], net828[47]}),
     .carry_out(net946), .vdd_cntl(vdd_cntl_l[127:0]),
     .sp12_h_r_04({net948[0], net948[1], net948[2], net948[3],
     net948[4], net948[5], net948[6], net948[7], net948[8], net948[9],
     net948[10], net948[11], net948[12], net948[13], net948[14],
     net948[15], net948[16], net948[17], net948[18], net948[19],
     net948[20], net948[21], net948[22], net948[23]}),
     .sp12_h_r_03({net949[0], net949[1], net949[2], net949[3],
     net949[4], net949[5], net949[6], net949[7], net949[8], net949[9],
     net949[10], net949[11], net949[12], net949[13], net949[14],
     net949[15], net949[16], net949[17], net949[18], net949[19],
     net949[20], net949[21], net949[22], net949[23]}),
     .sp12_h_r_02({net950[0], net950[1], net950[2], net950[3],
     net950[4], net950[5], net950[6], net950[7], net950[8], net950[9],
     net950[10], net950[11], net950[12], net950[13], net950[14],
     net950[15], net950[16], net950[17], net950[18], net950[19],
     net950[20], net950[21], net950[22], net950[23]}),
     .sp12_h_r_01({net951[0], net951[1], net951[2], net951[3],
     net951[4], net951[5], net951[6], net951[7], net951[8], net951[9],
     net951[10], net951[11], net951[12], net951[13], net951[14],
     net951[15], net951[16], net951[17], net951[18], net951[19],
     net951[20], net951[21], net951[22], net951[23]}),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_01_09[47:0]), .sp4_r_v_b_04({net954[0],
     net954[1], net954[2], net954[3], net954[4], net954[5], net954[6],
     net954[7], net954[8], net954[9], net954[10], net954[11],
     net954[12], net954[13], net954[14], net954[15], net954[16],
     net954[17], net954[18], net954[19], net954[20], net954[21],
     net954[22], net954[23], net954[24], net954[25], net954[26],
     net954[27], net954[28], net954[29], net954[30], net954[31],
     net954[32], net954[33], net954[34], net954[35], net954[36],
     net954[37], net954[38], net954[39], net954[40], net954[41],
     net954[42], net954[43], net954[44], net954[45], net954[46],
     net954[47]}), .sp4_r_v_b_03({net955[0], net955[1], net955[2],
     net955[3], net955[4], net955[5], net955[6], net955[7], net955[8],
     net955[9], net955[10], net955[11], net955[12], net955[13],
     net955[14], net955[15], net955[16], net955[17], net955[18],
     net955[19], net955[20], net955[21], net955[22], net955[23],
     net955[24], net955[25], net955[26], net955[27], net955[28],
     net955[29], net955[30], net955[31], net955[32], net955[33],
     net955[34], net955[35], net955[36], net955[37], net955[38],
     net955[39], net955[40], net955[41], net955[42], net955[43],
     net955[44], net955[45], net955[46], net955[47]}),
     .sp4_r_v_b_02({net956[0], net956[1], net956[2], net956[3],
     net956[4], net956[5], net956[6], net956[7], net956[8], net956[9],
     net956[10], net956[11], net956[12], net956[13], net956[14],
     net956[15], net956[16], net956[17], net956[18], net956[19],
     net956[20], net956[21], net956[22], net956[23], net956[24],
     net956[25], net956[26], net956[27], net956[28], net956[29],
     net956[30], net956[31], net956[32], net956[33], net956[34],
     net956[35], net956[36], net956[37], net956[38], net956[39],
     net956[40], net956[41], net956[42], net956[43], net956[44],
     net956[45], net956[46], net956[47]}),
     .sp4_r_v_b_01(sp4_v_b_02_09[47:0]), .sp4_h_r_04({net958[0],
     net958[1], net958[2], net958[3], net958[4], net958[5], net958[6],
     net958[7], net958[8], net958[9], net958[10], net958[11],
     net958[12], net958[13], net958[14], net958[15], net958[16],
     net958[17], net958[18], net958[19], net958[20], net958[21],
     net958[22], net958[23], net958[24], net958[25], net958[26],
     net958[27], net958[28], net958[29], net958[30], net958[31],
     net958[32], net958[33], net958[34], net958[35], net958[36],
     net958[37], net958[38], net958[39], net958[40], net958[41],
     net958[42], net958[43], net958[44], net958[45], net958[46],
     net958[47]}), .sp4_h_r_03({net959[0], net959[1], net959[2],
     net959[3], net959[4], net959[5], net959[6], net959[7], net959[8],
     net959[9], net959[10], net959[11], net959[12], net959[13],
     net959[14], net959[15], net959[16], net959[17], net959[18],
     net959[19], net959[20], net959[21], net959[22], net959[23],
     net959[24], net959[25], net959[26], net959[27], net959[28],
     net959[29], net959[30], net959[31], net959[32], net959[33],
     net959[34], net959[35], net959[36], net959[37], net959[38],
     net959[39], net959[40], net959[41], net959[42], net959[43],
     net959[44], net959[45], net959[46], net959[47]}),
     .sp4_h_r_02({net960[0], net960[1], net960[2], net960[3],
     net960[4], net960[5], net960[6], net960[7], net960[8], net960[9],
     net960[10], net960[11], net960[12], net960[13], net960[14],
     net960[15], net960[16], net960[17], net960[18], net960[19],
     net960[20], net960[21], net960[22], net960[23], net960[24],
     net960[25], net960[26], net960[27], net960[28], net960[29],
     net960[30], net960[31], net960[32], net960[33], net960[34],
     net960[35], net960[36], net960[37], net960[38], net960[39],
     net960[40], net960[41], net960[42], net960[43], net960[44],
     net960[45], net960[46], net960[47]}), .sp4_h_r_01({net961[0],
     net961[1], net961[2], net961[3], net961[4], net961[5], net961[6],
     net961[7], net961[8], net961[9], net961[10], net961[11],
     net961[12], net961[13], net961[14], net961[15], net961[16],
     net961[17], net961[18], net961[19], net961[20], net961[21],
     net961[22], net961[23], net961[24], net961[25], net961[26],
     net961[27], net961[28], net961[29], net961[30], net961[31],
     net961[32], net961[33], net961[34], net961[35], net961[36],
     net961[37], net961[38], net961[39], net961[40], net961[41],
     net961[42], net961[43], net961[44], net961[45], net961[46],
     net961[47]}), .sp4_h_l_03({net827[0], net827[1], net827[2],
     net827[3], net827[4], net827[5], net827[6], net827[7], net827[8],
     net827[9], net827[10], net827[11], net827[12], net827[13],
     net827[14], net827[15], net827[16], net827[17], net827[18],
     net827[19], net827[20], net827[21], net827[22], net827[23],
     net827[24], net827[25], net827[26], net827[27], net827[28],
     net827[29], net827[30], net827[31], net827[32], net827[33],
     net827[34], net827[35], net827[36], net827[37], net827[38],
     net827[39], net827[40], net827[41], net827[42], net827[43],
     net827[44], net827[45], net827[46], net827[47]}),
     .sp4_h_l_02({net829[0], net829[1], net829[2], net829[3],
     net829[4], net829[5], net829[6], net829[7], net829[8], net829[9],
     net829[10], net829[11], net829[12], net829[13], net829[14],
     net829[15], net829[16], net829[17], net829[18], net829[19],
     net829[20], net829[21], net829[22], net829[23], net829[24],
     net829[25], net829[26], net829[27], net829[28], net829[29],
     net829[30], net829[31], net829[32], net829[33], net829[34],
     net829[35], net829[36], net829[37], net829[38], net829[39],
     net829[40], net829[41], net829[42], net829[43], net829[44],
     net829[45], net829[46], net829[47]}), .sp4_h_l_01({net830[0],
     net830[1], net830[2], net830[3], net830[4], net830[5], net830[6],
     net830[7], net830[8], net830[9], net830[10], net830[11],
     net830[12], net830[13], net830[14], net830[15], net830[16],
     net830[17], net830[18], net830[19], net830[20], net830[21],
     net830[22], net830[23], net830[24], net830[25], net830[26],
     net830[27], net830[28], net830[29], net830[30], net830[31],
     net830[32], net830[33], net830[34], net830[35], net830[36],
     net830[37], net830[38], net830[39], net830[40], net830[41],
     net830[42], net830[43], net830[44], net830[45], net830[46],
     net830[47]}), .bl(bl[71:18]), .bot_op_01(bot_op_01_09[7:0]),
     .sp12_h_l_01({net855[0], net855[1], net855[2], net855[3],
     net855[4], net855[5], net855[6], net855[7], net855[8], net855[9],
     net855[10], net855[11], net855[12], net855[13], net855[14],
     net855[15], net855[16], net855[17], net855[18], net855[19],
     net855[20], net855[21], net855[22], net855[23]}),
     .sp12_h_l_02({net849[0], net849[1], net849[2], net849[3],
     net849[4], net849[5], net849[6], net849[7], net849[8], net849[9],
     net849[10], net849[11], net849[12], net849[13], net849[14],
     net849[15], net849[16], net849[17], net849[18], net849[19],
     net849[20], net849[21], net849[22], net849[23]}),
     .sp12_h_l_03({net856[0], net856[1], net856[2], net856[3],
     net856[4], net856[5], net856[6], net856[7], net856[8], net856[9],
     net856[10], net856[11], net856[12], net856[13], net856[14],
     net856[15], net856[16], net856[17], net856[18], net856[19],
     net856[20], net856[21], net856[22], net856[23]}),
     .sp12_h_l_04({net850[0], net850[1], net850[2], net850[3],
     net850[4], net850[5], net850[6], net850[7], net850[8], net850[9],
     net850[10], net850[11], net850[12], net850[13], net850[14],
     net850[15], net850[16], net850[17], net850[18], net850[19],
     net850[20], net850[21], net850[22], net850[23]}),
     .sp4_v_b_04({net1449[0], net1449[1], net1449[2], net1449[3],
     net1449[4], net1449[5], net1449[6], net1449[7], net1449[8],
     net1449[9], net1449[10], net1449[11], net1449[12], net1449[13],
     net1449[14], net1449[15], net1449[16], net1449[17], net1449[18],
     net1449[19], net1449[20], net1449[21], net1449[22], net1449[23],
     net1449[24], net1449[25], net1449[26], net1449[27], net1449[28],
     net1449[29], net1449[30], net1449[31], net1449[32], net1449[33],
     net1449[34], net1449[35], net1449[36], net1449[37], net1449[38],
     net1449[39], net1449[40], net1449[41], net1449[42], net1449[43],
     net1449[44], net1449[45], net1449[46], net1449[47]}),
     .sp4_v_b_03({net1450[0], net1450[1], net1450[2], net1450[3],
     net1450[4], net1450[5], net1450[6], net1450[7], net1450[8],
     net1450[9], net1450[10], net1450[11], net1450[12], net1450[13],
     net1450[14], net1450[15], net1450[16], net1450[17], net1450[18],
     net1450[19], net1450[20], net1450[21], net1450[22], net1450[23],
     net1450[24], net1450[25], net1450[26], net1450[27], net1450[28],
     net1450[29], net1450[30], net1450[31], net1450[32], net1450[33],
     net1450[34], net1450[35], net1450[36], net1450[37], net1450[38],
     net1450[39], net1450[40], net1450[41], net1450[42], net1450[43],
     net1450[44], net1450[45], net1450[46], net1450[47]}),
     .sp4_v_b_02({net1448[0], net1448[1], net1448[2], net1448[3],
     net1448[4], net1448[5], net1448[6], net1448[7], net1448[8],
     net1448[9], net1448[10], net1448[11], net1448[12], net1448[13],
     net1448[14], net1448[15], net1448[16], net1448[17], net1448[18],
     net1448[19], net1448[20], net1448[21], net1448[22], net1448[23],
     net1448[24], net1448[25], net1448[26], net1448[27], net1448[28],
     net1448[29], net1448[30], net1448[31], net1448[32], net1448[33],
     net1448[34], net1448[35], net1448[36], net1448[37], net1448[38],
     net1448[39], net1448[40], net1448[41], net1448[42], net1448[43],
     net1448[44], net1448[45], net1448[46], net1448[47]}),
     .bnr_op_01(bnr_op_01_09[7:0]), .sp4_h_l_05({net809[0], net809[1],
     net809[2], net809[3], net809[4], net809[5], net809[6], net809[7],
     net809[8], net809[9], net809[10], net809[11], net809[12],
     net809[13], net809[14], net809[15], net809[16], net809[17],
     net809[18], net809[19], net809[20], net809[21], net809[22],
     net809[23], net809[24], net809[25], net809[26], net809[27],
     net809[28], net809[29], net809[30], net809[31], net809[32],
     net809[33], net809[34], net809[35], net809[36], net809[37],
     net809[38], net809[39], net809[40], net809[41], net809[42],
     net809[43], net809[44], net809[45], net809[46], net809[47]}),
     .sp4_h_l_06({net819[0], net819[1], net819[2], net819[3],
     net819[4], net819[5], net819[6], net819[7], net819[8], net819[9],
     net819[10], net819[11], net819[12], net819[13], net819[14],
     net819[15], net819[16], net819[17], net819[18], net819[19],
     net819[20], net819[21], net819[22], net819[23], net819[24],
     net819[25], net819[26], net819[27], net819[28], net819[29],
     net819[30], net819[31], net819[32], net819[33], net819[34],
     net819[35], net819[36], net819[37], net819[38], net819[39],
     net819[40], net819[41], net819[42], net819[43], net819[44],
     net819[45], net819[46], net819[47]}), .sp4_h_l_07({net826[0],
     net826[1], net826[2], net826[3], net826[4], net826[5], net826[6],
     net826[7], net826[8], net826[9], net826[10], net826[11],
     net826[12], net826[13], net826[14], net826[15], net826[16],
     net826[17], net826[18], net826[19], net826[20], net826[21],
     net826[22], net826[23], net826[24], net826[25], net826[26],
     net826[27], net826[28], net826[29], net826[30], net826[31],
     net826[32], net826[33], net826[34], net826[35], net826[36],
     net826[37], net826[38], net826[39], net826[40], net826[41],
     net826[42], net826[43], net826[44], net826[45], net826[46],
     net826[47]}), .sp4_h_l_08({net825[0], net825[1], net825[2],
     net825[3], net825[4], net825[5], net825[6], net825[7], net825[8],
     net825[9], net825[10], net825[11], net825[12], net825[13],
     net825[14], net825[15], net825[16], net825[17], net825[18],
     net825[19], net825[20], net825[21], net825[22], net825[23],
     net825[24], net825[25], net825[26], net825[27], net825[28],
     net825[29], net825[30], net825[31], net825[32], net825[33],
     net825[34], net825[35], net825[36], net825[37], net825[38],
     net825[39], net825[40], net825[41], net825[42], net825[43],
     net825[44], net825[45], net825[46], net825[47]}),
     .sp4_h_r_08({net979[0], net979[1], net979[2], net979[3],
     net979[4], net979[5], net979[6], net979[7], net979[8], net979[9],
     net979[10], net979[11], net979[12], net979[13], net979[14],
     net979[15], net979[16], net979[17], net979[18], net979[19],
     net979[20], net979[21], net979[22], net979[23], net979[24],
     net979[25], net979[26], net979[27], net979[28], net979[29],
     net979[30], net979[31], net979[32], net979[33], net979[34],
     net979[35], net979[36], net979[37], net979[38], net979[39],
     net979[40], net979[41], net979[42], net979[43], net979[44],
     net979[45], net979[46], net979[47]}), .sp4_h_r_07({net980[0],
     net980[1], net980[2], net980[3], net980[4], net980[5], net980[6],
     net980[7], net980[8], net980[9], net980[10], net980[11],
     net980[12], net980[13], net980[14], net980[15], net980[16],
     net980[17], net980[18], net980[19], net980[20], net980[21],
     net980[22], net980[23], net980[24], net980[25], net980[26],
     net980[27], net980[28], net980[29], net980[30], net980[31],
     net980[32], net980[33], net980[34], net980[35], net980[36],
     net980[37], net980[38], net980[39], net980[40], net980[41],
     net980[42], net980[43], net980[44], net980[45], net980[46],
     net980[47]}), .sp4_h_r_06({net981[0], net981[1], net981[2],
     net981[3], net981[4], net981[5], net981[6], net981[7], net981[8],
     net981[9], net981[10], net981[11], net981[12], net981[13],
     net981[14], net981[15], net981[16], net981[17], net981[18],
     net981[19], net981[20], net981[21], net981[22], net981[23],
     net981[24], net981[25], net981[26], net981[27], net981[28],
     net981[29], net981[30], net981[31], net981[32], net981[33],
     net981[34], net981[35], net981[36], net981[37], net981[38],
     net981[39], net981[40], net981[41], net981[42], net981[43],
     net981[44], net981[45], net981[46], net981[47]}),
     .sp4_h_r_05({net982[0], net982[1], net982[2], net982[3],
     net982[4], net982[5], net982[6], net982[7], net982[8], net982[9],
     net982[10], net982[11], net982[12], net982[13], net982[14],
     net982[15], net982[16], net982[17], net982[18], net982[19],
     net982[20], net982[21], net982[22], net982[23], net982[24],
     net982[25], net982[26], net982[27], net982[28], net982[29],
     net982[30], net982[31], net982[32], net982[33], net982[34],
     net982[35], net982[36], net982[37], net982[38], net982[39],
     net982[40], net982[41], net982[42], net982[43], net982[44],
     net982[45], net982[46], net982[47]}), .slf_op_05({net833[0],
     net833[1], net833[2], net833[3], net833[4], net833[5], net833[6],
     net833[7]}), .slf_op_06({net832[0], net832[1], net832[2],
     net832[3], net832[4], net832[5], net832[6], net832[7]}),
     .slf_op_07({net831[0], net831[1], net831[2], net831[3], net831[4],
     net831[5], net831[6], net831[7]}), .slf_op_08({net836[0],
     net836[1], net836[2], net836[3], net836[4], net836[5], net836[6],
     net836[7]}), .rgt_op_08({net987[0], net987[1], net987[2],
     net987[3], net987[4], net987[5], net987[6], net987[7]}),
     .rgt_op_07({net988[0], net988[1], net988[2], net988[3], net988[4],
     net988[5], net988[6], net988[7]}), .rgt_op_06({net989[0],
     net989[1], net989[2], net989[3], net989[4], net989[5], net989[6],
     net989[7]}), .rgt_op_05({net990[0], net990[1], net990[2],
     net990[3], net990[4], net990[5], net990[6], net990[7]}),
     .lft_op_08({slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0], slf_op_00_16[3], slf_op_00_16[2],
     slf_op_00_16[1], slf_op_00_16[0]}), .lft_op_07({slf_op_00_15[3],
     slf_op_00_15[2], slf_op_00_15[1], slf_op_00_15[0],
     slf_op_00_15[3], slf_op_00_15[2], slf_op_00_15[1],
     slf_op_00_15[0]}), .lft_op_06({slf_op_00_14[3], slf_op_00_14[2],
     slf_op_00_14[1], slf_op_00_14[0], slf_op_00_14[3],
     slf_op_00_14[2], slf_op_00_14[1], slf_op_00_14[0]}),
     .lft_op_05({slf_op_00_13[3], slf_op_00_13[2], slf_op_00_13[1],
     slf_op_00_13[0], slf_op_00_13[3], slf_op_00_13[2],
     slf_op_00_13[1], slf_op_00_13[0]}), .sp12_h_l_08({net851[0],
     net851[1], net851[2], net851[3], net851[4], net851[5], net851[6],
     net851[7], net851[8], net851[9], net851[10], net851[11],
     net851[12], net851[13], net851[14], net851[15], net851[16],
     net851[17], net851[18], net851[19], net851[20], net851[21],
     net851[22], net851[23]}), .sp12_h_l_07({net857[0], net857[1],
     net857[2], net857[3], net857[4], net857[5], net857[6], net857[7],
     net857[8], net857[9], net857[10], net857[11], net857[12],
     net857[13], net857[14], net857[15], net857[16], net857[17],
     net857[18], net857[19], net857[20], net857[21], net857[22],
     net857[23]}), .sp12_h_l_06({net852[0], net852[1], net852[2],
     net852[3], net852[4], net852[5], net852[6], net852[7], net852[8],
     net852[9], net852[10], net852[11], net852[12], net852[13],
     net852[14], net852[15], net852[16], net852[17], net852[18],
     net852[19], net852[20], net852[21], net852[22], net852[23]}),
     .sp12_h_r_05({net998[0], net998[1], net998[2], net998[3],
     net998[4], net998[5], net998[6], net998[7], net998[8], net998[9],
     net998[10], net998[11], net998[12], net998[13], net998[14],
     net998[15], net998[16], net998[17], net998[18], net998[19],
     net998[20], net998[21], net998[22], net998[23]}),
     .sp12_h_r_06({net999[0], net999[1], net999[2], net999[3],
     net999[4], net999[5], net999[6], net999[7], net999[8], net999[9],
     net999[10], net999[11], net999[12], net999[13], net999[14],
     net999[15], net999[16], net999[17], net999[18], net999[19],
     net999[20], net999[21], net999[22], net999[23]}),
     .sp12_h_r_07({net1000[0], net1000[1], net1000[2], net1000[3],
     net1000[4], net1000[5], net1000[6], net1000[7], net1000[8],
     net1000[9], net1000[10], net1000[11], net1000[12], net1000[13],
     net1000[14], net1000[15], net1000[16], net1000[17], net1000[18],
     net1000[19], net1000[20], net1000[21], net1000[22], net1000[23]}),
     .sp12_h_r_08({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7], net1001[8],
     net1001[9], net1001[10], net1001[11], net1001[12], net1001[13],
     net1001[14], net1001[15], net1001[16], net1001[17], net1001[18],
     net1001[19], net1001[20], net1001[21], net1001[22], net1001[23]}),
     .sp12_h_l_05({net854[0], net854[1], net854[2], net854[3],
     net854[4], net854[5], net854[6], net854[7], net854[8], net854[9],
     net854[10], net854[11], net854[12], net854[13], net854[14],
     net854[15], net854[16], net854[17], net854[18], net854[19],
     net854[20], net854[21], net854[22], net854[23]}),
     .sp4_r_v_b_05({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7], net1003[8],
     net1003[9], net1003[10], net1003[11], net1003[12], net1003[13],
     net1003[14], net1003[15], net1003[16], net1003[17], net1003[18],
     net1003[19], net1003[20], net1003[21], net1003[22], net1003[23],
     net1003[24], net1003[25], net1003[26], net1003[27], net1003[28],
     net1003[29], net1003[30], net1003[31], net1003[32], net1003[33],
     net1003[34], net1003[35], net1003[36], net1003[37], net1003[38],
     net1003[39], net1003[40], net1003[41], net1003[42], net1003[43],
     net1003[44], net1003[45], net1003[46], net1003[47]}),
     .sp4_r_v_b_06({net1004[0], net1004[1], net1004[2], net1004[3],
     net1004[4], net1004[5], net1004[6], net1004[7], net1004[8],
     net1004[9], net1004[10], net1004[11], net1004[12], net1004[13],
     net1004[14], net1004[15], net1004[16], net1004[17], net1004[18],
     net1004[19], net1004[20], net1004[21], net1004[22], net1004[23],
     net1004[24], net1004[25], net1004[26], net1004[27], net1004[28],
     net1004[29], net1004[30], net1004[31], net1004[32], net1004[33],
     net1004[34], net1004[35], net1004[36], net1004[37], net1004[38],
     net1004[39], net1004[40], net1004[41], net1004[42], net1004[43],
     net1004[44], net1004[45], net1004[46], net1004[47]}),
     .sp4_r_v_b_07({net1005[0], net1005[1], net1005[2], net1005[3],
     net1005[4], net1005[5], net1005[6], net1005[7], net1005[8],
     net1005[9], net1005[10], net1005[11], net1005[12], net1005[13],
     net1005[14], net1005[15], net1005[16], net1005[17], net1005[18],
     net1005[19], net1005[20], net1005[21], net1005[22], net1005[23],
     net1005[24], net1005[25], net1005[26], net1005[27], net1005[28],
     net1005[29], net1005[30], net1005[31], net1005[32], net1005[33],
     net1005[34], net1005[35], net1005[36], net1005[37], net1005[38],
     net1005[39], net1005[40], net1005[41], net1005[42], net1005[43],
     net1005[44], net1005[45], net1005[46], net1005[47]}),
     .sp4_r_v_b_08({net1006[0], net1006[1], net1006[2], net1006[3],
     net1006[4], net1006[5], net1006[6], net1006[7], net1006[8],
     net1006[9], net1006[10], net1006[11], net1006[12], net1006[13],
     net1006[14], net1006[15], net1006[16], net1006[17], net1006[18],
     net1006[19], net1006[20], net1006[21], net1006[22], net1006[23],
     net1006[24], net1006[25], net1006[26], net1006[27], net1006[28],
     net1006[29], net1006[30], net1006[31], net1006[32], net1006[33],
     net1006[34], net1006[35], net1006[36], net1006[37], net1006[38],
     net1006[39], net1006[40], net1006[41], net1006[42], net1006[43],
     net1006[44], net1006[45], net1006[46], net1006[47]}),
     .sp4_v_b_08({net1443[0], net1443[1], net1443[2], net1443[3],
     net1443[4], net1443[5], net1443[6], net1443[7], net1443[8],
     net1443[9], net1443[10], net1443[11], net1443[12], net1443[13],
     net1443[14], net1443[15], net1443[16], net1443[17], net1443[18],
     net1443[19], net1443[20], net1443[21], net1443[22], net1443[23],
     net1443[24], net1443[25], net1443[26], net1443[27], net1443[28],
     net1443[29], net1443[30], net1443[31], net1443[32], net1443[33],
     net1443[34], net1443[35], net1443[36], net1443[37], net1443[38],
     net1443[39], net1443[40], net1443[41], net1443[42], net1443[43],
     net1443[44], net1443[45], net1443[46], net1443[47]}),
     .sp4_v_b_07({net1444[0], net1444[1], net1444[2], net1444[3],
     net1444[4], net1444[5], net1444[6], net1444[7], net1444[8],
     net1444[9], net1444[10], net1444[11], net1444[12], net1444[13],
     net1444[14], net1444[15], net1444[16], net1444[17], net1444[18],
     net1444[19], net1444[20], net1444[21], net1444[22], net1444[23],
     net1444[24], net1444[25], net1444[26], net1444[27], net1444[28],
     net1444[29], net1444[30], net1444[31], net1444[32], net1444[33],
     net1444[34], net1444[35], net1444[36], net1444[37], net1444[38],
     net1444[39], net1444[40], net1444[41], net1444[42], net1444[43],
     net1444[44], net1444[45], net1444[46], net1444[47]}),
     .sp4_v_b_06({net1445[0], net1445[1], net1445[2], net1445[3],
     net1445[4], net1445[5], net1445[6], net1445[7], net1445[8],
     net1445[9], net1445[10], net1445[11], net1445[12], net1445[13],
     net1445[14], net1445[15], net1445[16], net1445[17], net1445[18],
     net1445[19], net1445[20], net1445[21], net1445[22], net1445[23],
     net1445[24], net1445[25], net1445[26], net1445[27], net1445[28],
     net1445[29], net1445[30], net1445[31], net1445[32], net1445[33],
     net1445[34], net1445[35], net1445[36], net1445[37], net1445[38],
     net1445[39], net1445[40], net1445[41], net1445[42], net1445[43],
     net1445[44], net1445[45], net1445[46], net1445[47]}),
     .sp4_v_b_05({net1446[0], net1446[1], net1446[2], net1446[3],
     net1446[4], net1446[5], net1446[6], net1446[7], net1446[8],
     net1446[9], net1446[10], net1446[11], net1446[12], net1446[13],
     net1446[14], net1446[15], net1446[16], net1446[17], net1446[18],
     net1446[19], net1446[20], net1446[21], net1446[22], net1446[23],
     net1446[24], net1446[25], net1446[26], net1446[27], net1446[28],
     net1446[29], net1446[30], net1446[31], net1446[32], net1446[33],
     net1446[34], net1446[35], net1446[36], net1446[37], net1446[38],
     net1446[39], net1446[40], net1446[41], net1446[42], net1446[43],
     net1446[44], net1446[45], net1446[46], net1446[47]}),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .wl(wl_l[127:0]), .sp12_v_t_08({net1014[0], net1014[1],
     net1014[2], net1014[3], net1014[4], net1014[5], net1014[6],
     net1014[7], net1014[8], net1014[9], net1014[10], net1014[11],
     net1014[12], net1014[13], net1014[14], net1014[15], net1014[16],
     net1014[17], net1014[18], net1014[19], net1014[20], net1014[21],
     net1014[22], net1014[23]}), .tnr_op_08({slf_op_02_17[3],
     slf_op_02_17[2], slf_op_02_17[1], slf_op_02_17[0],
     slf_op_02_17[3], slf_op_02_17[2], slf_op_02_17[1],
     slf_op_02_17[0]}), .top_op_08({slf_op_01_17[3], slf_op_01_17[2],
     slf_op_01_17[1], slf_op_01_17[0], slf_op_01_17[3],
     slf_op_01_17[2], slf_op_01_17[1], slf_op_01_17[0]}),
     .tnl_op_08({tiegnd_qtl, tiegnd_qtl, tiegnd_qtl, tiegnd_qtl,
     tiegnd_qtl, tiegnd_qtl, tiegnd_qtl, tiegnd_qtl}),
     .sp4_v_t_08({net1018[0], net1018[1], net1018[2], net1018[3],
     net1018[4], net1018[5], net1018[6], net1018[7], net1018[8],
     net1018[9], net1018[10], net1018[11], net1018[12], net1018[13],
     net1018[14], net1018[15], net1018[16], net1018[17], net1018[18],
     net1018[19], net1018[20], net1018[21], net1018[22], net1018[23],
     net1018[24], net1018[25], net1018[26], net1018[27], net1018[28],
     net1018[29], net1018[30], net1018[31], net1018[32], net1018[33],
     net1018[34], net1018[35], net1018[36], net1018[37], net1018[38],
     net1018[39], net1018[40], net1018[41], net1018[42], net1018[43],
     net1018[44], net1018[45], net1018[46], net1018[47]}),
     .lc_bot(lc_bot_01_09), .op_vic(net1020),
     .sp12_v_b_01(sp12_v_b_01_09[23:0]), .glb_netwk_t({net1022[0],
     net1022[1], net1022[2], net1022[3], net1022[4], net1022[5],
     net1022[6], net1022[7]}));
lt_1x8_top_ice1f I_lt_col_t02 ( .glb_netwk_b({net1452[0], net1452[1],
     net1452[2], net1452[3], net1452[4], net1452[5], net1452[6],
     net1452[7]}), .rgt_op_03({net1024[0], net1024[1], net1024[2],
     net1024[3], net1024[4], net1024[5], net1024[6], net1024[7]}),
     .slf_op_02({net931[0], net931[1], net931[2], net931[3], net931[4],
     net931[5], net931[6], net931[7]}), .rgt_op_02({net1026[0],
     net1026[1], net1026[2], net1026[3], net1026[4], net1026[5],
     net1026[6], net1026[7]}), .rgt_op_01(slf_op_03_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04({net858[0], net858[1],
     net858[2], net858[3], net858[4], net858[5], net858[6],
     net858[7]}), .lft_op_03({net834[0], net834[1], net834[2],
     net834[3], net834[4], net834[5], net834[6], net834[7]}),
     .lft_op_02({net818[0], net818[1], net818[2], net818[3], net818[4],
     net818[5], net818[6], net818[7]}), .lft_op_01(slf_op_01_09[7:0]),
     .rgt_op_04({net1034[0], net1034[1], net1034[2], net1034[3],
     net1034[4], net1034[5], net1034[6], net1034[7]}),
     .carry_in(carry_in_02_09), .bnl_op_01(bnl_op_02_09[7:0]),
     .slf_op_04({net939[0], net939[1], net939[2], net939[3], net939[4],
     net939[5], net939[6], net939[7]}), .slf_op_03({net929[0],
     net929[1], net929[2], net929[3], net929[4], net929[5], net929[6],
     net929[7]}), .slf_op_01(slf_op_02_09[7:0]),
     .sp4_h_l_04({net958[0], net958[1], net958[2], net958[3],
     net958[4], net958[5], net958[6], net958[7], net958[8], net958[9],
     net958[10], net958[11], net958[12], net958[13], net958[14],
     net958[15], net958[16], net958[17], net958[18], net958[19],
     net958[20], net958[21], net958[22], net958[23], net958[24],
     net958[25], net958[26], net958[27], net958[28], net958[29],
     net958[30], net958[31], net958[32], net958[33], net958[34],
     net958[35], net958[36], net958[37], net958[38], net958[39],
     net958[40], net958[41], net958[42], net958[43], net958[44],
     net958[45], net958[46], net958[47]}), .carry_out(net1041),
     .vdd_cntl(vdd_cntl_l[127:0]), .sp12_h_r_04({net1043[0],
     net1043[1], net1043[2], net1043[3], net1043[4], net1043[5],
     net1043[6], net1043[7], net1043[8], net1043[9], net1043[10],
     net1043[11], net1043[12], net1043[13], net1043[14], net1043[15],
     net1043[16], net1043[17], net1043[18], net1043[19], net1043[20],
     net1043[21], net1043[22], net1043[23]}), .sp12_h_r_03({net1044[0],
     net1044[1], net1044[2], net1044[3], net1044[4], net1044[5],
     net1044[6], net1044[7], net1044[8], net1044[9], net1044[10],
     net1044[11], net1044[12], net1044[13], net1044[14], net1044[15],
     net1044[16], net1044[17], net1044[18], net1044[19], net1044[20],
     net1044[21], net1044[22], net1044[23]}), .sp12_h_r_02({net1045[0],
     net1045[1], net1045[2], net1045[3], net1045[4], net1045[5],
     net1045[6], net1045[7], net1045[8], net1045[9], net1045[10],
     net1045[11], net1045[12], net1045[13], net1045[14], net1045[15],
     net1045[16], net1045[17], net1045[18], net1045[19], net1045[20],
     net1045[21], net1045[22], net1045[23]}), .sp12_h_r_01({net1046[0],
     net1046[1], net1046[2], net1046[3], net1046[4], net1046[5],
     net1046[6], net1046[7], net1046[8], net1046[9], net1046[10],
     net1046[11], net1046[12], net1046[13], net1046[14], net1046[15],
     net1046[16], net1046[17], net1046[18], net1046[19], net1046[20],
     net1046[21], net1046[22], net1046[23]}),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_02_09[47:0]), .sp4_r_v_b_04({net1049[0],
     net1049[1], net1049[2], net1049[3], net1049[4], net1049[5],
     net1049[6], net1049[7], net1049[8], net1049[9], net1049[10],
     net1049[11], net1049[12], net1049[13], net1049[14], net1049[15],
     net1049[16], net1049[17], net1049[18], net1049[19], net1049[20],
     net1049[21], net1049[22], net1049[23], net1049[24], net1049[25],
     net1049[26], net1049[27], net1049[28], net1049[29], net1049[30],
     net1049[31], net1049[32], net1049[33], net1049[34], net1049[35],
     net1049[36], net1049[37], net1049[38], net1049[39], net1049[40],
     net1049[41], net1049[42], net1049[43], net1049[44], net1049[45],
     net1049[46], net1049[47]}), .sp4_r_v_b_03({net1050[0], net1050[1],
     net1050[2], net1050[3], net1050[4], net1050[5], net1050[6],
     net1050[7], net1050[8], net1050[9], net1050[10], net1050[11],
     net1050[12], net1050[13], net1050[14], net1050[15], net1050[16],
     net1050[17], net1050[18], net1050[19], net1050[20], net1050[21],
     net1050[22], net1050[23], net1050[24], net1050[25], net1050[26],
     net1050[27], net1050[28], net1050[29], net1050[30], net1050[31],
     net1050[32], net1050[33], net1050[34], net1050[35], net1050[36],
     net1050[37], net1050[38], net1050[39], net1050[40], net1050[41],
     net1050[42], net1050[43], net1050[44], net1050[45], net1050[46],
     net1050[47]}), .sp4_r_v_b_02({net1051[0], net1051[1], net1051[2],
     net1051[3], net1051[4], net1051[5], net1051[6], net1051[7],
     net1051[8], net1051[9], net1051[10], net1051[11], net1051[12],
     net1051[13], net1051[14], net1051[15], net1051[16], net1051[17],
     net1051[18], net1051[19], net1051[20], net1051[21], net1051[22],
     net1051[23], net1051[24], net1051[25], net1051[26], net1051[27],
     net1051[28], net1051[29], net1051[30], net1051[31], net1051[32],
     net1051[33], net1051[34], net1051[35], net1051[36], net1051[37],
     net1051[38], net1051[39], net1051[40], net1051[41], net1051[42],
     net1051[43], net1051[44], net1051[45], net1051[46], net1051[47]}),
     .sp4_r_v_b_01(sp4_v_b_03_09[47:0]), .sp4_h_r_04({net1053[0],
     net1053[1], net1053[2], net1053[3], net1053[4], net1053[5],
     net1053[6], net1053[7], net1053[8], net1053[9], net1053[10],
     net1053[11], net1053[12], net1053[13], net1053[14], net1053[15],
     net1053[16], net1053[17], net1053[18], net1053[19], net1053[20],
     net1053[21], net1053[22], net1053[23], net1053[24], net1053[25],
     net1053[26], net1053[27], net1053[28], net1053[29], net1053[30],
     net1053[31], net1053[32], net1053[33], net1053[34], net1053[35],
     net1053[36], net1053[37], net1053[38], net1053[39], net1053[40],
     net1053[41], net1053[42], net1053[43], net1053[44], net1053[45],
     net1053[46], net1053[47]}), .sp4_h_r_03({net1054[0], net1054[1],
     net1054[2], net1054[3], net1054[4], net1054[5], net1054[6],
     net1054[7], net1054[8], net1054[9], net1054[10], net1054[11],
     net1054[12], net1054[13], net1054[14], net1054[15], net1054[16],
     net1054[17], net1054[18], net1054[19], net1054[20], net1054[21],
     net1054[22], net1054[23], net1054[24], net1054[25], net1054[26],
     net1054[27], net1054[28], net1054[29], net1054[30], net1054[31],
     net1054[32], net1054[33], net1054[34], net1054[35], net1054[36],
     net1054[37], net1054[38], net1054[39], net1054[40], net1054[41],
     net1054[42], net1054[43], net1054[44], net1054[45], net1054[46],
     net1054[47]}), .sp4_h_r_02({net1055[0], net1055[1], net1055[2],
     net1055[3], net1055[4], net1055[5], net1055[6], net1055[7],
     net1055[8], net1055[9], net1055[10], net1055[11], net1055[12],
     net1055[13], net1055[14], net1055[15], net1055[16], net1055[17],
     net1055[18], net1055[19], net1055[20], net1055[21], net1055[22],
     net1055[23], net1055[24], net1055[25], net1055[26], net1055[27],
     net1055[28], net1055[29], net1055[30], net1055[31], net1055[32],
     net1055[33], net1055[34], net1055[35], net1055[36], net1055[37],
     net1055[38], net1055[39], net1055[40], net1055[41], net1055[42],
     net1055[43], net1055[44], net1055[45], net1055[46], net1055[47]}),
     .sp4_h_r_01({net1056[0], net1056[1], net1056[2], net1056[3],
     net1056[4], net1056[5], net1056[6], net1056[7], net1056[8],
     net1056[9], net1056[10], net1056[11], net1056[12], net1056[13],
     net1056[14], net1056[15], net1056[16], net1056[17], net1056[18],
     net1056[19], net1056[20], net1056[21], net1056[22], net1056[23],
     net1056[24], net1056[25], net1056[26], net1056[27], net1056[28],
     net1056[29], net1056[30], net1056[31], net1056[32], net1056[33],
     net1056[34], net1056[35], net1056[36], net1056[37], net1056[38],
     net1056[39], net1056[40], net1056[41], net1056[42], net1056[43],
     net1056[44], net1056[45], net1056[46], net1056[47]}),
     .sp4_h_l_03({net959[0], net959[1], net959[2], net959[3],
     net959[4], net959[5], net959[6], net959[7], net959[8], net959[9],
     net959[10], net959[11], net959[12], net959[13], net959[14],
     net959[15], net959[16], net959[17], net959[18], net959[19],
     net959[20], net959[21], net959[22], net959[23], net959[24],
     net959[25], net959[26], net959[27], net959[28], net959[29],
     net959[30], net959[31], net959[32], net959[33], net959[34],
     net959[35], net959[36], net959[37], net959[38], net959[39],
     net959[40], net959[41], net959[42], net959[43], net959[44],
     net959[45], net959[46], net959[47]}), .sp4_h_l_02({net960[0],
     net960[1], net960[2], net960[3], net960[4], net960[5], net960[6],
     net960[7], net960[8], net960[9], net960[10], net960[11],
     net960[12], net960[13], net960[14], net960[15], net960[16],
     net960[17], net960[18], net960[19], net960[20], net960[21],
     net960[22], net960[23], net960[24], net960[25], net960[26],
     net960[27], net960[28], net960[29], net960[30], net960[31],
     net960[32], net960[33], net960[34], net960[35], net960[36],
     net960[37], net960[38], net960[39], net960[40], net960[41],
     net960[42], net960[43], net960[44], net960[45], net960[46],
     net960[47]}), .sp4_h_l_01({net961[0], net961[1], net961[2],
     net961[3], net961[4], net961[5], net961[6], net961[7], net961[8],
     net961[9], net961[10], net961[11], net961[12], net961[13],
     net961[14], net961[15], net961[16], net961[17], net961[18],
     net961[19], net961[20], net961[21], net961[22], net961[23],
     net961[24], net961[25], net961[26], net961[27], net961[28],
     net961[29], net961[30], net961[31], net961[32], net961[33],
     net961[34], net961[35], net961[36], net961[37], net961[38],
     net961[39], net961[40], net961[41], net961[42], net961[43],
     net961[44], net961[45], net961[46], net961[47]}), .bl(bl[125:72]),
     .bot_op_01(bot_op_02_09[7:0]), .sp12_h_l_01({net951[0], net951[1],
     net951[2], net951[3], net951[4], net951[5], net951[6], net951[7],
     net951[8], net951[9], net951[10], net951[11], net951[12],
     net951[13], net951[14], net951[15], net951[16], net951[17],
     net951[18], net951[19], net951[20], net951[21], net951[22],
     net951[23]}), .sp12_h_l_02({net950[0], net950[1], net950[2],
     net950[3], net950[4], net950[5], net950[6], net950[7], net950[8],
     net950[9], net950[10], net950[11], net950[12], net950[13],
     net950[14], net950[15], net950[16], net950[17], net950[18],
     net950[19], net950[20], net950[21], net950[22], net950[23]}),
     .sp12_h_l_03({net949[0], net949[1], net949[2], net949[3],
     net949[4], net949[5], net949[6], net949[7], net949[8], net949[9],
     net949[10], net949[11], net949[12], net949[13], net949[14],
     net949[15], net949[16], net949[17], net949[18], net949[19],
     net949[20], net949[21], net949[22], net949[23]}),
     .sp12_h_l_04({net948[0], net948[1], net948[2], net948[3],
     net948[4], net948[5], net948[6], net948[7], net948[8], net948[9],
     net948[10], net948[11], net948[12], net948[13], net948[14],
     net948[15], net948[16], net948[17], net948[18], net948[19],
     net948[20], net948[21], net948[22], net948[23]}),
     .sp4_v_b_04({net954[0], net954[1], net954[2], net954[3],
     net954[4], net954[5], net954[6], net954[7], net954[8], net954[9],
     net954[10], net954[11], net954[12], net954[13], net954[14],
     net954[15], net954[16], net954[17], net954[18], net954[19],
     net954[20], net954[21], net954[22], net954[23], net954[24],
     net954[25], net954[26], net954[27], net954[28], net954[29],
     net954[30], net954[31], net954[32], net954[33], net954[34],
     net954[35], net954[36], net954[37], net954[38], net954[39],
     net954[40], net954[41], net954[42], net954[43], net954[44],
     net954[45], net954[46], net954[47]}), .sp4_v_b_03({net955[0],
     net955[1], net955[2], net955[3], net955[4], net955[5], net955[6],
     net955[7], net955[8], net955[9], net955[10], net955[11],
     net955[12], net955[13], net955[14], net955[15], net955[16],
     net955[17], net955[18], net955[19], net955[20], net955[21],
     net955[22], net955[23], net955[24], net955[25], net955[26],
     net955[27], net955[28], net955[29], net955[30], net955[31],
     net955[32], net955[33], net955[34], net955[35], net955[36],
     net955[37], net955[38], net955[39], net955[40], net955[41],
     net955[42], net955[43], net955[44], net955[45], net955[46],
     net955[47]}), .sp4_v_b_02({net956[0], net956[1], net956[2],
     net956[3], net956[4], net956[5], net956[6], net956[7], net956[8],
     net956[9], net956[10], net956[11], net956[12], net956[13],
     net956[14], net956[15], net956[16], net956[17], net956[18],
     net956[19], net956[20], net956[21], net956[22], net956[23],
     net956[24], net956[25], net956[26], net956[27], net956[28],
     net956[29], net956[30], net956[31], net956[32], net956[33],
     net956[34], net956[35], net956[36], net956[37], net956[38],
     net956[39], net956[40], net956[41], net956[42], net956[43],
     net956[44], net956[45], net956[46], net956[47]}),
     .bnr_op_01(bnr_op_02_09[7:0]), .sp4_h_l_05({net982[0], net982[1],
     net982[2], net982[3], net982[4], net982[5], net982[6], net982[7],
     net982[8], net982[9], net982[10], net982[11], net982[12],
     net982[13], net982[14], net982[15], net982[16], net982[17],
     net982[18], net982[19], net982[20], net982[21], net982[22],
     net982[23], net982[24], net982[25], net982[26], net982[27],
     net982[28], net982[29], net982[30], net982[31], net982[32],
     net982[33], net982[34], net982[35], net982[36], net982[37],
     net982[38], net982[39], net982[40], net982[41], net982[42],
     net982[43], net982[44], net982[45], net982[46], net982[47]}),
     .sp4_h_l_06({net981[0], net981[1], net981[2], net981[3],
     net981[4], net981[5], net981[6], net981[7], net981[8], net981[9],
     net981[10], net981[11], net981[12], net981[13], net981[14],
     net981[15], net981[16], net981[17], net981[18], net981[19],
     net981[20], net981[21], net981[22], net981[23], net981[24],
     net981[25], net981[26], net981[27], net981[28], net981[29],
     net981[30], net981[31], net981[32], net981[33], net981[34],
     net981[35], net981[36], net981[37], net981[38], net981[39],
     net981[40], net981[41], net981[42], net981[43], net981[44],
     net981[45], net981[46], net981[47]}), .sp4_h_l_07({net980[0],
     net980[1], net980[2], net980[3], net980[4], net980[5], net980[6],
     net980[7], net980[8], net980[9], net980[10], net980[11],
     net980[12], net980[13], net980[14], net980[15], net980[16],
     net980[17], net980[18], net980[19], net980[20], net980[21],
     net980[22], net980[23], net980[24], net980[25], net980[26],
     net980[27], net980[28], net980[29], net980[30], net980[31],
     net980[32], net980[33], net980[34], net980[35], net980[36],
     net980[37], net980[38], net980[39], net980[40], net980[41],
     net980[42], net980[43], net980[44], net980[45], net980[46],
     net980[47]}), .sp4_h_l_08({net979[0], net979[1], net979[2],
     net979[3], net979[4], net979[5], net979[6], net979[7], net979[8],
     net979[9], net979[10], net979[11], net979[12], net979[13],
     net979[14], net979[15], net979[16], net979[17], net979[18],
     net979[19], net979[20], net979[21], net979[22], net979[23],
     net979[24], net979[25], net979[26], net979[27], net979[28],
     net979[29], net979[30], net979[31], net979[32], net979[33],
     net979[34], net979[35], net979[36], net979[37], net979[38],
     net979[39], net979[40], net979[41], net979[42], net979[43],
     net979[44], net979[45], net979[46], net979[47]}),
     .sp4_h_r_08({net1074[0], net1074[1], net1074[2], net1074[3],
     net1074[4], net1074[5], net1074[6], net1074[7], net1074[8],
     net1074[9], net1074[10], net1074[11], net1074[12], net1074[13],
     net1074[14], net1074[15], net1074[16], net1074[17], net1074[18],
     net1074[19], net1074[20], net1074[21], net1074[22], net1074[23],
     net1074[24], net1074[25], net1074[26], net1074[27], net1074[28],
     net1074[29], net1074[30], net1074[31], net1074[32], net1074[33],
     net1074[34], net1074[35], net1074[36], net1074[37], net1074[38],
     net1074[39], net1074[40], net1074[41], net1074[42], net1074[43],
     net1074[44], net1074[45], net1074[46], net1074[47]}),
     .sp4_h_r_07({net1075[0], net1075[1], net1075[2], net1075[3],
     net1075[4], net1075[5], net1075[6], net1075[7], net1075[8],
     net1075[9], net1075[10], net1075[11], net1075[12], net1075[13],
     net1075[14], net1075[15], net1075[16], net1075[17], net1075[18],
     net1075[19], net1075[20], net1075[21], net1075[22], net1075[23],
     net1075[24], net1075[25], net1075[26], net1075[27], net1075[28],
     net1075[29], net1075[30], net1075[31], net1075[32], net1075[33],
     net1075[34], net1075[35], net1075[36], net1075[37], net1075[38],
     net1075[39], net1075[40], net1075[41], net1075[42], net1075[43],
     net1075[44], net1075[45], net1075[46], net1075[47]}),
     .sp4_h_r_06({net1076[0], net1076[1], net1076[2], net1076[3],
     net1076[4], net1076[5], net1076[6], net1076[7], net1076[8],
     net1076[9], net1076[10], net1076[11], net1076[12], net1076[13],
     net1076[14], net1076[15], net1076[16], net1076[17], net1076[18],
     net1076[19], net1076[20], net1076[21], net1076[22], net1076[23],
     net1076[24], net1076[25], net1076[26], net1076[27], net1076[28],
     net1076[29], net1076[30], net1076[31], net1076[32], net1076[33],
     net1076[34], net1076[35], net1076[36], net1076[37], net1076[38],
     net1076[39], net1076[40], net1076[41], net1076[42], net1076[43],
     net1076[44], net1076[45], net1076[46], net1076[47]}),
     .sp4_h_r_05({net1077[0], net1077[1], net1077[2], net1077[3],
     net1077[4], net1077[5], net1077[6], net1077[7], net1077[8],
     net1077[9], net1077[10], net1077[11], net1077[12], net1077[13],
     net1077[14], net1077[15], net1077[16], net1077[17], net1077[18],
     net1077[19], net1077[20], net1077[21], net1077[22], net1077[23],
     net1077[24], net1077[25], net1077[26], net1077[27], net1077[28],
     net1077[29], net1077[30], net1077[31], net1077[32], net1077[33],
     net1077[34], net1077[35], net1077[36], net1077[37], net1077[38],
     net1077[39], net1077[40], net1077[41], net1077[42], net1077[43],
     net1077[44], net1077[45], net1077[46], net1077[47]}),
     .slf_op_05({net990[0], net990[1], net990[2], net990[3], net990[4],
     net990[5], net990[6], net990[7]}), .slf_op_06({net989[0],
     net989[1], net989[2], net989[3], net989[4], net989[5], net989[6],
     net989[7]}), .slf_op_07({net988[0], net988[1], net988[2],
     net988[3], net988[4], net988[5], net988[6], net988[7]}),
     .slf_op_08({net987[0], net987[1], net987[2], net987[3], net987[4],
     net987[5], net987[6], net987[7]}), .rgt_op_08({net1082[0],
     net1082[1], net1082[2], net1082[3], net1082[4], net1082[5],
     net1082[6], net1082[7]}), .rgt_op_07({net1083[0], net1083[1],
     net1083[2], net1083[3], net1083[4], net1083[5], net1083[6],
     net1083[7]}), .rgt_op_06({net1084[0], net1084[1], net1084[2],
     net1084[3], net1084[4], net1084[5], net1084[6], net1084[7]}),
     .rgt_op_05({net1085[0], net1085[1], net1085[2], net1085[3],
     net1085[4], net1085[5], net1085[6], net1085[7]}),
     .lft_op_08({net836[0], net836[1], net836[2], net836[3], net836[4],
     net836[5], net836[6], net836[7]}), .lft_op_07({net831[0],
     net831[1], net831[2], net831[3], net831[4], net831[5], net831[6],
     net831[7]}), .lft_op_06({net832[0], net832[1], net832[2],
     net832[3], net832[4], net832[5], net832[6], net832[7]}),
     .lft_op_05({net833[0], net833[1], net833[2], net833[3], net833[4],
     net833[5], net833[6], net833[7]}), .sp12_h_l_08({net1001[0],
     net1001[1], net1001[2], net1001[3], net1001[4], net1001[5],
     net1001[6], net1001[7], net1001[8], net1001[9], net1001[10],
     net1001[11], net1001[12], net1001[13], net1001[14], net1001[15],
     net1001[16], net1001[17], net1001[18], net1001[19], net1001[20],
     net1001[21], net1001[22], net1001[23]}), .sp12_h_l_07({net1000[0],
     net1000[1], net1000[2], net1000[3], net1000[4], net1000[5],
     net1000[6], net1000[7], net1000[8], net1000[9], net1000[10],
     net1000[11], net1000[12], net1000[13], net1000[14], net1000[15],
     net1000[16], net1000[17], net1000[18], net1000[19], net1000[20],
     net1000[21], net1000[22], net1000[23]}), .sp12_h_l_06({net999[0],
     net999[1], net999[2], net999[3], net999[4], net999[5], net999[6],
     net999[7], net999[8], net999[9], net999[10], net999[11],
     net999[12], net999[13], net999[14], net999[15], net999[16],
     net999[17], net999[18], net999[19], net999[20], net999[21],
     net999[22], net999[23]}), .sp12_h_r_05({net1093[0], net1093[1],
     net1093[2], net1093[3], net1093[4], net1093[5], net1093[6],
     net1093[7], net1093[8], net1093[9], net1093[10], net1093[11],
     net1093[12], net1093[13], net1093[14], net1093[15], net1093[16],
     net1093[17], net1093[18], net1093[19], net1093[20], net1093[21],
     net1093[22], net1093[23]}), .sp12_h_r_06({net1094[0], net1094[1],
     net1094[2], net1094[3], net1094[4], net1094[5], net1094[6],
     net1094[7], net1094[8], net1094[9], net1094[10], net1094[11],
     net1094[12], net1094[13], net1094[14], net1094[15], net1094[16],
     net1094[17], net1094[18], net1094[19], net1094[20], net1094[21],
     net1094[22], net1094[23]}), .sp12_h_r_07({net1095[0], net1095[1],
     net1095[2], net1095[3], net1095[4], net1095[5], net1095[6],
     net1095[7], net1095[8], net1095[9], net1095[10], net1095[11],
     net1095[12], net1095[13], net1095[14], net1095[15], net1095[16],
     net1095[17], net1095[18], net1095[19], net1095[20], net1095[21],
     net1095[22], net1095[23]}), .sp12_h_r_08({net1096[0], net1096[1],
     net1096[2], net1096[3], net1096[4], net1096[5], net1096[6],
     net1096[7], net1096[8], net1096[9], net1096[10], net1096[11],
     net1096[12], net1096[13], net1096[14], net1096[15], net1096[16],
     net1096[17], net1096[18], net1096[19], net1096[20], net1096[21],
     net1096[22], net1096[23]}), .sp12_h_l_05({net998[0], net998[1],
     net998[2], net998[3], net998[4], net998[5], net998[6], net998[7],
     net998[8], net998[9], net998[10], net998[11], net998[12],
     net998[13], net998[14], net998[15], net998[16], net998[17],
     net998[18], net998[19], net998[20], net998[21], net998[22],
     net998[23]}), .sp4_r_v_b_05({net1098[0], net1098[1], net1098[2],
     net1098[3], net1098[4], net1098[5], net1098[6], net1098[7],
     net1098[8], net1098[9], net1098[10], net1098[11], net1098[12],
     net1098[13], net1098[14], net1098[15], net1098[16], net1098[17],
     net1098[18], net1098[19], net1098[20], net1098[21], net1098[22],
     net1098[23], net1098[24], net1098[25], net1098[26], net1098[27],
     net1098[28], net1098[29], net1098[30], net1098[31], net1098[32],
     net1098[33], net1098[34], net1098[35], net1098[36], net1098[37],
     net1098[38], net1098[39], net1098[40], net1098[41], net1098[42],
     net1098[43], net1098[44], net1098[45], net1098[46], net1098[47]}),
     .sp4_r_v_b_06({net1099[0], net1099[1], net1099[2], net1099[3],
     net1099[4], net1099[5], net1099[6], net1099[7], net1099[8],
     net1099[9], net1099[10], net1099[11], net1099[12], net1099[13],
     net1099[14], net1099[15], net1099[16], net1099[17], net1099[18],
     net1099[19], net1099[20], net1099[21], net1099[22], net1099[23],
     net1099[24], net1099[25], net1099[26], net1099[27], net1099[28],
     net1099[29], net1099[30], net1099[31], net1099[32], net1099[33],
     net1099[34], net1099[35], net1099[36], net1099[37], net1099[38],
     net1099[39], net1099[40], net1099[41], net1099[42], net1099[43],
     net1099[44], net1099[45], net1099[46], net1099[47]}),
     .sp4_r_v_b_07({net1100[0], net1100[1], net1100[2], net1100[3],
     net1100[4], net1100[5], net1100[6], net1100[7], net1100[8],
     net1100[9], net1100[10], net1100[11], net1100[12], net1100[13],
     net1100[14], net1100[15], net1100[16], net1100[17], net1100[18],
     net1100[19], net1100[20], net1100[21], net1100[22], net1100[23],
     net1100[24], net1100[25], net1100[26], net1100[27], net1100[28],
     net1100[29], net1100[30], net1100[31], net1100[32], net1100[33],
     net1100[34], net1100[35], net1100[36], net1100[37], net1100[38],
     net1100[39], net1100[40], net1100[41], net1100[42], net1100[43],
     net1100[44], net1100[45], net1100[46], net1100[47]}),
     .sp4_r_v_b_08({net1101[0], net1101[1], net1101[2], net1101[3],
     net1101[4], net1101[5], net1101[6], net1101[7], net1101[8],
     net1101[9], net1101[10], net1101[11], net1101[12], net1101[13],
     net1101[14], net1101[15], net1101[16], net1101[17], net1101[18],
     net1101[19], net1101[20], net1101[21], net1101[22], net1101[23],
     net1101[24], net1101[25], net1101[26], net1101[27], net1101[28],
     net1101[29], net1101[30], net1101[31], net1101[32], net1101[33],
     net1101[34], net1101[35], net1101[36], net1101[37], net1101[38],
     net1101[39], net1101[40], net1101[41], net1101[42], net1101[43],
     net1101[44], net1101[45], net1101[46], net1101[47]}),
     .sp4_v_b_08({net1006[0], net1006[1], net1006[2], net1006[3],
     net1006[4], net1006[5], net1006[6], net1006[7], net1006[8],
     net1006[9], net1006[10], net1006[11], net1006[12], net1006[13],
     net1006[14], net1006[15], net1006[16], net1006[17], net1006[18],
     net1006[19], net1006[20], net1006[21], net1006[22], net1006[23],
     net1006[24], net1006[25], net1006[26], net1006[27], net1006[28],
     net1006[29], net1006[30], net1006[31], net1006[32], net1006[33],
     net1006[34], net1006[35], net1006[36], net1006[37], net1006[38],
     net1006[39], net1006[40], net1006[41], net1006[42], net1006[43],
     net1006[44], net1006[45], net1006[46], net1006[47]}),
     .sp4_v_b_07({net1005[0], net1005[1], net1005[2], net1005[3],
     net1005[4], net1005[5], net1005[6], net1005[7], net1005[8],
     net1005[9], net1005[10], net1005[11], net1005[12], net1005[13],
     net1005[14], net1005[15], net1005[16], net1005[17], net1005[18],
     net1005[19], net1005[20], net1005[21], net1005[22], net1005[23],
     net1005[24], net1005[25], net1005[26], net1005[27], net1005[28],
     net1005[29], net1005[30], net1005[31], net1005[32], net1005[33],
     net1005[34], net1005[35], net1005[36], net1005[37], net1005[38],
     net1005[39], net1005[40], net1005[41], net1005[42], net1005[43],
     net1005[44], net1005[45], net1005[46], net1005[47]}),
     .sp4_v_b_06({net1004[0], net1004[1], net1004[2], net1004[3],
     net1004[4], net1004[5], net1004[6], net1004[7], net1004[8],
     net1004[9], net1004[10], net1004[11], net1004[12], net1004[13],
     net1004[14], net1004[15], net1004[16], net1004[17], net1004[18],
     net1004[19], net1004[20], net1004[21], net1004[22], net1004[23],
     net1004[24], net1004[25], net1004[26], net1004[27], net1004[28],
     net1004[29], net1004[30], net1004[31], net1004[32], net1004[33],
     net1004[34], net1004[35], net1004[36], net1004[37], net1004[38],
     net1004[39], net1004[40], net1004[41], net1004[42], net1004[43],
     net1004[44], net1004[45], net1004[46], net1004[47]}),
     .sp4_v_b_05({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7], net1003[8],
     net1003[9], net1003[10], net1003[11], net1003[12], net1003[13],
     net1003[14], net1003[15], net1003[16], net1003[17], net1003[18],
     net1003[19], net1003[20], net1003[21], net1003[22], net1003[23],
     net1003[24], net1003[25], net1003[26], net1003[27], net1003[28],
     net1003[29], net1003[30], net1003[31], net1003[32], net1003[33],
     net1003[34], net1003[35], net1003[36], net1003[37], net1003[38],
     net1003[39], net1003[40], net1003[41], net1003[42], net1003[43],
     net1003[44], net1003[45], net1003[46], net1003[47]}),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .wl(wl_l[127:0]), .sp12_v_t_08({net1109[0], net1109[1],
     net1109[2], net1109[3], net1109[4], net1109[5], net1109[6],
     net1109[7], net1109[8], net1109[9], net1109[10], net1109[11],
     net1109[12], net1109[13], net1109[14], net1109[15], net1109[16],
     net1109[17], net1109[18], net1109[19], net1109[20], net1109[21],
     net1109[22], net1109[23]}), .tnr_op_08({slf_op_08_17[3],
     slf_op_08_17[2], slf_op_08_17[1], slf_op_08_17[0],
     slf_op_08_17[3], slf_op_08_17[2], slf_op_08_17[1],
     slf_op_08_17[0]}), .top_op_08({slf_op_02_17[3], slf_op_02_17[2],
     slf_op_02_17[1], slf_op_02_17[0], slf_op_02_17[3],
     slf_op_02_17[2], slf_op_02_17[1], slf_op_02_17[0]}),
     .tnl_op_08({slf_op_01_17[3], slf_op_01_17[2], slf_op_01_17[1],
     slf_op_01_17[0], slf_op_01_17[3], slf_op_01_17[2],
     slf_op_01_17[1], slf_op_01_17[0]}), .sp4_v_t_08({net1113[0],
     net1113[1], net1113[2], net1113[3], net1113[4], net1113[5],
     net1113[6], net1113[7], net1113[8], net1113[9], net1113[10],
     net1113[11], net1113[12], net1113[13], net1113[14], net1113[15],
     net1113[16], net1113[17], net1113[18], net1113[19], net1113[20],
     net1113[21], net1113[22], net1113[23], net1113[24], net1113[25],
     net1113[26], net1113[27], net1113[28], net1113[29], net1113[30],
     net1113[31], net1113[32], net1113[33], net1113[34], net1113[35],
     net1113[36], net1113[37], net1113[38], net1113[39], net1113[40],
     net1113[41], net1113[42], net1113[43], net1113[44], net1113[45],
     net1113[46], net1113[47]}), .lc_bot(lc_bot_02_09),
     .op_vic(net1458), .sp12_v_b_01(sp12_v_b_02_09[23:0]),
     .glb_netwk_t({net1117[0], net1117[1], net1117[2], net1117[3],
     net1117[4], net1117[5], net1117[6], net1117[7]}));
lt_1x8_top_ice1f I_lt_col_t05 ( .glb_netwk_b({net1118[0], net1118[1],
     net1118[2], net1118[3], net1118[4], net1118[5], net1118[6],
     net1118[7]}), .rgt_op_03(slf_op_06_11[7:0]),
     .slf_op_02({net1216[0], net1216[1], net1216[2], net1216[3],
     net1216[4], net1216[5], net1216[6], net1216[7]}),
     .rgt_op_02(slf_op_06_10[7:0]), .rgt_op_01(slf_op_06_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04({net771[0], net771[1],
     net771[2], net771[3], net771[4], net771[5], net771[6],
     net771[7]}), .lft_op_03({net772[0], net772[1], net772[2],
     net772[3], net772[4], net772[5], net772[6], net772[7]}),
     .lft_op_02({net773[0], net773[1], net773[2], net773[3], net773[4],
     net773[5], net773[6], net773[7]}), .lft_op_01(slf_op_04_09[7:0]),
     .rgt_op_04(slf_op_06_12[7:0]), .carry_in(carry_in_05_09),
     .bnl_op_01(bnl_op_05_09[7:0]), .slf_op_04({net1224[0], net1224[1],
     net1224[2], net1224[3], net1224[4], net1224[5], net1224[6],
     net1224[7]}), .slf_op_03({net1214[0], net1214[1], net1214[2],
     net1214[3], net1214[4], net1214[5], net1214[6], net1214[7]}),
     .slf_op_01(slf_op_05_09[7:0]), .sp4_h_l_04({net1243[0],
     net1243[1], net1243[2], net1243[3], net1243[4], net1243[5],
     net1243[6], net1243[7], net1243[8], net1243[9], net1243[10],
     net1243[11], net1243[12], net1243[13], net1243[14], net1243[15],
     net1243[16], net1243[17], net1243[18], net1243[19], net1243[20],
     net1243[21], net1243[22], net1243[23], net1243[24], net1243[25],
     net1243[26], net1243[27], net1243[28], net1243[29], net1243[30],
     net1243[31], net1243[32], net1243[33], net1243[34], net1243[35],
     net1243[36], net1243[37], net1243[38], net1243[39], net1243[40],
     net1243[41], net1243[42], net1243[43], net1243[44], net1243[45],
     net1243[46], net1243[47]}), .carry_out(net1136),
     .vdd_cntl(vdd_cntl_l[127:0]), .sp12_h_r_04({net1138[0],
     net1138[1], net1138[2], net1138[3], net1138[4], net1138[5],
     net1138[6], net1138[7], net1138[8], net1138[9], net1138[10],
     net1138[11], net1138[12], net1138[13], net1138[14], net1138[15],
     net1138[16], net1138[17], net1138[18], net1138[19], net1138[20],
     net1138[21], net1138[22], net1138[23]}), .sp12_h_r_03({net1139[0],
     net1139[1], net1139[2], net1139[3], net1139[4], net1139[5],
     net1139[6], net1139[7], net1139[8], net1139[9], net1139[10],
     net1139[11], net1139[12], net1139[13], net1139[14], net1139[15],
     net1139[16], net1139[17], net1139[18], net1139[19], net1139[20],
     net1139[21], net1139[22], net1139[23]}), .sp12_h_r_02({net1140[0],
     net1140[1], net1140[2], net1140[3], net1140[4], net1140[5],
     net1140[6], net1140[7], net1140[8], net1140[9], net1140[10],
     net1140[11], net1140[12], net1140[13], net1140[14], net1140[15],
     net1140[16], net1140[17], net1140[18], net1140[19], net1140[20],
     net1140[21], net1140[22], net1140[23]}), .sp12_h_r_01({net1141[0],
     net1141[1], net1141[2], net1141[3], net1141[4], net1141[5],
     net1141[6], net1141[7], net1141[8], net1141[9], net1141[10],
     net1141[11], net1141[12], net1141[13], net1141[14], net1141[15],
     net1141[16], net1141[17], net1141[18], net1141[19], net1141[20],
     net1141[21], net1141[22], net1141[23]}),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_05_09[47:0]), .sp4_r_v_b_04({net1144[0],
     net1144[1], net1144[2], net1144[3], net1144[4], net1144[5],
     net1144[6], net1144[7], net1144[8], net1144[9], net1144[10],
     net1144[11], net1144[12], net1144[13], net1144[14], net1144[15],
     net1144[16], net1144[17], net1144[18], net1144[19], net1144[20],
     net1144[21], net1144[22], net1144[23], net1144[24], net1144[25],
     net1144[26], net1144[27], net1144[28], net1144[29], net1144[30],
     net1144[31], net1144[32], net1144[33], net1144[34], net1144[35],
     net1144[36], net1144[37], net1144[38], net1144[39], net1144[40],
     net1144[41], net1144[42], net1144[43], net1144[44], net1144[45],
     net1144[46], net1144[47]}), .sp4_r_v_b_03({net1145[0], net1145[1],
     net1145[2], net1145[3], net1145[4], net1145[5], net1145[6],
     net1145[7], net1145[8], net1145[9], net1145[10], net1145[11],
     net1145[12], net1145[13], net1145[14], net1145[15], net1145[16],
     net1145[17], net1145[18], net1145[19], net1145[20], net1145[21],
     net1145[22], net1145[23], net1145[24], net1145[25], net1145[26],
     net1145[27], net1145[28], net1145[29], net1145[30], net1145[31],
     net1145[32], net1145[33], net1145[34], net1145[35], net1145[36],
     net1145[37], net1145[38], net1145[39], net1145[40], net1145[41],
     net1145[42], net1145[43], net1145[44], net1145[45], net1145[46],
     net1145[47]}), .sp4_r_v_b_02({net1146[0], net1146[1], net1146[2],
     net1146[3], net1146[4], net1146[5], net1146[6], net1146[7],
     net1146[8], net1146[9], net1146[10], net1146[11], net1146[12],
     net1146[13], net1146[14], net1146[15], net1146[16], net1146[17],
     net1146[18], net1146[19], net1146[20], net1146[21], net1146[22],
     net1146[23], net1146[24], net1146[25], net1146[26], net1146[27],
     net1146[28], net1146[29], net1146[30], net1146[31], net1146[32],
     net1146[33], net1146[34], net1146[35], net1146[36], net1146[37],
     net1146[38], net1146[39], net1146[40], net1146[41], net1146[42],
     net1146[43], net1146[44], net1146[45], net1146[46], net1146[47]}),
     .sp4_r_v_b_01(sp4_v_b_06_09[47:0]), .sp4_h_r_04({net1148[0],
     net1148[1], net1148[2], net1148[3], net1148[4], net1148[5],
     net1148[6], net1148[7], net1148[8], net1148[9], net1148[10],
     net1148[11], net1148[12], net1148[13], net1148[14], net1148[15],
     net1148[16], net1148[17], net1148[18], net1148[19], net1148[20],
     net1148[21], net1148[22], net1148[23], net1148[24], net1148[25],
     net1148[26], net1148[27], net1148[28], net1148[29], net1148[30],
     net1148[31], net1148[32], net1148[33], net1148[34], net1148[35],
     net1148[36], net1148[37], net1148[38], net1148[39], net1148[40],
     net1148[41], net1148[42], net1148[43], net1148[44], net1148[45],
     net1148[46], net1148[47]}), .sp4_h_r_03({net1149[0], net1149[1],
     net1149[2], net1149[3], net1149[4], net1149[5], net1149[6],
     net1149[7], net1149[8], net1149[9], net1149[10], net1149[11],
     net1149[12], net1149[13], net1149[14], net1149[15], net1149[16],
     net1149[17], net1149[18], net1149[19], net1149[20], net1149[21],
     net1149[22], net1149[23], net1149[24], net1149[25], net1149[26],
     net1149[27], net1149[28], net1149[29], net1149[30], net1149[31],
     net1149[32], net1149[33], net1149[34], net1149[35], net1149[36],
     net1149[37], net1149[38], net1149[39], net1149[40], net1149[41],
     net1149[42], net1149[43], net1149[44], net1149[45], net1149[46],
     net1149[47]}), .sp4_h_r_02({net1150[0], net1150[1], net1150[2],
     net1150[3], net1150[4], net1150[5], net1150[6], net1150[7],
     net1150[8], net1150[9], net1150[10], net1150[11], net1150[12],
     net1150[13], net1150[14], net1150[15], net1150[16], net1150[17],
     net1150[18], net1150[19], net1150[20], net1150[21], net1150[22],
     net1150[23], net1150[24], net1150[25], net1150[26], net1150[27],
     net1150[28], net1150[29], net1150[30], net1150[31], net1150[32],
     net1150[33], net1150[34], net1150[35], net1150[36], net1150[37],
     net1150[38], net1150[39], net1150[40], net1150[41], net1150[42],
     net1150[43], net1150[44], net1150[45], net1150[46], net1150[47]}),
     .sp4_h_r_01({net1151[0], net1151[1], net1151[2], net1151[3],
     net1151[4], net1151[5], net1151[6], net1151[7], net1151[8],
     net1151[9], net1151[10], net1151[11], net1151[12], net1151[13],
     net1151[14], net1151[15], net1151[16], net1151[17], net1151[18],
     net1151[19], net1151[20], net1151[21], net1151[22], net1151[23],
     net1151[24], net1151[25], net1151[26], net1151[27], net1151[28],
     net1151[29], net1151[30], net1151[31], net1151[32], net1151[33],
     net1151[34], net1151[35], net1151[36], net1151[37], net1151[38],
     net1151[39], net1151[40], net1151[41], net1151[42], net1151[43],
     net1151[44], net1151[45], net1151[46], net1151[47]}),
     .sp4_h_l_03({net1244[0], net1244[1], net1244[2], net1244[3],
     net1244[4], net1244[5], net1244[6], net1244[7], net1244[8],
     net1244[9], net1244[10], net1244[11], net1244[12], net1244[13],
     net1244[14], net1244[15], net1244[16], net1244[17], net1244[18],
     net1244[19], net1244[20], net1244[21], net1244[22], net1244[23],
     net1244[24], net1244[25], net1244[26], net1244[27], net1244[28],
     net1244[29], net1244[30], net1244[31], net1244[32], net1244[33],
     net1244[34], net1244[35], net1244[36], net1244[37], net1244[38],
     net1244[39], net1244[40], net1244[41], net1244[42], net1244[43],
     net1244[44], net1244[45], net1244[46], net1244[47]}),
     .sp4_h_l_02({net1245[0], net1245[1], net1245[2], net1245[3],
     net1245[4], net1245[5], net1245[6], net1245[7], net1245[8],
     net1245[9], net1245[10], net1245[11], net1245[12], net1245[13],
     net1245[14], net1245[15], net1245[16], net1245[17], net1245[18],
     net1245[19], net1245[20], net1245[21], net1245[22], net1245[23],
     net1245[24], net1245[25], net1245[26], net1245[27], net1245[28],
     net1245[29], net1245[30], net1245[31], net1245[32], net1245[33],
     net1245[34], net1245[35], net1245[36], net1245[37], net1245[38],
     net1245[39], net1245[40], net1245[41], net1245[42], net1245[43],
     net1245[44], net1245[45], net1245[46], net1245[47]}),
     .sp4_h_l_01({net1246[0], net1246[1], net1246[2], net1246[3],
     net1246[4], net1246[5], net1246[6], net1246[7], net1246[8],
     net1246[9], net1246[10], net1246[11], net1246[12], net1246[13],
     net1246[14], net1246[15], net1246[16], net1246[17], net1246[18],
     net1246[19], net1246[20], net1246[21], net1246[22], net1246[23],
     net1246[24], net1246[25], net1246[26], net1246[27], net1246[28],
     net1246[29], net1246[30], net1246[31], net1246[32], net1246[33],
     net1246[34], net1246[35], net1246[36], net1246[37], net1246[38],
     net1246[39], net1246[40], net1246[41], net1246[42], net1246[43],
     net1246[44], net1246[45], net1246[46], net1246[47]}),
     .bl(bl[275:222]), .bot_op_01(bot_op_05_09[7:0]),
     .sp12_h_l_01({net1236[0], net1236[1], net1236[2], net1236[3],
     net1236[4], net1236[5], net1236[6], net1236[7], net1236[8],
     net1236[9], net1236[10], net1236[11], net1236[12], net1236[13],
     net1236[14], net1236[15], net1236[16], net1236[17], net1236[18],
     net1236[19], net1236[20], net1236[21], net1236[22], net1236[23]}),
     .sp12_h_l_02({net1235[0], net1235[1], net1235[2], net1235[3],
     net1235[4], net1235[5], net1235[6], net1235[7], net1235[8],
     net1235[9], net1235[10], net1235[11], net1235[12], net1235[13],
     net1235[14], net1235[15], net1235[16], net1235[17], net1235[18],
     net1235[19], net1235[20], net1235[21], net1235[22], net1235[23]}),
     .sp12_h_l_03({net1234[0], net1234[1], net1234[2], net1234[3],
     net1234[4], net1234[5], net1234[6], net1234[7], net1234[8],
     net1234[9], net1234[10], net1234[11], net1234[12], net1234[13],
     net1234[14], net1234[15], net1234[16], net1234[17], net1234[18],
     net1234[19], net1234[20], net1234[21], net1234[22], net1234[23]}),
     .sp12_h_l_04({net1233[0], net1233[1], net1233[2], net1233[3],
     net1233[4], net1233[5], net1233[6], net1233[7], net1233[8],
     net1233[9], net1233[10], net1233[11], net1233[12], net1233[13],
     net1233[14], net1233[15], net1233[16], net1233[17], net1233[18],
     net1233[19], net1233[20], net1233[21], net1233[22], net1233[23]}),
     .sp4_v_b_04({net1239[0], net1239[1], net1239[2], net1239[3],
     net1239[4], net1239[5], net1239[6], net1239[7], net1239[8],
     net1239[9], net1239[10], net1239[11], net1239[12], net1239[13],
     net1239[14], net1239[15], net1239[16], net1239[17], net1239[18],
     net1239[19], net1239[20], net1239[21], net1239[22], net1239[23],
     net1239[24], net1239[25], net1239[26], net1239[27], net1239[28],
     net1239[29], net1239[30], net1239[31], net1239[32], net1239[33],
     net1239[34], net1239[35], net1239[36], net1239[37], net1239[38],
     net1239[39], net1239[40], net1239[41], net1239[42], net1239[43],
     net1239[44], net1239[45], net1239[46], net1239[47]}),
     .sp4_v_b_03({net1240[0], net1240[1], net1240[2], net1240[3],
     net1240[4], net1240[5], net1240[6], net1240[7], net1240[8],
     net1240[9], net1240[10], net1240[11], net1240[12], net1240[13],
     net1240[14], net1240[15], net1240[16], net1240[17], net1240[18],
     net1240[19], net1240[20], net1240[21], net1240[22], net1240[23],
     net1240[24], net1240[25], net1240[26], net1240[27], net1240[28],
     net1240[29], net1240[30], net1240[31], net1240[32], net1240[33],
     net1240[34], net1240[35], net1240[36], net1240[37], net1240[38],
     net1240[39], net1240[40], net1240[41], net1240[42], net1240[43],
     net1240[44], net1240[45], net1240[46], net1240[47]}),
     .sp4_v_b_02({net1241[0], net1241[1], net1241[2], net1241[3],
     net1241[4], net1241[5], net1241[6], net1241[7], net1241[8],
     net1241[9], net1241[10], net1241[11], net1241[12], net1241[13],
     net1241[14], net1241[15], net1241[16], net1241[17], net1241[18],
     net1241[19], net1241[20], net1241[21], net1241[22], net1241[23],
     net1241[24], net1241[25], net1241[26], net1241[27], net1241[28],
     net1241[29], net1241[30], net1241[31], net1241[32], net1241[33],
     net1241[34], net1241[35], net1241[36], net1241[37], net1241[38],
     net1241[39], net1241[40], net1241[41], net1241[42], net1241[43],
     net1241[44], net1241[45], net1241[46], net1241[47]}),
     .bnr_op_01(bnr_op_05_09[7:0]), .sp4_h_l_05({net1267[0],
     net1267[1], net1267[2], net1267[3], net1267[4], net1267[5],
     net1267[6], net1267[7], net1267[8], net1267[9], net1267[10],
     net1267[11], net1267[12], net1267[13], net1267[14], net1267[15],
     net1267[16], net1267[17], net1267[18], net1267[19], net1267[20],
     net1267[21], net1267[22], net1267[23], net1267[24], net1267[25],
     net1267[26], net1267[27], net1267[28], net1267[29], net1267[30],
     net1267[31], net1267[32], net1267[33], net1267[34], net1267[35],
     net1267[36], net1267[37], net1267[38], net1267[39], net1267[40],
     net1267[41], net1267[42], net1267[43], net1267[44], net1267[45],
     net1267[46], net1267[47]}), .sp4_h_l_06({net1266[0], net1266[1],
     net1266[2], net1266[3], net1266[4], net1266[5], net1266[6],
     net1266[7], net1266[8], net1266[9], net1266[10], net1266[11],
     net1266[12], net1266[13], net1266[14], net1266[15], net1266[16],
     net1266[17], net1266[18], net1266[19], net1266[20], net1266[21],
     net1266[22], net1266[23], net1266[24], net1266[25], net1266[26],
     net1266[27], net1266[28], net1266[29], net1266[30], net1266[31],
     net1266[32], net1266[33], net1266[34], net1266[35], net1266[36],
     net1266[37], net1266[38], net1266[39], net1266[40], net1266[41],
     net1266[42], net1266[43], net1266[44], net1266[45], net1266[46],
     net1266[47]}), .sp4_h_l_07({net1265[0], net1265[1], net1265[2],
     net1265[3], net1265[4], net1265[5], net1265[6], net1265[7],
     net1265[8], net1265[9], net1265[10], net1265[11], net1265[12],
     net1265[13], net1265[14], net1265[15], net1265[16], net1265[17],
     net1265[18], net1265[19], net1265[20], net1265[21], net1265[22],
     net1265[23], net1265[24], net1265[25], net1265[26], net1265[27],
     net1265[28], net1265[29], net1265[30], net1265[31], net1265[32],
     net1265[33], net1265[34], net1265[35], net1265[36], net1265[37],
     net1265[38], net1265[39], net1265[40], net1265[41], net1265[42],
     net1265[43], net1265[44], net1265[45], net1265[46], net1265[47]}),
     .sp4_h_l_08({net1264[0], net1264[1], net1264[2], net1264[3],
     net1264[4], net1264[5], net1264[6], net1264[7], net1264[8],
     net1264[9], net1264[10], net1264[11], net1264[12], net1264[13],
     net1264[14], net1264[15], net1264[16], net1264[17], net1264[18],
     net1264[19], net1264[20], net1264[21], net1264[22], net1264[23],
     net1264[24], net1264[25], net1264[26], net1264[27], net1264[28],
     net1264[29], net1264[30], net1264[31], net1264[32], net1264[33],
     net1264[34], net1264[35], net1264[36], net1264[37], net1264[38],
     net1264[39], net1264[40], net1264[41], net1264[42], net1264[43],
     net1264[44], net1264[45], net1264[46], net1264[47]}),
     .sp4_h_r_08({net1169[0], net1169[1], net1169[2], net1169[3],
     net1169[4], net1169[5], net1169[6], net1169[7], net1169[8],
     net1169[9], net1169[10], net1169[11], net1169[12], net1169[13],
     net1169[14], net1169[15], net1169[16], net1169[17], net1169[18],
     net1169[19], net1169[20], net1169[21], net1169[22], net1169[23],
     net1169[24], net1169[25], net1169[26], net1169[27], net1169[28],
     net1169[29], net1169[30], net1169[31], net1169[32], net1169[33],
     net1169[34], net1169[35], net1169[36], net1169[37], net1169[38],
     net1169[39], net1169[40], net1169[41], net1169[42], net1169[43],
     net1169[44], net1169[45], net1169[46], net1169[47]}),
     .sp4_h_r_07({net1170[0], net1170[1], net1170[2], net1170[3],
     net1170[4], net1170[5], net1170[6], net1170[7], net1170[8],
     net1170[9], net1170[10], net1170[11], net1170[12], net1170[13],
     net1170[14], net1170[15], net1170[16], net1170[17], net1170[18],
     net1170[19], net1170[20], net1170[21], net1170[22], net1170[23],
     net1170[24], net1170[25], net1170[26], net1170[27], net1170[28],
     net1170[29], net1170[30], net1170[31], net1170[32], net1170[33],
     net1170[34], net1170[35], net1170[36], net1170[37], net1170[38],
     net1170[39], net1170[40], net1170[41], net1170[42], net1170[43],
     net1170[44], net1170[45], net1170[46], net1170[47]}),
     .sp4_h_r_06({net1171[0], net1171[1], net1171[2], net1171[3],
     net1171[4], net1171[5], net1171[6], net1171[7], net1171[8],
     net1171[9], net1171[10], net1171[11], net1171[12], net1171[13],
     net1171[14], net1171[15], net1171[16], net1171[17], net1171[18],
     net1171[19], net1171[20], net1171[21], net1171[22], net1171[23],
     net1171[24], net1171[25], net1171[26], net1171[27], net1171[28],
     net1171[29], net1171[30], net1171[31], net1171[32], net1171[33],
     net1171[34], net1171[35], net1171[36], net1171[37], net1171[38],
     net1171[39], net1171[40], net1171[41], net1171[42], net1171[43],
     net1171[44], net1171[45], net1171[46], net1171[47]}),
     .sp4_h_r_05({net1172[0], net1172[1], net1172[2], net1172[3],
     net1172[4], net1172[5], net1172[6], net1172[7], net1172[8],
     net1172[9], net1172[10], net1172[11], net1172[12], net1172[13],
     net1172[14], net1172[15], net1172[16], net1172[17], net1172[18],
     net1172[19], net1172[20], net1172[21], net1172[22], net1172[23],
     net1172[24], net1172[25], net1172[26], net1172[27], net1172[28],
     net1172[29], net1172[30], net1172[31], net1172[32], net1172[33],
     net1172[34], net1172[35], net1172[36], net1172[37], net1172[38],
     net1172[39], net1172[40], net1172[41], net1172[42], net1172[43],
     net1172[44], net1172[45], net1172[46], net1172[47]}),
     .slf_op_05({net1275[0], net1275[1], net1275[2], net1275[3],
     net1275[4], net1275[5], net1275[6], net1275[7]}),
     .slf_op_06({net1274[0], net1274[1], net1274[2], net1274[3],
     net1274[4], net1274[5], net1274[6], net1274[7]}),
     .slf_op_07({net1273[0], net1273[1], net1273[2], net1273[3],
     net1273[4], net1273[5], net1273[6], net1273[7]}),
     .slf_op_08({net1272[0], net1272[1], net1272[2], net1272[3],
     net1272[4], net1272[5], net1272[6], net1272[7]}),
     .rgt_op_08(slf_op_06_16[7:0]), .rgt_op_07(slf_op_06_15[7:0]),
     .rgt_op_06(slf_op_06_14[7:0]), .rgt_op_05(slf_op_06_13[7:0]),
     .lft_op_08({net767[0], net767[1], net767[2], net767[3], net767[4],
     net767[5], net767[6], net767[7]}), .lft_op_07({net768[0],
     net768[1], net768[2], net768[3], net768[4], net768[5], net768[6],
     net768[7]}), .lft_op_06({net769[0], net769[1], net769[2],
     net769[3], net769[4], net769[5], net769[6], net769[7]}),
     .lft_op_05({net770[0], net770[1], net770[2], net770[3], net770[4],
     net770[5], net770[6], net770[7]}), .sp12_h_l_08({net1286[0],
     net1286[1], net1286[2], net1286[3], net1286[4], net1286[5],
     net1286[6], net1286[7], net1286[8], net1286[9], net1286[10],
     net1286[11], net1286[12], net1286[13], net1286[14], net1286[15],
     net1286[16], net1286[17], net1286[18], net1286[19], net1286[20],
     net1286[21], net1286[22], net1286[23]}), .sp12_h_l_07({net1285[0],
     net1285[1], net1285[2], net1285[3], net1285[4], net1285[5],
     net1285[6], net1285[7], net1285[8], net1285[9], net1285[10],
     net1285[11], net1285[12], net1285[13], net1285[14], net1285[15],
     net1285[16], net1285[17], net1285[18], net1285[19], net1285[20],
     net1285[21], net1285[22], net1285[23]}), .sp12_h_l_06({net1284[0],
     net1284[1], net1284[2], net1284[3], net1284[4], net1284[5],
     net1284[6], net1284[7], net1284[8], net1284[9], net1284[10],
     net1284[11], net1284[12], net1284[13], net1284[14], net1284[15],
     net1284[16], net1284[17], net1284[18], net1284[19], net1284[20],
     net1284[21], net1284[22], net1284[23]}), .sp12_h_r_05({net1188[0],
     net1188[1], net1188[2], net1188[3], net1188[4], net1188[5],
     net1188[6], net1188[7], net1188[8], net1188[9], net1188[10],
     net1188[11], net1188[12], net1188[13], net1188[14], net1188[15],
     net1188[16], net1188[17], net1188[18], net1188[19], net1188[20],
     net1188[21], net1188[22], net1188[23]}), .sp12_h_r_06({net1189[0],
     net1189[1], net1189[2], net1189[3], net1189[4], net1189[5],
     net1189[6], net1189[7], net1189[8], net1189[9], net1189[10],
     net1189[11], net1189[12], net1189[13], net1189[14], net1189[15],
     net1189[16], net1189[17], net1189[18], net1189[19], net1189[20],
     net1189[21], net1189[22], net1189[23]}), .sp12_h_r_07({net1190[0],
     net1190[1], net1190[2], net1190[3], net1190[4], net1190[5],
     net1190[6], net1190[7], net1190[8], net1190[9], net1190[10],
     net1190[11], net1190[12], net1190[13], net1190[14], net1190[15],
     net1190[16], net1190[17], net1190[18], net1190[19], net1190[20],
     net1190[21], net1190[22], net1190[23]}), .sp12_h_r_08({net1191[0],
     net1191[1], net1191[2], net1191[3], net1191[4], net1191[5],
     net1191[6], net1191[7], net1191[8], net1191[9], net1191[10],
     net1191[11], net1191[12], net1191[13], net1191[14], net1191[15],
     net1191[16], net1191[17], net1191[18], net1191[19], net1191[20],
     net1191[21], net1191[22], net1191[23]}), .sp12_h_l_05({net1283[0],
     net1283[1], net1283[2], net1283[3], net1283[4], net1283[5],
     net1283[6], net1283[7], net1283[8], net1283[9], net1283[10],
     net1283[11], net1283[12], net1283[13], net1283[14], net1283[15],
     net1283[16], net1283[17], net1283[18], net1283[19], net1283[20],
     net1283[21], net1283[22], net1283[23]}),
     .sp4_r_v_b_05({net1193[0], net1193[1], net1193[2], net1193[3],
     net1193[4], net1193[5], net1193[6], net1193[7], net1193[8],
     net1193[9], net1193[10], net1193[11], net1193[12], net1193[13],
     net1193[14], net1193[15], net1193[16], net1193[17], net1193[18],
     net1193[19], net1193[20], net1193[21], net1193[22], net1193[23],
     net1193[24], net1193[25], net1193[26], net1193[27], net1193[28],
     net1193[29], net1193[30], net1193[31], net1193[32], net1193[33],
     net1193[34], net1193[35], net1193[36], net1193[37], net1193[38],
     net1193[39], net1193[40], net1193[41], net1193[42], net1193[43],
     net1193[44], net1193[45], net1193[46], net1193[47]}),
     .sp4_r_v_b_06({net1194[0], net1194[1], net1194[2], net1194[3],
     net1194[4], net1194[5], net1194[6], net1194[7], net1194[8],
     net1194[9], net1194[10], net1194[11], net1194[12], net1194[13],
     net1194[14], net1194[15], net1194[16], net1194[17], net1194[18],
     net1194[19], net1194[20], net1194[21], net1194[22], net1194[23],
     net1194[24], net1194[25], net1194[26], net1194[27], net1194[28],
     net1194[29], net1194[30], net1194[31], net1194[32], net1194[33],
     net1194[34], net1194[35], net1194[36], net1194[37], net1194[38],
     net1194[39], net1194[40], net1194[41], net1194[42], net1194[43],
     net1194[44], net1194[45], net1194[46], net1194[47]}),
     .sp4_r_v_b_07({net1195[0], net1195[1], net1195[2], net1195[3],
     net1195[4], net1195[5], net1195[6], net1195[7], net1195[8],
     net1195[9], net1195[10], net1195[11], net1195[12], net1195[13],
     net1195[14], net1195[15], net1195[16], net1195[17], net1195[18],
     net1195[19], net1195[20], net1195[21], net1195[22], net1195[23],
     net1195[24], net1195[25], net1195[26], net1195[27], net1195[28],
     net1195[29], net1195[30], net1195[31], net1195[32], net1195[33],
     net1195[34], net1195[35], net1195[36], net1195[37], net1195[38],
     net1195[39], net1195[40], net1195[41], net1195[42], net1195[43],
     net1195[44], net1195[45], net1195[46], net1195[47]}),
     .sp4_r_v_b_08({net1196[0], net1196[1], net1196[2], net1196[3],
     net1196[4], net1196[5], net1196[6], net1196[7], net1196[8],
     net1196[9], net1196[10], net1196[11], net1196[12], net1196[13],
     net1196[14], net1196[15], net1196[16], net1196[17], net1196[18],
     net1196[19], net1196[20], net1196[21], net1196[22], net1196[23],
     net1196[24], net1196[25], net1196[26], net1196[27], net1196[28],
     net1196[29], net1196[30], net1196[31], net1196[32], net1196[33],
     net1196[34], net1196[35], net1196[36], net1196[37], net1196[38],
     net1196[39], net1196[40], net1196[41], net1196[42], net1196[43],
     net1196[44], net1196[45], net1196[46], net1196[47]}),
     .sp4_v_b_08({net1291[0], net1291[1], net1291[2], net1291[3],
     net1291[4], net1291[5], net1291[6], net1291[7], net1291[8],
     net1291[9], net1291[10], net1291[11], net1291[12], net1291[13],
     net1291[14], net1291[15], net1291[16], net1291[17], net1291[18],
     net1291[19], net1291[20], net1291[21], net1291[22], net1291[23],
     net1291[24], net1291[25], net1291[26], net1291[27], net1291[28],
     net1291[29], net1291[30], net1291[31], net1291[32], net1291[33],
     net1291[34], net1291[35], net1291[36], net1291[37], net1291[38],
     net1291[39], net1291[40], net1291[41], net1291[42], net1291[43],
     net1291[44], net1291[45], net1291[46], net1291[47]}),
     .sp4_v_b_07({net1290[0], net1290[1], net1290[2], net1290[3],
     net1290[4], net1290[5], net1290[6], net1290[7], net1290[8],
     net1290[9], net1290[10], net1290[11], net1290[12], net1290[13],
     net1290[14], net1290[15], net1290[16], net1290[17], net1290[18],
     net1290[19], net1290[20], net1290[21], net1290[22], net1290[23],
     net1290[24], net1290[25], net1290[26], net1290[27], net1290[28],
     net1290[29], net1290[30], net1290[31], net1290[32], net1290[33],
     net1290[34], net1290[35], net1290[36], net1290[37], net1290[38],
     net1290[39], net1290[40], net1290[41], net1290[42], net1290[43],
     net1290[44], net1290[45], net1290[46], net1290[47]}),
     .sp4_v_b_06({net1289[0], net1289[1], net1289[2], net1289[3],
     net1289[4], net1289[5], net1289[6], net1289[7], net1289[8],
     net1289[9], net1289[10], net1289[11], net1289[12], net1289[13],
     net1289[14], net1289[15], net1289[16], net1289[17], net1289[18],
     net1289[19], net1289[20], net1289[21], net1289[22], net1289[23],
     net1289[24], net1289[25], net1289[26], net1289[27], net1289[28],
     net1289[29], net1289[30], net1289[31], net1289[32], net1289[33],
     net1289[34], net1289[35], net1289[36], net1289[37], net1289[38],
     net1289[39], net1289[40], net1289[41], net1289[42], net1289[43],
     net1289[44], net1289[45], net1289[46], net1289[47]}),
     .sp4_v_b_05({net1288[0], net1288[1], net1288[2], net1288[3],
     net1288[4], net1288[5], net1288[6], net1288[7], net1288[8],
     net1288[9], net1288[10], net1288[11], net1288[12], net1288[13],
     net1288[14], net1288[15], net1288[16], net1288[17], net1288[18],
     net1288[19], net1288[20], net1288[21], net1288[22], net1288[23],
     net1288[24], net1288[25], net1288[26], net1288[27], net1288[28],
     net1288[29], net1288[30], net1288[31], net1288[32], net1288[33],
     net1288[34], net1288[35], net1288[36], net1288[37], net1288[38],
     net1288[39], net1288[40], net1288[41], net1288[42], net1288[43],
     net1288[44], net1288[45], net1288[46], net1288[47]}),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .wl(wl_l[127:0]), .sp12_v_t_08({net1204[0], net1204[1],
     net1204[2], net1204[3], net1204[4], net1204[5], net1204[6],
     net1204[7], net1204[8], net1204[9], net1204[10], net1204[11],
     net1204[12], net1204[13], net1204[14], net1204[15], net1204[16],
     net1204[17], net1204[18], net1204[19], net1204[20], net1204[21],
     net1204[22], net1204[23]}), .tnr_op_08({slf_op_06_17[3],
     slf_op_06_17[2], slf_op_06_17[1], slf_op_06_17[0],
     slf_op_06_17[3], slf_op_06_17[2], slf_op_06_17[1],
     slf_op_06_17[0]}), .top_op_08({slf_op_05_17[3], slf_op_05_17[2],
     slf_op_05_17[1], slf_op_05_17[0], slf_op_05_17[3],
     slf_op_05_17[2], slf_op_05_17[1], slf_op_05_17[0]}),
     .tnl_op_08({slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0], slf_op_04_17[3], slf_op_04_17[2],
     slf_op_04_17[1], slf_op_04_17[0]}), .sp4_v_t_08({net1208[0],
     net1208[1], net1208[2], net1208[3], net1208[4], net1208[5],
     net1208[6], net1208[7], net1208[8], net1208[9], net1208[10],
     net1208[11], net1208[12], net1208[13], net1208[14], net1208[15],
     net1208[16], net1208[17], net1208[18], net1208[19], net1208[20],
     net1208[21], net1208[22], net1208[23], net1208[24], net1208[25],
     net1208[26], net1208[27], net1208[28], net1208[29], net1208[30],
     net1208[31], net1208[32], net1208[33], net1208[34], net1208[35],
     net1208[36], net1208[37], net1208[38], net1208[39], net1208[40],
     net1208[41], net1208[42], net1208[43], net1208[44], net1208[45],
     net1208[46], net1208[47]}), .lc_bot(lc_bot_05_09),
     .op_vic(net1462), .sp12_v_b_01(sp12_v_b_05_09[23:0]),
     .glb_netwk_t({net1212[0], net1212[1], net1212[2], net1212[3],
     net1212[4], net1212[5], net1212[6], net1212[7]}));
lt_1x8_top_ice1f I_lt_col_t04 ( .glb_netwk_b({net1213[0], net1213[1],
     net1213[2], net1213[3], net1213[4], net1213[5], net1213[6],
     net1213[7]}), .rgt_op_03({net1214[0], net1214[1], net1214[2],
     net1214[3], net1214[4], net1214[5], net1214[6], net1214[7]}),
     .slf_op_02({net773[0], net773[1], net773[2], net773[3], net773[4],
     net773[5], net773[6], net773[7]}), .rgt_op_02({net1216[0],
     net1216[1], net1216[2], net1216[3], net1216[4], net1216[5],
     net1216[6], net1216[7]}), .rgt_op_01(slf_op_05_09[7:0]),
     .purst(purst), .prog(prog), .lft_op_04({net1034[0], net1034[1],
     net1034[2], net1034[3], net1034[4], net1034[5], net1034[6],
     net1034[7]}), .lft_op_03({net1024[0], net1024[1], net1024[2],
     net1024[3], net1024[4], net1024[5], net1024[6], net1024[7]}),
     .lft_op_02({net1026[0], net1026[1], net1026[2], net1026[3],
     net1026[4], net1026[5], net1026[6], net1026[7]}),
     .lft_op_01(slf_op_03_09[7:0]), .rgt_op_04({net1224[0], net1224[1],
     net1224[2], net1224[3], net1224[4], net1224[5], net1224[6],
     net1224[7]}), .carry_in(carry_in_04_09),
     .bnl_op_01(bnl_op_04_09[7:0]), .slf_op_04({net771[0], net771[1],
     net771[2], net771[3], net771[4], net771[5], net771[6],
     net771[7]}), .slf_op_03({net772[0], net772[1], net772[2],
     net772[3], net772[4], net772[5], net772[6], net772[7]}),
     .slf_op_01(slf_op_04_09[7:0]), .sp4_h_l_04({net792[0], net792[1],
     net792[2], net792[3], net792[4], net792[5], net792[6], net792[7],
     net792[8], net792[9], net792[10], net792[11], net792[12],
     net792[13], net792[14], net792[15], net792[16], net792[17],
     net792[18], net792[19], net792[20], net792[21], net792[22],
     net792[23], net792[24], net792[25], net792[26], net792[27],
     net792[28], net792[29], net792[30], net792[31], net792[32],
     net792[33], net792[34], net792[35], net792[36], net792[37],
     net792[38], net792[39], net792[40], net792[41], net792[42],
     net792[43], net792[44], net792[45], net792[46], net792[47]}),
     .carry_out(net1231), .vdd_cntl(vdd_cntl_l[127:0]),
     .sp12_h_r_04({net1233[0], net1233[1], net1233[2], net1233[3],
     net1233[4], net1233[5], net1233[6], net1233[7], net1233[8],
     net1233[9], net1233[10], net1233[11], net1233[12], net1233[13],
     net1233[14], net1233[15], net1233[16], net1233[17], net1233[18],
     net1233[19], net1233[20], net1233[21], net1233[22], net1233[23]}),
     .sp12_h_r_03({net1234[0], net1234[1], net1234[2], net1234[3],
     net1234[4], net1234[5], net1234[6], net1234[7], net1234[8],
     net1234[9], net1234[10], net1234[11], net1234[12], net1234[13],
     net1234[14], net1234[15], net1234[16], net1234[17], net1234[18],
     net1234[19], net1234[20], net1234[21], net1234[22], net1234[23]}),
     .sp12_h_r_02({net1235[0], net1235[1], net1235[2], net1235[3],
     net1235[4], net1235[5], net1235[6], net1235[7], net1235[8],
     net1235[9], net1235[10], net1235[11], net1235[12], net1235[13],
     net1235[14], net1235[15], net1235[16], net1235[17], net1235[18],
     net1235[19], net1235[20], net1235[21], net1235[22], net1235[23]}),
     .sp12_h_r_01({net1236[0], net1236[1], net1236[2], net1236[3],
     net1236[4], net1236[5], net1236[6], net1236[7], net1236[8],
     net1236[9], net1236[10], net1236[11], net1236[12], net1236[13],
     net1236[14], net1236[15], net1236[16], net1236[17], net1236[18],
     net1236[19], net1236[20], net1236[21], net1236[22], net1236[23]}),
     .glb_netwk_col(clk_tree_drv_tl[7:0]),
     .sp4_v_b_01(sp4_v_b_04_09[47:0]), .sp4_r_v_b_04({net1239[0],
     net1239[1], net1239[2], net1239[3], net1239[4], net1239[5],
     net1239[6], net1239[7], net1239[8], net1239[9], net1239[10],
     net1239[11], net1239[12], net1239[13], net1239[14], net1239[15],
     net1239[16], net1239[17], net1239[18], net1239[19], net1239[20],
     net1239[21], net1239[22], net1239[23], net1239[24], net1239[25],
     net1239[26], net1239[27], net1239[28], net1239[29], net1239[30],
     net1239[31], net1239[32], net1239[33], net1239[34], net1239[35],
     net1239[36], net1239[37], net1239[38], net1239[39], net1239[40],
     net1239[41], net1239[42], net1239[43], net1239[44], net1239[45],
     net1239[46], net1239[47]}), .sp4_r_v_b_03({net1240[0], net1240[1],
     net1240[2], net1240[3], net1240[4], net1240[5], net1240[6],
     net1240[7], net1240[8], net1240[9], net1240[10], net1240[11],
     net1240[12], net1240[13], net1240[14], net1240[15], net1240[16],
     net1240[17], net1240[18], net1240[19], net1240[20], net1240[21],
     net1240[22], net1240[23], net1240[24], net1240[25], net1240[26],
     net1240[27], net1240[28], net1240[29], net1240[30], net1240[31],
     net1240[32], net1240[33], net1240[34], net1240[35], net1240[36],
     net1240[37], net1240[38], net1240[39], net1240[40], net1240[41],
     net1240[42], net1240[43], net1240[44], net1240[45], net1240[46],
     net1240[47]}), .sp4_r_v_b_02({net1241[0], net1241[1], net1241[2],
     net1241[3], net1241[4], net1241[5], net1241[6], net1241[7],
     net1241[8], net1241[9], net1241[10], net1241[11], net1241[12],
     net1241[13], net1241[14], net1241[15], net1241[16], net1241[17],
     net1241[18], net1241[19], net1241[20], net1241[21], net1241[22],
     net1241[23], net1241[24], net1241[25], net1241[26], net1241[27],
     net1241[28], net1241[29], net1241[30], net1241[31], net1241[32],
     net1241[33], net1241[34], net1241[35], net1241[36], net1241[37],
     net1241[38], net1241[39], net1241[40], net1241[41], net1241[42],
     net1241[43], net1241[44], net1241[45], net1241[46], net1241[47]}),
     .sp4_r_v_b_01(sp4_v_b_05_09[47:0]), .sp4_h_r_04({net1243[0],
     net1243[1], net1243[2], net1243[3], net1243[4], net1243[5],
     net1243[6], net1243[7], net1243[8], net1243[9], net1243[10],
     net1243[11], net1243[12], net1243[13], net1243[14], net1243[15],
     net1243[16], net1243[17], net1243[18], net1243[19], net1243[20],
     net1243[21], net1243[22], net1243[23], net1243[24], net1243[25],
     net1243[26], net1243[27], net1243[28], net1243[29], net1243[30],
     net1243[31], net1243[32], net1243[33], net1243[34], net1243[35],
     net1243[36], net1243[37], net1243[38], net1243[39], net1243[40],
     net1243[41], net1243[42], net1243[43], net1243[44], net1243[45],
     net1243[46], net1243[47]}), .sp4_h_r_03({net1244[0], net1244[1],
     net1244[2], net1244[3], net1244[4], net1244[5], net1244[6],
     net1244[7], net1244[8], net1244[9], net1244[10], net1244[11],
     net1244[12], net1244[13], net1244[14], net1244[15], net1244[16],
     net1244[17], net1244[18], net1244[19], net1244[20], net1244[21],
     net1244[22], net1244[23], net1244[24], net1244[25], net1244[26],
     net1244[27], net1244[28], net1244[29], net1244[30], net1244[31],
     net1244[32], net1244[33], net1244[34], net1244[35], net1244[36],
     net1244[37], net1244[38], net1244[39], net1244[40], net1244[41],
     net1244[42], net1244[43], net1244[44], net1244[45], net1244[46],
     net1244[47]}), .sp4_h_r_02({net1245[0], net1245[1], net1245[2],
     net1245[3], net1245[4], net1245[5], net1245[6], net1245[7],
     net1245[8], net1245[9], net1245[10], net1245[11], net1245[12],
     net1245[13], net1245[14], net1245[15], net1245[16], net1245[17],
     net1245[18], net1245[19], net1245[20], net1245[21], net1245[22],
     net1245[23], net1245[24], net1245[25], net1245[26], net1245[27],
     net1245[28], net1245[29], net1245[30], net1245[31], net1245[32],
     net1245[33], net1245[34], net1245[35], net1245[36], net1245[37],
     net1245[38], net1245[39], net1245[40], net1245[41], net1245[42],
     net1245[43], net1245[44], net1245[45], net1245[46], net1245[47]}),
     .sp4_h_r_01({net1246[0], net1246[1], net1246[2], net1246[3],
     net1246[4], net1246[5], net1246[6], net1246[7], net1246[8],
     net1246[9], net1246[10], net1246[11], net1246[12], net1246[13],
     net1246[14], net1246[15], net1246[16], net1246[17], net1246[18],
     net1246[19], net1246[20], net1246[21], net1246[22], net1246[23],
     net1246[24], net1246[25], net1246[26], net1246[27], net1246[28],
     net1246[29], net1246[30], net1246[31], net1246[32], net1246[33],
     net1246[34], net1246[35], net1246[36], net1246[37], net1246[38],
     net1246[39], net1246[40], net1246[41], net1246[42], net1246[43],
     net1246[44], net1246[45], net1246[46], net1246[47]}),
     .sp4_h_l_03({net791[0], net791[1], net791[2], net791[3],
     net791[4], net791[5], net791[6], net791[7], net791[8], net791[9],
     net791[10], net791[11], net791[12], net791[13], net791[14],
     net791[15], net791[16], net791[17], net791[18], net791[19],
     net791[20], net791[21], net791[22], net791[23], net791[24],
     net791[25], net791[26], net791[27], net791[28], net791[29],
     net791[30], net791[31], net791[32], net791[33], net791[34],
     net791[35], net791[36], net791[37], net791[38], net791[39],
     net791[40], net791[41], net791[42], net791[43], net791[44],
     net791[45], net791[46], net791[47]}), .sp4_h_l_02({net790[0],
     net790[1], net790[2], net790[3], net790[4], net790[5], net790[6],
     net790[7], net790[8], net790[9], net790[10], net790[11],
     net790[12], net790[13], net790[14], net790[15], net790[16],
     net790[17], net790[18], net790[19], net790[20], net790[21],
     net790[22], net790[23], net790[24], net790[25], net790[26],
     net790[27], net790[28], net790[29], net790[30], net790[31],
     net790[32], net790[33], net790[34], net790[35], net790[36],
     net790[37], net790[38], net790[39], net790[40], net790[41],
     net790[42], net790[43], net790[44], net790[45], net790[46],
     net790[47]}), .sp4_h_l_01({net746[0], net746[1], net746[2],
     net746[3], net746[4], net746[5], net746[6], net746[7], net746[8],
     net746[9], net746[10], net746[11], net746[12], net746[13],
     net746[14], net746[15], net746[16], net746[17], net746[18],
     net746[19], net746[20], net746[21], net746[22], net746[23],
     net746[24], net746[25], net746[26], net746[27], net746[28],
     net746[29], net746[30], net746[31], net746[32], net746[33],
     net746[34], net746[35], net746[36], net746[37], net746[38],
     net746[39], net746[40], net746[41], net746[42], net746[43],
     net746[44], net746[45], net746[46], net746[47]}),
     .bl(bl[221:168]), .bot_op_01(bot_op_04_09[7:0]),
     .sp12_h_l_01({net740[0], net740[1], net740[2], net740[3],
     net740[4], net740[5], net740[6], net740[7], net740[8], net740[9],
     net740[10], net740[11], net740[12], net740[13], net740[14],
     net740[15], net740[16], net740[17], net740[18], net740[19],
     net740[20], net740[21], net740[22], net740[23]}),
     .sp12_h_l_02({net748[0], net748[1], net748[2], net748[3],
     net748[4], net748[5], net748[6], net748[7], net748[8], net748[9],
     net748[10], net748[11], net748[12], net748[13], net748[14],
     net748[15], net748[16], net748[17], net748[18], net748[19],
     net748[20], net748[21], net748[22], net748[23]}),
     .sp12_h_l_03({net704[0], net704[1], net704[2], net704[3],
     net704[4], net704[5], net704[6], net704[7], net704[8], net704[9],
     net704[10], net704[11], net704[12], net704[13], net704[14],
     net704[15], net704[16], net704[17], net704[18], net704[19],
     net704[20], net704[21], net704[22], net704[23]}),
     .sp12_h_l_04({net749[0], net749[1], net749[2], net749[3],
     net749[4], net749[5], net749[6], net749[7], net749[8], net749[9],
     net749[10], net749[11], net749[12], net749[13], net749[14],
     net749[15], net749[16], net749[17], net749[18], net749[19],
     net749[20], net749[21], net749[22], net749[23]}),
     .sp4_v_b_04({net728[0], net728[1], net728[2], net728[3],
     net728[4], net728[5], net728[6], net728[7], net728[8], net728[9],
     net728[10], net728[11], net728[12], net728[13], net728[14],
     net728[15], net728[16], net728[17], net728[18], net728[19],
     net728[20], net728[21], net728[22], net728[23], net728[24],
     net728[25], net728[26], net728[27], net728[28], net728[29],
     net728[30], net728[31], net728[32], net728[33], net728[34],
     net728[35], net728[36], net728[37], net728[38], net728[39],
     net728[40], net728[41], net728[42], net728[43], net728[44],
     net728[45], net728[46], net728[47]}), .sp4_v_b_03({net724[0],
     net724[1], net724[2], net724[3], net724[4], net724[5], net724[6],
     net724[7], net724[8], net724[9], net724[10], net724[11],
     net724[12], net724[13], net724[14], net724[15], net724[16],
     net724[17], net724[18], net724[19], net724[20], net724[21],
     net724[22], net724[23], net724[24], net724[25], net724[26],
     net724[27], net724[28], net724[29], net724[30], net724[31],
     net724[32], net724[33], net724[34], net724[35], net724[36],
     net724[37], net724[38], net724[39], net724[40], net724[41],
     net724[42], net724[43], net724[44], net724[45], net724[46],
     net724[47]}), .sp4_v_b_02({net735[0], net735[1], net735[2],
     net735[3], net735[4], net735[5], net735[6], net735[7], net735[8],
     net735[9], net735[10], net735[11], net735[12], net735[13],
     net735[14], net735[15], net735[16], net735[17], net735[18],
     net735[19], net735[20], net735[21], net735[22], net735[23],
     net735[24], net735[25], net735[26], net735[27], net735[28],
     net735[29], net735[30], net735[31], net735[32], net735[33],
     net735[34], net735[35], net735[36], net735[37], net735[38],
     net735[39], net735[40], net735[41], net735[42], net735[43],
     net735[44], net735[45], net735[46], net735[47]}),
     .bnr_op_01(bnr_op_04_09[7:0]), .sp4_h_l_05({net793[0], net793[1],
     net793[2], net793[3], net793[4], net793[5], net793[6], net793[7],
     net793[8], net793[9], net793[10], net793[11], net793[12],
     net793[13], net793[14], net793[15], net793[16], net793[17],
     net793[18], net793[19], net793[20], net793[21], net793[22],
     net793[23], net793[24], net793[25], net793[26], net793[27],
     net793[28], net793[29], net793[30], net793[31], net793[32],
     net793[33], net793[34], net793[35], net793[36], net793[37],
     net793[38], net793[39], net793[40], net793[41], net793[42],
     net793[43], net793[44], net793[45], net793[46], net793[47]}),
     .sp4_h_l_06({net794[0], net794[1], net794[2], net794[3],
     net794[4], net794[5], net794[6], net794[7], net794[8], net794[9],
     net794[10], net794[11], net794[12], net794[13], net794[14],
     net794[15], net794[16], net794[17], net794[18], net794[19],
     net794[20], net794[21], net794[22], net794[23], net794[24],
     net794[25], net794[26], net794[27], net794[28], net794[29],
     net794[30], net794[31], net794[32], net794[33], net794[34],
     net794[35], net794[36], net794[37], net794[38], net794[39],
     net794[40], net794[41], net794[42], net794[43], net794[44],
     net794[45], net794[46], net794[47]}), .sp4_h_l_07({net795[0],
     net795[1], net795[2], net795[3], net795[4], net795[5], net795[6],
     net795[7], net795[8], net795[9], net795[10], net795[11],
     net795[12], net795[13], net795[14], net795[15], net795[16],
     net795[17], net795[18], net795[19], net795[20], net795[21],
     net795[22], net795[23], net795[24], net795[25], net795[26],
     net795[27], net795[28], net795[29], net795[30], net795[31],
     net795[32], net795[33], net795[34], net795[35], net795[36],
     net795[37], net795[38], net795[39], net795[40], net795[41],
     net795[42], net795[43], net795[44], net795[45], net795[46],
     net795[47]}), .sp4_h_l_08({net731[0], net731[1], net731[2],
     net731[3], net731[4], net731[5], net731[6], net731[7], net731[8],
     net731[9], net731[10], net731[11], net731[12], net731[13],
     net731[14], net731[15], net731[16], net731[17], net731[18],
     net731[19], net731[20], net731[21], net731[22], net731[23],
     net731[24], net731[25], net731[26], net731[27], net731[28],
     net731[29], net731[30], net731[31], net731[32], net731[33],
     net731[34], net731[35], net731[36], net731[37], net731[38],
     net731[39], net731[40], net731[41], net731[42], net731[43],
     net731[44], net731[45], net731[46], net731[47]}),
     .sp4_h_r_08({net1264[0], net1264[1], net1264[2], net1264[3],
     net1264[4], net1264[5], net1264[6], net1264[7], net1264[8],
     net1264[9], net1264[10], net1264[11], net1264[12], net1264[13],
     net1264[14], net1264[15], net1264[16], net1264[17], net1264[18],
     net1264[19], net1264[20], net1264[21], net1264[22], net1264[23],
     net1264[24], net1264[25], net1264[26], net1264[27], net1264[28],
     net1264[29], net1264[30], net1264[31], net1264[32], net1264[33],
     net1264[34], net1264[35], net1264[36], net1264[37], net1264[38],
     net1264[39], net1264[40], net1264[41], net1264[42], net1264[43],
     net1264[44], net1264[45], net1264[46], net1264[47]}),
     .sp4_h_r_07({net1265[0], net1265[1], net1265[2], net1265[3],
     net1265[4], net1265[5], net1265[6], net1265[7], net1265[8],
     net1265[9], net1265[10], net1265[11], net1265[12], net1265[13],
     net1265[14], net1265[15], net1265[16], net1265[17], net1265[18],
     net1265[19], net1265[20], net1265[21], net1265[22], net1265[23],
     net1265[24], net1265[25], net1265[26], net1265[27], net1265[28],
     net1265[29], net1265[30], net1265[31], net1265[32], net1265[33],
     net1265[34], net1265[35], net1265[36], net1265[37], net1265[38],
     net1265[39], net1265[40], net1265[41], net1265[42], net1265[43],
     net1265[44], net1265[45], net1265[46], net1265[47]}),
     .sp4_h_r_06({net1266[0], net1266[1], net1266[2], net1266[3],
     net1266[4], net1266[5], net1266[6], net1266[7], net1266[8],
     net1266[9], net1266[10], net1266[11], net1266[12], net1266[13],
     net1266[14], net1266[15], net1266[16], net1266[17], net1266[18],
     net1266[19], net1266[20], net1266[21], net1266[22], net1266[23],
     net1266[24], net1266[25], net1266[26], net1266[27], net1266[28],
     net1266[29], net1266[30], net1266[31], net1266[32], net1266[33],
     net1266[34], net1266[35], net1266[36], net1266[37], net1266[38],
     net1266[39], net1266[40], net1266[41], net1266[42], net1266[43],
     net1266[44], net1266[45], net1266[46], net1266[47]}),
     .sp4_h_r_05({net1267[0], net1267[1], net1267[2], net1267[3],
     net1267[4], net1267[5], net1267[6], net1267[7], net1267[8],
     net1267[9], net1267[10], net1267[11], net1267[12], net1267[13],
     net1267[14], net1267[15], net1267[16], net1267[17], net1267[18],
     net1267[19], net1267[20], net1267[21], net1267[22], net1267[23],
     net1267[24], net1267[25], net1267[26], net1267[27], net1267[28],
     net1267[29], net1267[30], net1267[31], net1267[32], net1267[33],
     net1267[34], net1267[35], net1267[36], net1267[37], net1267[38],
     net1267[39], net1267[40], net1267[41], net1267[42], net1267[43],
     net1267[44], net1267[45], net1267[46], net1267[47]}),
     .slf_op_05({net770[0], net770[1], net770[2], net770[3], net770[4],
     net770[5], net770[6], net770[7]}), .slf_op_06({net769[0],
     net769[1], net769[2], net769[3], net769[4], net769[5], net769[6],
     net769[7]}), .slf_op_07({net768[0], net768[1], net768[2],
     net768[3], net768[4], net768[5], net768[6], net768[7]}),
     .slf_op_08({net767[0], net767[1], net767[2], net767[3], net767[4],
     net767[5], net767[6], net767[7]}), .rgt_op_08({net1272[0],
     net1272[1], net1272[2], net1272[3], net1272[4], net1272[5],
     net1272[6], net1272[7]}), .rgt_op_07({net1273[0], net1273[1],
     net1273[2], net1273[3], net1273[4], net1273[5], net1273[6],
     net1273[7]}), .rgt_op_06({net1274[0], net1274[1], net1274[2],
     net1274[3], net1274[4], net1274[5], net1274[6], net1274[7]}),
     .rgt_op_05({net1275[0], net1275[1], net1275[2], net1275[3],
     net1275[4], net1275[5], net1275[6], net1275[7]}),
     .lft_op_08({net1082[0], net1082[1], net1082[2], net1082[3],
     net1082[4], net1082[5], net1082[6], net1082[7]}),
     .lft_op_07({net1083[0], net1083[1], net1083[2], net1083[3],
     net1083[4], net1083[5], net1083[6], net1083[7]}),
     .lft_op_06({net1084[0], net1084[1], net1084[2], net1084[3],
     net1084[4], net1084[5], net1084[6], net1084[7]}),
     .lft_op_05({net1085[0], net1085[1], net1085[2], net1085[3],
     net1085[4], net1085[5], net1085[6], net1085[7]}),
     .sp12_h_l_08({net721[0], net721[1], net721[2], net721[3],
     net721[4], net721[5], net721[6], net721[7], net721[8], net721[9],
     net721[10], net721[11], net721[12], net721[13], net721[14],
     net721[15], net721[16], net721[17], net721[18], net721[19],
     net721[20], net721[21], net721[22], net721[23]}),
     .sp12_h_l_07({net716[0], net716[1], net716[2], net716[3],
     net716[4], net716[5], net716[6], net716[7], net716[8], net716[9],
     net716[10], net716[11], net716[12], net716[13], net716[14],
     net716[15], net716[16], net716[17], net716[18], net716[19],
     net716[20], net716[21], net716[22], net716[23]}),
     .sp12_h_l_06({net718[0], net718[1], net718[2], net718[3],
     net718[4], net718[5], net718[6], net718[7], net718[8], net718[9],
     net718[10], net718[11], net718[12], net718[13], net718[14],
     net718[15], net718[16], net718[17], net718[18], net718[19],
     net718[20], net718[21], net718[22], net718[23]}),
     .sp12_h_r_05({net1283[0], net1283[1], net1283[2], net1283[3],
     net1283[4], net1283[5], net1283[6], net1283[7], net1283[8],
     net1283[9], net1283[10], net1283[11], net1283[12], net1283[13],
     net1283[14], net1283[15], net1283[16], net1283[17], net1283[18],
     net1283[19], net1283[20], net1283[21], net1283[22], net1283[23]}),
     .sp12_h_r_06({net1284[0], net1284[1], net1284[2], net1284[3],
     net1284[4], net1284[5], net1284[6], net1284[7], net1284[8],
     net1284[9], net1284[10], net1284[11], net1284[12], net1284[13],
     net1284[14], net1284[15], net1284[16], net1284[17], net1284[18],
     net1284[19], net1284[20], net1284[21], net1284[22], net1284[23]}),
     .sp12_h_r_07({net1285[0], net1285[1], net1285[2], net1285[3],
     net1285[4], net1285[5], net1285[6], net1285[7], net1285[8],
     net1285[9], net1285[10], net1285[11], net1285[12], net1285[13],
     net1285[14], net1285[15], net1285[16], net1285[17], net1285[18],
     net1285[19], net1285[20], net1285[21], net1285[22], net1285[23]}),
     .sp12_h_r_08({net1286[0], net1286[1], net1286[2], net1286[3],
     net1286[4], net1286[5], net1286[6], net1286[7], net1286[8],
     net1286[9], net1286[10], net1286[11], net1286[12], net1286[13],
     net1286[14], net1286[15], net1286[16], net1286[17], net1286[18],
     net1286[19], net1286[20], net1286[21], net1286[22], net1286[23]}),
     .sp12_h_l_05({net720[0], net720[1], net720[2], net720[3],
     net720[4], net720[5], net720[6], net720[7], net720[8], net720[9],
     net720[10], net720[11], net720[12], net720[13], net720[14],
     net720[15], net720[16], net720[17], net720[18], net720[19],
     net720[20], net720[21], net720[22], net720[23]}),
     .sp4_r_v_b_05({net1288[0], net1288[1], net1288[2], net1288[3],
     net1288[4], net1288[5], net1288[6], net1288[7], net1288[8],
     net1288[9], net1288[10], net1288[11], net1288[12], net1288[13],
     net1288[14], net1288[15], net1288[16], net1288[17], net1288[18],
     net1288[19], net1288[20], net1288[21], net1288[22], net1288[23],
     net1288[24], net1288[25], net1288[26], net1288[27], net1288[28],
     net1288[29], net1288[30], net1288[31], net1288[32], net1288[33],
     net1288[34], net1288[35], net1288[36], net1288[37], net1288[38],
     net1288[39], net1288[40], net1288[41], net1288[42], net1288[43],
     net1288[44], net1288[45], net1288[46], net1288[47]}),
     .sp4_r_v_b_06({net1289[0], net1289[1], net1289[2], net1289[3],
     net1289[4], net1289[5], net1289[6], net1289[7], net1289[8],
     net1289[9], net1289[10], net1289[11], net1289[12], net1289[13],
     net1289[14], net1289[15], net1289[16], net1289[17], net1289[18],
     net1289[19], net1289[20], net1289[21], net1289[22], net1289[23],
     net1289[24], net1289[25], net1289[26], net1289[27], net1289[28],
     net1289[29], net1289[30], net1289[31], net1289[32], net1289[33],
     net1289[34], net1289[35], net1289[36], net1289[37], net1289[38],
     net1289[39], net1289[40], net1289[41], net1289[42], net1289[43],
     net1289[44], net1289[45], net1289[46], net1289[47]}),
     .sp4_r_v_b_07({net1290[0], net1290[1], net1290[2], net1290[3],
     net1290[4], net1290[5], net1290[6], net1290[7], net1290[8],
     net1290[9], net1290[10], net1290[11], net1290[12], net1290[13],
     net1290[14], net1290[15], net1290[16], net1290[17], net1290[18],
     net1290[19], net1290[20], net1290[21], net1290[22], net1290[23],
     net1290[24], net1290[25], net1290[26], net1290[27], net1290[28],
     net1290[29], net1290[30], net1290[31], net1290[32], net1290[33],
     net1290[34], net1290[35], net1290[36], net1290[37], net1290[38],
     net1290[39], net1290[40], net1290[41], net1290[42], net1290[43],
     net1290[44], net1290[45], net1290[46], net1290[47]}),
     .sp4_r_v_b_08({net1291[0], net1291[1], net1291[2], net1291[3],
     net1291[4], net1291[5], net1291[6], net1291[7], net1291[8],
     net1291[9], net1291[10], net1291[11], net1291[12], net1291[13],
     net1291[14], net1291[15], net1291[16], net1291[17], net1291[18],
     net1291[19], net1291[20], net1291[21], net1291[22], net1291[23],
     net1291[24], net1291[25], net1291[26], net1291[27], net1291[28],
     net1291[29], net1291[30], net1291[31], net1291[32], net1291[33],
     net1291[34], net1291[35], net1291[36], net1291[37], net1291[38],
     net1291[39], net1291[40], net1291[41], net1291[42], net1291[43],
     net1291[44], net1291[45], net1291[46], net1291[47]}),
     .sp4_v_b_08({net763[0], net763[1], net763[2], net763[3],
     net763[4], net763[5], net763[6], net763[7], net763[8], net763[9],
     net763[10], net763[11], net763[12], net763[13], net763[14],
     net763[15], net763[16], net763[17], net763[18], net763[19],
     net763[20], net763[21], net763[22], net763[23], net763[24],
     net763[25], net763[26], net763[27], net763[28], net763[29],
     net763[30], net763[31], net763[32], net763[33], net763[34],
     net763[35], net763[36], net763[37], net763[38], net763[39],
     net763[40], net763[41], net763[42], net763[43], net763[44],
     net763[45], net763[46], net763[47]}), .sp4_v_b_07({net764[0],
     net764[1], net764[2], net764[3], net764[4], net764[5], net764[6],
     net764[7], net764[8], net764[9], net764[10], net764[11],
     net764[12], net764[13], net764[14], net764[15], net764[16],
     net764[17], net764[18], net764[19], net764[20], net764[21],
     net764[22], net764[23], net764[24], net764[25], net764[26],
     net764[27], net764[28], net764[29], net764[30], net764[31],
     net764[32], net764[33], net764[34], net764[35], net764[36],
     net764[37], net764[38], net764[39], net764[40], net764[41],
     net764[42], net764[43], net764[44], net764[45], net764[46],
     net764[47]}), .sp4_v_b_06({net765[0], net765[1], net765[2],
     net765[3], net765[4], net765[5], net765[6], net765[7], net765[8],
     net765[9], net765[10], net765[11], net765[12], net765[13],
     net765[14], net765[15], net765[16], net765[17], net765[18],
     net765[19], net765[20], net765[21], net765[22], net765[23],
     net765[24], net765[25], net765[26], net765[27], net765[28],
     net765[29], net765[30], net765[31], net765[32], net765[33],
     net765[34], net765[35], net765[36], net765[37], net765[38],
     net765[39], net765[40], net765[41], net765[42], net765[43],
     net765[44], net765[45], net765[46], net765[47]}),
     .sp4_v_b_05({net732[0], net732[1], net732[2], net732[3],
     net732[4], net732[5], net732[6], net732[7], net732[8], net732[9],
     net732[10], net732[11], net732[12], net732[13], net732[14],
     net732[15], net732[16], net732[17], net732[18], net732[19],
     net732[20], net732[21], net732[22], net732[23], net732[24],
     net732[25], net732[26], net732[27], net732[28], net732[29],
     net732[30], net732[31], net732[32], net732[33], net732[34],
     net732[35], net732[36], net732[37], net732[38], net732[39],
     net732[40], net732[41], net732[42], net732[43], net732[44],
     net732[45], net732[46], net732[47]}), .pgate(pgate_l[127:0]),
     .reset_b(reset_b_l[127:0]), .wl(wl_l[127:0]),
     .sp12_v_t_08({net1299[0], net1299[1], net1299[2], net1299[3],
     net1299[4], net1299[5], net1299[6], net1299[7], net1299[8],
     net1299[9], net1299[10], net1299[11], net1299[12], net1299[13],
     net1299[14], net1299[15], net1299[16], net1299[17], net1299[18],
     net1299[19], net1299[20], net1299[21], net1299[22], net1299[23]}),
     .tnr_op_08({slf_op_05_17[3], slf_op_05_17[2], slf_op_05_17[1],
     slf_op_05_17[0], slf_op_05_17[3], slf_op_05_17[2],
     slf_op_05_17[1], slf_op_05_17[0]}), .top_op_08({slf_op_04_17[3],
     slf_op_04_17[2], slf_op_04_17[1], slf_op_04_17[0],
     slf_op_04_17[3], slf_op_04_17[2], slf_op_04_17[1],
     slf_op_04_17[0]}), .tnl_op_08({slf_op_08_17[3], slf_op_08_17[2],
     slf_op_08_17[1], slf_op_08_17[0], slf_op_08_17[3],
     slf_op_08_17[2], slf_op_08_17[1], slf_op_08_17[0]}),
     .sp4_v_t_08({net1303[0], net1303[1], net1303[2], net1303[3],
     net1303[4], net1303[5], net1303[6], net1303[7], net1303[8],
     net1303[9], net1303[10], net1303[11], net1303[12], net1303[13],
     net1303[14], net1303[15], net1303[16], net1303[17], net1303[18],
     net1303[19], net1303[20], net1303[21], net1303[22], net1303[23],
     net1303[24], net1303[25], net1303[26], net1303[27], net1303[28],
     net1303[29], net1303[30], net1303[31], net1303[32], net1303[33],
     net1303[34], net1303[35], net1303[36], net1303[37], net1303[38],
     net1303[39], net1303[40], net1303[41], net1303[42], net1303[43],
     net1303[44], net1303[45], net1303[46], net1303[47]}),
     .lc_bot(lc_bot_04_09), .op_vic(net1459),
     .sp12_v_b_01(sp12_v_b_04_09[23:0]), .glb_netwk_t({net1307[0],
     net1307[1], net1307[2], net1307[3], net1307[4], net1307[5],
     net1307[6], net1307[7]}));
lt_1x8_top_ice1f I_lt_col_t06 ( .glb_netwk_b({net1460[0], net1460[1],
     net1460[2], net1460[3], net1460[4], net1460[5], net1460[6],
     net1460[7]}), .rgt_op_03(rgt_op_06_11[7:0]),
     .slf_op_02(slf_op_06_10[7:0]), .rgt_op_02(rgt_op_06_10[7:0]),
     .rgt_op_01(rgt_op_06_09[7:0]), .purst(purst), .prog(prog),
     .lft_op_04({net1224[0], net1224[1], net1224[2], net1224[3],
     net1224[4], net1224[5], net1224[6], net1224[7]}),
     .lft_op_03({net1214[0], net1214[1], net1214[2], net1214[3],
     net1214[4], net1214[5], net1214[6], net1214[7]}),
     .lft_op_02({net1216[0], net1216[1], net1216[2], net1216[3],
     net1216[4], net1216[5], net1216[6], net1216[7]}),
     .lft_op_01(slf_op_05_09[7:0]), .rgt_op_04(rgt_op_06_12[7:0]),
     .carry_in(carry_in_06_09), .bnl_op_01(bnl_op_06_09[7:0]),
     .slf_op_04(slf_op_06_12[7:0]), .slf_op_03(slf_op_06_11[7:0]),
     .slf_op_01(slf_op_06_09[7:0]), .sp4_h_l_04({net1148[0],
     net1148[1], net1148[2], net1148[3], net1148[4], net1148[5],
     net1148[6], net1148[7], net1148[8], net1148[9], net1148[10],
     net1148[11], net1148[12], net1148[13], net1148[14], net1148[15],
     net1148[16], net1148[17], net1148[18], net1148[19], net1148[20],
     net1148[21], net1148[22], net1148[23], net1148[24], net1148[25],
     net1148[26], net1148[27], net1148[28], net1148[29], net1148[30],
     net1148[31], net1148[32], net1148[33], net1148[34], net1148[35],
     net1148[36], net1148[37], net1148[38], net1148[39], net1148[40],
     net1148[41], net1148[42], net1148[43], net1148[44], net1148[45],
     net1148[46], net1148[47]}), .carry_out(net1326),
     .vdd_cntl(vdd_cntl_l[127:0]), .sp12_h_r_04(sp12_h_r_06_12[23:0]),
     .sp12_h_r_03(sp12_h_r_06_11[23:0]),
     .sp12_h_r_02(sp12_h_r_06_10[23:0]),
     .sp12_h_r_01(sp12_h_r_06_09[23:0]), .glb_netwk_col({net1332[0],
     net1332[1], net1332[2], net1332[3], net1332[4], net1332[5],
     net1332[6], net1332[7]}), .sp4_v_b_01(sp4_v_b_06_09[47:0]),
     .sp4_r_v_b_04(sp4_r_v_b_06_12[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_06_11[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_06_10[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_06_09[47:0]),
     .sp4_h_r_04(sp4_h_r_06_12[47:0]),
     .sp4_h_r_03(sp4_h_r_06_11[47:0]),
     .sp4_h_r_02(sp4_h_r_06_10[47:0]),
     .sp4_h_r_01(sp4_h_r_06_09[47:0]), .sp4_h_l_03({net1149[0],
     net1149[1], net1149[2], net1149[3], net1149[4], net1149[5],
     net1149[6], net1149[7], net1149[8], net1149[9], net1149[10],
     net1149[11], net1149[12], net1149[13], net1149[14], net1149[15],
     net1149[16], net1149[17], net1149[18], net1149[19], net1149[20],
     net1149[21], net1149[22], net1149[23], net1149[24], net1149[25],
     net1149[26], net1149[27], net1149[28], net1149[29], net1149[30],
     net1149[31], net1149[32], net1149[33], net1149[34], net1149[35],
     net1149[36], net1149[37], net1149[38], net1149[39], net1149[40],
     net1149[41], net1149[42], net1149[43], net1149[44], net1149[45],
     net1149[46], net1149[47]}), .sp4_h_l_02({net1150[0], net1150[1],
     net1150[2], net1150[3], net1150[4], net1150[5], net1150[6],
     net1150[7], net1150[8], net1150[9], net1150[10], net1150[11],
     net1150[12], net1150[13], net1150[14], net1150[15], net1150[16],
     net1150[17], net1150[18], net1150[19], net1150[20], net1150[21],
     net1150[22], net1150[23], net1150[24], net1150[25], net1150[26],
     net1150[27], net1150[28], net1150[29], net1150[30], net1150[31],
     net1150[32], net1150[33], net1150[34], net1150[35], net1150[36],
     net1150[37], net1150[38], net1150[39], net1150[40], net1150[41],
     net1150[42], net1150[43], net1150[44], net1150[45], net1150[46],
     net1150[47]}), .sp4_h_l_01({net1151[0], net1151[1], net1151[2],
     net1151[3], net1151[4], net1151[5], net1151[6], net1151[7],
     net1151[8], net1151[9], net1151[10], net1151[11], net1151[12],
     net1151[13], net1151[14], net1151[15], net1151[16], net1151[17],
     net1151[18], net1151[19], net1151[20], net1151[21], net1151[22],
     net1151[23], net1151[24], net1151[25], net1151[26], net1151[27],
     net1151[28], net1151[29], net1151[30], net1151[31], net1151[32],
     net1151[33], net1151[34], net1151[35], net1151[36], net1151[37],
     net1151[38], net1151[39], net1151[40], net1151[41], net1151[42],
     net1151[43], net1151[44], net1151[45], net1151[46], net1151[47]}),
     .bl(bl[329:276]), .bot_op_01(bot_op_06_09[7:0]),
     .sp12_h_l_01({net1141[0], net1141[1], net1141[2], net1141[3],
     net1141[4], net1141[5], net1141[6], net1141[7], net1141[8],
     net1141[9], net1141[10], net1141[11], net1141[12], net1141[13],
     net1141[14], net1141[15], net1141[16], net1141[17], net1141[18],
     net1141[19], net1141[20], net1141[21], net1141[22], net1141[23]}),
     .sp12_h_l_02({net1140[0], net1140[1], net1140[2], net1140[3],
     net1140[4], net1140[5], net1140[6], net1140[7], net1140[8],
     net1140[9], net1140[10], net1140[11], net1140[12], net1140[13],
     net1140[14], net1140[15], net1140[16], net1140[17], net1140[18],
     net1140[19], net1140[20], net1140[21], net1140[22], net1140[23]}),
     .sp12_h_l_03({net1139[0], net1139[1], net1139[2], net1139[3],
     net1139[4], net1139[5], net1139[6], net1139[7], net1139[8],
     net1139[9], net1139[10], net1139[11], net1139[12], net1139[13],
     net1139[14], net1139[15], net1139[16], net1139[17], net1139[18],
     net1139[19], net1139[20], net1139[21], net1139[22], net1139[23]}),
     .sp12_h_l_04({net1138[0], net1138[1], net1138[2], net1138[3],
     net1138[4], net1138[5], net1138[6], net1138[7], net1138[8],
     net1138[9], net1138[10], net1138[11], net1138[12], net1138[13],
     net1138[14], net1138[15], net1138[16], net1138[17], net1138[18],
     net1138[19], net1138[20], net1138[21], net1138[22], net1138[23]}),
     .sp4_v_b_04({net1144[0], net1144[1], net1144[2], net1144[3],
     net1144[4], net1144[5], net1144[6], net1144[7], net1144[8],
     net1144[9], net1144[10], net1144[11], net1144[12], net1144[13],
     net1144[14], net1144[15], net1144[16], net1144[17], net1144[18],
     net1144[19], net1144[20], net1144[21], net1144[22], net1144[23],
     net1144[24], net1144[25], net1144[26], net1144[27], net1144[28],
     net1144[29], net1144[30], net1144[31], net1144[32], net1144[33],
     net1144[34], net1144[35], net1144[36], net1144[37], net1144[38],
     net1144[39], net1144[40], net1144[41], net1144[42], net1144[43],
     net1144[44], net1144[45], net1144[46], net1144[47]}),
     .sp4_v_b_03({net1145[0], net1145[1], net1145[2], net1145[3],
     net1145[4], net1145[5], net1145[6], net1145[7], net1145[8],
     net1145[9], net1145[10], net1145[11], net1145[12], net1145[13],
     net1145[14], net1145[15], net1145[16], net1145[17], net1145[18],
     net1145[19], net1145[20], net1145[21], net1145[22], net1145[23],
     net1145[24], net1145[25], net1145[26], net1145[27], net1145[28],
     net1145[29], net1145[30], net1145[31], net1145[32], net1145[33],
     net1145[34], net1145[35], net1145[36], net1145[37], net1145[38],
     net1145[39], net1145[40], net1145[41], net1145[42], net1145[43],
     net1145[44], net1145[45], net1145[46], net1145[47]}),
     .sp4_v_b_02({net1146[0], net1146[1], net1146[2], net1146[3],
     net1146[4], net1146[5], net1146[6], net1146[7], net1146[8],
     net1146[9], net1146[10], net1146[11], net1146[12], net1146[13],
     net1146[14], net1146[15], net1146[16], net1146[17], net1146[18],
     net1146[19], net1146[20], net1146[21], net1146[22], net1146[23],
     net1146[24], net1146[25], net1146[26], net1146[27], net1146[28],
     net1146[29], net1146[30], net1146[31], net1146[32], net1146[33],
     net1146[34], net1146[35], net1146[36], net1146[37], net1146[38],
     net1146[39], net1146[40], net1146[41], net1146[42], net1146[43],
     net1146[44], net1146[45], net1146[46], net1146[47]}),
     .bnr_op_01(bnr_op_06_09[7:0]), .sp4_h_l_05({net1172[0],
     net1172[1], net1172[2], net1172[3], net1172[4], net1172[5],
     net1172[6], net1172[7], net1172[8], net1172[9], net1172[10],
     net1172[11], net1172[12], net1172[13], net1172[14], net1172[15],
     net1172[16], net1172[17], net1172[18], net1172[19], net1172[20],
     net1172[21], net1172[22], net1172[23], net1172[24], net1172[25],
     net1172[26], net1172[27], net1172[28], net1172[29], net1172[30],
     net1172[31], net1172[32], net1172[33], net1172[34], net1172[35],
     net1172[36], net1172[37], net1172[38], net1172[39], net1172[40],
     net1172[41], net1172[42], net1172[43], net1172[44], net1172[45],
     net1172[46], net1172[47]}), .sp4_h_l_06({net1171[0], net1171[1],
     net1171[2], net1171[3], net1171[4], net1171[5], net1171[6],
     net1171[7], net1171[8], net1171[9], net1171[10], net1171[11],
     net1171[12], net1171[13], net1171[14], net1171[15], net1171[16],
     net1171[17], net1171[18], net1171[19], net1171[20], net1171[21],
     net1171[22], net1171[23], net1171[24], net1171[25], net1171[26],
     net1171[27], net1171[28], net1171[29], net1171[30], net1171[31],
     net1171[32], net1171[33], net1171[34], net1171[35], net1171[36],
     net1171[37], net1171[38], net1171[39], net1171[40], net1171[41],
     net1171[42], net1171[43], net1171[44], net1171[45], net1171[46],
     net1171[47]}), .sp4_h_l_07({net1170[0], net1170[1], net1170[2],
     net1170[3], net1170[4], net1170[5], net1170[6], net1170[7],
     net1170[8], net1170[9], net1170[10], net1170[11], net1170[12],
     net1170[13], net1170[14], net1170[15], net1170[16], net1170[17],
     net1170[18], net1170[19], net1170[20], net1170[21], net1170[22],
     net1170[23], net1170[24], net1170[25], net1170[26], net1170[27],
     net1170[28], net1170[29], net1170[30], net1170[31], net1170[32],
     net1170[33], net1170[34], net1170[35], net1170[36], net1170[37],
     net1170[38], net1170[39], net1170[40], net1170[41], net1170[42],
     net1170[43], net1170[44], net1170[45], net1170[46], net1170[47]}),
     .sp4_h_l_08({net1169[0], net1169[1], net1169[2], net1169[3],
     net1169[4], net1169[5], net1169[6], net1169[7], net1169[8],
     net1169[9], net1169[10], net1169[11], net1169[12], net1169[13],
     net1169[14], net1169[15], net1169[16], net1169[17], net1169[18],
     net1169[19], net1169[20], net1169[21], net1169[22], net1169[23],
     net1169[24], net1169[25], net1169[26], net1169[27], net1169[28],
     net1169[29], net1169[30], net1169[31], net1169[32], net1169[33],
     net1169[34], net1169[35], net1169[36], net1169[37], net1169[38],
     net1169[39], net1169[40], net1169[41], net1169[42], net1169[43],
     net1169[44], net1169[45], net1169[46], net1169[47]}),
     .sp4_h_r_08(sp4_h_r_06_16[47:0]),
     .sp4_h_r_07(sp4_h_r_06_15[47:0]),
     .sp4_h_r_06(sp4_h_r_06_14[47:0]),
     .sp4_h_r_05(sp4_h_r_06_13[47:0]), .slf_op_05(slf_op_06_13[7:0]),
     .slf_op_06(slf_op_06_14[7:0]), .slf_op_07(slf_op_06_15[7:0]),
     .slf_op_08(slf_op_06_16[7:0]), .rgt_op_08(rgt_op_06_16[7:0]),
     .rgt_op_07(rgt_op_06_15[7:0]), .rgt_op_06(rgt_op_06_14[7:0]),
     .rgt_op_05(rgt_op_06_13[7:0]), .lft_op_08({net1272[0], net1272[1],
     net1272[2], net1272[3], net1272[4], net1272[5], net1272[6],
     net1272[7]}), .lft_op_07({net1273[0], net1273[1], net1273[2],
     net1273[3], net1273[4], net1273[5], net1273[6], net1273[7]}),
     .lft_op_06({net1274[0], net1274[1], net1274[2], net1274[3],
     net1274[4], net1274[5], net1274[6], net1274[7]}),
     .lft_op_05({net1275[0], net1275[1], net1275[2], net1275[3],
     net1275[4], net1275[5], net1275[6], net1275[7]}),
     .sp12_h_l_08({net1191[0], net1191[1], net1191[2], net1191[3],
     net1191[4], net1191[5], net1191[6], net1191[7], net1191[8],
     net1191[9], net1191[10], net1191[11], net1191[12], net1191[13],
     net1191[14], net1191[15], net1191[16], net1191[17], net1191[18],
     net1191[19], net1191[20], net1191[21], net1191[22], net1191[23]}),
     .sp12_h_l_07({net1190[0], net1190[1], net1190[2], net1190[3],
     net1190[4], net1190[5], net1190[6], net1190[7], net1190[8],
     net1190[9], net1190[10], net1190[11], net1190[12], net1190[13],
     net1190[14], net1190[15], net1190[16], net1190[17], net1190[18],
     net1190[19], net1190[20], net1190[21], net1190[22], net1190[23]}),
     .sp12_h_l_06({net1189[0], net1189[1], net1189[2], net1189[3],
     net1189[4], net1189[5], net1189[6], net1189[7], net1189[8],
     net1189[9], net1189[10], net1189[11], net1189[12], net1189[13],
     net1189[14], net1189[15], net1189[16], net1189[17], net1189[18],
     net1189[19], net1189[20], net1189[21], net1189[22], net1189[23]}),
     .sp12_h_r_05(sp12_h_r_06_13[23:0]),
     .sp12_h_r_06(sp12_h_r_06_14[23:0]),
     .sp12_h_r_07(sp12_h_r_06_15[23:0]),
     .sp12_h_r_08(sp12_h_r_06_16[23:0]), .sp12_h_l_05({net1188[0],
     net1188[1], net1188[2], net1188[3], net1188[4], net1188[5],
     net1188[6], net1188[7], net1188[8], net1188[9], net1188[10],
     net1188[11], net1188[12], net1188[13], net1188[14], net1188[15],
     net1188[16], net1188[17], net1188[18], net1188[19], net1188[20],
     net1188[21], net1188[22], net1188[23]}),
     .sp4_r_v_b_05(sp4_r_v_b_06_13[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_06_14[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_06_15[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_06_16[47:0]), .sp4_v_b_08({net1196[0],
     net1196[1], net1196[2], net1196[3], net1196[4], net1196[5],
     net1196[6], net1196[7], net1196[8], net1196[9], net1196[10],
     net1196[11], net1196[12], net1196[13], net1196[14], net1196[15],
     net1196[16], net1196[17], net1196[18], net1196[19], net1196[20],
     net1196[21], net1196[22], net1196[23], net1196[24], net1196[25],
     net1196[26], net1196[27], net1196[28], net1196[29], net1196[30],
     net1196[31], net1196[32], net1196[33], net1196[34], net1196[35],
     net1196[36], net1196[37], net1196[38], net1196[39], net1196[40],
     net1196[41], net1196[42], net1196[43], net1196[44], net1196[45],
     net1196[46], net1196[47]}), .sp4_v_b_07({net1195[0], net1195[1],
     net1195[2], net1195[3], net1195[4], net1195[5], net1195[6],
     net1195[7], net1195[8], net1195[9], net1195[10], net1195[11],
     net1195[12], net1195[13], net1195[14], net1195[15], net1195[16],
     net1195[17], net1195[18], net1195[19], net1195[20], net1195[21],
     net1195[22], net1195[23], net1195[24], net1195[25], net1195[26],
     net1195[27], net1195[28], net1195[29], net1195[30], net1195[31],
     net1195[32], net1195[33], net1195[34], net1195[35], net1195[36],
     net1195[37], net1195[38], net1195[39], net1195[40], net1195[41],
     net1195[42], net1195[43], net1195[44], net1195[45], net1195[46],
     net1195[47]}), .sp4_v_b_06({net1194[0], net1194[1], net1194[2],
     net1194[3], net1194[4], net1194[5], net1194[6], net1194[7],
     net1194[8], net1194[9], net1194[10], net1194[11], net1194[12],
     net1194[13], net1194[14], net1194[15], net1194[16], net1194[17],
     net1194[18], net1194[19], net1194[20], net1194[21], net1194[22],
     net1194[23], net1194[24], net1194[25], net1194[26], net1194[27],
     net1194[28], net1194[29], net1194[30], net1194[31], net1194[32],
     net1194[33], net1194[34], net1194[35], net1194[36], net1194[37],
     net1194[38], net1194[39], net1194[40], net1194[41], net1194[42],
     net1194[43], net1194[44], net1194[45], net1194[46], net1194[47]}),
     .sp4_v_b_05({net1193[0], net1193[1], net1193[2], net1193[3],
     net1193[4], net1193[5], net1193[6], net1193[7], net1193[8],
     net1193[9], net1193[10], net1193[11], net1193[12], net1193[13],
     net1193[14], net1193[15], net1193[16], net1193[17], net1193[18],
     net1193[19], net1193[20], net1193[21], net1193[22], net1193[23],
     net1193[24], net1193[25], net1193[26], net1193[27], net1193[28],
     net1193[29], net1193[30], net1193[31], net1193[32], net1193[33],
     net1193[34], net1193[35], net1193[36], net1193[37], net1193[38],
     net1193[39], net1193[40], net1193[41], net1193[42], net1193[43],
     net1193[44], net1193[45], net1193[46], net1193[47]}),
     .pgate(pgate_l[127:0]), .reset_b(reset_b_l[127:0]),
     .wl(wl_l[127:0]), .sp12_v_t_08({net1394[0], net1394[1],
     net1394[2], net1394[3], net1394[4], net1394[5], net1394[6],
     net1394[7], net1394[8], net1394[9], net1394[10], net1394[11],
     net1394[12], net1394[13], net1394[14], net1394[15], net1394[16],
     net1394[17], net1394[18], net1394[19], net1394[20], net1394[21],
     net1394[22], net1394[23]}), .tnr_op_08({tnr_op_06_16[3],
     tnr_op_06_16[2], tnr_op_06_16[1], tnr_op_06_16[0],
     tnr_op_06_16[3], tnr_op_06_16[2], tnr_op_06_16[1],
     tnr_op_06_16[0]}), .top_op_08({slf_op_06_17[3], slf_op_06_17[2],
     slf_op_06_17[1], slf_op_06_17[0], slf_op_06_17[3],
     slf_op_06_17[2], slf_op_06_17[1], slf_op_06_17[0]}),
     .tnl_op_08({slf_op_05_17[3], slf_op_05_17[2], slf_op_05_17[1],
     slf_op_05_17[0], slf_op_05_17[3], slf_op_05_17[2],
     slf_op_05_17[1], slf_op_05_17[0]}), .sp4_v_t_08({net1398[0],
     net1398[1], net1398[2], net1398[3], net1398[4], net1398[5],
     net1398[6], net1398[7], net1398[8], net1398[9], net1398[10],
     net1398[11], net1398[12], net1398[13], net1398[14], net1398[15],
     net1398[16], net1398[17], net1398[18], net1398[19], net1398[20],
     net1398[21], net1398[22], net1398[23], net1398[24], net1398[25],
     net1398[26], net1398[27], net1398[28], net1398[29], net1398[30],
     net1398[31], net1398[32], net1398[33], net1398[34], net1398[35],
     net1398[36], net1398[37], net1398[38], net1398[39], net1398[40],
     net1398[41], net1398[42], net1398[43], net1398[44], net1398[45],
     net1398[46], net1398[47]}), .lc_bot(lc_bot_06_09),
     .op_vic(net1465), .sp12_v_b_01(sp12_v_b_06_09[23:0]),
     .glb_netwk_t({net1402[0], net1402[1], net1402[2], net1402[3],
     net1402[4], net1402[5], net1402[6], net1402[7]}));
tielo I369 ( .tielo(tiegnd_qtl));
tielo I365 ( .tielo(tiegnd_bram_t));
scan_buf_ice8p I_scanbuf_8p_tl ( .update_i(net1405), .tclk_i(net1406),
     .shift_i(net1407), .sdi(net1408), .r_i(net1409), .mode_i(net1410),
     .hiz_b_i(net1411), .ceb_i(net1412), .bs_en_i(net1413),
     .update_o(update_o), .tclk_o(net816), .shift_o(shift_o),
     .sdo(net803), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
fabric_buf_ice8p I385 ( .f_in(net1423), .f_out(fabric_out_00_09));
fabric_buf_ice8p I390 ( .f_in(net675), .f_out(padin_06_17b));
fabric_buf_ice8p I391 ( .f_in(net1427), .f_out(padin_00_09a));
fabric_buf_ice8p I388 ( .f_in(net859), .f_out(fabric_out_06_17));
clk_quad_buf_x8_ice8p I_clk_qtl_center ( .clko(clk_tree_drv_tl[7:0]),
     .clki(clk_center[7:0]));
clk_quad_buf_x8_ice8p I_clktree_quad_drv_tl ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));

endmodule
// Library - leafcell, Cell - pinlatbuf12p_1, View - schematic
// LAST TIME SAVED: Dec 24 09:06:49 2010
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module pinlatbuf12p_1 ( cout, cbit, icegate, pad_in, prog );
output  cout;

input  cbit, icegate, pad_in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I_txgate_lvt_2 ( .in(cout), .out(net13), .pp(net046),
     .nn(net17));
txgate_lvt I_txgate_lvt_1 ( .in(pad_in), .out(net13), .pp(net17),
     .nn(net046));
inv_lvt I6 ( .A(net046), .Y(net17));
inv_lvt I24 ( .A(prog), .Y(net19));
inv_lvt I_inv_lvt ( .A(net044), .Y(cout));
nand2_lvt I_nand2_lvt ( .A(net19), .Y(net044), .B(net13));
nand2_lvt I5 ( .A(icegate), .Y(net046), .B(cbit));

endmodule
// Library - ice1chip, Cell - io_rgt_bot_1x8_ice1f, View - schematic
// LAST TIME SAVED: Mar 10 17:31:55 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module io_rgt_bot_1x8_ice1f ( cf_r[191:0], fabric_out_01,
     fabric_out_02, fabric_out_08, padeb[12:0], pado[12:0], sdo,
     slf_op_01[3:0], slf_op_02[3:0], slf_op_03[3:0], slf_op_04[3:0],
     slf_op_05[3:0], slf_op_06[3:0], slf_op_07[3:0], slf_op_08[3:0],
     tck_pad, tclk_o, tdi_pad, tms_pad, SP4_h_l_01[47:0],
     SP4_h_l_02[47:0], SP4_h_l_03[47:0], SP4_h_l_04[47:0],
     SP4_h_l_05[47:0], SP4_h_l_06[47:0], SP4_h_l_07[47:0],
     SP4_h_l_08[47:0], SP12_h_l_01[23:0], SP12_h_l_02[23:0],
     SP12_h_l_03[23:0], SP12_h_l_04[23:0], SP12_h_l_05[23:0],
     SP12_h_l_06[23:0], SP12_h_l_07[23:0], SP12_h_l_08[23:0], bl[17:0],
     pgate[127:0], reset_b[127:0], sp4_v_b_13_09[15:0],
     sp4_v_t_08[15:0], vdd_cntl[127:0], wl[127:0], bnl_op_13_09[7:0],
     bs_en, ceb, glb_netwk_col[7:0], hiz_b, hold,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[2],
     last_rsr[3], lft_op_01[7:0], lft_op_02[7:0], lft_op_03[7:0],
     lft_op_04[7:0], lft_op_05[7:0], lft_op_06[7:0], lft_op_07[7:0],
     lft_op_08[7:0], mode, mux_jtag_sel_b, padin[12:0], prog, r, sdi,
     sdo_enable, shift, tclk, tnl_op_08[7:0], totdopad, trstb_pad,
     update );
output  fabric_out_01, fabric_out_02, fabric_out_08, sdo, tck_pad,
     tclk_o, tdi_pad, tms_pad;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, mode, mux_jtag_sel_b, prog, r, sdi,
     sdo_enable, shift, tclk, totdopad, trstb_pad, update;

output [3:0]  slf_op_01;
output [3:0]  slf_op_08;
output [3:0]  slf_op_07;
output [3:0]  slf_op_02;
output [3:0]  slf_op_06;
output [12:0]  pado;
output [3:0]  slf_op_03;
output [191:0]  cf_r;
output [12:0]  padeb;
output [3:0]  slf_op_05;
output [3:0]  slf_op_04;

inout [23:0]  SP12_h_l_02;
inout [23:0]  SP12_h_l_06;
inout [23:0]  SP12_h_l_07;
inout [23:0]  SP12_h_l_03;
inout [47:0]  SP4_h_l_04;
inout [17:0]  bl;
inout [23:0]  SP12_h_l_04;
inout [47:0]  SP4_h_l_05;
inout [15:0]  sp4_v_t_08;
inout [47:0]  SP4_h_l_01;
inout [47:0]  SP4_h_l_06;
inout [47:0]  SP4_h_l_02;
inout [23:0]  SP12_h_l_05;
inout [47:0]  SP4_h_l_08;
inout [47:0]  SP4_h_l_03;
inout [15:0]  sp4_v_b_13_09;
inout [127:0]  reset_b;
inout [127:0]  vdd_cntl;
inout [127:0]  wl;
inout [23:0]  SP12_h_l_01;
inout [127:0]  pgate;
inout [23:0]  SP12_h_l_08;
inout [47:0]  SP4_h_l_07;

input [7:0]  lft_op_01;
input [7:0]  lft_op_06;
input [7:0]  lft_op_04;
input [7:0]  lft_op_03;
input [7:0]  lft_op_05;
input [7:0]  lft_op_07;
input [7:0]  lft_op_02;
input [7:0]  lft_op_08;
input [7:0]  tnl_op_08;
input [3:2]  last_rsr;
input [7:0]  bnl_op_13_09;
input [12:0]  padin;
input [7:0]  glb_netwk_col;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  net544;

wire  [15:0]  net400;

wire  [1:0]  net507;

wire  [7:0]  net584;

wire  [7:0]  glb_netwk_t;

wire  [36:11]  cf_rd;

wire  [1:0]  net345;

wire  [15:0]  net472;

wire  [7:0]  colbuf_cntl_t;

wire  [15:0]  net652;

wire  [1:0]  net350;

wire  [7:0]  net548;

wire  [7:0]  colbuf_cntl_b;

wire  [1:0]  net352;

wire  [15:0]  net580;

wire  [7:0]  net346;

wire  [1:0]  net344;

wire  [7:0]  net349;

wire  [15:0]  net616;

wire  [7:0]  net476;

wire  [1:0]  net360;

wire  [7:0]  glb_netwk_b;

wire  [1:0]  net363;

wire  [36:11]  cf_rp;

wire  [15:0]  net508;

wire  [1:0]  net361;

wire  [7:0]  net440;



mux2_hvt I_mux_jtagcf_2_ ( .in1(cf_rp[36]), .in0(vdd_),
     .out(cf_rd[36]), .sel(mux_jtag_sel_b));
mux2_hvt I_mux_jtagcf_1_ ( .in1(cf_rp[12]), .in0(vdd_),
     .out(cf_rd[12]), .sel(mux_jtag_sel_b));
mux2_hvt I_mux_jtagcf_0_ ( .in1(cf_rp[11]), .in0(vdd_),
     .out(cf_rd[11]), .sel(mux_jtag_sel_b));
bram_bufferx4 I_muxedjtagbuf_2_ ( .in(cf_rd[36]), .out(cf_r[36]));
bram_bufferx4 I_muxedjtagbuf_1_ ( .in(cf_rd[12]), .out(cf_r[12]));
bram_bufferx4 I_muxedjtagbuf_0_ ( .in(cf_rd[11]), .out(cf_r[11]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tiegnd));
tckbufx32_ice8p I_tmsbuf ( .in(tms), .out(tms_pad));
tckbufx32_ice8p I_tckbuf ( .in(tck), .out(tck_pad));
tckbufx32_ice8p I_tdibuf ( .in(tdi), .out(tdi_pad));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
io_col4_rgt_ice8p_v2 I_io_00_02 ( .slf_op(slf_op_02[3:0]),
     .cdone_in(trstb_pad), .spioeb({sdo_enable, tievdd}),
     .tnl_op(lft_op_03[7:0]), .spi_ss_in_b({nc_ss, tck}), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_02[23:0]),
     .spiout({totdopad, tiegnd}), .sp4_v_b({net580[0], net580[1],
     net580[2], net580[3], net580[4], net580[5], net580[6], net580[7],
     net580[8], net580[9], net580[10], net580[11], net580[12],
     net580[13], net580[14], net580[15]}), .prog(prog),
     .cf({cf_r[47:37], cf_rp[36], cf_r[35:24]}),
     .vdd_cntl(vdd_cntl[31:16]), .lft_op(lft_op_02[7:0]),
     .padin(padin[3:2]), .mode(mode), .wl(wl[31:16]), .pado(pado[3:2]),
     .sp4_v_t({net400[0], net400[1], net400[2], net400[3], net400[4],
     net400[5], net400[6], net400[7], net400[8], net400[9], net400[10],
     net400[11], net400[12], net400[13], net400[14], net400[15]}),
     .padeb(padeb[3:2]), .reset(reset_b[31:16]), .bl(bl[17:0]),
     .cbit_colcntl({net346[0], net346[1], net346[2], net346[3],
     net346[4], net346[5], net346[6], net346[7]}), .sdo(net405),
     .fabric_out(fabric_out_02), .glb_netwk(glb_netwk_b[7:0]),
     .pgate(pgate[31:16]), .sdi(net585), .sp4_h_l(SP4_h_l_02[47:0]),
     .bnl_op(lft_op_01[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_08 ( .slf_op(slf_op_08[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(tnl_op_08[7:0]), .spi_ss_in_b({net361[0], net361[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_08[23:0]), .spiout({tiegnd, tiegnd}),
     .sp4_v_b({net472[0], net472[1], net472[2], net472[3], net472[4],
     net472[5], net472[6], net472[7], net472[8], net472[9], net472[10],
     net472[11], net472[12], net472[13], net472[14], net472[15]}),
     .prog(prog), .cf(cf_r[191:168]), .vdd_cntl(vdd_cntl[127:112]),
     .lft_op(lft_op_08[7:0]), .padin(padin[12:11]), .mode(mode),
     .wl(wl[127:112]), .pado(pado[12:11]), .sp4_v_t(sp4_v_t_08[15:0]),
     .padeb(padeb[12:11]), .reset(reset_b[127:112]), .bl(bl[17:0]),
     .cbit_colcntl({net440[0], net440[1], net440[2], net440[3],
     net440[4], net440[5], net440[6], net440[7]}), .sdo(sdo),
     .fabric_out(fabric_out_08), .glb_netwk(glb_netwk_t[7:0]),
     .pgate(pgate[127:112]), .sdi(net477), .sp4_h_l(SP4_h_l_08[47:0]),
     .bnl_op(lft_op_07[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_07 ( .slf_op(slf_op_07[3:0]),
     .cdone_in(jtag_rowtest_mode_rowu3_b), .spioeb({tievdd, tiegnd}),
     .tnl_op(lft_op_08[7:0]), .spi_ss_in_b({net352[0], net352[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_07[23:0]), .spiout({tiegnd, last_rsr[3]}),
     .sp4_v_b({net544[0], net544[1], net544[2], net544[3], net544[4],
     net544[5], net544[6], net544[7], net544[8], net544[9], net544[10],
     net544[11], net544[12], net544[13], net544[14], net544[15]}),
     .prog(prog), .cf(cf_r[167:144]), .vdd_cntl(vdd_cntl[111:96]),
     .lft_op(lft_op_07[7:0]), .padin(padin[10:9]), .mode(mode),
     .wl(wl[111:96]), .pado(pado[10:9]), .sp4_v_t({net472[0],
     net472[1], net472[2], net472[3], net472[4], net472[5], net472[6],
     net472[7], net472[8], net472[9], net472[10], net472[11],
     net472[12], net472[13], net472[14], net472[15]}),
     .padeb(padeb[10:9]), .reset(reset_b[111:96]), .bl(bl[17:0]),
     .cbit_colcntl({net476[0], net476[1], net476[2], net476[3],
     net476[4], net476[5], net476[6], net476[7]}), .sdo(net477),
     .fabric_out(net478), .glb_netwk(glb_netwk_t[7:0]),
     .pgate(pgate[111:96]), .sdi(net549), .sp4_h_l(SP4_h_l_07[47:0]),
     .bnl_op(lft_op_06[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_05 ( .slf_op(slf_op_05[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_06[7:0]), .spi_ss_in_b({net345[0], net345[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_05[23:0]), .spiout({tiegnd, tiegnd}),
     .sp4_v_b({net652[0], net652[1], net652[2], net652[3], net652[4],
     net652[5], net652[6], net652[7], net652[8], net652[9], net652[10],
     net652[11], net652[12], net652[13], net652[14], net652[15]}),
     .prog(prog), .cf(cf_r[119:96]), .vdd_cntl(vdd_cntl[79:64]),
     .lft_op(lft_op_05[7:0]), .padin({net507[0], net507[1]}),
     .mode(mode), .wl(wl[79:64]), .pado({net507[0], net507[1]}),
     .sp4_v_t({net508[0], net508[1], net508[2], net508[3], net508[4],
     net508[5], net508[6], net508[7], net508[8], net508[9], net508[10],
     net508[11], net508[12], net508[13], net508[14], net508[15]}),
     .padeb({net363[0], net363[1]}), .reset(reset_b[79:64]),
     .bl(bl[17:0]), .cbit_colcntl(colbuf_cntl_t[7:0]), .sdo(net513),
     .fabric_out(net514), .glb_netwk(glb_netwk_t[7:0]),
     .pgate(pgate[79:64]), .sdi(net657), .sp4_h_l(SP4_h_l_05[47:0]),
     .bnl_op(lft_op_04[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_06 ( .slf_op(slf_op_06[3:0]),
     .cdone_in(jtag_rowtest_mode_rowu2_b), .spioeb({tievdd, tiegnd}),
     .tnl_op(lft_op_07[7:0]), .spi_ss_in_b({net360[0], net360[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_06[23:0]), .spiout({tiegnd, last_rsr[2]}),
     .sp4_v_b({net508[0], net508[1], net508[2], net508[3], net508[4],
     net508[5], net508[6], net508[7], net508[8], net508[9], net508[10],
     net508[11], net508[12], net508[13], net508[14], net508[15]}),
     .prog(prog), .cf(cf_r[143:120]), .vdd_cntl(vdd_cntl[95:80]),
     .lft_op(lft_op_06[7:0]), .padin(padin[8:7]), .mode(mode),
     .wl(wl[95:80]), .pado(pado[8:7]), .sp4_v_t({net544[0], net544[1],
     net544[2], net544[3], net544[4], net544[5], net544[6], net544[7],
     net544[8], net544[9], net544[10], net544[11], net544[12],
     net544[13], net544[14], net544[15]}), .padeb(padeb[8:7]),
     .reset(reset_b[95:80]), .bl(bl[17:0]), .cbit_colcntl({net548[0],
     net548[1], net548[2], net548[3], net548[4], net548[5], net548[6],
     net548[7]}), .sdo(net549), .fabric_out(net550),
     .glb_netwk(glb_netwk_t[7:0]), .pgate(pgate[95:80]), .sdi(net513),
     .sp4_h_l(SP4_h_l_06[47:0]), .bnl_op(lft_op_05[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_01 ( .slf_op(slf_op_01[3:0]),
     .cdone_in(mux_jtag_sel_b), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_02[7:0]), .spi_ss_in_b({tms, tdi}), .hold(hold),
     .update(update), .shift(shift), .hiz_b(hiz_b), .bs_en(bs_en),
     .r(r), .tclk(tclk_o), .ceb(ceb), .sp12_h_l(SP12_h_l_01[23:0]),
     .spiout({tiegnd, tiegnd}), .sp4_v_b(sp4_v_b_13_09[15:0]),
     .prog(prog), .cf({cf_r[23:13], cf_rp[12], cf_rp[11], cf_r[10:0]}),
     .vdd_cntl(vdd_cntl[15:0]), .lft_op(lft_op_01[7:0]),
     .padin(padin[1:0]), .mode(mode), .wl(wl[15:0]), .pado(pado[1:0]),
     .sp4_v_t({net580[0], net580[1], net580[2], net580[3], net580[4],
     net580[5], net580[6], net580[7], net580[8], net580[9], net580[10],
     net580[11], net580[12], net580[13], net580[14], net580[15]}),
     .padeb(padeb[1:0]), .reset(reset_b[15:0]), .bl(bl[17:0]),
     .cbit_colcntl({net584[0], net584[1], net584[2], net584[3],
     net584[4], net584[5], net584[6], net584[7]}), .sdo(net585),
     .fabric_out(fabric_out_01), .glb_netwk(glb_netwk_b[7:0]),
     .pgate(pgate[15:0]), .sdi(sdi), .sp4_h_l(SP4_h_l_01[47:0]),
     .bnl_op(bnl_op_13_09[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_03 ( .slf_op(slf_op_03[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_04[7:0]), .spi_ss_in_b({net350[0], net350[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_03[23:0]), .spiout({tiegnd, tiegnd}),
     .sp4_v_b({net400[0], net400[1], net400[2], net400[3], net400[4],
     net400[5], net400[6], net400[7], net400[8], net400[9], net400[10],
     net400[11], net400[12], net400[13], net400[14], net400[15]}),
     .prog(prog), .cf(cf_r[71:48]), .vdd_cntl(vdd_cntl[47:32]),
     .lft_op(lft_op_03[7:0]), .padin({padin[4], padin_nc}),
     .mode(mode), .wl(wl[47:32]), .pado({pado[4], pado_nc}),
     .sp4_v_t({net616[0], net616[1], net616[2], net616[3], net616[4],
     net616[5], net616[6], net616[7], net616[8], net616[9], net616[10],
     net616[11], net616[12], net616[13], net616[14], net616[15]}),
     .padeb({padeb[4], padeb_nc}), .reset(reset_b[47:32]),
     .bl(bl[17:0]), .cbit_colcntl({net349[0], net349[1], net349[2],
     net349[3], net349[4], net349[5], net349[6], net349[7]}),
     .sdo(net621), .fabric_out(net622), .glb_netwk(glb_netwk_b[7:0]),
     .pgate(pgate[47:32]), .sdi(net405), .sp4_h_l(SP4_h_l_03[47:0]),
     .bnl_op(lft_op_02[7:0]));
io_col4_rgt_ice8p_v2 I_io_00_04 ( .slf_op(slf_op_04[3:0]),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .tnl_op(lft_op_05[7:0]), .spi_ss_in_b({net344[0], net344[1]}),
     .hold(hold), .update(update), .shift(shift), .hiz_b(hiz_b),
     .bs_en(bs_en), .r(r), .tclk(tclk_o), .ceb(ceb),
     .sp12_h_l(SP12_h_l_04[23:0]), .spiout({tiegnd, tiegnd}),
     .sp4_v_b({net616[0], net616[1], net616[2], net616[3], net616[4],
     net616[5], net616[6], net616[7], net616[8], net616[9], net616[10],
     net616[11], net616[12], net616[13], net616[14], net616[15]}),
     .prog(prog), .cf(cf_r[95:72]), .vdd_cntl(vdd_cntl[63:48]),
     .lft_op(lft_op_04[7:0]), .padin(padin[6:5]), .mode(mode),
     .wl(wl[63:48]), .pado(pado[6:5]), .sp4_v_t({net652[0], net652[1],
     net652[2], net652[3], net652[4], net652[5], net652[6], net652[7],
     net652[8], net652[9], net652[10], net652[11], net652[12],
     net652[13], net652[14], net652[15]}), .padeb(padeb[6:5]),
     .reset(reset_b[63:48]), .bl(bl[17:0]),
     .cbit_colcntl(colbuf_cntl_b[7:0]), .sdo(net657),
     .fabric_out(net658), .glb_netwk(glb_netwk_b[7:0]),
     .pgate(pgate[63:48]), .sdi(net621), .sp4_h_l(SP4_h_l_04[47:0]),
     .bnl_op(lft_op_03[7:0]));

endmodule
// Library - ice8chip, Cell - io_col4_bot_ice8p, View - schematic
// LAST TIME SAVED: Jan 12 14:58:38 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module io_col4_bot_ice8p ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [23:0]  cf;
output [1:0]  pado;
output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [3:0]  slf_op;

inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;

input [1:0]  padin;
input [1:0]  spiout;
input [15:0]  reset;
input [15:0]  pgate;
input [7:0]  glb_netwk;
input [1:0]  spioeb;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [15:0]  wl;
input [15:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [7:0]  net225;



inv_lvt I_inv1 ( .A(prog), .Y(progb));
inv_lvt I_inv2 ( .A(progb), .Y(progd));
io_gmux_x16bare_v3 I_io_gmux_x16bare_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .lc_trk_g0(lc_trk_g0[7:0]), .bl(bl[9:4]),
     .prog(progd), .lc_trk_g1(lc_trk_g1[7:0]), .min7({sp4_h_l[47],
     sp4_h_l[39], sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7],
     sp12_h_l[23], sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7],
     bnl_op[7], lft_op[7], tnl_op[7], gnd_, gnd_}), .min6({sp4_h_l[46],
     sp4_h_l[38], sp4_h_l[30], sp4_h_l[22], sp4_h_l[14], sp4_h_l[6],
     sp12_h_l[22], sp12_h_l[14], sp12_h_l[6], sp4_v_b[14], sp4_v_b[6],
     bnl_op[6], lft_op[6], tnl_op[6], gnd_, gnd_}),
     .cbitb_colcntl({net225[0], net225[1], net225[2], net225[3],
     net225[4], net225[5], net225[6], net225[7]}),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .min5({sp4_h_l[45], sp4_h_l[37],
     sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5], sp12_h_l[21],
     sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5], bnl_op[5],
     lft_op[5], tnl_op[5], gnd_, gnd_}), .min4({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}), .min3({sp4_h_l[43],
     sp4_h_l[35], sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3],
     sp12_h_l[19], sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3],
     bnl_op[3], lft_op[3], tnl_op[3], gnd_, gnd_}), .min2({sp4_h_l[42],
     sp4_h_l[34], sp4_h_l[26], sp4_h_l[18], sp4_h_l[10], sp4_h_l[2],
     sp12_h_l[18], sp12_h_l[10], sp12_h_l[2], sp4_v_b[10], sp4_v_b[2],
     bnl_op[2], lft_op[2], tnl_op[2], gnd_, gnd_}), .min1({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}), .min0({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min8({sp4_h_l[40],
     sp4_h_l[32], sp4_h_l[24], sp4_h_l[16], sp4_h_l[8], sp4_h_l[0],
     sp12_h_l[16], sp12_h_l[8], sp12_h_l[0], sp4_v_b[8], sp4_v_b[0],
     bnl_op[0], lft_op[0], tnl_op[0], gnd_, gnd_}), .min9({sp4_h_l[41],
     sp4_h_l[33], sp4_h_l[25], sp4_h_l[17], sp4_h_l[9], sp4_h_l[1],
     sp12_h_l[17], sp12_h_l[9], sp12_h_l[1], sp4_v_b[9], sp4_v_b[1],
     bnl_op[1], lft_op[1], tnl_op[1], gnd_, gnd_}),
     .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min11({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27],
     sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11],
     sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3],
     tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44], sp4_h_l[36],
     sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4], sp12_h_l[20],
     sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4], bnl_op[4],
     lft_op[4], tnl_op[4], gnd_, gnd_}), .min13({sp4_h_l[45],
     sp4_h_l[37], sp4_h_l[29], sp4_h_l[21], sp4_h_l[13], sp4_h_l[5],
     sp12_h_l[21], sp12_h_l[13], sp12_h_l[5], sp4_v_b[13], sp4_v_b[5],
     bnl_op[5], lft_op[5], tnl_op[5], gnd_, gnd_}),
     .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min15({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31],
     sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15],
     sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7],
     tnl_op[7], gnd_, gnd_}));
io_col_odrv4_x40bare_v3 I_io_col_odrv4_x40bare_v3 ( cf[23:0], bl[3:0],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}, progd,
     {reset[14], reset[15], reset[12], reset[13], reset[10], reset[11],
     reset[8], reset[9], reset[6], reset[7], reset[4], reset[5],
     reset[2], reset[3], reset[0], reset[1]}, {vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}, {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11],
     wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0],
     wl[1]});
sbox1_colbdlc_v3 I_sbox1_colbdlc_v3 ( .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .reset({reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}), .prog(progd), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .outclk(outclk),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .fabric_out(fabric_out), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}));
ioe_col2_v3 I_ioe_col2_v3 ( .update(enable_update), .ti(ti[5:0]),
     .tclk(tclk), .shift(shift), .sdi(sdi), .prog(progd),
     .padin(padin[1:0]), .mode(mode), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .inclk(inclk), .outclk(outclk),
     .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo),
     .pado(om[1:0]), .padeb(oenm[1:0]), .ceb(ceb),
     .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12], vdd_cntl[13],
     vdd_cntl[10], vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6],
     vdd_cntl[7], vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3],
     vdd_cntl[0], vdd_cntl[1]}), .pgate({pgate[14], pgate[15],
     pgate[12], pgate[13], pgate[10], pgate[11], pgate[8], pgate[9],
     pgate[6], pgate[7], pgate[4], pgate[5], pgate[2], pgate[3],
     pgate[0], pgate[1]}), .bl(bl[17:16]), .dout(slf_op[3:0]),
     .hold(hold), .hiz_b(hiz_b), .rstio(r));
rm6w  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6w  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6w  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6w  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6w  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6w  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6w  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6w  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6w  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6w  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6w  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6w  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6w  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6w  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6w  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6w  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));

endmodule
// Library - ice1chip, Cell - io_bot_rgt_1x6_ice1f, View - schematic
// LAST TIME SAVED: May  3 12:10:20 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module io_bot_rgt_1x6_ice1f ( cf_b_r[143:0], fabric_out_07_00,
     fabric_out_12_00, padeb_b_r[11], padeb_b_r[23:13], pado_b_r[11],
     pado_b_r[23:13], sdo_pad, slf_op_01_00[3:0], slf_op_02_00[3:0],
     slf_op_03_00[3:0], slf_op_04_00[3:0], slf_op_05_00[3:0],
     slf_op_06_00[3:0], spi_ss_in_bbank[4:0], bl_01[53:0], bl_02[53:0],
     bl_03[53:0], bl_04[41:0], bl_05[53:0], bl_06[53:0],
     sp4_h_l_07_00[15:0], sp4_h_r_12_17[15:0], sp4_v_b_01_00[47:0],
     sp4_v_b_02_00[47:0], sp4_v_b_03_00[47:0], sp4_v_b_04_00[47:0],
     sp4_v_b_05_00[47:0], sp4_v_b_06_00[47:0], sp12_v_b_01_00[23:0],
     sp12_v_b_02_00[23:0], sp12_v_b_03_00[23:0], sp12_v_b_04_00[23:0],
     sp12_v_b_05_00[23:0], sp12_v_b_06_00[23:0], bnl_op_01_00[7:0],
     bs_en_i, ceb_i, end_of_startup, glb_net_01[7:0], glb_net_02[7:0],
     glb_net_03[7:0], glb_net_04[7:0], glb_net_05[7:0],
     glb_net_06[7:0], hiz_b_i, hold_b_r, lft_op_01_00[7:0],
     lft_op_02_00[7:0], lft_op_03_00[7:0], lft_op_04_00[7:0],
     lft_op_05_00[7:0], lft_op_06_00[7:0], md_spi_b, mode_i,
     padin_b_r[11], padin_b_r[23:13], pgate_l[15:0], prog, r_i,
     reset_l[15:0], sdi, shift_i, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk_i, tnr_op_06_00[7:0], update_i, vdd_cntl_l[15:0],
     wl_l[15:0] );
output  fabric_out_07_00, fabric_out_12_00, sdo_pad;


input  bs_en_i, ceb_i, end_of_startup, hiz_b_i, hold_b_r, md_spi_b,
     mode_i, prog, r_i, sdi, shift_i, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk_i, update_i;

output [3:0]  slf_op_05_00;
output [3:0]  slf_op_03_00;
output [3:0]  slf_op_06_00;
output [3:0]  slf_op_01_00;
output [3:0]  slf_op_04_00;
output [3:0]  slf_op_02_00;
output [4:0]  spi_ss_in_bbank;
output [23:11]  padeb_b_r;
output [143:0]  cf_b_r;
output [23:11]  pado_b_r;

inout [47:0]  sp4_v_b_01_00;
inout [47:0]  sp4_v_b_02_00;
inout [15:0]  sp4_h_r_12_17;
inout [47:0]  sp4_v_b_04_00;
inout [47:0]  sp4_v_b_06_00;
inout [23:0]  sp12_v_b_05_00;
inout [23:0]  sp12_v_b_02_00;
inout [23:0]  sp12_v_b_03_00;
inout [41:0]  bl_04;
inout [23:0]  sp12_v_b_01_00;
inout [47:0]  sp4_v_b_05_00;
inout [23:0]  sp12_v_b_06_00;
inout [53:0]  bl_02;
inout [53:0]  bl_03;
inout [53:0]  bl_05;
inout [53:0]  bl_06;
inout [23:0]  sp12_v_b_04_00;
inout [47:0]  sp4_v_b_03_00;
inout [15:0]  sp4_h_l_07_00;
inout [53:0]  bl_01;

input [15:0]  pgate_l;
input [7:0]  glb_net_02;
input [7:0]  lft_op_05_00;
input [7:0]  glb_net_03;
input [7:0]  glb_net_06;
input [15:0]  wl_l;
input [7:0]  glb_net_05;
input [7:0]  glb_net_01;
input [7:0]  lft_op_02_00;
input [7:0]  lft_op_01_00;
input [7:0]  bnl_op_01_00;
input [15:0]  reset_l;
input [7:0]  lft_op_03_00;
input [7:0]  glb_net_04;
input [7:0]  lft_op_04_00;
input [7:0]  lft_op_06_00;
input [23:11]  padin_b_r;
input [15:0]  vdd_cntl_l;
input [7:0]  tnr_op_06_00;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net543;

wire  [15:0]  net514;

wire  [1:0]  net545;

wire  [15:0]  net374;

wire  [1:0]  net546;

wire  [15:0]  net409;

wire  [132:83]  cf_b_r_pd;

wire  [15:0]  net444;

wire  [132:83]  cf_b_r_p;

wire  [15:0]  net339;



bram_bufferx4 I_cfbuf_spiss_ck_1_ ( .in(cf_b_r_pd[132]),
     .out(cf_b_r[132]));
bram_bufferx4 I_cfbuf_spiss_ck_0_ ( .in(cf_b_r_pd[131]),
     .out(cf_b_r[131]));
bram_bufferx4 I_buf_spisdi ( .in(cf_b_r_pd[107]), .out(cf_b_r[107]));
bram_bufferx4 I_buf_coldboot_1_ ( .in(cf_b_r_pd[84]),
     .out(cf_b_r[84]));
bram_bufferx4 I_buf_coldboot_0_ ( .in(cf_b_r_pd[83]),
     .out(cf_b_r[83]));
mux2_hvt I_cfmux_spiss_ck_1_ ( .in1(cf_b_r_p[132]), .in0(vdd_),
     .out(cf_b_r_pd[132]), .sel(end_of_startup));
mux2_hvt I_cfmux_spiss_ck_0_ ( .in1(cf_b_r_p[131]), .in0(vdd_),
     .out(cf_b_r_pd[131]), .sel(end_of_startup));
mux2_hvt I_cfmux_spisdi ( .in1(cf_b_r_p[107]), .in0(vdd_),
     .out(cf_b_r_pd[107]), .sel(end_of_startup));
mux2_hvt I_cfmux_coldboot_1_ ( .in1(cf_b_r_p[84]), .in0(vdd_),
     .out(cf_b_r_pd[84]), .sel(end_of_startup));
mux2_hvt I_cfmux_coldboot_0_ ( .in1(cf_b_r_p[83]), .in0(vdd_),
     .out(cf_b_r_pd[83]), .sel(end_of_startup));
bram_bufferx4x6 I_bram_bufferx4x6 ( .in(net463), .out(net301));
lowla_modified I_lowla_modified ( .clk(endtck), .min(net301),
     .lao(sdo_pad));
scan_buf_ice8p I_scanbuf_8p_mb ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net314), .tclk_o(net315), .shift_o(net316),
     .sdo(net317), .r_o(net318), .mode_o(net319), .hiz_b_o(net320),
     .ceb_o(net321), .bs_en_o(net322));
io_col4_bot_ice8p I_IO_08_00 ( .sdo(net323), .sdi(net393),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net409[0], net409[1], net409[2], net409[3],
     net409[4], net409[5], net409[6], net409[7], net409[8], net409[9],
     net409[10], net409[11], net409[12], net409[13], net409[14],
     net409[15]}), .mode(net319), .shift(net316), .hiz_b(net320),
     .r(net318), .bs_en(net322), .tclk(endtck), .update(net314),
     .padin(padin_b_r[15:14]), .pado(pado_b_r[15:14]),
     .padeb(padeb_b_r[15:14]), .sp4_v_b({net339[0], net339[1],
     net339[2], net339[3], net339[4], net339[5], net339[6], net339[7],
     net339[8], net339[9], net339[10], net339[11], net339[12],
     net339[13], net339[14], net339[15]}),
     .sp4_h_l(sp4_v_b_02_00[47:0]), .sp12_h_l(sp12_v_b_02_00[23:0]),
     .prog(prog), .spi_ss_in_b({net545[0], net545[1]}),
     .tnl_op(lft_op_01_00[7:0]), .lft_op(lft_op_02_00[7:0]),
     .bnl_op(lft_op_03_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_02[5], bl_02[4], bl_02[37],
     bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32], bl_02[14],
     bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16], bl_02[27],
     bl_02[26], bl_02[25], bl_02[23]}), .wl(wl_l[15:0]),
     .cf(cf_b_r[47:24]), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_00[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_b_r), .fabric_out(net357));
io_col4_bot_ice8p I_IO_10_00_bram ( .sdo(net358), .sdi(net498),
     .spiout({tielow, tielow}), .cdone_in(end_of_startup),
     .spioeb({tievdd, tievdd}), .sp4_v_t({net514[0], net514[1],
     net514[2], net514[3], net514[4], net514[5], net514[6], net514[7],
     net514[8], net514[9], net514[10], net514[11], net514[12],
     net514[13], net514[14], net514[15]}), .mode(net319),
     .shift(net316), .hiz_b(net320), .r(net318), .bs_en(net322),
     .tclk(endtck), .update(net314), .padin(padin_b_r[19:18]),
     .pado(pado_b_r[19:18]), .padeb(padeb_b_r[19:18]),
     .sp4_v_b({net374[0], net374[1], net374[2], net374[3], net374[4],
     net374[5], net374[6], net374[7], net374[8], net374[9], net374[10],
     net374[11], net374[12], net374[13], net374[14], net374[15]}),
     .sp4_h_l(sp4_v_b_04_00[47:0]), .sp12_h_l(sp12_v_b_04_00[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_bbank[1:0]),
     .tnl_op(lft_op_03_00[7:0]), .lft_op(lft_op_04_00[7:0]),
     .bnl_op(lft_op_05_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_04[5], bl_04[4], bl_04[37],
     bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32], bl_04[14],
     bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16], bl_04[27],
     bl_04[26], bl_04[25], bl_04[23]}), .wl(wl_l[15:0]),
     .cf({cf_b_r[95:85], cf_b_r_p[84:83], cf_b_r[82:72]}),
     .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_00[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_b_r), .fabric_out(net392));
io_col4_bot_ice8p I_IO_07_00 ( .sdo(net393), .sdi(net317),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_07_00[15:0]), .mode(net319),
     .shift(net316), .hiz_b(net320), .r(net318), .bs_en(net322),
     .tclk(endtck), .update(net314), .padin({padin_b_r[13],
     padin_b_r[11]}), .pado({pado_b_r[13], pado_b_r[11]}),
     .padeb({padeb_b_r[13], padeb_b_r[11]}), .sp4_v_b({net409[0],
     net409[1], net409[2], net409[3], net409[4], net409[5], net409[6],
     net409[7], net409[8], net409[9], net409[10], net409[11],
     net409[12], net409[13], net409[14], net409[15]}),
     .sp4_h_l(sp4_v_b_01_00[47:0]), .sp12_h_l(sp12_v_b_01_00[23:0]),
     .prog(prog), .spi_ss_in_b({net546[0], net546[1]}),
     .tnl_op(bnl_op_01_00[7:0]), .lft_op(lft_op_01_00[7:0]),
     .bnl_op(lft_op_02_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_b_r[23:0]), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_00[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_b_r), .fabric_out(fabric_out_07_00));
io_col4_bot_ice8p I_IO_11_00 ( .sdo(net428), .sdi(net358),
     .spiout({tielow, spi_sdo}), .cdone_in(end_of_startup),
     .spioeb({tievdd, spi_sdo_oe_b}), .sp4_v_t({net374[0], net374[1],
     net374[2], net374[3], net374[4], net374[5], net374[6], net374[7],
     net374[8], net374[9], net374[10], net374[11], net374[12],
     net374[13], net374[14], net374[15]}), .mode(net319),
     .shift(net316), .hiz_b(net320), .r(net318), .bs_en(net322),
     .tclk(endtck), .update(net314), .padin(padin_b_r[21:20]),
     .pado(pado_b_r[21:20]), .padeb(padeb_b_r[21:20]),
     .sp4_v_b({net444[0], net444[1], net444[2], net444[3], net444[4],
     net444[5], net444[6], net444[7], net444[8], net444[9], net444[10],
     net444[11], net444[12], net444[13], net444[14], net444[15]}),
     .sp4_h_l(sp4_v_b_05_00[47:0]), .sp12_h_l(sp12_v_b_05_00[23:0]),
     .prog(prog), .spi_ss_in_b({spi_ss_in_bbank[2], spi_ss_nc}),
     .tnl_op(lft_op_04_00[7:0]), .lft_op(lft_op_05_00[7:0]),
     .bnl_op(lft_op_06_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_05[5], bl_05[4], bl_05[37],
     bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32], bl_05[14],
     bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16], bl_05[27],
     bl_05[26], bl_05[25], bl_05[23]}), .wl(wl_l[15:0]),
     .cf({cf_b_r[119:108], cf_b_r_p[107], cf_b_r[106:96]}),
     .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_00[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_b_r), .fabric_out(net462));
io_col4_bot_ice8p I_IO_12_00 ( .sdo(net463), .sdi(net428),
     .spiout({spi_ss_out, spi_clk_out}), .cdone_in(end_of_startup),
     .spioeb({md_spi_b, md_spi_b}), .sp4_v_t({net444[0], net444[1],
     net444[2], net444[3], net444[4], net444[5], net444[6], net444[7],
     net444[8], net444[9], net444[10], net444[11], net444[12],
     net444[13], net444[14], net444[15]}), .mode(net319),
     .shift(net316), .hiz_b(net320), .r(net318), .bs_en(net322),
     .tclk(endtck), .update(net314), .padin(padin_b_r[23:22]),
     .pado(pado_b_r[23:22]), .padeb(padeb_b_r[23:22]),
     .sp4_v_b(sp4_h_r_12_17[15:0]), .sp4_h_l(sp4_v_b_06_00[47:0]),
     .sp12_h_l(sp12_v_b_06_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_bbank[4:3]), .tnl_op(lft_op_05_00[7:0]),
     .lft_op(lft_op_06_00[7:0]), .bnl_op(tnr_op_06_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_l[15:0]), .cf({cf_b_r[143:133], cf_b_r_p[132:131],
     cf_b_r[130:120]}), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_00[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_b_r), .fabric_out(fabric_out_12_00));
io_col4_bot_ice8p I_IO_09_00 ( .sdo(net498), .sdi(net323),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net339[0], net339[1], net339[2], net339[3],
     net339[4], net339[5], net339[6], net339[7], net339[8], net339[9],
     net339[10], net339[11], net339[12], net339[13], net339[14],
     net339[15]}), .mode(net319), .shift(net316), .hiz_b(net320),
     .r(net318), .bs_en(net322), .tclk(endtck), .update(net314),
     .padin(padin_b_r[17:16]), .pado(pado_b_r[17:16]),
     .padeb(padeb_b_r[17:16]), .sp4_v_b({net514[0], net514[1],
     net514[2], net514[3], net514[4], net514[5], net514[6], net514[7],
     net514[8], net514[9], net514[10], net514[11], net514[12],
     net514[13], net514[14], net514[15]}),
     .sp4_h_l(sp4_v_b_03_00[47:0]), .sp12_h_l(sp12_v_b_03_00[23:0]),
     .prog(prog), .spi_ss_in_b({net543[0], net543[1]}),
     .tnl_op(lft_op_02_00[7:0]), .lft_op(lft_op_03_00[7:0]),
     .bnl_op(lft_op_04_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_03[5], bl_03[4], bl_03[37],
     bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32], bl_03[14],
     bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16], bl_03[27],
     bl_03[26], bl_03[25], bl_03[23]}), .wl(wl_l[15:0]),
     .cf(cf_b_r[71:48]), .ceb(net321), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_00[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_b_r), .fabric_out(net544));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(net315), .out(endtck));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));

endmodule
// Library - ice1chip, Cell - lt_1x8_bot_ice1f, View - schematic
// LAST TIME SAVED: Mar  9 14:57:57 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module lt_1x8_bot_ice1f ( carry_out, glb_netwk_bot, op_vic, slf_op_01,
     slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07,
     slf_op_08, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02, sp4_h_l_03,
     sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07, sp4_h_l_08,
     sp4_h_r_01, sp4_h_r_02, sp4_h_r_03, sp4_h_r_04, sp4_h_r_05,
     sp4_h_r_06, sp4_h_r_07, sp4_h_r_08, sp4_r_v_b_01, sp4_r_v_b_02,
     sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05, sp4_r_v_b_06,
     sp4_r_v_b_07, sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03,
     sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07, sp4_v_b_08,
     sp4_v_t_08, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04,
     sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_r_01,
     sp12_h_r_02, sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06,
     sp12_h_r_07, sp12_h_r_08, sp12_v_b_01, sp12_v_t_08, vdd_cntl, wl,
     bnl_op_01, bnr_op_01, bot_op_01, carry_in, glb_netwk_col, lc_bot,
     lft_op_01, lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06,
     lft_op_07, lft_op_08, prog, purst, rgt_op_01, rgt_op_02,
     rgt_op_03, rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08,
     tnl_op_08, tnr_op_08, top_op_08 );
output  carry_out, op_vic;


input  carry_in, lc_bot, prog, purst;

output [7:0]  slf_op_07;
output [7:0]  slf_op_02;
output [7:0]  slf_op_08;
output [7:0]  slf_op_06;
output [7:0]  slf_op_05;
output [7:0]  slf_op_01;
output [7:0]  glb_netwk_bot;
output [7:0]  slf_op_04;
output [7:0]  slf_op_03;

inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_r_v_b_04;
inout [23:0]  sp12_h_l_05;
inout [23:0]  sp12_h_r_01;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_v_b_06;
inout [47:0]  sp4_h_l_07;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_r_v_b_05;
inout [47:0]  sp4_h_l_04;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_h_l_02;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_h_r_03;
inout [23:0]  sp12_h_r_08;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_v_t_08;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_v_b_03;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_r_v_b_08;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_v_b_05;
inout [23:0]  sp12_h_l_04;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_h_l_06;
inout [127:0]  pgate;
inout [127:0]  wl;
inout [127:0]  vdd_cntl;
inout [127:0]  reset_b;
inout [47:0]  sp4_v_b_07;
inout [23:0]  sp12_h_r_02;
inout [23:0]  sp12_v_t_08;
inout [23:0]  sp12_v_b_01;
inout [23:0]  sp12_h_l_08;
inout [53:0]  bl;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_h_r_08;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_r_v_b_06;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_h_r_05;
inout [23:0]  sp12_h_r_03;

input [7:0]  rgt_op_08;
input [7:0]  lft_op_01;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_07;
input [7:0]  lft_op_05;
input [7:0]  glb_netwk_col;
input [7:0]  top_op_08;
input [7:0]  lft_op_02;
input [7:0]  lft_op_08;
input [7:0]  lft_op_07;
input [7:0]  lft_op_06;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_06;
input [7:0]  bot_op_01;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_02;
input [7:0]  tnl_op_08;
input [7:0]  rgt_op_04;
input [7:0]  lft_op_03;
input [7:0]  lft_op_04;
input [7:0]  bnr_op_01;
input [7:0]  bnl_op_01;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  net944;

wire  [7:0]  colbuf_cntl_bot;

wire  [7:0]  colbuf_cntl_top;

wire  [7:0]  glb_netwk_top;

wire  [7:0]  net1118;

wire  [7:0]  net0755;

wire  [23:0]  net1006;

wire  [7:0]  net932;

wire  [7:0]  net963;

wire  [7:0]  net1056;

wire  [23:0]  net1130;

wire  [23:0]  net975;

wire  [7:0]  net1087;

wire  [23:0]  net1037;

wire  [23:0]  net1068;

wire  [23:0]  net1099;



ltile4_ice8p_v1 I_LT06 ( .cntl_cbit({net963[0], net963[1], net963[2],
     net963[3], net963[4], net963[5], net963[6], net963[7]}),
     .op_bot(net996), .op_vic(net965), .prog(prog), .carry_out(net967),
     .lft_op(lft_op_06[7:0]), .sp12_h_l(sp12_h_l_06[23:0]),
     .sp4_h_l(sp4_h_l_06[47:0]), .sp4_v_b(sp4_v_b_06[47:0]),
     .sp12_v_b({net1006[0], net1006[1], net1006[2], net1006[3],
     net1006[4], net1006[5], net1006[6], net1006[7], net1006[8],
     net1006[9], net1006[10], net1006[11], net1006[12], net1006[13],
     net1006[14], net1006[15], net1006[16], net1006[17], net1006[18],
     net1006[19], net1006[20], net1006[21], net1006[22], net1006[23]}),
     .sp12_h_r(sp12_h_r_06[23:0]), .sp4_h_r(sp4_h_r_06[47:0]),
     .sp12_v_t({net975[0], net975[1], net975[2], net975[3], net975[4],
     net975[5], net975[6], net975[7], net975[8], net975[9], net975[10],
     net975[11], net975[12], net975[13], net975[14], net975[15],
     net975[16], net975[17], net975[18], net975[19], net975[20],
     net975[21], net975[22], net975[23]}), .sp4_v_t(sp4_v_b_07[47:0]),
     .sp4_r_v_b(sp4_r_v_b_06[47:0]), .wl(wl[95:80]),
     .top_op(slf_op_07[7:0]), .rgt_op(rgt_op_06[7:0]),
     .bot_op(slf_op_05[7:0]), .bl(bl[53:0]), .reset_b(reset_b[95:80]),
     .vdd_cntl(vdd_cntl[95:80]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net998), .purst(purst), .slf_op(slf_op_06[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_05[7:0]),
     .bnl_op(lft_op_05[7:0]), .tnr_op(rgt_op_07[7:0]),
     .tnl_op(lft_op_07[7:0]));
ltile4_ice8p_v1 I_LT03 ( .cntl_cbit({net1056[0], net1056[1],
     net1056[2], net1056[3], net1056[4], net1056[5], net1056[6],
     net1056[7]}), .op_bot(net1089), .op_vic(net1058), .prog(prog),
     .carry_out(net1060), .lft_op(lft_op_03[7:0]),
     .sp12_h_l(sp12_h_l_03[23:0]), .sp4_h_l(sp4_h_l_03[47:0]),
     .sp4_v_b(sp4_v_b_03[47:0]), .sp12_v_b({net1099[0], net1099[1],
     net1099[2], net1099[3], net1099[4], net1099[5], net1099[6],
     net1099[7], net1099[8], net1099[9], net1099[10], net1099[11],
     net1099[12], net1099[13], net1099[14], net1099[15], net1099[16],
     net1099[17], net1099[18], net1099[19], net1099[20], net1099[21],
     net1099[22], net1099[23]}), .sp12_h_r(sp12_h_r_03[23:0]),
     .sp4_h_r(sp4_h_r_03[47:0]), .sp12_v_t({net1068[0], net1068[1],
     net1068[2], net1068[3], net1068[4], net1068[5], net1068[6],
     net1068[7], net1068[8], net1068[9], net1068[10], net1068[11],
     net1068[12], net1068[13], net1068[14], net1068[15], net1068[16],
     net1068[17], net1068[18], net1068[19], net1068[20], net1068[21],
     net1068[22], net1068[23]}), .sp4_v_t(sp4_v_b_04[47:0]),
     .sp4_r_v_b(sp4_r_v_b_03[47:0]), .wl(wl[47:32]),
     .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net1091), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4_ice8p_v1 I_LT04 ( .cntl_cbit(colbuf_cntl_bot[7:0]),
     .op_bot(net1058), .op_vic(net1027), .prog(prog),
     .carry_out(net1029), .lft_op(lft_op_04[7:0]),
     .sp12_h_l(sp12_h_l_04[23:0]), .sp4_h_l(sp4_h_l_04[47:0]),
     .sp4_v_b(sp4_v_b_04[47:0]), .sp12_v_b({net1068[0], net1068[1],
     net1068[2], net1068[3], net1068[4], net1068[5], net1068[6],
     net1068[7], net1068[8], net1068[9], net1068[10], net1068[11],
     net1068[12], net1068[13], net1068[14], net1068[15], net1068[16],
     net1068[17], net1068[18], net1068[19], net1068[20], net1068[21],
     net1068[22], net1068[23]}), .sp12_h_r(sp12_h_r_04[23:0]),
     .sp4_h_r(sp4_h_r_04[47:0]), .sp12_v_t({net1037[0], net1037[1],
     net1037[2], net1037[3], net1037[4], net1037[5], net1037[6],
     net1037[7], net1037[8], net1037[9], net1037[10], net1037[11],
     net1037[12], net1037[13], net1037[14], net1037[15], net1037[16],
     net1037[17], net1037[18], net1037[19], net1037[20], net1037[21],
     net1037[22], net1037[23]}), .sp4_v_t(sp4_v_b_05[47:0]),
     .sp4_r_v_b(sp4_r_v_b_04[47:0]), .wl(wl[63:48]),
     .top_op(slf_op_05[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net1060), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(rgt_op_05[7:0]),
     .tnl_op(lft_op_05[7:0]));
ltile4_ice8p_v1 I_LT05 ( .cntl_cbit(colbuf_cntl_top[7:0]),
     .op_bot(net1027), .op_vic(net996), .prog(prog),
     .carry_out(net998), .lft_op(lft_op_05[7:0]),
     .sp12_h_l(sp12_h_l_05[23:0]), .sp4_h_l(sp4_h_l_05[47:0]),
     .sp4_v_b(sp4_v_b_05[47:0]), .sp12_v_b({net1037[0], net1037[1],
     net1037[2], net1037[3], net1037[4], net1037[5], net1037[6],
     net1037[7], net1037[8], net1037[9], net1037[10], net1037[11],
     net1037[12], net1037[13], net1037[14], net1037[15], net1037[16],
     net1037[17], net1037[18], net1037[19], net1037[20], net1037[21],
     net1037[22], net1037[23]}), .sp12_h_r(sp12_h_r_05[23:0]),
     .sp4_h_r(sp4_h_r_05[47:0]), .sp12_v_t({net1006[0], net1006[1],
     net1006[2], net1006[3], net1006[4], net1006[5], net1006[6],
     net1006[7], net1006[8], net1006[9], net1006[10], net1006[11],
     net1006[12], net1006[13], net1006[14], net1006[15], net1006[16],
     net1006[17], net1006[18], net1006[19], net1006[20], net1006[21],
     net1006[22], net1006[23]}), .sp4_v_t(sp4_v_b_06[47:0]),
     .sp4_r_v_b(sp4_r_v_b_05[47:0]), .wl(wl[79:64]),
     .top_op(slf_op_06[7:0]), .rgt_op(rgt_op_05[7:0]),
     .bot_op(slf_op_04[7:0]), .bl(bl[53:0]), .reset_b(reset_b[79:64]),
     .vdd_cntl(vdd_cntl[79:64]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net1029), .purst(purst), .slf_op(slf_op_05[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_04[7:0]),
     .bnl_op(lft_op_04[7:0]), .tnr_op(rgt_op_06[7:0]),
     .tnl_op(lft_op_06[7:0]));
ltile4_ice8p_v1 I_LT01 ( .cntl_cbit({net1118[0], net1118[1],
     net1118[2], net1118[3], net1118[4], net1118[5], net1118[6],
     net1118[7]}), .op_bot(lc_bot), .op_vic(net1120), .prog(prog),
     .carry_out(net1122), .lft_op(lft_op_01[7:0]),
     .sp12_h_l(sp12_h_l_01[23:0]), .sp4_h_l(sp4_h_l_01[47:0]),
     .sp4_v_b(sp4_v_b_01[47:0]), .sp12_v_b(sp12_v_b_01[23:0]),
     .sp12_h_r(sp12_h_r_01[23:0]), .sp4_h_r(sp4_h_r_01[47:0]),
     .sp12_v_t({net1130[0], net1130[1], net1130[2], net1130[3],
     net1130[4], net1130[5], net1130[6], net1130[7], net1130[8],
     net1130[9], net1130[10], net1130[11], net1130[12], net1130[13],
     net1130[14], net1130[15], net1130[16], net1130[17], net1130[18],
     net1130[19], net1130[20], net1130[21], net1130[22], net1130[23]}),
     .sp4_v_t(sp4_v_b_02[47:0]), .sp4_r_v_b(sp4_r_v_b_01[47:0]),
     .wl(wl[15:0]), .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4_ice8p_v1 I_LT02 ( .cntl_cbit({net1087[0], net1087[1],
     net1087[2], net1087[3], net1087[4], net1087[5], net1087[6],
     net1087[7]}), .op_bot(net1120), .op_vic(net1089), .prog(prog),
     .carry_out(net1091), .lft_op(lft_op_02[7:0]),
     .sp12_h_l(sp12_h_l_02[23:0]), .sp4_h_l(sp4_h_l_02[47:0]),
     .sp4_v_b(sp4_v_b_02[47:0]), .sp12_v_b({net1130[0], net1130[1],
     net1130[2], net1130[3], net1130[4], net1130[5], net1130[6],
     net1130[7], net1130[8], net1130[9], net1130[10], net1130[11],
     net1130[12], net1130[13], net1130[14], net1130[15], net1130[16],
     net1130[17], net1130[18], net1130[19], net1130[20], net1130[21],
     net1130[22], net1130[23]}), .sp12_h_r(sp12_h_r_02[23:0]),
     .sp4_h_r(sp4_h_r_02[47:0]), .sp12_v_t({net1099[0], net1099[1],
     net1099[2], net1099[3], net1099[4], net1099[5], net1099[6],
     net1099[7], net1099[8], net1099[9], net1099[10], net1099[11],
     net1099[12], net1099[13], net1099[14], net1099[15], net1099[16],
     net1099[17], net1099[18], net1099[19], net1099[20], net1099[21],
     net1099[22], net1099[23]}), .sp4_v_t(sp4_v_b_03[47:0]),
     .sp4_r_v_b(sp4_r_v_b_02[47:0]), .wl(wl[31:16]),
     .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk_bot[7:0]),
     .carry_in(net1122), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));
ltile4_ice8p_v1 I_LT08 ( .cntl_cbit({net0755[0], net0755[1],
     net0755[2], net0755[3], net0755[4], net0755[5], net0755[6],
     net0755[7]}), .op_bot(net934), .op_vic(op_vic), .prog(prog),
     .carry_out(carry_out), .lft_op(lft_op_08[7:0]),
     .sp12_h_l(sp12_h_l_08[23:0]), .sp4_h_l(sp4_h_l_08[47:0]),
     .sp4_v_b(sp4_v_b_08[47:0]), .sp12_v_b({net944[0], net944[1],
     net944[2], net944[3], net944[4], net944[5], net944[6], net944[7],
     net944[8], net944[9], net944[10], net944[11], net944[12],
     net944[13], net944[14], net944[15], net944[16], net944[17],
     net944[18], net944[19], net944[20], net944[21], net944[22],
     net944[23]}), .sp12_h_r(sp12_h_r_08[23:0]),
     .sp4_h_r(sp4_h_r_08[47:0]), .sp12_v_t(sp12_v_t_08[23:0]),
     .sp4_v_t(sp4_v_t_08[47:0]), .sp4_r_v_b(sp4_r_v_b_08[47:0]),
     .wl(wl[127:112]), .top_op(top_op_08[7:0]),
     .rgt_op(rgt_op_08[7:0]), .bot_op(slf_op_07[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[127:112]), .vdd_cntl(vdd_cntl[127:112]),
     .glb_netwk(glb_netwk_top[7:0]), .carry_in(net936), .purst(purst),
     .slf_op(slf_op_08[7:0]), .pgate(pgate[127:112]),
     .bnr_op(rgt_op_07[7:0]), .bnl_op(lft_op_07[7:0]),
     .tnr_op(tnr_op_08[7:0]), .tnl_op(tnl_op_08[7:0]));
ltile4_ice8p_v1 I_LT07 ( .cntl_cbit({net932[0], net932[1], net932[2],
     net932[3], net932[4], net932[5], net932[6], net932[7]}),
     .op_bot(net965), .op_vic(net934), .prog(prog), .carry_out(net936),
     .lft_op(lft_op_07[7:0]), .sp12_h_l(sp12_h_l_07[23:0]),
     .sp4_h_l(sp4_h_l_07[47:0]), .sp4_v_b(sp4_v_b_07[47:0]),
     .sp12_v_b({net975[0], net975[1], net975[2], net975[3], net975[4],
     net975[5], net975[6], net975[7], net975[8], net975[9], net975[10],
     net975[11], net975[12], net975[13], net975[14], net975[15],
     net975[16], net975[17], net975[18], net975[19], net975[20],
     net975[21], net975[22], net975[23]}),
     .sp12_h_r(sp12_h_r_07[23:0]), .sp4_h_r(sp4_h_r_07[47:0]),
     .sp12_v_t({net944[0], net944[1], net944[2], net944[3], net944[4],
     net944[5], net944[6], net944[7], net944[8], net944[9], net944[10],
     net944[11], net944[12], net944[13], net944[14], net944[15],
     net944[16], net944[17], net944[18], net944[19], net944[20],
     net944[21], net944[22], net944[23]}), .sp4_v_t(sp4_v_b_08[47:0]),
     .sp4_r_v_b(sp4_r_v_b_07[47:0]), .wl(wl[111:96]),
     .top_op(slf_op_08[7:0]), .rgt_op(rgt_op_07[7:0]),
     .bot_op(slf_op_06[7:0]), .bl(bl[53:0]), .reset_b(reset_b[111:96]),
     .vdd_cntl(vdd_cntl[111:96]), .glb_netwk(glb_netwk_top[7:0]),
     .carry_in(net967), .purst(purst), .slf_op(slf_op_07[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_06[7:0]),
     .bnl_op(lft_op_06[7:0]), .tnr_op(rgt_op_08[7:0]),
     .tnl_op(lft_op_08[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_bot (
     .colbuf_cntl(colbuf_cntl_bot[7:0]), .col_clk(glb_netwk_bot[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_top (
     .colbuf_cntl(colbuf_cntl_top[7:0]), .col_clk(glb_netwk_top[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - clkbuffer200u, View - schematic
// LAST TIME SAVED: Jun 30 10:54:26 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module clkbuffer200u ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - ice1chip, Cell - quad_br_ice1, View - schematic
// LAST TIME SAVED: May  3 12:05:59 2011
// NETLIST TIME: May  5 11:56:43 2011
`timescale 1ns / 1ns 

module quad_br_ice1 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o[7:0],
     bm_sclk_o, bm_sclkrw_o[1:0], bm_sdi_o[1:0], bm_sdo_o[1:0],
     bm_sreb_o, bm_sweb_o[1:0], bm_wdummymux_en_o, bs_en_o,
     carry_out_07_08, carry_out_08_08, carry_out_09_08,
     carry_out_11_08, carry_out_12_08, ceb_o, cf_b_r[143:0],
     cf_r[191:0], fabric_out_07_00, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fabric_out_13_08, hiz_b_o, mode_o, op_vic_07_08,
     op_vic_08_08, op_vic_09_08, op_vic_11_08, op_vic_12_08,
     padeb_b_r[11], padeb_b_r[23:13], padeb_r[12:0], padin_07_00a,
     padin_13_08b, pado_b_r[11], pado_b_r[23:13], pado_r[12:0], r_o,
     sdo, sdo_pad, shift_o, slf_op_07_00[3:0], slf_op_07_01[7:0],
     slf_op_07_02[7:0], slf_op_07_03[7:0], slf_op_07_04[7:0],
     slf_op_07_05[7:0], slf_op_07_06[7:0], slf_op_07_07[7:0],
     slf_op_07_08[7:0], slf_op_08_08[7:0], slf_op_09_08[7:0],
     slf_op_10_08[7:0], slf_op_11_08[7:0], slf_op_12_08[7:0],
     slf_op_13_08[3:0], spi_ss_in_bbank[4:0], tck_pad, tclk_o, tdi_pad,
     tms_pad, update_o, bl[329:0], pgate_r[143:0], reset_b_r[143:0],
     sp4_h_l_07_00[15:0], sp4_h_l_07_01[47:0], sp4_h_l_07_02[47:0],
     sp4_h_l_07_03[47:0], sp4_h_l_07_04[47:0], sp4_h_l_07_05[47:0],
     sp4_h_l_07_06[47:0], sp4_h_l_07_07[47:0], sp4_h_l_07_08[47:0],
     sp4_v_b_07_01[47:0], sp4_v_b_07_02[47:0], sp4_v_b_07_03[47:0],
     sp4_v_b_07_04[47:0], sp4_v_b_07_05[47:0], sp4_v_b_07_06[47:0],
     sp4_v_b_07_07[47:0], sp4_v_b_07_08[47:0], sp4_v_t_07_08[47:0],
     sp4_v_t_08_08[47:0], sp4_v_t_09_08[47:0], sp4_v_t_10_08[47:0],
     sp4_v_t_11_08[47:0], sp4_v_t_12_08[47:0], sp4_v_t_13_08[15:0],
     sp12_h_l_07_01[23:0], sp12_h_l_07_02[23:0], sp12_h_l_07_03[23:0],
     sp12_h_l_07_04[23:0], sp12_h_l_07_05[23:0], sp12_h_l_07_06[23:0],
     sp12_h_l_07_07[23:0], sp12_h_l_07_08[23:0], sp12_v_t_07_08[23:0],
     sp12_v_t_08_08[23:0], sp12_v_t_09_08[23:0], sp12_v_t_10_08[23:0],
     sp12_v_t_11_08[23:0], sp12_v_t_12_08[23:0], vdd_cntl_r[143:0],
     wl_r[143:0], bm_aa_top[10:0], bm_ab_top[10:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i[1:0],
     bm_sdi_i[1:0], bm_sdo_i[1:0], bm_sreb_i, bm_sweb_i[1:0],
     bm_wdummymux_en_i, bnl_op_07_01[3:0], bs_en_i, bs_en_mi, ceb_i,
     ceb_mi, end_of_startup, glb_in[7:0], hiz_b_i, hiz_b_mi, hold_b_r,
     hold_r_b, jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     last_rsr[2], last_rsr[3], lft_op_07_01[7:0], lft_op_07_02[7:0],
     lft_op_07_03[7:0], lft_op_07_04[7:0], lft_op_07_05[7:0],
     lft_op_07_06[7:0], lft_op_07_07[7:0], lft_op_07_08[7:0], md_spi_b,
     mode_i, mode_mi, mux_jtag_sel_b, padin_b_r[11], padin_b_r[23:13],
     padin_r[12:0], pll_sdo, prog, purst, r_i, r_mi, sdi, sdi_pad,
     sdo_enable, shift_i, shift_mi, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk_i, tclk_mi, tnl_op_07_08[7:0], tnl_op_08_08[7:0],
     tnl_op_09_08[7:0], tnl_op_10_08[7:0], tnl_op_11_08[7:0],
     tnl_op_12_08[7:0], tnl_op_13_08[7:0], tnr_op_07_08[7:0],
     tnr_op_08_08[7:0], tnr_op_09_08[7:0], tnr_op_10_08[7:0],
     tnr_op_11_08[7:0], tnr_op_12_08[7:0], top_op_07_08[7:0],
     top_op_08_08[7:0], top_op_09_08[7:0], top_op_10_08[7:0],
     top_op_11_08[7:0], top_op_12_08[7:0], totdopad, trstb_pad,
     update_i, update_mi );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_07_08, carry_out_08_08,
     carry_out_09_08, carry_out_11_08, carry_out_12_08, ceb_o,
     fabric_out_07_00, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fabric_out_13_08, hiz_b_o, mode_o, op_vic_07_08,
     op_vic_08_08, op_vic_09_08, op_vic_11_08, op_vic_12_08,
     padin_07_00a, padin_13_08b, r_o, sdo, sdo_pad, shift_o, tck_pad,
     tclk_o, tdi_pad, tms_pad, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, bs_en_mi, ceb_i, ceb_mi,
     end_of_startup, hiz_b_i, hiz_b_mi, hold_b_r, hold_r_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode_i, mode_mi, mux_jtag_sel_b, pll_sdo, prog, purst, r_i, r_mi,
     sdi, sdi_pad, sdo_enable, shift_i, shift_mi, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out, tclk_i, tclk_mi, totdopad, trstb_pad,
     update_i, update_mi;

output [1:0]  bm_sdo_o;
output [7:0]  slf_op_07_04;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_07_08;
output [7:0]  slf_op_07_05;
output [4:0]  spi_ss_in_bbank;
output [7:0]  slf_op_07_03;
output [7:0]  slf_op_12_08;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_07_07;
output [3:0]  slf_op_13_08;
output [143:0]  cf_b_r;
output [7:0]  slf_op_11_08;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_08_08;
output [7:0]  slf_op_07_01;
output [23:11]  padeb_b_r;
output [191:0]  cf_r;
output [12:0]  padeb_r;
output [23:11]  pado_b_r;
output [3:0]  slf_op_07_00;
output [12:0]  pado_r;
output [7:0]  slf_op_07_02;
output [7:0]  slf_op_07_06;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_10_08;
output [7:0]  slf_op_09_08;

inout [47:0]  sp4_v_b_07_06;
inout [47:0]  sp4_v_t_12_08;
inout [23:0]  sp12_v_t_07_08;
inout [47:0]  sp4_h_l_07_07;
inout [47:0]  sp4_h_l_07_03;
inout [23:0]  sp12_v_t_10_08;
inout [47:0]  sp4_v_b_07_08;
inout [23:0]  sp12_h_l_07_08;
inout [23:0]  sp12_h_l_07_01;
inout [15:0]  sp4_h_l_07_00;
inout [15:0]  sp4_v_t_13_08;
inout [47:0]  sp4_h_l_07_08;
inout [47:0]  sp4_h_l_07_04;
inout [47:0]  sp4_h_l_07_01;
inout [47:0]  sp4_v_b_07_02;
inout [47:0]  sp4_h_l_07_02;
inout [47:0]  sp4_v_t_08_08;
inout [23:0]  sp12_v_t_11_08;
inout [23:0]  sp12_h_l_07_04;
inout [23:0]  sp12_v_t_08_08;
inout [23:0]  sp12_h_l_07_06;
inout [47:0]  sp4_v_t_09_08;
inout [23:0]  sp12_v_t_12_08;
inout [47:0]  sp4_h_l_07_05;
inout [47:0]  sp4_v_b_07_04;
inout [23:0]  sp12_h_l_07_05;
inout [47:0]  sp4_v_b_07_03;
inout [47:0]  sp4_v_t_11_08;
inout [47:0]  sp4_v_t_07_08;
inout [47:0]  sp4_h_l_07_06;
inout [47:0]  sp4_v_b_07_05;
inout [143:0]  wl_r;
inout [143:0]  pgate_r;
inout [23:0]  sp12_h_l_07_07;
inout [47:0]  sp4_v_t_10_08;
inout [47:0]  sp4_v_b_07_07;
inout [143:0]  vdd_cntl_r;
inout [329:0]  bl;
inout [23:0]  sp12_h_l_07_02;
inout [47:0]  sp4_v_b_07_01;
inout [23:0]  sp12_v_t_09_08;
inout [23:0]  sp12_h_l_07_03;
inout [143:0]  reset_b_r;

input [1:0]  bm_sweb_i;
input [7:0]  tnr_op_08_08;
input [7:0]  lft_op_07_03;
input [7:0]  top_op_11_08;
input [7:0]  lft_op_07_07;
input [7:0]  lft_op_07_01;
input [7:0]  glb_in;
input [7:0]  top_op_10_08;
input [23:11]  padin_b_r;
input [7:0]  tnl_op_11_08;
input [7:0]  lft_op_07_08;
input [7:0]  tnr_op_12_08;
input [7:0]  tnl_op_13_08;
input [7:0]  lft_op_07_02;
input [1:0]  bm_sclkrw_i;
input [3:2]  last_rsr;
input [10:0]  bm_aa_top;
input [1:0]  bm_sdi_i;
input [7:0]  tnl_op_08_08;
input [7:0]  tnr_op_09_08;
input [7:0]  tnl_op_07_08;
input [7:0]  top_op_09_08;
input [7:0]  lft_op_07_04;
input [3:0]  bnl_op_07_01;
input [12:0]  padin_r;
input [7:0]  top_op_07_08;
input [7:0]  top_op_08_08;
input [7:0]  lft_op_07_05;
input [7:0]  tnl_op_10_08;
input [1:0]  bm_sdo_i;
input [10:0]  bm_ab_top;
input [7:0]  top_op_12_08;
input [7:0]  tnl_op_12_08;
input [7:0]  tnl_op_09_08;
input [7:0]  tnr_op_07_08;
input [7:0]  lft_op_07_06;
input [7:0]  bm_sa_i;
input [7:0]  tnr_op_11_08;
input [7:0]  tnr_op_10_08;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [47:0]  net1288;

wire  [47:0]  net1383;

wire  [47:0]  net1484;

wire  [23:0]  net1478;

wire  [23:0]  net1509;

wire  [47:0]  net1192;

wire  [7:0]  net1389;

wire  [47:0]  net907;

wire  [23:0]  net1212;

wire  [7:0]  net784;

wire  [7:0]  net913;

wire  [47:0]  net1119;

wire  [23:0]  net901;

wire  [47:0]  net976;

wire  [47:0]  net1169;

wire  [47:0]  net1264;

wire  [23:0]  net1305;

wire  [47:0]  net1492;

wire  [23:0]  net1464;

wire  [23:0]  net911;

wire  [23:0]  net1210;

wire  [7:0]  net1104;

wire  [23:0]  net1209;

wire  [23:0]  net1480;

wire  [47:0]  net980;

wire  [47:0]  net979;

wire  [47:0]  net1551;

wire  [23:0]  net1500;

wire  [47:0]  net1309;

wire  [47:0]  net1000;

wire  [47:0]  net1310;

wire  [23:0]  net1402;

wire  [47:0]  net1360;

wire  [47:0]  net1550;

wire  [7:0]  net1390;

wire  [47:0]  net1262;

wire  [23:0]  net1020;

wire  [7:0]  net936;

wire  [23:0]  net894;

wire  [7:0]  net1045;

wire  [47:0]  net1261;

wire  [47:0]  net889;

wire  [23:0]  net1022;

wire  [23:0]  net1400;

wire  [47:0]  net1382;

wire  [23:0]  net1114;

wire  [47:0]  net1095;

wire  [47:0]  net1003;

wire  [7:0]  clk_center;

wire  [3:0]  slf_op_13_04;

wire  [3:0]  slf_op_12_00;

wire  [47:0]  net1266;

wire  [47:0]  net1076;

wire  [3:0]  slf_op_13_01;

wire  [3:0]  slf_op_13_03;

wire  [7:0]  net1340;

wire  [23:0]  net1257;

wire  [3:0]  slf_op_13_05;

wire  [3:0]  slf_op_08_00;

wire  [23:0]  net1255;

wire  [7:0]  net934;

wire  [7:0]  net1200;

wire  [3:0]  slf_op_13_06;

wire  [23:0]  net1211;

wire  [23:0]  net1019;

wire  [47:0]  net1495;

wire  [23:0]  net1352;

wire  [7:0]  net910;

wire  [47:0]  net1286;

wire  [47:0]  net1171;

wire  [47:0]  net1071;

wire  [10:0]  net792;

wire  [7:0]  net1105;

wire  [7:0]  net1047;

wire  [7:0]  net01436;

wire  [47:0]  net916;

wire  [23:0]  net1350;

wire  [7:0]  net1199;

wire  [3:0]  slf_op_11_00;

wire  [23:0]  net1306;

wire  [47:0]  net1098;

wire  [7:0]  net1531;

wire  [47:0]  net1191;

wire  [47:0]  net1287;

wire  [23:0]  net1476;

wire  [47:0]  net802;

wire  [23:0]  net1021;

wire  [47:0]  net1096;

wire  [7:0]  net1142;

wire  [23:0]  net1508;

wire  [47:0]  net1193;

wire  [47:0]  net1025;

wire  [47:0]  net805;

wire  [23:0]  net1115;

wire  [23:0]  net1160;

wire  [47:0]  net1122;

wire  [47:0]  net1312;

wire  [47:0]  net977;

wire  [47:0]  net1167;

wire  [15:0]  net948;

wire  [47:0]  net1121;

wire  [47:0]  net1380;

wire  [47:0]  net1120;

wire  [47:0]  net1555;

wire  [3:0]  slf_op_09_00;

wire  [23:0]  net970;

wire  [23:0]  net1162;

wire  [23:0]  net1256;

wire  [47:0]  net1405;

wire  [23:0]  net1399;

wire  [47:0]  net1406;

wire  [23:0]  net903;

wire  [7:0]  net1245;

wire  [47:0]  net1267;

wire  [7:0]  net1529;

wire  [23:0]  net1066;

wire  [47:0]  net1166;

wire  [47:0]  net1072;

wire  [7:0]  net938;

wire  [7:0]  net1106;

wire  [23:0]  net1304;

wire  [47:0]  net1554;

wire  [47:0]  net1214;

wire  [47:0]  net982;

wire  [7:0]  net935;

wire  [47:0]  net1001;

wire  [23:0]  net971;

wire  [7:0]  net1295;

wire  [23:0]  net1067;

wire  [47:0]  net1381;

wire  [47:0]  net1404;

wire  [23:0]  net1064;

wire  [7:0]  net937;

wire  [23:0]  net1117;

wire  [47:0]  net1525;

wire  [47:0]  net1260;

wire  [47:0]  net1172;

wire  [7:0]  net1055;

wire  [47:0]  net1524;

wire  [7:0]  net1391;

wire  [47:0]  net1488;

wire  [7:0]  net1530;

wire  [47:0]  net1027;

wire  [7:0]  net939;

wire  [23:0]  net1254;

wire  [47:0]  net1361;

wire  [7:0]  net1528;

wire  [47:0]  net1362;

wire  [47:0]  net1491;

wire  [23:0]  net1159;

wire  [7:0]  net782;

wire  [7:0]  net1533;

wire  [7:0]  net1532;

wire  [10:0]  net791;

wire  [7:0]  net1237;

wire  [47:0]  net1002;

wire  [47:0]  net1506;

wire  [47:0]  net1215;

wire  [47:0]  net1216;

wire  [47:0]  net1311;

wire  [47:0]  net1285;

wire  [47:0]  net1355;

wire  [7:0]  clk_tree_drv_br;

wire  [23:0]  net1065;

wire  [47:0]  net1190;

wire  [23:0]  net972;

wire  [47:0]  net1407;

wire  [3:0]  slf_op_13_07;

wire  [3:0]  slf_op_10_00;

wire  [23:0]  net1161;

wire  [47:0]  net800;

wire  [7:0]  net1296;

wire  [11:11]  padinlat_b_r;

wire  [23:0]  net899;

wire  [23:0]  net969;

wire  [47:0]  net1359;

wire  [7:0]  net1235;

wire  [47:0]  net1170;

wire  [7:0]  net1150;

wire  [7:0]  net1332;

wire  [23:0]  net898;

wire  [23:0]  net1401;

wire  [47:0]  net1553;

wire  [47:0]  net1077;

wire  [47:0]  net1075;

wire  [7:0]  net1330;

wire  [23:0]  net1351;

wire  [47:0]  net1168;

wire  [47:0]  net799;

wire  [23:0]  net1116;

wire  [47:0]  net1357;

wire  [7:0]  net1294;

wire  [47:0]  net896;

wire  [47:0]  net1070;

wire  [47:0]  net1165;

wire  [23:0]  net1307;

wire  [23:0]  net1349;

wire  [47:0]  net1552;

wire  [47:0]  net1356;

wire  [47:0]  net1265;

wire  [47:0]  net981;

wire  [23:0]  net1481;

wire  [7:0]  net793;

wire  [47:0]  net1523;

wire  [47:0]  net1097;

wire  [7:0]  net1140;

wire  [3:0]  slf_op_13_02;

wire  [47:0]  net1217;

wire  [7:0]  net1201;

wire  [47:0]  net1074;



bram1x4_ice1f I_bram_col_b10 ( .glb_netwk_top({net01436[0],
     net01436[1], net01436[2], net01436[3], net01436[4], net01436[5],
     net01436[6], net01436[7]}), .prog(prog),
     .glb_netwk_col(clk_tree_drv_br[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .reset_b(reset_b_r[143:16]),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sreb_o(bm_sreb_o),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .lft_op_05({net1296[0], net1296[1],
     net1296[2], net1296[3], net1296[4], net1296[5], net1296[6],
     net1296[7]}), .bl(bl[203:162]), .sp4_h_l_06({net1097[0],
     net1097[1], net1097[2], net1097[3], net1097[4], net1097[5],
     net1097[6], net1097[7], net1097[8], net1097[9], net1097[10],
     net1097[11], net1097[12], net1097[13], net1097[14], net1097[15],
     net1097[16], net1097[17], net1097[18], net1097[19], net1097[20],
     net1097[21], net1097[22], net1097[23], net1097[24], net1097[25],
     net1097[26], net1097[27], net1097[28], net1097[29], net1097[30],
     net1097[31], net1097[32], net1097[33], net1097[34], net1097[35],
     net1097[36], net1097[37], net1097[38], net1097[39], net1097[40],
     net1097[41], net1097[42], net1097[43], net1097[44], net1097[45],
     net1097[46], net1097[47]}), .sp12_h_l_02({net1066[0], net1066[1],
     net1066[2], net1066[3], net1066[4], net1066[5], net1066[6],
     net1066[7], net1066[8], net1066[9], net1066[10], net1066[11],
     net1066[12], net1066[13], net1066[14], net1066[15], net1066[16],
     net1066[17], net1066[18], net1066[19], net1066[20], net1066[21],
     net1066[22], net1066[23]}), .lft_op_06({net1295[0], net1295[1],
     net1295[2], net1295[3], net1295[4], net1295[5], net1295[6],
     net1295[7]}), .sp12_h_l_03({net1065[0], net1065[1], net1065[2],
     net1065[3], net1065[4], net1065[5], net1065[6], net1065[7],
     net1065[8], net1065[9], net1065[10], net1065[11], net1065[12],
     net1065[13], net1065[14], net1065[15], net1065[16], net1065[17],
     net1065[18], net1065[19], net1065[20], net1065[21], net1065[22],
     net1065[23]}), .sp12_h_r_03({net1464[0], net1464[1], net1464[2],
     net1464[3], net1464[4], net1464[5], net1464[6], net1464[7],
     net1464[8], net1464[9], net1464[10], net1464[11], net1464[12],
     net1464[13], net1464[14], net1464[15], net1464[16], net1464[17],
     net1464[18], net1464[19], net1464[20], net1464[21], net1464[22],
     net1464[23]}), .sp12_h_l_01({net1067[0], net1067[1], net1067[2],
     net1067[3], net1067[4], net1067[5], net1067[6], net1067[7],
     net1067[8], net1067[9], net1067[10], net1067[11], net1067[12],
     net1067[13], net1067[14], net1067[15], net1067[16], net1067[17],
     net1067[18], net1067[19], net1067[20], net1067[21], net1067[22],
     net1067[23]}), .sp4_v_b_04({net1070[0], net1070[1], net1070[2],
     net1070[3], net1070[4], net1070[5], net1070[6], net1070[7],
     net1070[8], net1070[9], net1070[10], net1070[11], net1070[12],
     net1070[13], net1070[14], net1070[15], net1070[16], net1070[17],
     net1070[18], net1070[19], net1070[20], net1070[21], net1070[22],
     net1070[23], net1070[24], net1070[25], net1070[26], net1070[27],
     net1070[28], net1070[29], net1070[30], net1070[31], net1070[32],
     net1070[33], net1070[34], net1070[35], net1070[36], net1070[37],
     net1070[38], net1070[39], net1070[40], net1070[41], net1070[42],
     net1070[43], net1070[44], net1070[45], net1070[46], net1070[47]}),
     .sp4_v_b_05({net1119[0], net1119[1], net1119[2], net1119[3],
     net1119[4], net1119[5], net1119[6], net1119[7], net1119[8],
     net1119[9], net1119[10], net1119[11], net1119[12], net1119[13],
     net1119[14], net1119[15], net1119[16], net1119[17], net1119[18],
     net1119[19], net1119[20], net1119[21], net1119[22], net1119[23],
     net1119[24], net1119[25], net1119[26], net1119[27], net1119[28],
     net1119[29], net1119[30], net1119[31], net1119[32], net1119[33],
     net1119[34], net1119[35], net1119[36], net1119[37], net1119[38],
     net1119[39], net1119[40], net1119[41], net1119[42], net1119[43],
     net1119[44], net1119[45], net1119[46], net1119[47]}),
     .lft_op_07({net1294[0], net1294[1], net1294[2], net1294[3],
     net1294[4], net1294[5], net1294[6], net1294[7]}),
     .sp4_v_b_06({net1120[0], net1120[1], net1120[2], net1120[3],
     net1120[4], net1120[5], net1120[6], net1120[7], net1120[8],
     net1120[9], net1120[10], net1120[11], net1120[12], net1120[13],
     net1120[14], net1120[15], net1120[16], net1120[17], net1120[18],
     net1120[19], net1120[20], net1120[21], net1120[22], net1120[23],
     net1120[24], net1120[25], net1120[26], net1120[27], net1120[28],
     net1120[29], net1120[30], net1120[31], net1120[32], net1120[33],
     net1120[34], net1120[35], net1120[36], net1120[37], net1120[38],
     net1120[39], net1120[40], net1120[41], net1120[42], net1120[43],
     net1120[44], net1120[45], net1120[46], net1120[47]}),
     .sp4_v_b_08({net1122[0], net1122[1], net1122[2], net1122[3],
     net1122[4], net1122[5], net1122[6], net1122[7], net1122[8],
     net1122[9], net1122[10], net1122[11], net1122[12], net1122[13],
     net1122[14], net1122[15], net1122[16], net1122[17], net1122[18],
     net1122[19], net1122[20], net1122[21], net1122[22], net1122[23],
     net1122[24], net1122[25], net1122[26], net1122[27], net1122[28],
     net1122[29], net1122[30], net1122[31], net1122[32], net1122[33],
     net1122[34], net1122[35], net1122[36], net1122[37], net1122[38],
     net1122[39], net1122[40], net1122[41], net1122[42], net1122[43],
     net1122[44], net1122[45], net1122[46], net1122[47]}),
     .sp4_v_b_07({net1121[0], net1121[1], net1121[2], net1121[3],
     net1121[4], net1121[5], net1121[6], net1121[7], net1121[8],
     net1121[9], net1121[10], net1121[11], net1121[12], net1121[13],
     net1121[14], net1121[15], net1121[16], net1121[17], net1121[18],
     net1121[19], net1121[20], net1121[21], net1121[22], net1121[23],
     net1121[24], net1121[25], net1121[26], net1121[27], net1121[28],
     net1121[29], net1121[30], net1121[31], net1121[32], net1121[33],
     net1121[34], net1121[35], net1121[36], net1121[37], net1121[38],
     net1121[39], net1121[40], net1121[41], net1121[42], net1121[43],
     net1121[44], net1121[45], net1121[46], net1121[47]}),
     .lft_op_03({net1235[0], net1235[1], net1235[2], net1235[3],
     net1235[4], net1235[5], net1235[6], net1235[7]}),
     .lft_op_01({net910[0], net910[1], net910[2], net910[3], net910[4],
     net910[5], net910[6], net910[7]}), .sp4_h_l_02({net1076[0],
     net1076[1], net1076[2], net1076[3], net1076[4], net1076[5],
     net1076[6], net1076[7], net1076[8], net1076[9], net1076[10],
     net1076[11], net1076[12], net1076[13], net1076[14], net1076[15],
     net1076[16], net1076[17], net1076[18], net1076[19], net1076[20],
     net1076[21], net1076[22], net1076[23], net1076[24], net1076[25],
     net1076[26], net1076[27], net1076[28], net1076[29], net1076[30],
     net1076[31], net1076[32], net1076[33], net1076[34], net1076[35],
     net1076[36], net1076[37], net1076[38], net1076[39], net1076[40],
     net1076[41], net1076[42], net1076[43], net1076[44], net1076[45],
     net1076[46], net1076[47]}), .sp12_h_l_06({net1115[0], net1115[1],
     net1115[2], net1115[3], net1115[4], net1115[5], net1115[6],
     net1115[7], net1115[8], net1115[9], net1115[10], net1115[11],
     net1115[12], net1115[13], net1115[14], net1115[15], net1115[16],
     net1115[17], net1115[18], net1115[19], net1115[20], net1115[21],
     net1115[22], net1115[23]}), .sp12_h_r_07({net1476[0], net1476[1],
     net1476[2], net1476[3], net1476[4], net1476[5], net1476[6],
     net1476[7], net1476[8], net1476[9], net1476[10], net1476[11],
     net1476[12], net1476[13], net1476[14], net1476[15], net1476[16],
     net1476[17], net1476[18], net1476[19], net1476[20], net1476[21],
     net1476[22], net1476[23]}), .sp12_h_l_05({net1114[0], net1114[1],
     net1114[2], net1114[3], net1114[4], net1114[5], net1114[6],
     net1114[7], net1114[8], net1114[9], net1114[10], net1114[11],
     net1114[12], net1114[13], net1114[14], net1114[15], net1114[16],
     net1114[17], net1114[18], net1114[19], net1114[20], net1114[21],
     net1114[22], net1114[23]}), .sp12_h_r_06({net1478[0], net1478[1],
     net1478[2], net1478[3], net1478[4], net1478[5], net1478[6],
     net1478[7], net1478[8], net1478[9], net1478[10], net1478[11],
     net1478[12], net1478[13], net1478[14], net1478[15], net1478[16],
     net1478[17], net1478[18], net1478[19], net1478[20], net1478[21],
     net1478[22], net1478[23]}), .sp12_h_l_04({net1064[0], net1064[1],
     net1064[2], net1064[3], net1064[4], net1064[5], net1064[6],
     net1064[7], net1064[8], net1064[9], net1064[10], net1064[11],
     net1064[12], net1064[13], net1064[14], net1064[15], net1064[16],
     net1064[17], net1064[18], net1064[19], net1064[20], net1064[21],
     net1064[22], net1064[23]}), .sp12_h_r_05({net1480[0], net1480[1],
     net1480[2], net1480[3], net1480[4], net1480[5], net1480[6],
     net1480[7], net1480[8], net1480[9], net1480[10], net1480[11],
     net1480[12], net1480[13], net1480[14], net1480[15], net1480[16],
     net1480[17], net1480[18], net1480[19], net1480[20], net1480[21],
     net1480[22], net1480[23]}), .sp12_h_r_08({net1481[0], net1481[1],
     net1481[2], net1481[3], net1481[4], net1481[5], net1481[6],
     net1481[7], net1481[8], net1481[9], net1481[10], net1481[11],
     net1481[12], net1481[13], net1481[14], net1481[15], net1481[16],
     net1481[17], net1481[18], net1481[19], net1481[20], net1481[21],
     net1481[22], net1481[23]}), .sp12_h_l_07({net1116[0], net1116[1],
     net1116[2], net1116[3], net1116[4], net1116[5], net1116[6],
     net1116[7], net1116[8], net1116[9], net1116[10], net1116[11],
     net1116[12], net1116[13], net1116[14], net1116[15], net1116[16],
     net1116[17], net1116[18], net1116[19], net1116[20], net1116[21],
     net1116[22], net1116[23]}), .sp12_h_l_08({net1117[0], net1117[1],
     net1117[2], net1117[3], net1117[4], net1117[5], net1117[6],
     net1117[7], net1117[8], net1117[9], net1117[10], net1117[11],
     net1117[12], net1117[13], net1117[14], net1117[15], net1117[16],
     net1117[17], net1117[18], net1117[19], net1117[20], net1117[21],
     net1117[22], net1117[23]}), .sp4_r_v_b_03({net1484[0], net1484[1],
     net1484[2], net1484[3], net1484[4], net1484[5], net1484[6],
     net1484[7], net1484[8], net1484[9], net1484[10], net1484[11],
     net1484[12], net1484[13], net1484[14], net1484[15], net1484[16],
     net1484[17], net1484[18], net1484[19], net1484[20], net1484[21],
     net1484[22], net1484[23], net1484[24], net1484[25], net1484[26],
     net1484[27], net1484[28], net1484[29], net1484[30], net1484[31],
     net1484[32], net1484[33], net1484[34], net1484[35], net1484[36],
     net1484[37], net1484[38], net1484[39], net1484[40], net1484[41],
     net1484[42], net1484[43], net1484[44], net1484[45], net1484[46],
     net1484[47]}), .vdd_cntl(vdd_cntl_r[143:16]),
     .pgate(pgate_r[143:16]), .bot_op_01({slf_op_10_00[3],
     slf_op_10_00[2], slf_op_10_00[1], slf_op_10_00[0],
     slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0]}), .sp4_r_v_b_04({net1488[0], net1488[1],
     net1488[2], net1488[3], net1488[4], net1488[5], net1488[6],
     net1488[7], net1488[8], net1488[9], net1488[10], net1488[11],
     net1488[12], net1488[13], net1488[14], net1488[15], net1488[16],
     net1488[17], net1488[18], net1488[19], net1488[20], net1488[21],
     net1488[22], net1488[23], net1488[24], net1488[25], net1488[26],
     net1488[27], net1488[28], net1488[29], net1488[30], net1488[31],
     net1488[32], net1488[33], net1488[34], net1488[35], net1488[36],
     net1488[37], net1488[38], net1488[39], net1488[40], net1488[41],
     net1488[42], net1488[43], net1488[44], net1488[45], net1488[46],
     net1488[47]}), .sp4_v_b_01({net907[0], net907[1], net907[2],
     net907[3], net907[4], net907[5], net907[6], net907[7], net907[8],
     net907[9], net907[10], net907[11], net907[12], net907[13],
     net907[14], net907[15], net907[16], net907[17], net907[18],
     net907[19], net907[20], net907[21], net907[22], net907[23],
     net907[24], net907[25], net907[26], net907[27], net907[28],
     net907[29], net907[30], net907[31], net907[32], net907[33],
     net907[34], net907[35], net907[36], net907[37], net907[38],
     net907[39], net907[40], net907[41], net907[42], net907[43],
     net907[44], net907[45], net907[46], net907[47]}),
     .sp4_v_b_03({net1071[0], net1071[1], net1071[2], net1071[3],
     net1071[4], net1071[5], net1071[6], net1071[7], net1071[8],
     net1071[9], net1071[10], net1071[11], net1071[12], net1071[13],
     net1071[14], net1071[15], net1071[16], net1071[17], net1071[18],
     net1071[19], net1071[20], net1071[21], net1071[22], net1071[23],
     net1071[24], net1071[25], net1071[26], net1071[27], net1071[28],
     net1071[29], net1071[30], net1071[31], net1071[32], net1071[33],
     net1071[34], net1071[35], net1071[36], net1071[37], net1071[38],
     net1071[39], net1071[40], net1071[41], net1071[42], net1071[43],
     net1071[44], net1071[45], net1071[46], net1071[47]}),
     .sp4_h_r_08({net1491[0], net1491[1], net1491[2], net1491[3],
     net1491[4], net1491[5], net1491[6], net1491[7], net1491[8],
     net1491[9], net1491[10], net1491[11], net1491[12], net1491[13],
     net1491[14], net1491[15], net1491[16], net1491[17], net1491[18],
     net1491[19], net1491[20], net1491[21], net1491[22], net1491[23],
     net1491[24], net1491[25], net1491[26], net1491[27], net1491[28],
     net1491[29], net1491[30], net1491[31], net1491[32], net1491[33],
     net1491[34], net1491[35], net1491[36], net1491[37], net1491[38],
     net1491[39], net1491[40], net1491[41], net1491[42], net1491[43],
     net1491[44], net1491[45], net1491[46], net1491[47]}),
     .sp4_r_v_b_05({net1492[0], net1492[1], net1492[2], net1492[3],
     net1492[4], net1492[5], net1492[6], net1492[7], net1492[8],
     net1492[9], net1492[10], net1492[11], net1492[12], net1492[13],
     net1492[14], net1492[15], net1492[16], net1492[17], net1492[18],
     net1492[19], net1492[20], net1492[21], net1492[22], net1492[23],
     net1492[24], net1492[25], net1492[26], net1492[27], net1492[28],
     net1492[29], net1492[30], net1492[31], net1492[32], net1492[33],
     net1492[34], net1492[35], net1492[36], net1492[37], net1492[38],
     net1492[39], net1492[40], net1492[41], net1492[42], net1492[43],
     net1492[44], net1492[45], net1492[46], net1492[47]}),
     .sp4_v_b_02({net1072[0], net1072[1], net1072[2], net1072[3],
     net1072[4], net1072[5], net1072[6], net1072[7], net1072[8],
     net1072[9], net1072[10], net1072[11], net1072[12], net1072[13],
     net1072[14], net1072[15], net1072[16], net1072[17], net1072[18],
     net1072[19], net1072[20], net1072[21], net1072[22], net1072[23],
     net1072[24], net1072[25], net1072[26], net1072[27], net1072[28],
     net1072[29], net1072[30], net1072[31], net1072[32], net1072[33],
     net1072[34], net1072[35], net1072[36], net1072[37], net1072[38],
     net1072[39], net1072[40], net1072[41], net1072[42], net1072[43],
     net1072[44], net1072[45], net1072[46], net1072[47]}),
     .sp4_v_t_08(sp4_v_t_10_08[47:0]), .sp4_r_v_b_02({net1495[0],
     net1495[1], net1495[2], net1495[3], net1495[4], net1495[5],
     net1495[6], net1495[7], net1495[8], net1495[9], net1495[10],
     net1495[11], net1495[12], net1495[13], net1495[14], net1495[15],
     net1495[16], net1495[17], net1495[18], net1495[19], net1495[20],
     net1495[21], net1495[22], net1495[23], net1495[24], net1495[25],
     net1495[26], net1495[27], net1495[28], net1495[29], net1495[30],
     net1495[31], net1495[32], net1495[33], net1495[34], net1495[35],
     net1495[36], net1495[37], net1495[38], net1495[39], net1495[40],
     net1495[41], net1495[42], net1495[43], net1495[44], net1495[45],
     net1495[46], net1495[47]}), .bnr_op_01({slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0],
     slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0]}), .bm_sdi_o(bm_sdi_o[1:0]),
     .sp4_h_l_04({net1074[0], net1074[1], net1074[2], net1074[3],
     net1074[4], net1074[5], net1074[6], net1074[7], net1074[8],
     net1074[9], net1074[10], net1074[11], net1074[12], net1074[13],
     net1074[14], net1074[15], net1074[16], net1074[17], net1074[18],
     net1074[19], net1074[20], net1074[21], net1074[22], net1074[23],
     net1074[24], net1074[25], net1074[26], net1074[27], net1074[28],
     net1074[29], net1074[30], net1074[31], net1074[32], net1074[33],
     net1074[34], net1074[35], net1074[36], net1074[37], net1074[38],
     net1074[39], net1074[40], net1074[41], net1074[42], net1074[43],
     net1074[44], net1074[45], net1074[46], net1074[47]}),
     .lft_op_08(slf_op_09_08[7:0]), .sp12_h_r_01({net1500[0],
     net1500[1], net1500[2], net1500[3], net1500[4], net1500[5],
     net1500[6], net1500[7], net1500[8], net1500[9], net1500[10],
     net1500[11], net1500[12], net1500[13], net1500[14], net1500[15],
     net1500[16], net1500[17], net1500[18], net1500[19], net1500[20],
     net1500[21], net1500[22], net1500[23]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .sp4_h_l_03({net1075[0], net1075[1], net1075[2], net1075[3],
     net1075[4], net1075[5], net1075[6], net1075[7], net1075[8],
     net1075[9], net1075[10], net1075[11], net1075[12], net1075[13],
     net1075[14], net1075[15], net1075[16], net1075[17], net1075[18],
     net1075[19], net1075[20], net1075[21], net1075[22], net1075[23],
     net1075[24], net1075[25], net1075[26], net1075[27], net1075[28],
     net1075[29], net1075[30], net1075[31], net1075[32], net1075[33],
     net1075[34], net1075[35], net1075[36], net1075[37], net1075[38],
     net1075[39], net1075[40], net1075[41], net1075[42], net1075[43],
     net1075[44], net1075[45], net1075[46], net1075[47]}),
     .sp4_h_l_01({net1077[0], net1077[1], net1077[2], net1077[3],
     net1077[4], net1077[5], net1077[6], net1077[7], net1077[8],
     net1077[9], net1077[10], net1077[11], net1077[12], net1077[13],
     net1077[14], net1077[15], net1077[16], net1077[17], net1077[18],
     net1077[19], net1077[20], net1077[21], net1077[22], net1077[23],
     net1077[24], net1077[25], net1077[26], net1077[27], net1077[28],
     net1077[29], net1077[30], net1077[31], net1077[32], net1077[33],
     net1077[34], net1077[35], net1077[36], net1077[37], net1077[38],
     net1077[39], net1077[40], net1077[41], net1077[42], net1077[43],
     net1077[44], net1077[45], net1077[46], net1077[47]}),
     .sp4_h_r_01({net1506[0], net1506[1], net1506[2], net1506[3],
     net1506[4], net1506[5], net1506[6], net1506[7], net1506[8],
     net1506[9], net1506[10], net1506[11], net1506[12], net1506[13],
     net1506[14], net1506[15], net1506[16], net1506[17], net1506[18],
     net1506[19], net1506[20], net1506[21], net1506[22], net1506[23],
     net1506[24], net1506[25], net1506[26], net1506[27], net1506[28],
     net1506[29], net1506[30], net1506[31], net1506[32], net1506[33],
     net1506[34], net1506[35], net1506[36], net1506[37], net1506[38],
     net1506[39], net1506[40], net1506[41], net1506[42], net1506[43],
     net1506[44], net1506[45], net1506[46], net1506[47]}),
     .tnr_op_08(tnr_op_10_08[7:0]), .sp12_h_r_02({net1508[0],
     net1508[1], net1508[2], net1508[3], net1508[4], net1508[5],
     net1508[6], net1508[7], net1508[8], net1508[9], net1508[10],
     net1508[11], net1508[12], net1508[13], net1508[14], net1508[15],
     net1508[16], net1508[17], net1508[18], net1508[19], net1508[20],
     net1508[21], net1508[22], net1508[23]}), .sp12_h_r_04({net1509[0],
     net1509[1], net1509[2], net1509[3], net1509[4], net1509[5],
     net1509[6], net1509[7], net1509[8], net1509[9], net1509[10],
     net1509[11], net1509[12], net1509[13], net1509[14], net1509[15],
     net1509[16], net1509[17], net1509[18], net1509[19], net1509[20],
     net1509[21], net1509[22], net1509[23]}),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .lft_op_02({net1237[0], net1237[1], net1237[2], net1237[3],
     net1237[4], net1237[5], net1237[6], net1237[7]}),
     .lft_op_04({net1245[0], net1245[1], net1245[2], net1245[3],
     net1245[4], net1245[5], net1245[6], net1245[7]}),
     .bm_sweb_i(bm_sweb_i[1:0]), .bnl_op_01({slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0],
     slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0]}), .sp12_v_t_08(sp12_v_t_10_08[23:0]),
     .wl(wl_r[143:16]), .tnl_op_08(tnl_op_10_08[7:0]),
     .top_op_08(top_op_10_08[7:0]), .bm_ab_2bot({net792[0], net792[1],
     net792[2], net792[3], net792[4], net792[5], net792[6], net792[7],
     net792[8], net792[9], net792[10]}), .bm_aa_2bot({net791[0],
     net791[1], net791[2], net791[3], net791[4], net791[5], net791[6],
     net791[7], net791[8], net791[9], net791[10]}),
     .sp12_v_b_01({net899[0], net899[1], net899[2], net899[3],
     net899[4], net899[5], net899[6], net899[7], net899[8], net899[9],
     net899[10], net899[11], net899[12], net899[13], net899[14],
     net899[15], net899[16], net899[17], net899[18], net899[19],
     net899[20], net899[21], net899[22], net899[23]}),
     .sp4_r_v_b_08({net1523[0], net1523[1], net1523[2], net1523[3],
     net1523[4], net1523[5], net1523[6], net1523[7], net1523[8],
     net1523[9], net1523[10], net1523[11], net1523[12], net1523[13],
     net1523[14], net1523[15], net1523[16], net1523[17], net1523[18],
     net1523[19], net1523[20], net1523[21], net1523[22], net1523[23],
     net1523[24], net1523[25], net1523[26], net1523[27], net1523[28],
     net1523[29], net1523[30], net1523[31], net1523[32], net1523[33],
     net1523[34], net1523[35], net1523[36], net1523[37], net1523[38],
     net1523[39], net1523[40], net1523[41], net1523[42], net1523[43],
     net1523[44], net1523[45], net1523[46], net1523[47]}),
     .sp4_r_v_b_07({net1524[0], net1524[1], net1524[2], net1524[3],
     net1524[4], net1524[5], net1524[6], net1524[7], net1524[8],
     net1524[9], net1524[10], net1524[11], net1524[12], net1524[13],
     net1524[14], net1524[15], net1524[16], net1524[17], net1524[18],
     net1524[19], net1524[20], net1524[21], net1524[22], net1524[23],
     net1524[24], net1524[25], net1524[26], net1524[27], net1524[28],
     net1524[29], net1524[30], net1524[31], net1524[32], net1524[33],
     net1524[34], net1524[35], net1524[36], net1524[37], net1524[38],
     net1524[39], net1524[40], net1524[41], net1524[42], net1524[43],
     net1524[44], net1524[45], net1524[46], net1524[47]}),
     .sp4_r_v_b_06({net1525[0], net1525[1], net1525[2], net1525[3],
     net1525[4], net1525[5], net1525[6], net1525[7], net1525[8],
     net1525[9], net1525[10], net1525[11], net1525[12], net1525[13],
     net1525[14], net1525[15], net1525[16], net1525[17], net1525[18],
     net1525[19], net1525[20], net1525[21], net1525[22], net1525[23],
     net1525[24], net1525[25], net1525[26], net1525[27], net1525[28],
     net1525[29], net1525[30], net1525[31], net1525[32], net1525[33],
     net1525[34], net1525[35], net1525[36], net1525[37], net1525[38],
     net1525[39], net1525[40], net1525[41], net1525[42], net1525[43],
     net1525[44], net1525[45], net1525[46], net1525[47]}),
     .sp4_r_v_b_01({net896[0], net896[1], net896[2], net896[3],
     net896[4], net896[5], net896[6], net896[7], net896[8], net896[9],
     net896[10], net896[11], net896[12], net896[13], net896[14],
     net896[15], net896[16], net896[17], net896[18], net896[19],
     net896[20], net896[21], net896[22], net896[23], net896[24],
     net896[25], net896[26], net896[27], net896[28], net896[29],
     net896[30], net896[31], net896[32], net896[33], net896[34],
     net896[35], net896[36], net896[37], net896[38], net896[39],
     net896[40], net896[41], net896[42], net896[43], net896[44],
     net896[45], net896[46], net896[47]}),
     .rgt_op_08(slf_op_11_08[7:0]), .rgt_op_07({net1528[0], net1528[1],
     net1528[2], net1528[3], net1528[4], net1528[5], net1528[6],
     net1528[7]}), .rgt_op_06({net1529[0], net1529[1], net1529[2],
     net1529[3], net1529[4], net1529[5], net1529[6], net1529[7]}),
     .rgt_op_05({net1530[0], net1530[1], net1530[2], net1530[3],
     net1530[4], net1530[5], net1530[6], net1530[7]}),
     .rgt_op_04({net1531[0], net1531[1], net1531[2], net1531[3],
     net1531[4], net1531[5], net1531[6], net1531[7]}),
     .rgt_op_03({net1532[0], net1532[1], net1532[2], net1532[3],
     net1532[4], net1532[5], net1532[6], net1532[7]}),
     .rgt_op_02({net1533[0], net1533[1], net1533[2], net1533[3],
     net1533[4], net1533[5], net1533[6], net1533[7]}),
     .rgt_op_01({net782[0], net782[1], net782[2], net782[3], net782[4],
     net782[5], net782[6], net782[7]}), .slf_op_02({net1047[0],
     net1047[1], net1047[2], net1047[3], net1047[4], net1047[5],
     net1047[6], net1047[7]}), .slf_op_01({net784[0], net784[1],
     net784[2], net784[3], net784[4], net784[5], net784[6],
     net784[7]}), .slf_op_03({net1045[0], net1045[1], net1045[2],
     net1045[3], net1045[4], net1045[5], net1045[6], net1045[7]}),
     .slf_op_04({net1055[0], net1055[1], net1055[2], net1055[3],
     net1055[4], net1055[5], net1055[6], net1055[7]}),
     .slf_op_05({net1106[0], net1106[1], net1106[2], net1106[3],
     net1106[4], net1106[5], net1106[6], net1106[7]}),
     .slf_op_06({net1105[0], net1105[1], net1105[2], net1105[3],
     net1105[4], net1105[5], net1105[6], net1105[7]}),
     .slf_op_07({net1104[0], net1104[1], net1104[2], net1104[3],
     net1104[4], net1104[5], net1104[6], net1104[7]}),
     .slf_op_08(slf_op_10_08[7:0]), .bm_ab_top(bm_ab_top[10:0]),
     .bm_aa_top(bm_aa_top[10:0]), .glb_netwk_bot({net936[0], net936[1],
     net936[2], net936[3], net936[4], net936[5], net936[6],
     net936[7]}), .sp4_h_l_08({net1095[0], net1095[1], net1095[2],
     net1095[3], net1095[4], net1095[5], net1095[6], net1095[7],
     net1095[8], net1095[9], net1095[10], net1095[11], net1095[12],
     net1095[13], net1095[14], net1095[15], net1095[16], net1095[17],
     net1095[18], net1095[19], net1095[20], net1095[21], net1095[22],
     net1095[23], net1095[24], net1095[25], net1095[26], net1095[27],
     net1095[28], net1095[29], net1095[30], net1095[31], net1095[32],
     net1095[33], net1095[34], net1095[35], net1095[36], net1095[37],
     net1095[38], net1095[39], net1095[40], net1095[41], net1095[42],
     net1095[43], net1095[44], net1095[45], net1095[46], net1095[47]}),
     .sp4_h_l_07({net1096[0], net1096[1], net1096[2], net1096[3],
     net1096[4], net1096[5], net1096[6], net1096[7], net1096[8],
     net1096[9], net1096[10], net1096[11], net1096[12], net1096[13],
     net1096[14], net1096[15], net1096[16], net1096[17], net1096[18],
     net1096[19], net1096[20], net1096[21], net1096[22], net1096[23],
     net1096[24], net1096[25], net1096[26], net1096[27], net1096[28],
     net1096[29], net1096[30], net1096[31], net1096[32], net1096[33],
     net1096[34], net1096[35], net1096[36], net1096[37], net1096[38],
     net1096[39], net1096[40], net1096[41], net1096[42], net1096[43],
     net1096[44], net1096[45], net1096[46], net1096[47]}),
     .sp4_h_l_05({net1098[0], net1098[1], net1098[2], net1098[3],
     net1098[4], net1098[5], net1098[6], net1098[7], net1098[8],
     net1098[9], net1098[10], net1098[11], net1098[12], net1098[13],
     net1098[14], net1098[15], net1098[16], net1098[17], net1098[18],
     net1098[19], net1098[20], net1098[21], net1098[22], net1098[23],
     net1098[24], net1098[25], net1098[26], net1098[27], net1098[28],
     net1098[29], net1098[30], net1098[31], net1098[32], net1098[33],
     net1098[34], net1098[35], net1098[36], net1098[37], net1098[38],
     net1098[39], net1098[40], net1098[41], net1098[42], net1098[43],
     net1098[44], net1098[45], net1098[46], net1098[47]}),
     .sp4_h_r_02({net1550[0], net1550[1], net1550[2], net1550[3],
     net1550[4], net1550[5], net1550[6], net1550[7], net1550[8],
     net1550[9], net1550[10], net1550[11], net1550[12], net1550[13],
     net1550[14], net1550[15], net1550[16], net1550[17], net1550[18],
     net1550[19], net1550[20], net1550[21], net1550[22], net1550[23],
     net1550[24], net1550[25], net1550[26], net1550[27], net1550[28],
     net1550[29], net1550[30], net1550[31], net1550[32], net1550[33],
     net1550[34], net1550[35], net1550[36], net1550[37], net1550[38],
     net1550[39], net1550[40], net1550[41], net1550[42], net1550[43],
     net1550[44], net1550[45], net1550[46], net1550[47]}),
     .sp4_h_r_03({net1551[0], net1551[1], net1551[2], net1551[3],
     net1551[4], net1551[5], net1551[6], net1551[7], net1551[8],
     net1551[9], net1551[10], net1551[11], net1551[12], net1551[13],
     net1551[14], net1551[15], net1551[16], net1551[17], net1551[18],
     net1551[19], net1551[20], net1551[21], net1551[22], net1551[23],
     net1551[24], net1551[25], net1551[26], net1551[27], net1551[28],
     net1551[29], net1551[30], net1551[31], net1551[32], net1551[33],
     net1551[34], net1551[35], net1551[36], net1551[37], net1551[38],
     net1551[39], net1551[40], net1551[41], net1551[42], net1551[43],
     net1551[44], net1551[45], net1551[46], net1551[47]}),
     .sp4_h_r_04({net1552[0], net1552[1], net1552[2], net1552[3],
     net1552[4], net1552[5], net1552[6], net1552[7], net1552[8],
     net1552[9], net1552[10], net1552[11], net1552[12], net1552[13],
     net1552[14], net1552[15], net1552[16], net1552[17], net1552[18],
     net1552[19], net1552[20], net1552[21], net1552[22], net1552[23],
     net1552[24], net1552[25], net1552[26], net1552[27], net1552[28],
     net1552[29], net1552[30], net1552[31], net1552[32], net1552[33],
     net1552[34], net1552[35], net1552[36], net1552[37], net1552[38],
     net1552[39], net1552[40], net1552[41], net1552[42], net1552[43],
     net1552[44], net1552[45], net1552[46], net1552[47]}),
     .sp4_h_r_05({net1553[0], net1553[1], net1553[2], net1553[3],
     net1553[4], net1553[5], net1553[6], net1553[7], net1553[8],
     net1553[9], net1553[10], net1553[11], net1553[12], net1553[13],
     net1553[14], net1553[15], net1553[16], net1553[17], net1553[18],
     net1553[19], net1553[20], net1553[21], net1553[22], net1553[23],
     net1553[24], net1553[25], net1553[26], net1553[27], net1553[28],
     net1553[29], net1553[30], net1553[31], net1553[32], net1553[33],
     net1553[34], net1553[35], net1553[36], net1553[37], net1553[38],
     net1553[39], net1553[40], net1553[41], net1553[42], net1553[43],
     net1553[44], net1553[45], net1553[46], net1553[47]}),
     .sp4_h_r_06({net1554[0], net1554[1], net1554[2], net1554[3],
     net1554[4], net1554[5], net1554[6], net1554[7], net1554[8],
     net1554[9], net1554[10], net1554[11], net1554[12], net1554[13],
     net1554[14], net1554[15], net1554[16], net1554[17], net1554[18],
     net1554[19], net1554[20], net1554[21], net1554[22], net1554[23],
     net1554[24], net1554[25], net1554[26], net1554[27], net1554[28],
     net1554[29], net1554[30], net1554[31], net1554[32], net1554[33],
     net1554[34], net1554[35], net1554[36], net1554[37], net1554[38],
     net1554[39], net1554[40], net1554[41], net1554[42], net1554[43],
     net1554[44], net1554[45], net1554[46], net1554[47]}),
     .sp4_h_r_07({net1555[0], net1555[1], net1555[2], net1555[3],
     net1555[4], net1555[5], net1555[6], net1555[7], net1555[8],
     net1555[9], net1555[10], net1555[11], net1555[12], net1555[13],
     net1555[14], net1555[15], net1555[16], net1555[17], net1555[18],
     net1555[19], net1555[20], net1555[21], net1555[22], net1555[23],
     net1555[24], net1555[25], net1555[26], net1555[27], net1555[28],
     net1555[29], net1555[30], net1555[31], net1555[32], net1555[33],
     net1555[34], net1555[35], net1555[36], net1555[37], net1555[38],
     net1555[39], net1555[40], net1555[41], net1555[42], net1555[43],
     net1555[44], net1555[45], net1555[46], net1555[47]}));
pinlatbuf12p_1 I484 ( .pad_in(padin_r[12]), .icegate(hold_r_b),
     .cbit(cf_r[183]), .cout(net0731), .prog(prog));
pinlatbuf12p_1 I486 ( .pad_in(padin_b_r[11]), .icegate(hold_b_r),
     .cbit(cf_b_r[15]), .cout(padinlat_b_r[11]), .prog(prog));
tielo I369 ( .tielo(tgnd_br_q));
scan_buf_ice8p I_scanbuf_8p_br ( .update_i(update_mi),
     .tclk_i(tclk_mi), .shift_i(shift_mi), .sdi(sdi_pad), .r_i(r_mi),
     .mode_i(mode_mi), .hiz_b_i(hiz_b_mi), .ceb_i(ceb_mi),
     .bs_en_i(bs_en_mi), .update_o(update_o), .tclk_o(net774),
     .shift_o(shift_o), .sdo(net776), .r_o(r_o), .mode_o(mode_o),
     .hiz_b_o(hiz_b_o), .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_rgt_bot_1x8_ice1f I_preio_rgt_b ( cf_r[191:0], net808, net807,
     net809, padeb_r[12:0], pado_r[12:0], sdo, slf_op_13_01[3:0],
     slf_op_13_02[3:0], slf_op_13_03[3:0], slf_op_13_04[3:0],
     slf_op_13_05[3:0], slf_op_13_06[3:0], slf_op_13_07[3:0],
     slf_op_13_08[3:0], tck_pad, tclk_o, tdi_pad, tms_pad, {net982[0],
     net982[1], net982[2], net982[3], net982[4], net982[5], net982[6],
     net982[7], net982[8], net982[9], net982[10], net982[11],
     net982[12], net982[13], net982[14], net982[15], net982[16],
     net982[17], net982[18], net982[19], net982[20], net982[21],
     net982[22], net982[23], net982[24], net982[25], net982[26],
     net982[27], net982[28], net982[29], net982[30], net982[31],
     net982[32], net982[33], net982[34], net982[35], net982[36],
     net982[37], net982[38], net982[39], net982[40], net982[41],
     net982[42], net982[43], net982[44], net982[45], net982[46],
     net982[47]}, {net981[0], net981[1], net981[2], net981[3],
     net981[4], net981[5], net981[6], net981[7], net981[8], net981[9],
     net981[10], net981[11], net981[12], net981[13], net981[14],
     net981[15], net981[16], net981[17], net981[18], net981[19],
     net981[20], net981[21], net981[22], net981[23], net981[24],
     net981[25], net981[26], net981[27], net981[28], net981[29],
     net981[30], net981[31], net981[32], net981[33], net981[34],
     net981[35], net981[36], net981[37], net981[38], net981[39],
     net981[40], net981[41], net981[42], net981[43], net981[44],
     net981[45], net981[46], net981[47]}, {net980[0], net980[1],
     net980[2], net980[3], net980[4], net980[5], net980[6], net980[7],
     net980[8], net980[9], net980[10], net980[11], net980[12],
     net980[13], net980[14], net980[15], net980[16], net980[17],
     net980[18], net980[19], net980[20], net980[21], net980[22],
     net980[23], net980[24], net980[25], net980[26], net980[27],
     net980[28], net980[29], net980[30], net980[31], net980[32],
     net980[33], net980[34], net980[35], net980[36], net980[37],
     net980[38], net980[39], net980[40], net980[41], net980[42],
     net980[43], net980[44], net980[45], net980[46], net980[47]},
     {net979[0], net979[1], net979[2], net979[3], net979[4], net979[5],
     net979[6], net979[7], net979[8], net979[9], net979[10],
     net979[11], net979[12], net979[13], net979[14], net979[15],
     net979[16], net979[17], net979[18], net979[19], net979[20],
     net979[21], net979[22], net979[23], net979[24], net979[25],
     net979[26], net979[27], net979[28], net979[29], net979[30],
     net979[31], net979[32], net979[33], net979[34], net979[35],
     net979[36], net979[37], net979[38], net979[39], net979[40],
     net979[41], net979[42], net979[43], net979[44], net979[45],
     net979[46], net979[47]}, {net1003[0], net1003[1], net1003[2],
     net1003[3], net1003[4], net1003[5], net1003[6], net1003[7],
     net1003[8], net1003[9], net1003[10], net1003[11], net1003[12],
     net1003[13], net1003[14], net1003[15], net1003[16], net1003[17],
     net1003[18], net1003[19], net1003[20], net1003[21], net1003[22],
     net1003[23], net1003[24], net1003[25], net1003[26], net1003[27],
     net1003[28], net1003[29], net1003[30], net1003[31], net1003[32],
     net1003[33], net1003[34], net1003[35], net1003[36], net1003[37],
     net1003[38], net1003[39], net1003[40], net1003[41], net1003[42],
     net1003[43], net1003[44], net1003[45], net1003[46], net1003[47]},
     {net1002[0], net1002[1], net1002[2], net1002[3], net1002[4],
     net1002[5], net1002[6], net1002[7], net1002[8], net1002[9],
     net1002[10], net1002[11], net1002[12], net1002[13], net1002[14],
     net1002[15], net1002[16], net1002[17], net1002[18], net1002[19],
     net1002[20], net1002[21], net1002[22], net1002[23], net1002[24],
     net1002[25], net1002[26], net1002[27], net1002[28], net1002[29],
     net1002[30], net1002[31], net1002[32], net1002[33], net1002[34],
     net1002[35], net1002[36], net1002[37], net1002[38], net1002[39],
     net1002[40], net1002[41], net1002[42], net1002[43], net1002[44],
     net1002[45], net1002[46], net1002[47]}, {net1001[0], net1001[1],
     net1001[2], net1001[3], net1001[4], net1001[5], net1001[6],
     net1001[7], net1001[8], net1001[9], net1001[10], net1001[11],
     net1001[12], net1001[13], net1001[14], net1001[15], net1001[16],
     net1001[17], net1001[18], net1001[19], net1001[20], net1001[21],
     net1001[22], net1001[23], net1001[24], net1001[25], net1001[26],
     net1001[27], net1001[28], net1001[29], net1001[30], net1001[31],
     net1001[32], net1001[33], net1001[34], net1001[35], net1001[36],
     net1001[37], net1001[38], net1001[39], net1001[40], net1001[41],
     net1001[42], net1001[43], net1001[44], net1001[45], net1001[46],
     net1001[47]}, {net1000[0], net1000[1], net1000[2], net1000[3],
     net1000[4], net1000[5], net1000[6], net1000[7], net1000[8],
     net1000[9], net1000[10], net1000[11], net1000[12], net1000[13],
     net1000[14], net1000[15], net1000[16], net1000[17], net1000[18],
     net1000[19], net1000[20], net1000[21], net1000[22], net1000[23],
     net1000[24], net1000[25], net1000[26], net1000[27], net1000[28],
     net1000[29], net1000[30], net1000[31], net1000[32], net1000[33],
     net1000[34], net1000[35], net1000[36], net1000[37], net1000[38],
     net1000[39], net1000[40], net1000[41], net1000[42], net1000[43],
     net1000[44], net1000[45], net1000[46], net1000[47]}, {net972[0],
     net972[1], net972[2], net972[3], net972[4], net972[5], net972[6],
     net972[7], net972[8], net972[9], net972[10], net972[11],
     net972[12], net972[13], net972[14], net972[15], net972[16],
     net972[17], net972[18], net972[19], net972[20], net972[21],
     net972[22], net972[23]}, {net971[0], net971[1], net971[2],
     net971[3], net971[4], net971[5], net971[6], net971[7], net971[8],
     net971[9], net971[10], net971[11], net971[12], net971[13],
     net971[14], net971[15], net971[16], net971[17], net971[18],
     net971[19], net971[20], net971[21], net971[22], net971[23]},
     {net970[0], net970[1], net970[2], net970[3], net970[4], net970[5],
     net970[6], net970[7], net970[8], net970[9], net970[10],
     net970[11], net970[12], net970[13], net970[14], net970[15],
     net970[16], net970[17], net970[18], net970[19], net970[20],
     net970[21], net970[22], net970[23]}, {net969[0], net969[1],
     net969[2], net969[3], net969[4], net969[5], net969[6], net969[7],
     net969[8], net969[9], net969[10], net969[11], net969[12],
     net969[13], net969[14], net969[15], net969[16], net969[17],
     net969[18], net969[19], net969[20], net969[21], net969[22],
     net969[23]}, {net1019[0], net1019[1], net1019[2], net1019[3],
     net1019[4], net1019[5], net1019[6], net1019[7], net1019[8],
     net1019[9], net1019[10], net1019[11], net1019[12], net1019[13],
     net1019[14], net1019[15], net1019[16], net1019[17], net1019[18],
     net1019[19], net1019[20], net1019[21], net1019[22], net1019[23]},
     {net1020[0], net1020[1], net1020[2], net1020[3], net1020[4],
     net1020[5], net1020[6], net1020[7], net1020[8], net1020[9],
     net1020[10], net1020[11], net1020[12], net1020[13], net1020[14],
     net1020[15], net1020[16], net1020[17], net1020[18], net1020[19],
     net1020[20], net1020[21], net1020[22], net1020[23]}, {net1021[0],
     net1021[1], net1021[2], net1021[3], net1021[4], net1021[5],
     net1021[6], net1021[7], net1021[8], net1021[9], net1021[10],
     net1021[11], net1021[12], net1021[13], net1021[14], net1021[15],
     net1021[16], net1021[17], net1021[18], net1021[19], net1021[20],
     net1021[21], net1021[22], net1021[23]}, {net1022[0], net1022[1],
     net1022[2], net1022[3], net1022[4], net1022[5], net1022[6],
     net1022[7], net1022[8], net1022[9], net1022[10], net1022[11],
     net1022[12], net1022[13], net1022[14], net1022[15], net1022[16],
     net1022[17], net1022[18], net1022[19], net1022[20], net1022[21],
     net1022[22], net1022[23]}, bl[329:312], pgate_r[143:16],
     reset_b_r[143:16], {net948[0], net948[1], net948[2], net948[3],
     net948[4], net948[5], net948[6], net948[7], net948[8], net948[9],
     net948[10], net948[11], net948[12], net948[13], net948[14],
     net948[15]}, sp4_v_t_13_08[15:0], vdd_cntl_r[143:16],
     wl_r[143:16], {slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0], slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0]}, bs_en_o, ceb_o,
     clk_tree_drv_br[7:0], hiz_b_o, hold_r_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[2],
     last_rsr[3], {net913[0], net913[1], net913[2], net913[3],
     net913[4], net913[5], net913[6], net913[7]}, {net1142[0],
     net1142[1], net1142[2], net1142[3], net1142[4], net1142[5],
     net1142[6], net1142[7]}, {net1140[0], net1140[1], net1140[2],
     net1140[3], net1140[4], net1140[5], net1140[6], net1140[7]},
     {net1150[0], net1150[1], net1150[2], net1150[3], net1150[4],
     net1150[5], net1150[6], net1150[7]}, {net1201[0], net1201[1],
     net1201[2], net1201[3], net1201[4], net1201[5], net1201[6],
     net1201[7]}, {net1200[0], net1200[1], net1200[2], net1200[3],
     net1200[4], net1200[5], net1200[6], net1200[7]}, {net1199[0],
     net1199[1], net1199[2], net1199[3], net1199[4], net1199[5],
     net1199[6], net1199[7]}, slf_op_12_08[7:0], mode_o,
     mux_jtag_sel_b, padin_r[12:0], prog, r_o, net776, sdo_enable,
     shift_o, net774, tnl_op_13_08[7:0], totdopad, trstb_pad,
     update_o);
io_bot_rgt_1x6_ice1f I_preio_bot_r ( cf_b_r[143:0], net1437, net912,
     padeb_b_r[11], padeb_b_r[23:13], pado_b_r[11], pado_b_r[23:13],
     sdo_pad, slf_op_07_00[3:0], slf_op_08_00[3:0], slf_op_09_00[3:0],
     slf_op_10_00[3:0], slf_op_11_00[3:0], slf_op_12_00[3:0],
     spi_ss_in_bbank[4:0], bl[53:0], bl[107:54], bl[161:108],
     bl[203:162], bl[257:204], bl[311:258], sp4_h_l_07_00[15:0],
     {net948[0], net948[1], net948[2], net948[3], net948[4], net948[5],
     net948[6], net948[7], net948[8], net948[9], net948[10],
     net948[11], net948[12], net948[13], net948[14], net948[15]},
     sp4_v_b_07_01[47:0], {net889[0], net889[1], net889[2], net889[3],
     net889[4], net889[5], net889[6], net889[7], net889[8], net889[9],
     net889[10], net889[11], net889[12], net889[13], net889[14],
     net889[15], net889[16], net889[17], net889[18], net889[19],
     net889[20], net889[21], net889[22], net889[23], net889[24],
     net889[25], net889[26], net889[27], net889[28], net889[29],
     net889[30], net889[31], net889[32], net889[33], net889[34],
     net889[35], net889[36], net889[37], net889[38], net889[39],
     net889[40], net889[41], net889[42], net889[43], net889[44],
     net889[45], net889[46], net889[47]}, {net916[0], net916[1],
     net916[2], net916[3], net916[4], net916[5], net916[6], net916[7],
     net916[8], net916[9], net916[10], net916[11], net916[12],
     net916[13], net916[14], net916[15], net916[16], net916[17],
     net916[18], net916[19], net916[20], net916[21], net916[22],
     net916[23], net916[24], net916[25], net916[26], net916[27],
     net916[28], net916[29], net916[30], net916[31], net916[32],
     net916[33], net916[34], net916[35], net916[36], net916[37],
     net916[38], net916[39], net916[40], net916[41], net916[42],
     net916[43], net916[44], net916[45], net916[46], net916[47]},
     {net907[0], net907[1], net907[2], net907[3], net907[4], net907[5],
     net907[6], net907[7], net907[8], net907[9], net907[10],
     net907[11], net907[12], net907[13], net907[14], net907[15],
     net907[16], net907[17], net907[18], net907[19], net907[20],
     net907[21], net907[22], net907[23], net907[24], net907[25],
     net907[26], net907[27], net907[28], net907[29], net907[30],
     net907[31], net907[32], net907[33], net907[34], net907[35],
     net907[36], net907[37], net907[38], net907[39], net907[40],
     net907[41], net907[42], net907[43], net907[44], net907[45],
     net907[46], net907[47]}, {net896[0], net896[1], net896[2],
     net896[3], net896[4], net896[5], net896[6], net896[7], net896[8],
     net896[9], net896[10], net896[11], net896[12], net896[13],
     net896[14], net896[15], net896[16], net896[17], net896[18],
     net896[19], net896[20], net896[21], net896[22], net896[23],
     net896[24], net896[25], net896[26], net896[27], net896[28],
     net896[29], net896[30], net896[31], net896[32], net896[33],
     net896[34], net896[35], net896[36], net896[37], net896[38],
     net896[39], net896[40], net896[41], net896[42], net896[43],
     net896[44], net896[45], net896[46], net896[47]}, {net1168[0],
     net1168[1], net1168[2], net1168[3], net1168[4], net1168[5],
     net1168[6], net1168[7], net1168[8], net1168[9], net1168[10],
     net1168[11], net1168[12], net1168[13], net1168[14], net1168[15],
     net1168[16], net1168[17], net1168[18], net1168[19], net1168[20],
     net1168[21], net1168[22], net1168[23], net1168[24], net1168[25],
     net1168[26], net1168[27], net1168[28], net1168[29], net1168[30],
     net1168[31], net1168[32], net1168[33], net1168[34], net1168[35],
     net1168[36], net1168[37], net1168[38], net1168[39], net1168[40],
     net1168[41], net1168[42], net1168[43], net1168[44], net1168[45],
     net1168[46], net1168[47]}, {net903[0], net903[1], net903[2],
     net903[3], net903[4], net903[5], net903[6], net903[7], net903[8],
     net903[9], net903[10], net903[11], net903[12], net903[13],
     net903[14], net903[15], net903[16], net903[17], net903[18],
     net903[19], net903[20], net903[21], net903[22], net903[23]},
     {net901[0], net901[1], net901[2], net901[3], net901[4], net901[5],
     net901[6], net901[7], net901[8], net901[9], net901[10],
     net901[11], net901[12], net901[13], net901[14], net901[15],
     net901[16], net901[17], net901[18], net901[19], net901[20],
     net901[21], net901[22], net901[23]}, {net911[0], net911[1],
     net911[2], net911[3], net911[4], net911[5], net911[6], net911[7],
     net911[8], net911[9], net911[10], net911[11], net911[12],
     net911[13], net911[14], net911[15], net911[16], net911[17],
     net911[18], net911[19], net911[20], net911[21], net911[22],
     net911[23]}, {net899[0], net899[1], net899[2], net899[3],
     net899[4], net899[5], net899[6], net899[7], net899[8], net899[9],
     net899[10], net899[11], net899[12], net899[13], net899[14],
     net899[15], net899[16], net899[17], net899[18], net899[19],
     net899[20], net899[21], net899[22], net899[23]}, {net894[0],
     net894[1], net894[2], net894[3], net894[4], net894[5], net894[6],
     net894[7], net894[8], net894[9], net894[10], net894[11],
     net894[12], net894[13], net894[14], net894[15], net894[16],
     net894[17], net894[18], net894[19], net894[20], net894[21],
     net894[22], net894[23]}, {net898[0], net898[1], net898[2],
     net898[3], net898[4], net898[5], net898[6], net898[7], net898[8],
     net898[9], net898[10], net898[11], net898[12], net898[13],
     net898[14], net898[15], net898[16], net898[17], net898[18],
     net898[19], net898[20], net898[21], net898[22], net898[23]},
     lft_op_07_01[7:0], bs_en_i, ceb_i, end_of_startup, {net939[0],
     net939[1], net939[2], net939[3], net939[4], net939[5], net939[6],
     net939[7]}, {net938[0], net938[1], net938[2], net938[3],
     net938[4], net938[5], net938[6], net938[7]}, {net937[0],
     net937[1], net937[2], net937[3], net937[4], net937[5], net937[6],
     net937[7]}, {net936[0], net936[1], net936[2], net936[3],
     net936[4], net936[5], net936[6], net936[7]}, {net935[0],
     net935[1], net935[2], net935[3], net935[4], net935[5], net935[6],
     net935[7]}, {net934[0], net934[1], net934[2], net934[3],
     net934[4], net934[5], net934[6], net934[7]}, hiz_b_i, hold_b_r,
     slf_op_07_01[7:0], {net793[0], net793[1], net793[2], net793[3],
     net793[4], net793[5], net793[6], net793[7]}, {net910[0],
     net910[1], net910[2], net910[3], net910[4], net910[5], net910[6],
     net910[7]}, {net784[0], net784[1], net784[2], net784[3],
     net784[4], net784[5], net784[6], net784[7]}, {net782[0],
     net782[1], net782[2], net782[3], net782[4], net782[5], net782[6],
     net782[7]}, {net913[0], net913[1], net913[2], net913[3],
     net913[4], net913[5], net913[6], net913[7]}, md_spi_b, mode_i,
     padin_b_r[11], padin_b_r[23:13], {pgate_r[1], pgate_r[0],
     pgate_r[2], pgate_r[3], pgate_r[5], pgate_r[4], pgate_r[6],
     pgate_r[7], pgate_r[9], pgate_r[8], pgate_r[10], pgate_r[11],
     pgate_r[13], pgate_r[12], pgate_r[14], pgate_r[15]}, prog, r_i,
     {reset_b_r[1], reset_b_r[0], reset_b_r[2], reset_b_r[3],
     reset_b_r[5], reset_b_r[4], reset_b_r[6], reset_b_r[7],
     reset_b_r[9], reset_b_r[8], reset_b_r[10], reset_b_r[11],
     reset_b_r[13], reset_b_r[12], reset_b_r[14], reset_b_r[15]}, sdi,
     shift_i, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out, tclk_i,
     {slf_op_13_01[3], slf_op_13_01[2], slf_op_13_01[1],
     slf_op_13_01[0], slf_op_13_01[3], slf_op_13_01[2],
     slf_op_13_01[1], slf_op_13_01[0]}, update_i, {vdd_cntl_r[1],
     vdd_cntl_r[0], vdd_cntl_r[2], vdd_cntl_r[3], vdd_cntl_r[5],
     vdd_cntl_r[4], vdd_cntl_r[6], vdd_cntl_r[7], vdd_cntl_r[9],
     vdd_cntl_r[8], vdd_cntl_r[10], vdd_cntl_r[11], vdd_cntl_r[13],
     vdd_cntl_r[12], vdd_cntl_r[14], vdd_cntl_r[15]}, {wl_r[1],
     wl_r[0], wl_r[2], wl_r[3], wl_r[5], wl_r[4], wl_r[6], wl_r[7],
     wl_r[9], wl_r[8], wl_r[10], wl_r[11], wl_r[13], wl_r[12],
     wl_r[14], wl_r[15]});
lt_1x8_bot_ice1f I_lt_col_b12 ( .glb_netwk_bot({net934[0], net934[1],
     net934[2], net934[3], net934[4], net934[5], net934[6],
     net934[7]}), .rgt_op_03({slf_op_13_03[3], slf_op_13_03[2],
     slf_op_13_03[1], slf_op_13_03[0], slf_op_13_03[3],
     slf_op_13_03[2], slf_op_13_03[1], slf_op_13_03[0]}),
     .slf_op_02({net1142[0], net1142[1], net1142[2], net1142[3],
     net1142[4], net1142[5], net1142[6], net1142[7]}),
     .rgt_op_02({slf_op_13_02[3], slf_op_13_02[2], slf_op_13_02[1],
     slf_op_13_02[0], slf_op_13_02[3], slf_op_13_02[2],
     slf_op_13_02[1], slf_op_13_02[0]}), .rgt_op_01({slf_op_13_01[3],
     slf_op_13_01[2], slf_op_13_01[1], slf_op_13_01[0],
     slf_op_13_01[3], slf_op_13_01[2], slf_op_13_01[1],
     slf_op_13_01[0]}), .purst(purst), .prog(prog),
     .lft_op_04({net1531[0], net1531[1], net1531[2], net1531[3],
     net1531[4], net1531[5], net1531[6], net1531[7]}),
     .lft_op_03({net1532[0], net1532[1], net1532[2], net1532[3],
     net1532[4], net1532[5], net1532[6], net1532[7]}),
     .lft_op_02({net1533[0], net1533[1], net1533[2], net1533[3],
     net1533[4], net1533[5], net1533[6], net1533[7]}),
     .lft_op_01({net782[0], net782[1], net782[2], net782[3], net782[4],
     net782[5], net782[6], net782[7]}), .rgt_op_04({slf_op_13_04[3],
     slf_op_13_04[2], slf_op_13_04[1], slf_op_13_04[0],
     slf_op_13_04[3], slf_op_13_04[2], slf_op_13_04[1],
     slf_op_13_04[0]}), .carry_in(tgnd_br_q),
     .bnl_op_01({slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0], slf_op_11_00[3], slf_op_11_00[2],
     slf_op_11_00[1], slf_op_11_00[0]}), .slf_op_04({net1150[0],
     net1150[1], net1150[2], net1150[3], net1150[4], net1150[5],
     net1150[6], net1150[7]}), .slf_op_03({net1140[0], net1140[1],
     net1140[2], net1140[3], net1140[4], net1140[5], net1140[6],
     net1140[7]}), .slf_op_01({net913[0], net913[1], net913[2],
     net913[3], net913[4], net913[5], net913[6], net913[7]}),
     .sp4_h_l_04({net1169[0], net1169[1], net1169[2], net1169[3],
     net1169[4], net1169[5], net1169[6], net1169[7], net1169[8],
     net1169[9], net1169[10], net1169[11], net1169[12], net1169[13],
     net1169[14], net1169[15], net1169[16], net1169[17], net1169[18],
     net1169[19], net1169[20], net1169[21], net1169[22], net1169[23],
     net1169[24], net1169[25], net1169[26], net1169[27], net1169[28],
     net1169[29], net1169[30], net1169[31], net1169[32], net1169[33],
     net1169[34], net1169[35], net1169[36], net1169[37], net1169[38],
     net1169[39], net1169[40], net1169[41], net1169[42], net1169[43],
     net1169[44], net1169[45], net1169[46], net1169[47]}),
     .carry_out(carry_out_12_08), .vdd_cntl(vdd_cntl_r[143:16]),
     .sp12_h_r_04({net969[0], net969[1], net969[2], net969[3],
     net969[4], net969[5], net969[6], net969[7], net969[8], net969[9],
     net969[10], net969[11], net969[12], net969[13], net969[14],
     net969[15], net969[16], net969[17], net969[18], net969[19],
     net969[20], net969[21], net969[22], net969[23]}),
     .sp12_h_r_03({net970[0], net970[1], net970[2], net970[3],
     net970[4], net970[5], net970[6], net970[7], net970[8], net970[9],
     net970[10], net970[11], net970[12], net970[13], net970[14],
     net970[15], net970[16], net970[17], net970[18], net970[19],
     net970[20], net970[21], net970[22], net970[23]}),
     .sp12_h_r_02({net971[0], net971[1], net971[2], net971[3],
     net971[4], net971[5], net971[6], net971[7], net971[8], net971[9],
     net971[10], net971[11], net971[12], net971[13], net971[14],
     net971[15], net971[16], net971[17], net971[18], net971[19],
     net971[20], net971[21], net971[22], net971[23]}),
     .sp12_h_r_01({net972[0], net972[1], net972[2], net972[3],
     net972[4], net972[5], net972[6], net972[7], net972[8], net972[9],
     net972[10], net972[11], net972[12], net972[13], net972[14],
     net972[15], net972[16], net972[17], net972[18], net972[19],
     net972[20], net972[21], net972[22], net972[23]}),
     .glb_netwk_col(clk_tree_drv_br[7:0]), .sp4_v_b_01({net1168[0],
     net1168[1], net1168[2], net1168[3], net1168[4], net1168[5],
     net1168[6], net1168[7], net1168[8], net1168[9], net1168[10],
     net1168[11], net1168[12], net1168[13], net1168[14], net1168[15],
     net1168[16], net1168[17], net1168[18], net1168[19], net1168[20],
     net1168[21], net1168[22], net1168[23], net1168[24], net1168[25],
     net1168[26], net1168[27], net1168[28], net1168[29], net1168[30],
     net1168[31], net1168[32], net1168[33], net1168[34], net1168[35],
     net1168[36], net1168[37], net1168[38], net1168[39], net1168[40],
     net1168[41], net1168[42], net1168[43], net1168[44], net1168[45],
     net1168[46], net1168[47]}), .sp4_r_v_b_04({net799[0], net799[1],
     net799[2], net799[3], net799[4], net799[5], net799[6], net799[7],
     net799[8], net799[9], net799[10], net799[11], net799[12],
     net799[13], net799[14], net799[15], net799[16], net799[17],
     net799[18], net799[19], net799[20], net799[21], net799[22],
     net799[23], net799[24], net799[25], net799[26], net799[27],
     net799[28], net799[29], net799[30], net799[31], net799[32],
     net799[33], net799[34], net799[35], net799[36], net799[37],
     net799[38], net799[39], net799[40], net799[41], net799[42],
     net799[43], net799[44], net799[45], net799[46], net799[47]}),
     .sp4_r_v_b_03({net976[0], net976[1], net976[2], net976[3],
     net976[4], net976[5], net976[6], net976[7], net976[8], net976[9],
     net976[10], net976[11], net976[12], net976[13], net976[14],
     net976[15], net976[16], net976[17], net976[18], net976[19],
     net976[20], net976[21], net976[22], net976[23], net976[24],
     net976[25], net976[26], net976[27], net976[28], net976[29],
     net976[30], net976[31], net976[32], net976[33], net976[34],
     net976[35], net976[36], net976[37], net976[38], net976[39],
     net976[40], net976[41], net976[42], net976[43], net976[44],
     net976[45], net976[46], net976[47]}), .sp4_r_v_b_02({net977[0],
     net977[1], net977[2], net977[3], net977[4], net977[5], net977[6],
     net977[7], net977[8], net977[9], net977[10], net977[11],
     net977[12], net977[13], net977[14], net977[15], net977[16],
     net977[17], net977[18], net977[19], net977[20], net977[21],
     net977[22], net977[23], net977[24], net977[25], net977[26],
     net977[27], net977[28], net977[29], net977[30], net977[31],
     net977[32], net977[33], net977[34], net977[35], net977[36],
     net977[37], net977[38], net977[39], net977[40], net977[41],
     net977[42], net977[43], net977[44], net977[45], net977[46],
     net977[47]}), .sp4_r_v_b_01({net805[0], net805[1], net805[2],
     net805[3], net805[4], net805[5], net805[6], net805[7], net805[8],
     net805[9], net805[10], net805[11], net805[12], net805[13],
     net805[14], net805[15], net805[16], net805[17], net805[18],
     net805[19], net805[20], net805[21], net805[22], net805[23],
     net805[24], net805[25], net805[26], net805[27], net805[28],
     net805[29], net805[30], net805[31], net805[32], net805[33],
     net805[34], net805[35], net805[36], net805[37], net805[38],
     net805[39], net805[40], net805[41], net805[42], net805[43],
     net805[44], net805[45], net805[46], net805[47]}),
     .sp4_h_r_04({net979[0], net979[1], net979[2], net979[3],
     net979[4], net979[5], net979[6], net979[7], net979[8], net979[9],
     net979[10], net979[11], net979[12], net979[13], net979[14],
     net979[15], net979[16], net979[17], net979[18], net979[19],
     net979[20], net979[21], net979[22], net979[23], net979[24],
     net979[25], net979[26], net979[27], net979[28], net979[29],
     net979[30], net979[31], net979[32], net979[33], net979[34],
     net979[35], net979[36], net979[37], net979[38], net979[39],
     net979[40], net979[41], net979[42], net979[43], net979[44],
     net979[45], net979[46], net979[47]}), .sp4_h_r_03({net980[0],
     net980[1], net980[2], net980[3], net980[4], net980[5], net980[6],
     net980[7], net980[8], net980[9], net980[10], net980[11],
     net980[12], net980[13], net980[14], net980[15], net980[16],
     net980[17], net980[18], net980[19], net980[20], net980[21],
     net980[22], net980[23], net980[24], net980[25], net980[26],
     net980[27], net980[28], net980[29], net980[30], net980[31],
     net980[32], net980[33], net980[34], net980[35], net980[36],
     net980[37], net980[38], net980[39], net980[40], net980[41],
     net980[42], net980[43], net980[44], net980[45], net980[46],
     net980[47]}), .sp4_h_r_02({net981[0], net981[1], net981[2],
     net981[3], net981[4], net981[5], net981[6], net981[7], net981[8],
     net981[9], net981[10], net981[11], net981[12], net981[13],
     net981[14], net981[15], net981[16], net981[17], net981[18],
     net981[19], net981[20], net981[21], net981[22], net981[23],
     net981[24], net981[25], net981[26], net981[27], net981[28],
     net981[29], net981[30], net981[31], net981[32], net981[33],
     net981[34], net981[35], net981[36], net981[37], net981[38],
     net981[39], net981[40], net981[41], net981[42], net981[43],
     net981[44], net981[45], net981[46], net981[47]}),
     .sp4_h_r_01({net982[0], net982[1], net982[2], net982[3],
     net982[4], net982[5], net982[6], net982[7], net982[8], net982[9],
     net982[10], net982[11], net982[12], net982[13], net982[14],
     net982[15], net982[16], net982[17], net982[18], net982[19],
     net982[20], net982[21], net982[22], net982[23], net982[24],
     net982[25], net982[26], net982[27], net982[28], net982[29],
     net982[30], net982[31], net982[32], net982[33], net982[34],
     net982[35], net982[36], net982[37], net982[38], net982[39],
     net982[40], net982[41], net982[42], net982[43], net982[44],
     net982[45], net982[46], net982[47]}), .sp4_h_l_03({net1170[0],
     net1170[1], net1170[2], net1170[3], net1170[4], net1170[5],
     net1170[6], net1170[7], net1170[8], net1170[9], net1170[10],
     net1170[11], net1170[12], net1170[13], net1170[14], net1170[15],
     net1170[16], net1170[17], net1170[18], net1170[19], net1170[20],
     net1170[21], net1170[22], net1170[23], net1170[24], net1170[25],
     net1170[26], net1170[27], net1170[28], net1170[29], net1170[30],
     net1170[31], net1170[32], net1170[33], net1170[34], net1170[35],
     net1170[36], net1170[37], net1170[38], net1170[39], net1170[40],
     net1170[41], net1170[42], net1170[43], net1170[44], net1170[45],
     net1170[46], net1170[47]}), .sp4_h_l_02({net1171[0], net1171[1],
     net1171[2], net1171[3], net1171[4], net1171[5], net1171[6],
     net1171[7], net1171[8], net1171[9], net1171[10], net1171[11],
     net1171[12], net1171[13], net1171[14], net1171[15], net1171[16],
     net1171[17], net1171[18], net1171[19], net1171[20], net1171[21],
     net1171[22], net1171[23], net1171[24], net1171[25], net1171[26],
     net1171[27], net1171[28], net1171[29], net1171[30], net1171[31],
     net1171[32], net1171[33], net1171[34], net1171[35], net1171[36],
     net1171[37], net1171[38], net1171[39], net1171[40], net1171[41],
     net1171[42], net1171[43], net1171[44], net1171[45], net1171[46],
     net1171[47]}), .sp4_h_l_01({net1172[0], net1172[1], net1172[2],
     net1172[3], net1172[4], net1172[5], net1172[6], net1172[7],
     net1172[8], net1172[9], net1172[10], net1172[11], net1172[12],
     net1172[13], net1172[14], net1172[15], net1172[16], net1172[17],
     net1172[18], net1172[19], net1172[20], net1172[21], net1172[22],
     net1172[23], net1172[24], net1172[25], net1172[26], net1172[27],
     net1172[28], net1172[29], net1172[30], net1172[31], net1172[32],
     net1172[33], net1172[34], net1172[35], net1172[36], net1172[37],
     net1172[38], net1172[39], net1172[40], net1172[41], net1172[42],
     net1172[43], net1172[44], net1172[45], net1172[46], net1172[47]}),
     .bl(bl[311:258]), .bot_op_01({slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0], slf_op_12_00[3],
     slf_op_12_00[2], slf_op_12_00[1], slf_op_12_00[0]}),
     .sp12_h_l_01({net1162[0], net1162[1], net1162[2], net1162[3],
     net1162[4], net1162[5], net1162[6], net1162[7], net1162[8],
     net1162[9], net1162[10], net1162[11], net1162[12], net1162[13],
     net1162[14], net1162[15], net1162[16], net1162[17], net1162[18],
     net1162[19], net1162[20], net1162[21], net1162[22], net1162[23]}),
     .sp12_h_l_02({net1161[0], net1161[1], net1161[2], net1161[3],
     net1161[4], net1161[5], net1161[6], net1161[7], net1161[8],
     net1161[9], net1161[10], net1161[11], net1161[12], net1161[13],
     net1161[14], net1161[15], net1161[16], net1161[17], net1161[18],
     net1161[19], net1161[20], net1161[21], net1161[22], net1161[23]}),
     .sp12_h_l_03({net1160[0], net1160[1], net1160[2], net1160[3],
     net1160[4], net1160[5], net1160[6], net1160[7], net1160[8],
     net1160[9], net1160[10], net1160[11], net1160[12], net1160[13],
     net1160[14], net1160[15], net1160[16], net1160[17], net1160[18],
     net1160[19], net1160[20], net1160[21], net1160[22], net1160[23]}),
     .sp12_h_l_04({net1159[0], net1159[1], net1159[2], net1159[3],
     net1159[4], net1159[5], net1159[6], net1159[7], net1159[8],
     net1159[9], net1159[10], net1159[11], net1159[12], net1159[13],
     net1159[14], net1159[15], net1159[16], net1159[17], net1159[18],
     net1159[19], net1159[20], net1159[21], net1159[22], net1159[23]}),
     .sp4_v_b_04({net1165[0], net1165[1], net1165[2], net1165[3],
     net1165[4], net1165[5], net1165[6], net1165[7], net1165[8],
     net1165[9], net1165[10], net1165[11], net1165[12], net1165[13],
     net1165[14], net1165[15], net1165[16], net1165[17], net1165[18],
     net1165[19], net1165[20], net1165[21], net1165[22], net1165[23],
     net1165[24], net1165[25], net1165[26], net1165[27], net1165[28],
     net1165[29], net1165[30], net1165[31], net1165[32], net1165[33],
     net1165[34], net1165[35], net1165[36], net1165[37], net1165[38],
     net1165[39], net1165[40], net1165[41], net1165[42], net1165[43],
     net1165[44], net1165[45], net1165[46], net1165[47]}),
     .sp4_v_b_03({net1166[0], net1166[1], net1166[2], net1166[3],
     net1166[4], net1166[5], net1166[6], net1166[7], net1166[8],
     net1166[9], net1166[10], net1166[11], net1166[12], net1166[13],
     net1166[14], net1166[15], net1166[16], net1166[17], net1166[18],
     net1166[19], net1166[20], net1166[21], net1166[22], net1166[23],
     net1166[24], net1166[25], net1166[26], net1166[27], net1166[28],
     net1166[29], net1166[30], net1166[31], net1166[32], net1166[33],
     net1166[34], net1166[35], net1166[36], net1166[37], net1166[38],
     net1166[39], net1166[40], net1166[41], net1166[42], net1166[43],
     net1166[44], net1166[45], net1166[46], net1166[47]}),
     .sp4_v_b_02({net1167[0], net1167[1], net1167[2], net1167[3],
     net1167[4], net1167[5], net1167[6], net1167[7], net1167[8],
     net1167[9], net1167[10], net1167[11], net1167[12], net1167[13],
     net1167[14], net1167[15], net1167[16], net1167[17], net1167[18],
     net1167[19], net1167[20], net1167[21], net1167[22], net1167[23],
     net1167[24], net1167[25], net1167[26], net1167[27], net1167[28],
     net1167[29], net1167[30], net1167[31], net1167[32], net1167[33],
     net1167[34], net1167[35], net1167[36], net1167[37], net1167[38],
     net1167[39], net1167[40], net1167[41], net1167[42], net1167[43],
     net1167[44], net1167[45], net1167[46], net1167[47]}),
     .bnr_op_01({pll_sdo, pll_sdo, pll_sdo, pll_sdo, pll_sdo, pll_sdo,
     pll_sdo, pll_sdo}), .sp4_h_l_05({net1193[0], net1193[1],
     net1193[2], net1193[3], net1193[4], net1193[5], net1193[6],
     net1193[7], net1193[8], net1193[9], net1193[10], net1193[11],
     net1193[12], net1193[13], net1193[14], net1193[15], net1193[16],
     net1193[17], net1193[18], net1193[19], net1193[20], net1193[21],
     net1193[22], net1193[23], net1193[24], net1193[25], net1193[26],
     net1193[27], net1193[28], net1193[29], net1193[30], net1193[31],
     net1193[32], net1193[33], net1193[34], net1193[35], net1193[36],
     net1193[37], net1193[38], net1193[39], net1193[40], net1193[41],
     net1193[42], net1193[43], net1193[44], net1193[45], net1193[46],
     net1193[47]}), .sp4_h_l_06({net1192[0], net1192[1], net1192[2],
     net1192[3], net1192[4], net1192[5], net1192[6], net1192[7],
     net1192[8], net1192[9], net1192[10], net1192[11], net1192[12],
     net1192[13], net1192[14], net1192[15], net1192[16], net1192[17],
     net1192[18], net1192[19], net1192[20], net1192[21], net1192[22],
     net1192[23], net1192[24], net1192[25], net1192[26], net1192[27],
     net1192[28], net1192[29], net1192[30], net1192[31], net1192[32],
     net1192[33], net1192[34], net1192[35], net1192[36], net1192[37],
     net1192[38], net1192[39], net1192[40], net1192[41], net1192[42],
     net1192[43], net1192[44], net1192[45], net1192[46], net1192[47]}),
     .sp4_h_l_07({net1191[0], net1191[1], net1191[2], net1191[3],
     net1191[4], net1191[5], net1191[6], net1191[7], net1191[8],
     net1191[9], net1191[10], net1191[11], net1191[12], net1191[13],
     net1191[14], net1191[15], net1191[16], net1191[17], net1191[18],
     net1191[19], net1191[20], net1191[21], net1191[22], net1191[23],
     net1191[24], net1191[25], net1191[26], net1191[27], net1191[28],
     net1191[29], net1191[30], net1191[31], net1191[32], net1191[33],
     net1191[34], net1191[35], net1191[36], net1191[37], net1191[38],
     net1191[39], net1191[40], net1191[41], net1191[42], net1191[43],
     net1191[44], net1191[45], net1191[46], net1191[47]}),
     .sp4_h_l_08({net1190[0], net1190[1], net1190[2], net1190[3],
     net1190[4], net1190[5], net1190[6], net1190[7], net1190[8],
     net1190[9], net1190[10], net1190[11], net1190[12], net1190[13],
     net1190[14], net1190[15], net1190[16], net1190[17], net1190[18],
     net1190[19], net1190[20], net1190[21], net1190[22], net1190[23],
     net1190[24], net1190[25], net1190[26], net1190[27], net1190[28],
     net1190[29], net1190[30], net1190[31], net1190[32], net1190[33],
     net1190[34], net1190[35], net1190[36], net1190[37], net1190[38],
     net1190[39], net1190[40], net1190[41], net1190[42], net1190[43],
     net1190[44], net1190[45], net1190[46], net1190[47]}),
     .sp4_h_r_08({net1000[0], net1000[1], net1000[2], net1000[3],
     net1000[4], net1000[5], net1000[6], net1000[7], net1000[8],
     net1000[9], net1000[10], net1000[11], net1000[12], net1000[13],
     net1000[14], net1000[15], net1000[16], net1000[17], net1000[18],
     net1000[19], net1000[20], net1000[21], net1000[22], net1000[23],
     net1000[24], net1000[25], net1000[26], net1000[27], net1000[28],
     net1000[29], net1000[30], net1000[31], net1000[32], net1000[33],
     net1000[34], net1000[35], net1000[36], net1000[37], net1000[38],
     net1000[39], net1000[40], net1000[41], net1000[42], net1000[43],
     net1000[44], net1000[45], net1000[46], net1000[47]}),
     .sp4_h_r_07({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7], net1001[8],
     net1001[9], net1001[10], net1001[11], net1001[12], net1001[13],
     net1001[14], net1001[15], net1001[16], net1001[17], net1001[18],
     net1001[19], net1001[20], net1001[21], net1001[22], net1001[23],
     net1001[24], net1001[25], net1001[26], net1001[27], net1001[28],
     net1001[29], net1001[30], net1001[31], net1001[32], net1001[33],
     net1001[34], net1001[35], net1001[36], net1001[37], net1001[38],
     net1001[39], net1001[40], net1001[41], net1001[42], net1001[43],
     net1001[44], net1001[45], net1001[46], net1001[47]}),
     .sp4_h_r_06({net1002[0], net1002[1], net1002[2], net1002[3],
     net1002[4], net1002[5], net1002[6], net1002[7], net1002[8],
     net1002[9], net1002[10], net1002[11], net1002[12], net1002[13],
     net1002[14], net1002[15], net1002[16], net1002[17], net1002[18],
     net1002[19], net1002[20], net1002[21], net1002[22], net1002[23],
     net1002[24], net1002[25], net1002[26], net1002[27], net1002[28],
     net1002[29], net1002[30], net1002[31], net1002[32], net1002[33],
     net1002[34], net1002[35], net1002[36], net1002[37], net1002[38],
     net1002[39], net1002[40], net1002[41], net1002[42], net1002[43],
     net1002[44], net1002[45], net1002[46], net1002[47]}),
     .sp4_h_r_05({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7], net1003[8],
     net1003[9], net1003[10], net1003[11], net1003[12], net1003[13],
     net1003[14], net1003[15], net1003[16], net1003[17], net1003[18],
     net1003[19], net1003[20], net1003[21], net1003[22], net1003[23],
     net1003[24], net1003[25], net1003[26], net1003[27], net1003[28],
     net1003[29], net1003[30], net1003[31], net1003[32], net1003[33],
     net1003[34], net1003[35], net1003[36], net1003[37], net1003[38],
     net1003[39], net1003[40], net1003[41], net1003[42], net1003[43],
     net1003[44], net1003[45], net1003[46], net1003[47]}),
     .slf_op_05({net1201[0], net1201[1], net1201[2], net1201[3],
     net1201[4], net1201[5], net1201[6], net1201[7]}),
     .slf_op_06({net1200[0], net1200[1], net1200[2], net1200[3],
     net1200[4], net1200[5], net1200[6], net1200[7]}),
     .slf_op_07({net1199[0], net1199[1], net1199[2], net1199[3],
     net1199[4], net1199[5], net1199[6], net1199[7]}),
     .slf_op_08(slf_op_12_08[7:0]), .rgt_op_08({slf_op_13_08[3],
     slf_op_13_08[2], slf_op_13_08[1], slf_op_13_08[0],
     slf_op_13_08[3], slf_op_13_08[2], slf_op_13_08[1],
     slf_op_13_08[0]}), .rgt_op_07({slf_op_13_07[3], slf_op_13_07[2],
     slf_op_13_07[1], slf_op_13_07[0], slf_op_13_07[3],
     slf_op_13_07[2], slf_op_13_07[1], slf_op_13_07[0]}),
     .rgt_op_06({slf_op_13_06[3], slf_op_13_06[2], slf_op_13_06[1],
     slf_op_13_06[0], slf_op_13_06[3], slf_op_13_06[2],
     slf_op_13_06[1], slf_op_13_06[0]}), .rgt_op_05({slf_op_13_05[3],
     slf_op_13_05[2], slf_op_13_05[1], slf_op_13_05[0],
     slf_op_13_05[3], slf_op_13_05[2], slf_op_13_05[1],
     slf_op_13_05[0]}), .lft_op_08(slf_op_11_08[7:0]),
     .lft_op_07({net1528[0], net1528[1], net1528[2], net1528[3],
     net1528[4], net1528[5], net1528[6], net1528[7]}),
     .lft_op_06({net1529[0], net1529[1], net1529[2], net1529[3],
     net1529[4], net1529[5], net1529[6], net1529[7]}),
     .lft_op_05({net1530[0], net1530[1], net1530[2], net1530[3],
     net1530[4], net1530[5], net1530[6], net1530[7]}),
     .sp12_h_l_08({net1212[0], net1212[1], net1212[2], net1212[3],
     net1212[4], net1212[5], net1212[6], net1212[7], net1212[8],
     net1212[9], net1212[10], net1212[11], net1212[12], net1212[13],
     net1212[14], net1212[15], net1212[16], net1212[17], net1212[18],
     net1212[19], net1212[20], net1212[21], net1212[22], net1212[23]}),
     .sp12_h_l_07({net1211[0], net1211[1], net1211[2], net1211[3],
     net1211[4], net1211[5], net1211[6], net1211[7], net1211[8],
     net1211[9], net1211[10], net1211[11], net1211[12], net1211[13],
     net1211[14], net1211[15], net1211[16], net1211[17], net1211[18],
     net1211[19], net1211[20], net1211[21], net1211[22], net1211[23]}),
     .sp12_h_l_06({net1210[0], net1210[1], net1210[2], net1210[3],
     net1210[4], net1210[5], net1210[6], net1210[7], net1210[8],
     net1210[9], net1210[10], net1210[11], net1210[12], net1210[13],
     net1210[14], net1210[15], net1210[16], net1210[17], net1210[18],
     net1210[19], net1210[20], net1210[21], net1210[22], net1210[23]}),
     .sp12_h_r_05({net1019[0], net1019[1], net1019[2], net1019[3],
     net1019[4], net1019[5], net1019[6], net1019[7], net1019[8],
     net1019[9], net1019[10], net1019[11], net1019[12], net1019[13],
     net1019[14], net1019[15], net1019[16], net1019[17], net1019[18],
     net1019[19], net1019[20], net1019[21], net1019[22], net1019[23]}),
     .sp12_h_r_06({net1020[0], net1020[1], net1020[2], net1020[3],
     net1020[4], net1020[5], net1020[6], net1020[7], net1020[8],
     net1020[9], net1020[10], net1020[11], net1020[12], net1020[13],
     net1020[14], net1020[15], net1020[16], net1020[17], net1020[18],
     net1020[19], net1020[20], net1020[21], net1020[22], net1020[23]}),
     .sp12_h_r_07({net1021[0], net1021[1], net1021[2], net1021[3],
     net1021[4], net1021[5], net1021[6], net1021[7], net1021[8],
     net1021[9], net1021[10], net1021[11], net1021[12], net1021[13],
     net1021[14], net1021[15], net1021[16], net1021[17], net1021[18],
     net1021[19], net1021[20], net1021[21], net1021[22], net1021[23]}),
     .sp12_h_r_08({net1022[0], net1022[1], net1022[2], net1022[3],
     net1022[4], net1022[5], net1022[6], net1022[7], net1022[8],
     net1022[9], net1022[10], net1022[11], net1022[12], net1022[13],
     net1022[14], net1022[15], net1022[16], net1022[17], net1022[18],
     net1022[19], net1022[20], net1022[21], net1022[22], net1022[23]}),
     .sp12_h_l_05({net1209[0], net1209[1], net1209[2], net1209[3],
     net1209[4], net1209[5], net1209[6], net1209[7], net1209[8],
     net1209[9], net1209[10], net1209[11], net1209[12], net1209[13],
     net1209[14], net1209[15], net1209[16], net1209[17], net1209[18],
     net1209[19], net1209[20], net1209[21], net1209[22], net1209[23]}),
     .sp4_r_v_b_05({net802[0], net802[1], net802[2], net802[3],
     net802[4], net802[5], net802[6], net802[7], net802[8], net802[9],
     net802[10], net802[11], net802[12], net802[13], net802[14],
     net802[15], net802[16], net802[17], net802[18], net802[19],
     net802[20], net802[21], net802[22], net802[23], net802[24],
     net802[25], net802[26], net802[27], net802[28], net802[29],
     net802[30], net802[31], net802[32], net802[33], net802[34],
     net802[35], net802[36], net802[37], net802[38], net802[39],
     net802[40], net802[41], net802[42], net802[43], net802[44],
     net802[45], net802[46], net802[47]}), .sp4_r_v_b_06({net1025[0],
     net1025[1], net1025[2], net1025[3], net1025[4], net1025[5],
     net1025[6], net1025[7], net1025[8], net1025[9], net1025[10],
     net1025[11], net1025[12], net1025[13], net1025[14], net1025[15],
     net1025[16], net1025[17], net1025[18], net1025[19], net1025[20],
     net1025[21], net1025[22], net1025[23], net1025[24], net1025[25],
     net1025[26], net1025[27], net1025[28], net1025[29], net1025[30],
     net1025[31], net1025[32], net1025[33], net1025[34], net1025[35],
     net1025[36], net1025[37], net1025[38], net1025[39], net1025[40],
     net1025[41], net1025[42], net1025[43], net1025[44], net1025[45],
     net1025[46], net1025[47]}), .sp4_r_v_b_07({net800[0], net800[1],
     net800[2], net800[3], net800[4], net800[5], net800[6], net800[7],
     net800[8], net800[9], net800[10], net800[11], net800[12],
     net800[13], net800[14], net800[15], net800[16], net800[17],
     net800[18], net800[19], net800[20], net800[21], net800[22],
     net800[23], net800[24], net800[25], net800[26], net800[27],
     net800[28], net800[29], net800[30], net800[31], net800[32],
     net800[33], net800[34], net800[35], net800[36], net800[37],
     net800[38], net800[39], net800[40], net800[41], net800[42],
     net800[43], net800[44], net800[45], net800[46], net800[47]}),
     .sp4_r_v_b_08({net1027[0], net1027[1], net1027[2], net1027[3],
     net1027[4], net1027[5], net1027[6], net1027[7], net1027[8],
     net1027[9], net1027[10], net1027[11], net1027[12], net1027[13],
     net1027[14], net1027[15], net1027[16], net1027[17], net1027[18],
     net1027[19], net1027[20], net1027[21], net1027[22], net1027[23],
     net1027[24], net1027[25], net1027[26], net1027[27], net1027[28],
     net1027[29], net1027[30], net1027[31], net1027[32], net1027[33],
     net1027[34], net1027[35], net1027[36], net1027[37], net1027[38],
     net1027[39], net1027[40], net1027[41], net1027[42], net1027[43],
     net1027[44], net1027[45], net1027[46], net1027[47]}),
     .sp4_v_b_08({net1217[0], net1217[1], net1217[2], net1217[3],
     net1217[4], net1217[5], net1217[6], net1217[7], net1217[8],
     net1217[9], net1217[10], net1217[11], net1217[12], net1217[13],
     net1217[14], net1217[15], net1217[16], net1217[17], net1217[18],
     net1217[19], net1217[20], net1217[21], net1217[22], net1217[23],
     net1217[24], net1217[25], net1217[26], net1217[27], net1217[28],
     net1217[29], net1217[30], net1217[31], net1217[32], net1217[33],
     net1217[34], net1217[35], net1217[36], net1217[37], net1217[38],
     net1217[39], net1217[40], net1217[41], net1217[42], net1217[43],
     net1217[44], net1217[45], net1217[46], net1217[47]}),
     .sp4_v_b_07({net1216[0], net1216[1], net1216[2], net1216[3],
     net1216[4], net1216[5], net1216[6], net1216[7], net1216[8],
     net1216[9], net1216[10], net1216[11], net1216[12], net1216[13],
     net1216[14], net1216[15], net1216[16], net1216[17], net1216[18],
     net1216[19], net1216[20], net1216[21], net1216[22], net1216[23],
     net1216[24], net1216[25], net1216[26], net1216[27], net1216[28],
     net1216[29], net1216[30], net1216[31], net1216[32], net1216[33],
     net1216[34], net1216[35], net1216[36], net1216[37], net1216[38],
     net1216[39], net1216[40], net1216[41], net1216[42], net1216[43],
     net1216[44], net1216[45], net1216[46], net1216[47]}),
     .sp4_v_b_06({net1215[0], net1215[1], net1215[2], net1215[3],
     net1215[4], net1215[5], net1215[6], net1215[7], net1215[8],
     net1215[9], net1215[10], net1215[11], net1215[12], net1215[13],
     net1215[14], net1215[15], net1215[16], net1215[17], net1215[18],
     net1215[19], net1215[20], net1215[21], net1215[22], net1215[23],
     net1215[24], net1215[25], net1215[26], net1215[27], net1215[28],
     net1215[29], net1215[30], net1215[31], net1215[32], net1215[33],
     net1215[34], net1215[35], net1215[36], net1215[37], net1215[38],
     net1215[39], net1215[40], net1215[41], net1215[42], net1215[43],
     net1215[44], net1215[45], net1215[46], net1215[47]}),
     .sp4_v_b_05({net1214[0], net1214[1], net1214[2], net1214[3],
     net1214[4], net1214[5], net1214[6], net1214[7], net1214[8],
     net1214[9], net1214[10], net1214[11], net1214[12], net1214[13],
     net1214[14], net1214[15], net1214[16], net1214[17], net1214[18],
     net1214[19], net1214[20], net1214[21], net1214[22], net1214[23],
     net1214[24], net1214[25], net1214[26], net1214[27], net1214[28],
     net1214[29], net1214[30], net1214[31], net1214[32], net1214[33],
     net1214[34], net1214[35], net1214[36], net1214[37], net1214[38],
     net1214[39], net1214[40], net1214[41], net1214[42], net1214[43],
     net1214[44], net1214[45], net1214[46], net1214[47]}),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .wl(wl_r[143:16]), .sp12_v_t_08(sp12_v_t_12_08[23:0]),
     .tnr_op_08(tnr_op_12_08[7:0]), .top_op_08(top_op_12_08[7:0]),
     .tnl_op_08(tnl_op_12_08[7:0]), .sp4_v_t_08(sp4_v_t_12_08[47:0]),
     .lc_bot(tgnd_br_q), .op_vic(op_vic_12_08),
     .sp12_v_b_01({net898[0], net898[1], net898[2], net898[3],
     net898[4], net898[5], net898[6], net898[7], net898[8], net898[9],
     net898[10], net898[11], net898[12], net898[13], net898[14],
     net898[15], net898[16], net898[17], net898[18], net898[19],
     net898[20], net898[21], net898[22], net898[23]}));
lt_1x8_bot_ice1f I_lt_col_b09 ( .glb_netwk_bot({net937[0], net937[1],
     net937[2], net937[3], net937[4], net937[5], net937[6],
     net937[7]}), .rgt_op_03({net1045[0], net1045[1], net1045[2],
     net1045[3], net1045[4], net1045[5], net1045[6], net1045[7]}),
     .slf_op_02({net1237[0], net1237[1], net1237[2], net1237[3],
     net1237[4], net1237[5], net1237[6], net1237[7]}),
     .rgt_op_02({net1047[0], net1047[1], net1047[2], net1047[3],
     net1047[4], net1047[5], net1047[6], net1047[7]}),
     .rgt_op_01({net784[0], net784[1], net784[2], net784[3], net784[4],
     net784[5], net784[6], net784[7]}), .purst(purst), .prog(prog),
     .lft_op_04({net1340[0], net1340[1], net1340[2], net1340[3],
     net1340[4], net1340[5], net1340[6], net1340[7]}),
     .lft_op_03({net1330[0], net1330[1], net1330[2], net1330[3],
     net1330[4], net1330[5], net1330[6], net1330[7]}),
     .lft_op_02({net1332[0], net1332[1], net1332[2], net1332[3],
     net1332[4], net1332[5], net1332[6], net1332[7]}),
     .lft_op_01({net793[0], net793[1], net793[2], net793[3], net793[4],
     net793[5], net793[6], net793[7]}), .rgt_op_04({net1055[0],
     net1055[1], net1055[2], net1055[3], net1055[4], net1055[5],
     net1055[6], net1055[7]}), .carry_in(tgnd_br_q),
     .bnl_op_01({slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0], slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0]}), .slf_op_04({net1245[0],
     net1245[1], net1245[2], net1245[3], net1245[4], net1245[5],
     net1245[6], net1245[7]}), .slf_op_03({net1235[0], net1235[1],
     net1235[2], net1235[3], net1235[4], net1235[5], net1235[6],
     net1235[7]}), .slf_op_01({net910[0], net910[1], net910[2],
     net910[3], net910[4], net910[5], net910[6], net910[7]}),
     .sp4_h_l_04({net1264[0], net1264[1], net1264[2], net1264[3],
     net1264[4], net1264[5], net1264[6], net1264[7], net1264[8],
     net1264[9], net1264[10], net1264[11], net1264[12], net1264[13],
     net1264[14], net1264[15], net1264[16], net1264[17], net1264[18],
     net1264[19], net1264[20], net1264[21], net1264[22], net1264[23],
     net1264[24], net1264[25], net1264[26], net1264[27], net1264[28],
     net1264[29], net1264[30], net1264[31], net1264[32], net1264[33],
     net1264[34], net1264[35], net1264[36], net1264[37], net1264[38],
     net1264[39], net1264[40], net1264[41], net1264[42], net1264[43],
     net1264[44], net1264[45], net1264[46], net1264[47]}),
     .carry_out(carry_out_09_08), .vdd_cntl(vdd_cntl_r[143:16]),
     .sp12_h_r_04({net1064[0], net1064[1], net1064[2], net1064[3],
     net1064[4], net1064[5], net1064[6], net1064[7], net1064[8],
     net1064[9], net1064[10], net1064[11], net1064[12], net1064[13],
     net1064[14], net1064[15], net1064[16], net1064[17], net1064[18],
     net1064[19], net1064[20], net1064[21], net1064[22], net1064[23]}),
     .sp12_h_r_03({net1065[0], net1065[1], net1065[2], net1065[3],
     net1065[4], net1065[5], net1065[6], net1065[7], net1065[8],
     net1065[9], net1065[10], net1065[11], net1065[12], net1065[13],
     net1065[14], net1065[15], net1065[16], net1065[17], net1065[18],
     net1065[19], net1065[20], net1065[21], net1065[22], net1065[23]}),
     .sp12_h_r_02({net1066[0], net1066[1], net1066[2], net1066[3],
     net1066[4], net1066[5], net1066[6], net1066[7], net1066[8],
     net1066[9], net1066[10], net1066[11], net1066[12], net1066[13],
     net1066[14], net1066[15], net1066[16], net1066[17], net1066[18],
     net1066[19], net1066[20], net1066[21], net1066[22], net1066[23]}),
     .sp12_h_r_01({net1067[0], net1067[1], net1067[2], net1067[3],
     net1067[4], net1067[5], net1067[6], net1067[7], net1067[8],
     net1067[9], net1067[10], net1067[11], net1067[12], net1067[13],
     net1067[14], net1067[15], net1067[16], net1067[17], net1067[18],
     net1067[19], net1067[20], net1067[21], net1067[22], net1067[23]}),
     .glb_netwk_col(clk_tree_drv_br[7:0]), .sp4_v_b_01({net916[0],
     net916[1], net916[2], net916[3], net916[4], net916[5], net916[6],
     net916[7], net916[8], net916[9], net916[10], net916[11],
     net916[12], net916[13], net916[14], net916[15], net916[16],
     net916[17], net916[18], net916[19], net916[20], net916[21],
     net916[22], net916[23], net916[24], net916[25], net916[26],
     net916[27], net916[28], net916[29], net916[30], net916[31],
     net916[32], net916[33], net916[34], net916[35], net916[36],
     net916[37], net916[38], net916[39], net916[40], net916[41],
     net916[42], net916[43], net916[44], net916[45], net916[46],
     net916[47]}), .sp4_r_v_b_04({net1070[0], net1070[1], net1070[2],
     net1070[3], net1070[4], net1070[5], net1070[6], net1070[7],
     net1070[8], net1070[9], net1070[10], net1070[11], net1070[12],
     net1070[13], net1070[14], net1070[15], net1070[16], net1070[17],
     net1070[18], net1070[19], net1070[20], net1070[21], net1070[22],
     net1070[23], net1070[24], net1070[25], net1070[26], net1070[27],
     net1070[28], net1070[29], net1070[30], net1070[31], net1070[32],
     net1070[33], net1070[34], net1070[35], net1070[36], net1070[37],
     net1070[38], net1070[39], net1070[40], net1070[41], net1070[42],
     net1070[43], net1070[44], net1070[45], net1070[46], net1070[47]}),
     .sp4_r_v_b_03({net1071[0], net1071[1], net1071[2], net1071[3],
     net1071[4], net1071[5], net1071[6], net1071[7], net1071[8],
     net1071[9], net1071[10], net1071[11], net1071[12], net1071[13],
     net1071[14], net1071[15], net1071[16], net1071[17], net1071[18],
     net1071[19], net1071[20], net1071[21], net1071[22], net1071[23],
     net1071[24], net1071[25], net1071[26], net1071[27], net1071[28],
     net1071[29], net1071[30], net1071[31], net1071[32], net1071[33],
     net1071[34], net1071[35], net1071[36], net1071[37], net1071[38],
     net1071[39], net1071[40], net1071[41], net1071[42], net1071[43],
     net1071[44], net1071[45], net1071[46], net1071[47]}),
     .sp4_r_v_b_02({net1072[0], net1072[1], net1072[2], net1072[3],
     net1072[4], net1072[5], net1072[6], net1072[7], net1072[8],
     net1072[9], net1072[10], net1072[11], net1072[12], net1072[13],
     net1072[14], net1072[15], net1072[16], net1072[17], net1072[18],
     net1072[19], net1072[20], net1072[21], net1072[22], net1072[23],
     net1072[24], net1072[25], net1072[26], net1072[27], net1072[28],
     net1072[29], net1072[30], net1072[31], net1072[32], net1072[33],
     net1072[34], net1072[35], net1072[36], net1072[37], net1072[38],
     net1072[39], net1072[40], net1072[41], net1072[42], net1072[43],
     net1072[44], net1072[45], net1072[46], net1072[47]}),
     .sp4_r_v_b_01({net907[0], net907[1], net907[2], net907[3],
     net907[4], net907[5], net907[6], net907[7], net907[8], net907[9],
     net907[10], net907[11], net907[12], net907[13], net907[14],
     net907[15], net907[16], net907[17], net907[18], net907[19],
     net907[20], net907[21], net907[22], net907[23], net907[24],
     net907[25], net907[26], net907[27], net907[28], net907[29],
     net907[30], net907[31], net907[32], net907[33], net907[34],
     net907[35], net907[36], net907[37], net907[38], net907[39],
     net907[40], net907[41], net907[42], net907[43], net907[44],
     net907[45], net907[46], net907[47]}), .sp4_h_r_04({net1074[0],
     net1074[1], net1074[2], net1074[3], net1074[4], net1074[5],
     net1074[6], net1074[7], net1074[8], net1074[9], net1074[10],
     net1074[11], net1074[12], net1074[13], net1074[14], net1074[15],
     net1074[16], net1074[17], net1074[18], net1074[19], net1074[20],
     net1074[21], net1074[22], net1074[23], net1074[24], net1074[25],
     net1074[26], net1074[27], net1074[28], net1074[29], net1074[30],
     net1074[31], net1074[32], net1074[33], net1074[34], net1074[35],
     net1074[36], net1074[37], net1074[38], net1074[39], net1074[40],
     net1074[41], net1074[42], net1074[43], net1074[44], net1074[45],
     net1074[46], net1074[47]}), .sp4_h_r_03({net1075[0], net1075[1],
     net1075[2], net1075[3], net1075[4], net1075[5], net1075[6],
     net1075[7], net1075[8], net1075[9], net1075[10], net1075[11],
     net1075[12], net1075[13], net1075[14], net1075[15], net1075[16],
     net1075[17], net1075[18], net1075[19], net1075[20], net1075[21],
     net1075[22], net1075[23], net1075[24], net1075[25], net1075[26],
     net1075[27], net1075[28], net1075[29], net1075[30], net1075[31],
     net1075[32], net1075[33], net1075[34], net1075[35], net1075[36],
     net1075[37], net1075[38], net1075[39], net1075[40], net1075[41],
     net1075[42], net1075[43], net1075[44], net1075[45], net1075[46],
     net1075[47]}), .sp4_h_r_02({net1076[0], net1076[1], net1076[2],
     net1076[3], net1076[4], net1076[5], net1076[6], net1076[7],
     net1076[8], net1076[9], net1076[10], net1076[11], net1076[12],
     net1076[13], net1076[14], net1076[15], net1076[16], net1076[17],
     net1076[18], net1076[19], net1076[20], net1076[21], net1076[22],
     net1076[23], net1076[24], net1076[25], net1076[26], net1076[27],
     net1076[28], net1076[29], net1076[30], net1076[31], net1076[32],
     net1076[33], net1076[34], net1076[35], net1076[36], net1076[37],
     net1076[38], net1076[39], net1076[40], net1076[41], net1076[42],
     net1076[43], net1076[44], net1076[45], net1076[46], net1076[47]}),
     .sp4_h_r_01({net1077[0], net1077[1], net1077[2], net1077[3],
     net1077[4], net1077[5], net1077[6], net1077[7], net1077[8],
     net1077[9], net1077[10], net1077[11], net1077[12], net1077[13],
     net1077[14], net1077[15], net1077[16], net1077[17], net1077[18],
     net1077[19], net1077[20], net1077[21], net1077[22], net1077[23],
     net1077[24], net1077[25], net1077[26], net1077[27], net1077[28],
     net1077[29], net1077[30], net1077[31], net1077[32], net1077[33],
     net1077[34], net1077[35], net1077[36], net1077[37], net1077[38],
     net1077[39], net1077[40], net1077[41], net1077[42], net1077[43],
     net1077[44], net1077[45], net1077[46], net1077[47]}),
     .sp4_h_l_03({net1265[0], net1265[1], net1265[2], net1265[3],
     net1265[4], net1265[5], net1265[6], net1265[7], net1265[8],
     net1265[9], net1265[10], net1265[11], net1265[12], net1265[13],
     net1265[14], net1265[15], net1265[16], net1265[17], net1265[18],
     net1265[19], net1265[20], net1265[21], net1265[22], net1265[23],
     net1265[24], net1265[25], net1265[26], net1265[27], net1265[28],
     net1265[29], net1265[30], net1265[31], net1265[32], net1265[33],
     net1265[34], net1265[35], net1265[36], net1265[37], net1265[38],
     net1265[39], net1265[40], net1265[41], net1265[42], net1265[43],
     net1265[44], net1265[45], net1265[46], net1265[47]}),
     .sp4_h_l_02({net1266[0], net1266[1], net1266[2], net1266[3],
     net1266[4], net1266[5], net1266[6], net1266[7], net1266[8],
     net1266[9], net1266[10], net1266[11], net1266[12], net1266[13],
     net1266[14], net1266[15], net1266[16], net1266[17], net1266[18],
     net1266[19], net1266[20], net1266[21], net1266[22], net1266[23],
     net1266[24], net1266[25], net1266[26], net1266[27], net1266[28],
     net1266[29], net1266[30], net1266[31], net1266[32], net1266[33],
     net1266[34], net1266[35], net1266[36], net1266[37], net1266[38],
     net1266[39], net1266[40], net1266[41], net1266[42], net1266[43],
     net1266[44], net1266[45], net1266[46], net1266[47]}),
     .sp4_h_l_01({net1267[0], net1267[1], net1267[2], net1267[3],
     net1267[4], net1267[5], net1267[6], net1267[7], net1267[8],
     net1267[9], net1267[10], net1267[11], net1267[12], net1267[13],
     net1267[14], net1267[15], net1267[16], net1267[17], net1267[18],
     net1267[19], net1267[20], net1267[21], net1267[22], net1267[23],
     net1267[24], net1267[25], net1267[26], net1267[27], net1267[28],
     net1267[29], net1267[30], net1267[31], net1267[32], net1267[33],
     net1267[34], net1267[35], net1267[36], net1267[37], net1267[38],
     net1267[39], net1267[40], net1267[41], net1267[42], net1267[43],
     net1267[44], net1267[45], net1267[46], net1267[47]}),
     .bl(bl[161:108]), .bot_op_01({slf_op_09_00[3], slf_op_09_00[2],
     slf_op_09_00[1], slf_op_09_00[0], slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0]}),
     .sp12_h_l_01({net1257[0], net1257[1], net1257[2], net1257[3],
     net1257[4], net1257[5], net1257[6], net1257[7], net1257[8],
     net1257[9], net1257[10], net1257[11], net1257[12], net1257[13],
     net1257[14], net1257[15], net1257[16], net1257[17], net1257[18],
     net1257[19], net1257[20], net1257[21], net1257[22], net1257[23]}),
     .sp12_h_l_02({net1256[0], net1256[1], net1256[2], net1256[3],
     net1256[4], net1256[5], net1256[6], net1256[7], net1256[8],
     net1256[9], net1256[10], net1256[11], net1256[12], net1256[13],
     net1256[14], net1256[15], net1256[16], net1256[17], net1256[18],
     net1256[19], net1256[20], net1256[21], net1256[22], net1256[23]}),
     .sp12_h_l_03({net1255[0], net1255[1], net1255[2], net1255[3],
     net1255[4], net1255[5], net1255[6], net1255[7], net1255[8],
     net1255[9], net1255[10], net1255[11], net1255[12], net1255[13],
     net1255[14], net1255[15], net1255[16], net1255[17], net1255[18],
     net1255[19], net1255[20], net1255[21], net1255[22], net1255[23]}),
     .sp12_h_l_04({net1254[0], net1254[1], net1254[2], net1254[3],
     net1254[4], net1254[5], net1254[6], net1254[7], net1254[8],
     net1254[9], net1254[10], net1254[11], net1254[12], net1254[13],
     net1254[14], net1254[15], net1254[16], net1254[17], net1254[18],
     net1254[19], net1254[20], net1254[21], net1254[22], net1254[23]}),
     .sp4_v_b_04({net1260[0], net1260[1], net1260[2], net1260[3],
     net1260[4], net1260[5], net1260[6], net1260[7], net1260[8],
     net1260[9], net1260[10], net1260[11], net1260[12], net1260[13],
     net1260[14], net1260[15], net1260[16], net1260[17], net1260[18],
     net1260[19], net1260[20], net1260[21], net1260[22], net1260[23],
     net1260[24], net1260[25], net1260[26], net1260[27], net1260[28],
     net1260[29], net1260[30], net1260[31], net1260[32], net1260[33],
     net1260[34], net1260[35], net1260[36], net1260[37], net1260[38],
     net1260[39], net1260[40], net1260[41], net1260[42], net1260[43],
     net1260[44], net1260[45], net1260[46], net1260[47]}),
     .sp4_v_b_03({net1261[0], net1261[1], net1261[2], net1261[3],
     net1261[4], net1261[5], net1261[6], net1261[7], net1261[8],
     net1261[9], net1261[10], net1261[11], net1261[12], net1261[13],
     net1261[14], net1261[15], net1261[16], net1261[17], net1261[18],
     net1261[19], net1261[20], net1261[21], net1261[22], net1261[23],
     net1261[24], net1261[25], net1261[26], net1261[27], net1261[28],
     net1261[29], net1261[30], net1261[31], net1261[32], net1261[33],
     net1261[34], net1261[35], net1261[36], net1261[37], net1261[38],
     net1261[39], net1261[40], net1261[41], net1261[42], net1261[43],
     net1261[44], net1261[45], net1261[46], net1261[47]}),
     .sp4_v_b_02({net1262[0], net1262[1], net1262[2], net1262[3],
     net1262[4], net1262[5], net1262[6], net1262[7], net1262[8],
     net1262[9], net1262[10], net1262[11], net1262[12], net1262[13],
     net1262[14], net1262[15], net1262[16], net1262[17], net1262[18],
     net1262[19], net1262[20], net1262[21], net1262[22], net1262[23],
     net1262[24], net1262[25], net1262[26], net1262[27], net1262[28],
     net1262[29], net1262[30], net1262[31], net1262[32], net1262[33],
     net1262[34], net1262[35], net1262[36], net1262[37], net1262[38],
     net1262[39], net1262[40], net1262[41], net1262[42], net1262[43],
     net1262[44], net1262[45], net1262[46], net1262[47]}),
     .bnr_op_01({slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0], slf_op_10_00[3], slf_op_10_00[2],
     slf_op_10_00[1], slf_op_10_00[0]}), .sp4_h_l_05({net1288[0],
     net1288[1], net1288[2], net1288[3], net1288[4], net1288[5],
     net1288[6], net1288[7], net1288[8], net1288[9], net1288[10],
     net1288[11], net1288[12], net1288[13], net1288[14], net1288[15],
     net1288[16], net1288[17], net1288[18], net1288[19], net1288[20],
     net1288[21], net1288[22], net1288[23], net1288[24], net1288[25],
     net1288[26], net1288[27], net1288[28], net1288[29], net1288[30],
     net1288[31], net1288[32], net1288[33], net1288[34], net1288[35],
     net1288[36], net1288[37], net1288[38], net1288[39], net1288[40],
     net1288[41], net1288[42], net1288[43], net1288[44], net1288[45],
     net1288[46], net1288[47]}), .sp4_h_l_06({net1287[0], net1287[1],
     net1287[2], net1287[3], net1287[4], net1287[5], net1287[6],
     net1287[7], net1287[8], net1287[9], net1287[10], net1287[11],
     net1287[12], net1287[13], net1287[14], net1287[15], net1287[16],
     net1287[17], net1287[18], net1287[19], net1287[20], net1287[21],
     net1287[22], net1287[23], net1287[24], net1287[25], net1287[26],
     net1287[27], net1287[28], net1287[29], net1287[30], net1287[31],
     net1287[32], net1287[33], net1287[34], net1287[35], net1287[36],
     net1287[37], net1287[38], net1287[39], net1287[40], net1287[41],
     net1287[42], net1287[43], net1287[44], net1287[45], net1287[46],
     net1287[47]}), .sp4_h_l_07({net1286[0], net1286[1], net1286[2],
     net1286[3], net1286[4], net1286[5], net1286[6], net1286[7],
     net1286[8], net1286[9], net1286[10], net1286[11], net1286[12],
     net1286[13], net1286[14], net1286[15], net1286[16], net1286[17],
     net1286[18], net1286[19], net1286[20], net1286[21], net1286[22],
     net1286[23], net1286[24], net1286[25], net1286[26], net1286[27],
     net1286[28], net1286[29], net1286[30], net1286[31], net1286[32],
     net1286[33], net1286[34], net1286[35], net1286[36], net1286[37],
     net1286[38], net1286[39], net1286[40], net1286[41], net1286[42],
     net1286[43], net1286[44], net1286[45], net1286[46], net1286[47]}),
     .sp4_h_l_08({net1285[0], net1285[1], net1285[2], net1285[3],
     net1285[4], net1285[5], net1285[6], net1285[7], net1285[8],
     net1285[9], net1285[10], net1285[11], net1285[12], net1285[13],
     net1285[14], net1285[15], net1285[16], net1285[17], net1285[18],
     net1285[19], net1285[20], net1285[21], net1285[22], net1285[23],
     net1285[24], net1285[25], net1285[26], net1285[27], net1285[28],
     net1285[29], net1285[30], net1285[31], net1285[32], net1285[33],
     net1285[34], net1285[35], net1285[36], net1285[37], net1285[38],
     net1285[39], net1285[40], net1285[41], net1285[42], net1285[43],
     net1285[44], net1285[45], net1285[46], net1285[47]}),
     .sp4_h_r_08({net1095[0], net1095[1], net1095[2], net1095[3],
     net1095[4], net1095[5], net1095[6], net1095[7], net1095[8],
     net1095[9], net1095[10], net1095[11], net1095[12], net1095[13],
     net1095[14], net1095[15], net1095[16], net1095[17], net1095[18],
     net1095[19], net1095[20], net1095[21], net1095[22], net1095[23],
     net1095[24], net1095[25], net1095[26], net1095[27], net1095[28],
     net1095[29], net1095[30], net1095[31], net1095[32], net1095[33],
     net1095[34], net1095[35], net1095[36], net1095[37], net1095[38],
     net1095[39], net1095[40], net1095[41], net1095[42], net1095[43],
     net1095[44], net1095[45], net1095[46], net1095[47]}),
     .sp4_h_r_07({net1096[0], net1096[1], net1096[2], net1096[3],
     net1096[4], net1096[5], net1096[6], net1096[7], net1096[8],
     net1096[9], net1096[10], net1096[11], net1096[12], net1096[13],
     net1096[14], net1096[15], net1096[16], net1096[17], net1096[18],
     net1096[19], net1096[20], net1096[21], net1096[22], net1096[23],
     net1096[24], net1096[25], net1096[26], net1096[27], net1096[28],
     net1096[29], net1096[30], net1096[31], net1096[32], net1096[33],
     net1096[34], net1096[35], net1096[36], net1096[37], net1096[38],
     net1096[39], net1096[40], net1096[41], net1096[42], net1096[43],
     net1096[44], net1096[45], net1096[46], net1096[47]}),
     .sp4_h_r_06({net1097[0], net1097[1], net1097[2], net1097[3],
     net1097[4], net1097[5], net1097[6], net1097[7], net1097[8],
     net1097[9], net1097[10], net1097[11], net1097[12], net1097[13],
     net1097[14], net1097[15], net1097[16], net1097[17], net1097[18],
     net1097[19], net1097[20], net1097[21], net1097[22], net1097[23],
     net1097[24], net1097[25], net1097[26], net1097[27], net1097[28],
     net1097[29], net1097[30], net1097[31], net1097[32], net1097[33],
     net1097[34], net1097[35], net1097[36], net1097[37], net1097[38],
     net1097[39], net1097[40], net1097[41], net1097[42], net1097[43],
     net1097[44], net1097[45], net1097[46], net1097[47]}),
     .sp4_h_r_05({net1098[0], net1098[1], net1098[2], net1098[3],
     net1098[4], net1098[5], net1098[6], net1098[7], net1098[8],
     net1098[9], net1098[10], net1098[11], net1098[12], net1098[13],
     net1098[14], net1098[15], net1098[16], net1098[17], net1098[18],
     net1098[19], net1098[20], net1098[21], net1098[22], net1098[23],
     net1098[24], net1098[25], net1098[26], net1098[27], net1098[28],
     net1098[29], net1098[30], net1098[31], net1098[32], net1098[33],
     net1098[34], net1098[35], net1098[36], net1098[37], net1098[38],
     net1098[39], net1098[40], net1098[41], net1098[42], net1098[43],
     net1098[44], net1098[45], net1098[46], net1098[47]}),
     .slf_op_05({net1296[0], net1296[1], net1296[2], net1296[3],
     net1296[4], net1296[5], net1296[6], net1296[7]}),
     .slf_op_06({net1295[0], net1295[1], net1295[2], net1295[3],
     net1295[4], net1295[5], net1295[6], net1295[7]}),
     .slf_op_07({net1294[0], net1294[1], net1294[2], net1294[3],
     net1294[4], net1294[5], net1294[6], net1294[7]}),
     .slf_op_08(slf_op_09_08[7:0]), .rgt_op_08(slf_op_10_08[7:0]),
     .rgt_op_07({net1104[0], net1104[1], net1104[2], net1104[3],
     net1104[4], net1104[5], net1104[6], net1104[7]}),
     .rgt_op_06({net1105[0], net1105[1], net1105[2], net1105[3],
     net1105[4], net1105[5], net1105[6], net1105[7]}),
     .rgt_op_05({net1106[0], net1106[1], net1106[2], net1106[3],
     net1106[4], net1106[5], net1106[6], net1106[7]}),
     .lft_op_08(slf_op_08_08[7:0]), .lft_op_07({net1389[0], net1389[1],
     net1389[2], net1389[3], net1389[4], net1389[5], net1389[6],
     net1389[7]}), .lft_op_06({net1390[0], net1390[1], net1390[2],
     net1390[3], net1390[4], net1390[5], net1390[6], net1390[7]}),
     .lft_op_05({net1391[0], net1391[1], net1391[2], net1391[3],
     net1391[4], net1391[5], net1391[6], net1391[7]}),
     .sp12_h_l_08({net1307[0], net1307[1], net1307[2], net1307[3],
     net1307[4], net1307[5], net1307[6], net1307[7], net1307[8],
     net1307[9], net1307[10], net1307[11], net1307[12], net1307[13],
     net1307[14], net1307[15], net1307[16], net1307[17], net1307[18],
     net1307[19], net1307[20], net1307[21], net1307[22], net1307[23]}),
     .sp12_h_l_07({net1306[0], net1306[1], net1306[2], net1306[3],
     net1306[4], net1306[5], net1306[6], net1306[7], net1306[8],
     net1306[9], net1306[10], net1306[11], net1306[12], net1306[13],
     net1306[14], net1306[15], net1306[16], net1306[17], net1306[18],
     net1306[19], net1306[20], net1306[21], net1306[22], net1306[23]}),
     .sp12_h_l_06({net1305[0], net1305[1], net1305[2], net1305[3],
     net1305[4], net1305[5], net1305[6], net1305[7], net1305[8],
     net1305[9], net1305[10], net1305[11], net1305[12], net1305[13],
     net1305[14], net1305[15], net1305[16], net1305[17], net1305[18],
     net1305[19], net1305[20], net1305[21], net1305[22], net1305[23]}),
     .sp12_h_r_05({net1114[0], net1114[1], net1114[2], net1114[3],
     net1114[4], net1114[5], net1114[6], net1114[7], net1114[8],
     net1114[9], net1114[10], net1114[11], net1114[12], net1114[13],
     net1114[14], net1114[15], net1114[16], net1114[17], net1114[18],
     net1114[19], net1114[20], net1114[21], net1114[22], net1114[23]}),
     .sp12_h_r_06({net1115[0], net1115[1], net1115[2], net1115[3],
     net1115[4], net1115[5], net1115[6], net1115[7], net1115[8],
     net1115[9], net1115[10], net1115[11], net1115[12], net1115[13],
     net1115[14], net1115[15], net1115[16], net1115[17], net1115[18],
     net1115[19], net1115[20], net1115[21], net1115[22], net1115[23]}),
     .sp12_h_r_07({net1116[0], net1116[1], net1116[2], net1116[3],
     net1116[4], net1116[5], net1116[6], net1116[7], net1116[8],
     net1116[9], net1116[10], net1116[11], net1116[12], net1116[13],
     net1116[14], net1116[15], net1116[16], net1116[17], net1116[18],
     net1116[19], net1116[20], net1116[21], net1116[22], net1116[23]}),
     .sp12_h_r_08({net1117[0], net1117[1], net1117[2], net1117[3],
     net1117[4], net1117[5], net1117[6], net1117[7], net1117[8],
     net1117[9], net1117[10], net1117[11], net1117[12], net1117[13],
     net1117[14], net1117[15], net1117[16], net1117[17], net1117[18],
     net1117[19], net1117[20], net1117[21], net1117[22], net1117[23]}),
     .sp12_h_l_05({net1304[0], net1304[1], net1304[2], net1304[3],
     net1304[4], net1304[5], net1304[6], net1304[7], net1304[8],
     net1304[9], net1304[10], net1304[11], net1304[12], net1304[13],
     net1304[14], net1304[15], net1304[16], net1304[17], net1304[18],
     net1304[19], net1304[20], net1304[21], net1304[22], net1304[23]}),
     .sp4_r_v_b_05({net1119[0], net1119[1], net1119[2], net1119[3],
     net1119[4], net1119[5], net1119[6], net1119[7], net1119[8],
     net1119[9], net1119[10], net1119[11], net1119[12], net1119[13],
     net1119[14], net1119[15], net1119[16], net1119[17], net1119[18],
     net1119[19], net1119[20], net1119[21], net1119[22], net1119[23],
     net1119[24], net1119[25], net1119[26], net1119[27], net1119[28],
     net1119[29], net1119[30], net1119[31], net1119[32], net1119[33],
     net1119[34], net1119[35], net1119[36], net1119[37], net1119[38],
     net1119[39], net1119[40], net1119[41], net1119[42], net1119[43],
     net1119[44], net1119[45], net1119[46], net1119[47]}),
     .sp4_r_v_b_06({net1120[0], net1120[1], net1120[2], net1120[3],
     net1120[4], net1120[5], net1120[6], net1120[7], net1120[8],
     net1120[9], net1120[10], net1120[11], net1120[12], net1120[13],
     net1120[14], net1120[15], net1120[16], net1120[17], net1120[18],
     net1120[19], net1120[20], net1120[21], net1120[22], net1120[23],
     net1120[24], net1120[25], net1120[26], net1120[27], net1120[28],
     net1120[29], net1120[30], net1120[31], net1120[32], net1120[33],
     net1120[34], net1120[35], net1120[36], net1120[37], net1120[38],
     net1120[39], net1120[40], net1120[41], net1120[42], net1120[43],
     net1120[44], net1120[45], net1120[46], net1120[47]}),
     .sp4_r_v_b_07({net1121[0], net1121[1], net1121[2], net1121[3],
     net1121[4], net1121[5], net1121[6], net1121[7], net1121[8],
     net1121[9], net1121[10], net1121[11], net1121[12], net1121[13],
     net1121[14], net1121[15], net1121[16], net1121[17], net1121[18],
     net1121[19], net1121[20], net1121[21], net1121[22], net1121[23],
     net1121[24], net1121[25], net1121[26], net1121[27], net1121[28],
     net1121[29], net1121[30], net1121[31], net1121[32], net1121[33],
     net1121[34], net1121[35], net1121[36], net1121[37], net1121[38],
     net1121[39], net1121[40], net1121[41], net1121[42], net1121[43],
     net1121[44], net1121[45], net1121[46], net1121[47]}),
     .sp4_r_v_b_08({net1122[0], net1122[1], net1122[2], net1122[3],
     net1122[4], net1122[5], net1122[6], net1122[7], net1122[8],
     net1122[9], net1122[10], net1122[11], net1122[12], net1122[13],
     net1122[14], net1122[15], net1122[16], net1122[17], net1122[18],
     net1122[19], net1122[20], net1122[21], net1122[22], net1122[23],
     net1122[24], net1122[25], net1122[26], net1122[27], net1122[28],
     net1122[29], net1122[30], net1122[31], net1122[32], net1122[33],
     net1122[34], net1122[35], net1122[36], net1122[37], net1122[38],
     net1122[39], net1122[40], net1122[41], net1122[42], net1122[43],
     net1122[44], net1122[45], net1122[46], net1122[47]}),
     .sp4_v_b_08({net1312[0], net1312[1], net1312[2], net1312[3],
     net1312[4], net1312[5], net1312[6], net1312[7], net1312[8],
     net1312[9], net1312[10], net1312[11], net1312[12], net1312[13],
     net1312[14], net1312[15], net1312[16], net1312[17], net1312[18],
     net1312[19], net1312[20], net1312[21], net1312[22], net1312[23],
     net1312[24], net1312[25], net1312[26], net1312[27], net1312[28],
     net1312[29], net1312[30], net1312[31], net1312[32], net1312[33],
     net1312[34], net1312[35], net1312[36], net1312[37], net1312[38],
     net1312[39], net1312[40], net1312[41], net1312[42], net1312[43],
     net1312[44], net1312[45], net1312[46], net1312[47]}),
     .sp4_v_b_07({net1311[0], net1311[1], net1311[2], net1311[3],
     net1311[4], net1311[5], net1311[6], net1311[7], net1311[8],
     net1311[9], net1311[10], net1311[11], net1311[12], net1311[13],
     net1311[14], net1311[15], net1311[16], net1311[17], net1311[18],
     net1311[19], net1311[20], net1311[21], net1311[22], net1311[23],
     net1311[24], net1311[25], net1311[26], net1311[27], net1311[28],
     net1311[29], net1311[30], net1311[31], net1311[32], net1311[33],
     net1311[34], net1311[35], net1311[36], net1311[37], net1311[38],
     net1311[39], net1311[40], net1311[41], net1311[42], net1311[43],
     net1311[44], net1311[45], net1311[46], net1311[47]}),
     .sp4_v_b_06({net1310[0], net1310[1], net1310[2], net1310[3],
     net1310[4], net1310[5], net1310[6], net1310[7], net1310[8],
     net1310[9], net1310[10], net1310[11], net1310[12], net1310[13],
     net1310[14], net1310[15], net1310[16], net1310[17], net1310[18],
     net1310[19], net1310[20], net1310[21], net1310[22], net1310[23],
     net1310[24], net1310[25], net1310[26], net1310[27], net1310[28],
     net1310[29], net1310[30], net1310[31], net1310[32], net1310[33],
     net1310[34], net1310[35], net1310[36], net1310[37], net1310[38],
     net1310[39], net1310[40], net1310[41], net1310[42], net1310[43],
     net1310[44], net1310[45], net1310[46], net1310[47]}),
     .sp4_v_b_05({net1309[0], net1309[1], net1309[2], net1309[3],
     net1309[4], net1309[5], net1309[6], net1309[7], net1309[8],
     net1309[9], net1309[10], net1309[11], net1309[12], net1309[13],
     net1309[14], net1309[15], net1309[16], net1309[17], net1309[18],
     net1309[19], net1309[20], net1309[21], net1309[22], net1309[23],
     net1309[24], net1309[25], net1309[26], net1309[27], net1309[28],
     net1309[29], net1309[30], net1309[31], net1309[32], net1309[33],
     net1309[34], net1309[35], net1309[36], net1309[37], net1309[38],
     net1309[39], net1309[40], net1309[41], net1309[42], net1309[43],
     net1309[44], net1309[45], net1309[46], net1309[47]}),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .wl(wl_r[143:16]), .sp12_v_t_08(sp12_v_t_09_08[23:0]),
     .tnr_op_08(tnr_op_09_08[7:0]), .top_op_08(top_op_09_08[7:0]),
     .tnl_op_08(tnl_op_09_08[7:0]), .sp4_v_t_08(sp4_v_t_09_08[47:0]),
     .lc_bot(tgnd_br_q), .op_vic(op_vic_09_08),
     .sp12_v_b_01({net911[0], net911[1], net911[2], net911[3],
     net911[4], net911[5], net911[6], net911[7], net911[8], net911[9],
     net911[10], net911[11], net911[12], net911[13], net911[14],
     net911[15], net911[16], net911[17], net911[18], net911[19],
     net911[20], net911[21], net911[22], net911[23]}));
lt_1x8_bot_ice1f I_lt_col_b11 ( .glb_netwk_bot({net935[0], net935[1],
     net935[2], net935[3], net935[4], net935[5], net935[6],
     net935[7]}), .rgt_op_03({net1140[0], net1140[1], net1140[2],
     net1140[3], net1140[4], net1140[5], net1140[6], net1140[7]}),
     .slf_op_02({net1533[0], net1533[1], net1533[2], net1533[3],
     net1533[4], net1533[5], net1533[6], net1533[7]}),
     .rgt_op_02({net1142[0], net1142[1], net1142[2], net1142[3],
     net1142[4], net1142[5], net1142[6], net1142[7]}),
     .rgt_op_01({net913[0], net913[1], net913[2], net913[3], net913[4],
     net913[5], net913[6], net913[7]}), .purst(purst), .prog(prog),
     .lft_op_04({net1055[0], net1055[1], net1055[2], net1055[3],
     net1055[4], net1055[5], net1055[6], net1055[7]}),
     .lft_op_03({net1045[0], net1045[1], net1045[2], net1045[3],
     net1045[4], net1045[5], net1045[6], net1045[7]}),
     .lft_op_02({net1047[0], net1047[1], net1047[2], net1047[3],
     net1047[4], net1047[5], net1047[6], net1047[7]}),
     .lft_op_01({net784[0], net784[1], net784[2], net784[3], net784[4],
     net784[5], net784[6], net784[7]}), .rgt_op_04({net1150[0],
     net1150[1], net1150[2], net1150[3], net1150[4], net1150[5],
     net1150[6], net1150[7]}), .carry_in(tgnd_br_q),
     .bnl_op_01({slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0], slf_op_10_00[3], slf_op_10_00[2],
     slf_op_10_00[1], slf_op_10_00[0]}), .slf_op_04({net1531[0],
     net1531[1], net1531[2], net1531[3], net1531[4], net1531[5],
     net1531[6], net1531[7]}), .slf_op_03({net1532[0], net1532[1],
     net1532[2], net1532[3], net1532[4], net1532[5], net1532[6],
     net1532[7]}), .slf_op_01({net782[0], net782[1], net782[2],
     net782[3], net782[4], net782[5], net782[6], net782[7]}),
     .sp4_h_l_04({net1552[0], net1552[1], net1552[2], net1552[3],
     net1552[4], net1552[5], net1552[6], net1552[7], net1552[8],
     net1552[9], net1552[10], net1552[11], net1552[12], net1552[13],
     net1552[14], net1552[15], net1552[16], net1552[17], net1552[18],
     net1552[19], net1552[20], net1552[21], net1552[22], net1552[23],
     net1552[24], net1552[25], net1552[26], net1552[27], net1552[28],
     net1552[29], net1552[30], net1552[31], net1552[32], net1552[33],
     net1552[34], net1552[35], net1552[36], net1552[37], net1552[38],
     net1552[39], net1552[40], net1552[41], net1552[42], net1552[43],
     net1552[44], net1552[45], net1552[46], net1552[47]}),
     .carry_out(carry_out_11_08), .vdd_cntl(vdd_cntl_r[143:16]),
     .sp12_h_r_04({net1159[0], net1159[1], net1159[2], net1159[3],
     net1159[4], net1159[5], net1159[6], net1159[7], net1159[8],
     net1159[9], net1159[10], net1159[11], net1159[12], net1159[13],
     net1159[14], net1159[15], net1159[16], net1159[17], net1159[18],
     net1159[19], net1159[20], net1159[21], net1159[22], net1159[23]}),
     .sp12_h_r_03({net1160[0], net1160[1], net1160[2], net1160[3],
     net1160[4], net1160[5], net1160[6], net1160[7], net1160[8],
     net1160[9], net1160[10], net1160[11], net1160[12], net1160[13],
     net1160[14], net1160[15], net1160[16], net1160[17], net1160[18],
     net1160[19], net1160[20], net1160[21], net1160[22], net1160[23]}),
     .sp12_h_r_02({net1161[0], net1161[1], net1161[2], net1161[3],
     net1161[4], net1161[5], net1161[6], net1161[7], net1161[8],
     net1161[9], net1161[10], net1161[11], net1161[12], net1161[13],
     net1161[14], net1161[15], net1161[16], net1161[17], net1161[18],
     net1161[19], net1161[20], net1161[21], net1161[22], net1161[23]}),
     .sp12_h_r_01({net1162[0], net1162[1], net1162[2], net1162[3],
     net1162[4], net1162[5], net1162[6], net1162[7], net1162[8],
     net1162[9], net1162[10], net1162[11], net1162[12], net1162[13],
     net1162[14], net1162[15], net1162[16], net1162[17], net1162[18],
     net1162[19], net1162[20], net1162[21], net1162[22], net1162[23]}),
     .glb_netwk_col(clk_tree_drv_br[7:0]), .sp4_v_b_01({net896[0],
     net896[1], net896[2], net896[3], net896[4], net896[5], net896[6],
     net896[7], net896[8], net896[9], net896[10], net896[11],
     net896[12], net896[13], net896[14], net896[15], net896[16],
     net896[17], net896[18], net896[19], net896[20], net896[21],
     net896[22], net896[23], net896[24], net896[25], net896[26],
     net896[27], net896[28], net896[29], net896[30], net896[31],
     net896[32], net896[33], net896[34], net896[35], net896[36],
     net896[37], net896[38], net896[39], net896[40], net896[41],
     net896[42], net896[43], net896[44], net896[45], net896[46],
     net896[47]}), .sp4_r_v_b_04({net1165[0], net1165[1], net1165[2],
     net1165[3], net1165[4], net1165[5], net1165[6], net1165[7],
     net1165[8], net1165[9], net1165[10], net1165[11], net1165[12],
     net1165[13], net1165[14], net1165[15], net1165[16], net1165[17],
     net1165[18], net1165[19], net1165[20], net1165[21], net1165[22],
     net1165[23], net1165[24], net1165[25], net1165[26], net1165[27],
     net1165[28], net1165[29], net1165[30], net1165[31], net1165[32],
     net1165[33], net1165[34], net1165[35], net1165[36], net1165[37],
     net1165[38], net1165[39], net1165[40], net1165[41], net1165[42],
     net1165[43], net1165[44], net1165[45], net1165[46], net1165[47]}),
     .sp4_r_v_b_03({net1166[0], net1166[1], net1166[2], net1166[3],
     net1166[4], net1166[5], net1166[6], net1166[7], net1166[8],
     net1166[9], net1166[10], net1166[11], net1166[12], net1166[13],
     net1166[14], net1166[15], net1166[16], net1166[17], net1166[18],
     net1166[19], net1166[20], net1166[21], net1166[22], net1166[23],
     net1166[24], net1166[25], net1166[26], net1166[27], net1166[28],
     net1166[29], net1166[30], net1166[31], net1166[32], net1166[33],
     net1166[34], net1166[35], net1166[36], net1166[37], net1166[38],
     net1166[39], net1166[40], net1166[41], net1166[42], net1166[43],
     net1166[44], net1166[45], net1166[46], net1166[47]}),
     .sp4_r_v_b_02({net1167[0], net1167[1], net1167[2], net1167[3],
     net1167[4], net1167[5], net1167[6], net1167[7], net1167[8],
     net1167[9], net1167[10], net1167[11], net1167[12], net1167[13],
     net1167[14], net1167[15], net1167[16], net1167[17], net1167[18],
     net1167[19], net1167[20], net1167[21], net1167[22], net1167[23],
     net1167[24], net1167[25], net1167[26], net1167[27], net1167[28],
     net1167[29], net1167[30], net1167[31], net1167[32], net1167[33],
     net1167[34], net1167[35], net1167[36], net1167[37], net1167[38],
     net1167[39], net1167[40], net1167[41], net1167[42], net1167[43],
     net1167[44], net1167[45], net1167[46], net1167[47]}),
     .sp4_r_v_b_01({net1168[0], net1168[1], net1168[2], net1168[3],
     net1168[4], net1168[5], net1168[6], net1168[7], net1168[8],
     net1168[9], net1168[10], net1168[11], net1168[12], net1168[13],
     net1168[14], net1168[15], net1168[16], net1168[17], net1168[18],
     net1168[19], net1168[20], net1168[21], net1168[22], net1168[23],
     net1168[24], net1168[25], net1168[26], net1168[27], net1168[28],
     net1168[29], net1168[30], net1168[31], net1168[32], net1168[33],
     net1168[34], net1168[35], net1168[36], net1168[37], net1168[38],
     net1168[39], net1168[40], net1168[41], net1168[42], net1168[43],
     net1168[44], net1168[45], net1168[46], net1168[47]}),
     .sp4_h_r_04({net1169[0], net1169[1], net1169[2], net1169[3],
     net1169[4], net1169[5], net1169[6], net1169[7], net1169[8],
     net1169[9], net1169[10], net1169[11], net1169[12], net1169[13],
     net1169[14], net1169[15], net1169[16], net1169[17], net1169[18],
     net1169[19], net1169[20], net1169[21], net1169[22], net1169[23],
     net1169[24], net1169[25], net1169[26], net1169[27], net1169[28],
     net1169[29], net1169[30], net1169[31], net1169[32], net1169[33],
     net1169[34], net1169[35], net1169[36], net1169[37], net1169[38],
     net1169[39], net1169[40], net1169[41], net1169[42], net1169[43],
     net1169[44], net1169[45], net1169[46], net1169[47]}),
     .sp4_h_r_03({net1170[0], net1170[1], net1170[2], net1170[3],
     net1170[4], net1170[5], net1170[6], net1170[7], net1170[8],
     net1170[9], net1170[10], net1170[11], net1170[12], net1170[13],
     net1170[14], net1170[15], net1170[16], net1170[17], net1170[18],
     net1170[19], net1170[20], net1170[21], net1170[22], net1170[23],
     net1170[24], net1170[25], net1170[26], net1170[27], net1170[28],
     net1170[29], net1170[30], net1170[31], net1170[32], net1170[33],
     net1170[34], net1170[35], net1170[36], net1170[37], net1170[38],
     net1170[39], net1170[40], net1170[41], net1170[42], net1170[43],
     net1170[44], net1170[45], net1170[46], net1170[47]}),
     .sp4_h_r_02({net1171[0], net1171[1], net1171[2], net1171[3],
     net1171[4], net1171[5], net1171[6], net1171[7], net1171[8],
     net1171[9], net1171[10], net1171[11], net1171[12], net1171[13],
     net1171[14], net1171[15], net1171[16], net1171[17], net1171[18],
     net1171[19], net1171[20], net1171[21], net1171[22], net1171[23],
     net1171[24], net1171[25], net1171[26], net1171[27], net1171[28],
     net1171[29], net1171[30], net1171[31], net1171[32], net1171[33],
     net1171[34], net1171[35], net1171[36], net1171[37], net1171[38],
     net1171[39], net1171[40], net1171[41], net1171[42], net1171[43],
     net1171[44], net1171[45], net1171[46], net1171[47]}),
     .sp4_h_r_01({net1172[0], net1172[1], net1172[2], net1172[3],
     net1172[4], net1172[5], net1172[6], net1172[7], net1172[8],
     net1172[9], net1172[10], net1172[11], net1172[12], net1172[13],
     net1172[14], net1172[15], net1172[16], net1172[17], net1172[18],
     net1172[19], net1172[20], net1172[21], net1172[22], net1172[23],
     net1172[24], net1172[25], net1172[26], net1172[27], net1172[28],
     net1172[29], net1172[30], net1172[31], net1172[32], net1172[33],
     net1172[34], net1172[35], net1172[36], net1172[37], net1172[38],
     net1172[39], net1172[40], net1172[41], net1172[42], net1172[43],
     net1172[44], net1172[45], net1172[46], net1172[47]}),
     .sp4_h_l_03({net1551[0], net1551[1], net1551[2], net1551[3],
     net1551[4], net1551[5], net1551[6], net1551[7], net1551[8],
     net1551[9], net1551[10], net1551[11], net1551[12], net1551[13],
     net1551[14], net1551[15], net1551[16], net1551[17], net1551[18],
     net1551[19], net1551[20], net1551[21], net1551[22], net1551[23],
     net1551[24], net1551[25], net1551[26], net1551[27], net1551[28],
     net1551[29], net1551[30], net1551[31], net1551[32], net1551[33],
     net1551[34], net1551[35], net1551[36], net1551[37], net1551[38],
     net1551[39], net1551[40], net1551[41], net1551[42], net1551[43],
     net1551[44], net1551[45], net1551[46], net1551[47]}),
     .sp4_h_l_02({net1550[0], net1550[1], net1550[2], net1550[3],
     net1550[4], net1550[5], net1550[6], net1550[7], net1550[8],
     net1550[9], net1550[10], net1550[11], net1550[12], net1550[13],
     net1550[14], net1550[15], net1550[16], net1550[17], net1550[18],
     net1550[19], net1550[20], net1550[21], net1550[22], net1550[23],
     net1550[24], net1550[25], net1550[26], net1550[27], net1550[28],
     net1550[29], net1550[30], net1550[31], net1550[32], net1550[33],
     net1550[34], net1550[35], net1550[36], net1550[37], net1550[38],
     net1550[39], net1550[40], net1550[41], net1550[42], net1550[43],
     net1550[44], net1550[45], net1550[46], net1550[47]}),
     .sp4_h_l_01({net1506[0], net1506[1], net1506[2], net1506[3],
     net1506[4], net1506[5], net1506[6], net1506[7], net1506[8],
     net1506[9], net1506[10], net1506[11], net1506[12], net1506[13],
     net1506[14], net1506[15], net1506[16], net1506[17], net1506[18],
     net1506[19], net1506[20], net1506[21], net1506[22], net1506[23],
     net1506[24], net1506[25], net1506[26], net1506[27], net1506[28],
     net1506[29], net1506[30], net1506[31], net1506[32], net1506[33],
     net1506[34], net1506[35], net1506[36], net1506[37], net1506[38],
     net1506[39], net1506[40], net1506[41], net1506[42], net1506[43],
     net1506[44], net1506[45], net1506[46], net1506[47]}),
     .bl(bl[257:204]), .bot_op_01({slf_op_11_00[3], slf_op_11_00[2],
     slf_op_11_00[1], slf_op_11_00[0], slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0]}),
     .sp12_h_l_01({net1500[0], net1500[1], net1500[2], net1500[3],
     net1500[4], net1500[5], net1500[6], net1500[7], net1500[8],
     net1500[9], net1500[10], net1500[11], net1500[12], net1500[13],
     net1500[14], net1500[15], net1500[16], net1500[17], net1500[18],
     net1500[19], net1500[20], net1500[21], net1500[22], net1500[23]}),
     .sp12_h_l_02({net1508[0], net1508[1], net1508[2], net1508[3],
     net1508[4], net1508[5], net1508[6], net1508[7], net1508[8],
     net1508[9], net1508[10], net1508[11], net1508[12], net1508[13],
     net1508[14], net1508[15], net1508[16], net1508[17], net1508[18],
     net1508[19], net1508[20], net1508[21], net1508[22], net1508[23]}),
     .sp12_h_l_03({net1464[0], net1464[1], net1464[2], net1464[3],
     net1464[4], net1464[5], net1464[6], net1464[7], net1464[8],
     net1464[9], net1464[10], net1464[11], net1464[12], net1464[13],
     net1464[14], net1464[15], net1464[16], net1464[17], net1464[18],
     net1464[19], net1464[20], net1464[21], net1464[22], net1464[23]}),
     .sp12_h_l_04({net1509[0], net1509[1], net1509[2], net1509[3],
     net1509[4], net1509[5], net1509[6], net1509[7], net1509[8],
     net1509[9], net1509[10], net1509[11], net1509[12], net1509[13],
     net1509[14], net1509[15], net1509[16], net1509[17], net1509[18],
     net1509[19], net1509[20], net1509[21], net1509[22], net1509[23]}),
     .sp4_v_b_04({net1488[0], net1488[1], net1488[2], net1488[3],
     net1488[4], net1488[5], net1488[6], net1488[7], net1488[8],
     net1488[9], net1488[10], net1488[11], net1488[12], net1488[13],
     net1488[14], net1488[15], net1488[16], net1488[17], net1488[18],
     net1488[19], net1488[20], net1488[21], net1488[22], net1488[23],
     net1488[24], net1488[25], net1488[26], net1488[27], net1488[28],
     net1488[29], net1488[30], net1488[31], net1488[32], net1488[33],
     net1488[34], net1488[35], net1488[36], net1488[37], net1488[38],
     net1488[39], net1488[40], net1488[41], net1488[42], net1488[43],
     net1488[44], net1488[45], net1488[46], net1488[47]}),
     .sp4_v_b_03({net1484[0], net1484[1], net1484[2], net1484[3],
     net1484[4], net1484[5], net1484[6], net1484[7], net1484[8],
     net1484[9], net1484[10], net1484[11], net1484[12], net1484[13],
     net1484[14], net1484[15], net1484[16], net1484[17], net1484[18],
     net1484[19], net1484[20], net1484[21], net1484[22], net1484[23],
     net1484[24], net1484[25], net1484[26], net1484[27], net1484[28],
     net1484[29], net1484[30], net1484[31], net1484[32], net1484[33],
     net1484[34], net1484[35], net1484[36], net1484[37], net1484[38],
     net1484[39], net1484[40], net1484[41], net1484[42], net1484[43],
     net1484[44], net1484[45], net1484[46], net1484[47]}),
     .sp4_v_b_02({net1495[0], net1495[1], net1495[2], net1495[3],
     net1495[4], net1495[5], net1495[6], net1495[7], net1495[8],
     net1495[9], net1495[10], net1495[11], net1495[12], net1495[13],
     net1495[14], net1495[15], net1495[16], net1495[17], net1495[18],
     net1495[19], net1495[20], net1495[21], net1495[22], net1495[23],
     net1495[24], net1495[25], net1495[26], net1495[27], net1495[28],
     net1495[29], net1495[30], net1495[31], net1495[32], net1495[33],
     net1495[34], net1495[35], net1495[36], net1495[37], net1495[38],
     net1495[39], net1495[40], net1495[41], net1495[42], net1495[43],
     net1495[44], net1495[45], net1495[46], net1495[47]}),
     .bnr_op_01({slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0], slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0]}), .sp4_h_l_05({net1553[0],
     net1553[1], net1553[2], net1553[3], net1553[4], net1553[5],
     net1553[6], net1553[7], net1553[8], net1553[9], net1553[10],
     net1553[11], net1553[12], net1553[13], net1553[14], net1553[15],
     net1553[16], net1553[17], net1553[18], net1553[19], net1553[20],
     net1553[21], net1553[22], net1553[23], net1553[24], net1553[25],
     net1553[26], net1553[27], net1553[28], net1553[29], net1553[30],
     net1553[31], net1553[32], net1553[33], net1553[34], net1553[35],
     net1553[36], net1553[37], net1553[38], net1553[39], net1553[40],
     net1553[41], net1553[42], net1553[43], net1553[44], net1553[45],
     net1553[46], net1553[47]}), .sp4_h_l_06({net1554[0], net1554[1],
     net1554[2], net1554[3], net1554[4], net1554[5], net1554[6],
     net1554[7], net1554[8], net1554[9], net1554[10], net1554[11],
     net1554[12], net1554[13], net1554[14], net1554[15], net1554[16],
     net1554[17], net1554[18], net1554[19], net1554[20], net1554[21],
     net1554[22], net1554[23], net1554[24], net1554[25], net1554[26],
     net1554[27], net1554[28], net1554[29], net1554[30], net1554[31],
     net1554[32], net1554[33], net1554[34], net1554[35], net1554[36],
     net1554[37], net1554[38], net1554[39], net1554[40], net1554[41],
     net1554[42], net1554[43], net1554[44], net1554[45], net1554[46],
     net1554[47]}), .sp4_h_l_07({net1555[0], net1555[1], net1555[2],
     net1555[3], net1555[4], net1555[5], net1555[6], net1555[7],
     net1555[8], net1555[9], net1555[10], net1555[11], net1555[12],
     net1555[13], net1555[14], net1555[15], net1555[16], net1555[17],
     net1555[18], net1555[19], net1555[20], net1555[21], net1555[22],
     net1555[23], net1555[24], net1555[25], net1555[26], net1555[27],
     net1555[28], net1555[29], net1555[30], net1555[31], net1555[32],
     net1555[33], net1555[34], net1555[35], net1555[36], net1555[37],
     net1555[38], net1555[39], net1555[40], net1555[41], net1555[42],
     net1555[43], net1555[44], net1555[45], net1555[46], net1555[47]}),
     .sp4_h_l_08({net1491[0], net1491[1], net1491[2], net1491[3],
     net1491[4], net1491[5], net1491[6], net1491[7], net1491[8],
     net1491[9], net1491[10], net1491[11], net1491[12], net1491[13],
     net1491[14], net1491[15], net1491[16], net1491[17], net1491[18],
     net1491[19], net1491[20], net1491[21], net1491[22], net1491[23],
     net1491[24], net1491[25], net1491[26], net1491[27], net1491[28],
     net1491[29], net1491[30], net1491[31], net1491[32], net1491[33],
     net1491[34], net1491[35], net1491[36], net1491[37], net1491[38],
     net1491[39], net1491[40], net1491[41], net1491[42], net1491[43],
     net1491[44], net1491[45], net1491[46], net1491[47]}),
     .sp4_h_r_08({net1190[0], net1190[1], net1190[2], net1190[3],
     net1190[4], net1190[5], net1190[6], net1190[7], net1190[8],
     net1190[9], net1190[10], net1190[11], net1190[12], net1190[13],
     net1190[14], net1190[15], net1190[16], net1190[17], net1190[18],
     net1190[19], net1190[20], net1190[21], net1190[22], net1190[23],
     net1190[24], net1190[25], net1190[26], net1190[27], net1190[28],
     net1190[29], net1190[30], net1190[31], net1190[32], net1190[33],
     net1190[34], net1190[35], net1190[36], net1190[37], net1190[38],
     net1190[39], net1190[40], net1190[41], net1190[42], net1190[43],
     net1190[44], net1190[45], net1190[46], net1190[47]}),
     .sp4_h_r_07({net1191[0], net1191[1], net1191[2], net1191[3],
     net1191[4], net1191[5], net1191[6], net1191[7], net1191[8],
     net1191[9], net1191[10], net1191[11], net1191[12], net1191[13],
     net1191[14], net1191[15], net1191[16], net1191[17], net1191[18],
     net1191[19], net1191[20], net1191[21], net1191[22], net1191[23],
     net1191[24], net1191[25], net1191[26], net1191[27], net1191[28],
     net1191[29], net1191[30], net1191[31], net1191[32], net1191[33],
     net1191[34], net1191[35], net1191[36], net1191[37], net1191[38],
     net1191[39], net1191[40], net1191[41], net1191[42], net1191[43],
     net1191[44], net1191[45], net1191[46], net1191[47]}),
     .sp4_h_r_06({net1192[0], net1192[1], net1192[2], net1192[3],
     net1192[4], net1192[5], net1192[6], net1192[7], net1192[8],
     net1192[9], net1192[10], net1192[11], net1192[12], net1192[13],
     net1192[14], net1192[15], net1192[16], net1192[17], net1192[18],
     net1192[19], net1192[20], net1192[21], net1192[22], net1192[23],
     net1192[24], net1192[25], net1192[26], net1192[27], net1192[28],
     net1192[29], net1192[30], net1192[31], net1192[32], net1192[33],
     net1192[34], net1192[35], net1192[36], net1192[37], net1192[38],
     net1192[39], net1192[40], net1192[41], net1192[42], net1192[43],
     net1192[44], net1192[45], net1192[46], net1192[47]}),
     .sp4_h_r_05({net1193[0], net1193[1], net1193[2], net1193[3],
     net1193[4], net1193[5], net1193[6], net1193[7], net1193[8],
     net1193[9], net1193[10], net1193[11], net1193[12], net1193[13],
     net1193[14], net1193[15], net1193[16], net1193[17], net1193[18],
     net1193[19], net1193[20], net1193[21], net1193[22], net1193[23],
     net1193[24], net1193[25], net1193[26], net1193[27], net1193[28],
     net1193[29], net1193[30], net1193[31], net1193[32], net1193[33],
     net1193[34], net1193[35], net1193[36], net1193[37], net1193[38],
     net1193[39], net1193[40], net1193[41], net1193[42], net1193[43],
     net1193[44], net1193[45], net1193[46], net1193[47]}),
     .slf_op_05({net1530[0], net1530[1], net1530[2], net1530[3],
     net1530[4], net1530[5], net1530[6], net1530[7]}),
     .slf_op_06({net1529[0], net1529[1], net1529[2], net1529[3],
     net1529[4], net1529[5], net1529[6], net1529[7]}),
     .slf_op_07({net1528[0], net1528[1], net1528[2], net1528[3],
     net1528[4], net1528[5], net1528[6], net1528[7]}),
     .slf_op_08(slf_op_11_08[7:0]), .rgt_op_08(slf_op_12_08[7:0]),
     .rgt_op_07({net1199[0], net1199[1], net1199[2], net1199[3],
     net1199[4], net1199[5], net1199[6], net1199[7]}),
     .rgt_op_06({net1200[0], net1200[1], net1200[2], net1200[3],
     net1200[4], net1200[5], net1200[6], net1200[7]}),
     .rgt_op_05({net1201[0], net1201[1], net1201[2], net1201[3],
     net1201[4], net1201[5], net1201[6], net1201[7]}),
     .lft_op_08(slf_op_10_08[7:0]), .lft_op_07({net1104[0], net1104[1],
     net1104[2], net1104[3], net1104[4], net1104[5], net1104[6],
     net1104[7]}), .lft_op_06({net1105[0], net1105[1], net1105[2],
     net1105[3], net1105[4], net1105[5], net1105[6], net1105[7]}),
     .lft_op_05({net1106[0], net1106[1], net1106[2], net1106[3],
     net1106[4], net1106[5], net1106[6], net1106[7]}),
     .sp12_h_l_08({net1481[0], net1481[1], net1481[2], net1481[3],
     net1481[4], net1481[5], net1481[6], net1481[7], net1481[8],
     net1481[9], net1481[10], net1481[11], net1481[12], net1481[13],
     net1481[14], net1481[15], net1481[16], net1481[17], net1481[18],
     net1481[19], net1481[20], net1481[21], net1481[22], net1481[23]}),
     .sp12_h_l_07({net1476[0], net1476[1], net1476[2], net1476[3],
     net1476[4], net1476[5], net1476[6], net1476[7], net1476[8],
     net1476[9], net1476[10], net1476[11], net1476[12], net1476[13],
     net1476[14], net1476[15], net1476[16], net1476[17], net1476[18],
     net1476[19], net1476[20], net1476[21], net1476[22], net1476[23]}),
     .sp12_h_l_06({net1478[0], net1478[1], net1478[2], net1478[3],
     net1478[4], net1478[5], net1478[6], net1478[7], net1478[8],
     net1478[9], net1478[10], net1478[11], net1478[12], net1478[13],
     net1478[14], net1478[15], net1478[16], net1478[17], net1478[18],
     net1478[19], net1478[20], net1478[21], net1478[22], net1478[23]}),
     .sp12_h_r_05({net1209[0], net1209[1], net1209[2], net1209[3],
     net1209[4], net1209[5], net1209[6], net1209[7], net1209[8],
     net1209[9], net1209[10], net1209[11], net1209[12], net1209[13],
     net1209[14], net1209[15], net1209[16], net1209[17], net1209[18],
     net1209[19], net1209[20], net1209[21], net1209[22], net1209[23]}),
     .sp12_h_r_06({net1210[0], net1210[1], net1210[2], net1210[3],
     net1210[4], net1210[5], net1210[6], net1210[7], net1210[8],
     net1210[9], net1210[10], net1210[11], net1210[12], net1210[13],
     net1210[14], net1210[15], net1210[16], net1210[17], net1210[18],
     net1210[19], net1210[20], net1210[21], net1210[22], net1210[23]}),
     .sp12_h_r_07({net1211[0], net1211[1], net1211[2], net1211[3],
     net1211[4], net1211[5], net1211[6], net1211[7], net1211[8],
     net1211[9], net1211[10], net1211[11], net1211[12], net1211[13],
     net1211[14], net1211[15], net1211[16], net1211[17], net1211[18],
     net1211[19], net1211[20], net1211[21], net1211[22], net1211[23]}),
     .sp12_h_r_08({net1212[0], net1212[1], net1212[2], net1212[3],
     net1212[4], net1212[5], net1212[6], net1212[7], net1212[8],
     net1212[9], net1212[10], net1212[11], net1212[12], net1212[13],
     net1212[14], net1212[15], net1212[16], net1212[17], net1212[18],
     net1212[19], net1212[20], net1212[21], net1212[22], net1212[23]}),
     .sp12_h_l_05({net1480[0], net1480[1], net1480[2], net1480[3],
     net1480[4], net1480[5], net1480[6], net1480[7], net1480[8],
     net1480[9], net1480[10], net1480[11], net1480[12], net1480[13],
     net1480[14], net1480[15], net1480[16], net1480[17], net1480[18],
     net1480[19], net1480[20], net1480[21], net1480[22], net1480[23]}),
     .sp4_r_v_b_05({net1214[0], net1214[1], net1214[2], net1214[3],
     net1214[4], net1214[5], net1214[6], net1214[7], net1214[8],
     net1214[9], net1214[10], net1214[11], net1214[12], net1214[13],
     net1214[14], net1214[15], net1214[16], net1214[17], net1214[18],
     net1214[19], net1214[20], net1214[21], net1214[22], net1214[23],
     net1214[24], net1214[25], net1214[26], net1214[27], net1214[28],
     net1214[29], net1214[30], net1214[31], net1214[32], net1214[33],
     net1214[34], net1214[35], net1214[36], net1214[37], net1214[38],
     net1214[39], net1214[40], net1214[41], net1214[42], net1214[43],
     net1214[44], net1214[45], net1214[46], net1214[47]}),
     .sp4_r_v_b_06({net1215[0], net1215[1], net1215[2], net1215[3],
     net1215[4], net1215[5], net1215[6], net1215[7], net1215[8],
     net1215[9], net1215[10], net1215[11], net1215[12], net1215[13],
     net1215[14], net1215[15], net1215[16], net1215[17], net1215[18],
     net1215[19], net1215[20], net1215[21], net1215[22], net1215[23],
     net1215[24], net1215[25], net1215[26], net1215[27], net1215[28],
     net1215[29], net1215[30], net1215[31], net1215[32], net1215[33],
     net1215[34], net1215[35], net1215[36], net1215[37], net1215[38],
     net1215[39], net1215[40], net1215[41], net1215[42], net1215[43],
     net1215[44], net1215[45], net1215[46], net1215[47]}),
     .sp4_r_v_b_07({net1216[0], net1216[1], net1216[2], net1216[3],
     net1216[4], net1216[5], net1216[6], net1216[7], net1216[8],
     net1216[9], net1216[10], net1216[11], net1216[12], net1216[13],
     net1216[14], net1216[15], net1216[16], net1216[17], net1216[18],
     net1216[19], net1216[20], net1216[21], net1216[22], net1216[23],
     net1216[24], net1216[25], net1216[26], net1216[27], net1216[28],
     net1216[29], net1216[30], net1216[31], net1216[32], net1216[33],
     net1216[34], net1216[35], net1216[36], net1216[37], net1216[38],
     net1216[39], net1216[40], net1216[41], net1216[42], net1216[43],
     net1216[44], net1216[45], net1216[46], net1216[47]}),
     .sp4_r_v_b_08({net1217[0], net1217[1], net1217[2], net1217[3],
     net1217[4], net1217[5], net1217[6], net1217[7], net1217[8],
     net1217[9], net1217[10], net1217[11], net1217[12], net1217[13],
     net1217[14], net1217[15], net1217[16], net1217[17], net1217[18],
     net1217[19], net1217[20], net1217[21], net1217[22], net1217[23],
     net1217[24], net1217[25], net1217[26], net1217[27], net1217[28],
     net1217[29], net1217[30], net1217[31], net1217[32], net1217[33],
     net1217[34], net1217[35], net1217[36], net1217[37], net1217[38],
     net1217[39], net1217[40], net1217[41], net1217[42], net1217[43],
     net1217[44], net1217[45], net1217[46], net1217[47]}),
     .sp4_v_b_08({net1523[0], net1523[1], net1523[2], net1523[3],
     net1523[4], net1523[5], net1523[6], net1523[7], net1523[8],
     net1523[9], net1523[10], net1523[11], net1523[12], net1523[13],
     net1523[14], net1523[15], net1523[16], net1523[17], net1523[18],
     net1523[19], net1523[20], net1523[21], net1523[22], net1523[23],
     net1523[24], net1523[25], net1523[26], net1523[27], net1523[28],
     net1523[29], net1523[30], net1523[31], net1523[32], net1523[33],
     net1523[34], net1523[35], net1523[36], net1523[37], net1523[38],
     net1523[39], net1523[40], net1523[41], net1523[42], net1523[43],
     net1523[44], net1523[45], net1523[46], net1523[47]}),
     .sp4_v_b_07({net1524[0], net1524[1], net1524[2], net1524[3],
     net1524[4], net1524[5], net1524[6], net1524[7], net1524[8],
     net1524[9], net1524[10], net1524[11], net1524[12], net1524[13],
     net1524[14], net1524[15], net1524[16], net1524[17], net1524[18],
     net1524[19], net1524[20], net1524[21], net1524[22], net1524[23],
     net1524[24], net1524[25], net1524[26], net1524[27], net1524[28],
     net1524[29], net1524[30], net1524[31], net1524[32], net1524[33],
     net1524[34], net1524[35], net1524[36], net1524[37], net1524[38],
     net1524[39], net1524[40], net1524[41], net1524[42], net1524[43],
     net1524[44], net1524[45], net1524[46], net1524[47]}),
     .sp4_v_b_06({net1525[0], net1525[1], net1525[2], net1525[3],
     net1525[4], net1525[5], net1525[6], net1525[7], net1525[8],
     net1525[9], net1525[10], net1525[11], net1525[12], net1525[13],
     net1525[14], net1525[15], net1525[16], net1525[17], net1525[18],
     net1525[19], net1525[20], net1525[21], net1525[22], net1525[23],
     net1525[24], net1525[25], net1525[26], net1525[27], net1525[28],
     net1525[29], net1525[30], net1525[31], net1525[32], net1525[33],
     net1525[34], net1525[35], net1525[36], net1525[37], net1525[38],
     net1525[39], net1525[40], net1525[41], net1525[42], net1525[43],
     net1525[44], net1525[45], net1525[46], net1525[47]}),
     .sp4_v_b_05({net1492[0], net1492[1], net1492[2], net1492[3],
     net1492[4], net1492[5], net1492[6], net1492[7], net1492[8],
     net1492[9], net1492[10], net1492[11], net1492[12], net1492[13],
     net1492[14], net1492[15], net1492[16], net1492[17], net1492[18],
     net1492[19], net1492[20], net1492[21], net1492[22], net1492[23],
     net1492[24], net1492[25], net1492[26], net1492[27], net1492[28],
     net1492[29], net1492[30], net1492[31], net1492[32], net1492[33],
     net1492[34], net1492[35], net1492[36], net1492[37], net1492[38],
     net1492[39], net1492[40], net1492[41], net1492[42], net1492[43],
     net1492[44], net1492[45], net1492[46], net1492[47]}),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .wl(wl_r[143:16]), .sp12_v_t_08(sp12_v_t_11_08[23:0]),
     .tnr_op_08(tnr_op_11_08[7:0]), .top_op_08(top_op_11_08[7:0]),
     .tnl_op_08(tnl_op_11_08[7:0]), .sp4_v_t_08(sp4_v_t_11_08[47:0]),
     .lc_bot(tgnd_br_q), .op_vic(op_vic_11_08),
     .sp12_v_b_01({net894[0], net894[1], net894[2], net894[3],
     net894[4], net894[5], net894[6], net894[7], net894[8], net894[9],
     net894[10], net894[11], net894[12], net894[13], net894[14],
     net894[15], net894[16], net894[17], net894[18], net894[19],
     net894[20], net894[21], net894[22], net894[23]}));
lt_1x8_bot_ice1f I_lt_col_b08 ( .glb_netwk_bot({net938[0], net938[1],
     net938[2], net938[3], net938[4], net938[5], net938[6],
     net938[7]}), .rgt_op_03({net1235[0], net1235[1], net1235[2],
     net1235[3], net1235[4], net1235[5], net1235[6], net1235[7]}),
     .slf_op_02({net1332[0], net1332[1], net1332[2], net1332[3],
     net1332[4], net1332[5], net1332[6], net1332[7]}),
     .rgt_op_02({net1237[0], net1237[1], net1237[2], net1237[3],
     net1237[4], net1237[5], net1237[6], net1237[7]}),
     .rgt_op_01({net910[0], net910[1], net910[2], net910[3], net910[4],
     net910[5], net910[6], net910[7]}), .purst(purst), .prog(prog),
     .lft_op_04(slf_op_07_04[7:0]), .lft_op_03(slf_op_07_03[7:0]),
     .lft_op_02(slf_op_07_02[7:0]), .lft_op_01(slf_op_07_01[7:0]),
     .rgt_op_04({net1245[0], net1245[1], net1245[2], net1245[3],
     net1245[4], net1245[5], net1245[6], net1245[7]}),
     .carry_in(tgnd_br_q), .bnl_op_01({slf_op_07_00[3],
     slf_op_07_00[2], slf_op_07_00[1], slf_op_07_00[0],
     slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0]}), .slf_op_04({net1340[0], net1340[1], net1340[2],
     net1340[3], net1340[4], net1340[5], net1340[6], net1340[7]}),
     .slf_op_03({net1330[0], net1330[1], net1330[2], net1330[3],
     net1330[4], net1330[5], net1330[6], net1330[7]}),
     .slf_op_01({net793[0], net793[1], net793[2], net793[3], net793[4],
     net793[5], net793[6], net793[7]}), .sp4_h_l_04({net1359[0],
     net1359[1], net1359[2], net1359[3], net1359[4], net1359[5],
     net1359[6], net1359[7], net1359[8], net1359[9], net1359[10],
     net1359[11], net1359[12], net1359[13], net1359[14], net1359[15],
     net1359[16], net1359[17], net1359[18], net1359[19], net1359[20],
     net1359[21], net1359[22], net1359[23], net1359[24], net1359[25],
     net1359[26], net1359[27], net1359[28], net1359[29], net1359[30],
     net1359[31], net1359[32], net1359[33], net1359[34], net1359[35],
     net1359[36], net1359[37], net1359[38], net1359[39], net1359[40],
     net1359[41], net1359[42], net1359[43], net1359[44], net1359[45],
     net1359[46], net1359[47]}), .carry_out(carry_out_08_08),
     .vdd_cntl(vdd_cntl_r[143:16]), .sp12_h_r_04({net1254[0],
     net1254[1], net1254[2], net1254[3], net1254[4], net1254[5],
     net1254[6], net1254[7], net1254[8], net1254[9], net1254[10],
     net1254[11], net1254[12], net1254[13], net1254[14], net1254[15],
     net1254[16], net1254[17], net1254[18], net1254[19], net1254[20],
     net1254[21], net1254[22], net1254[23]}), .sp12_h_r_03({net1255[0],
     net1255[1], net1255[2], net1255[3], net1255[4], net1255[5],
     net1255[6], net1255[7], net1255[8], net1255[9], net1255[10],
     net1255[11], net1255[12], net1255[13], net1255[14], net1255[15],
     net1255[16], net1255[17], net1255[18], net1255[19], net1255[20],
     net1255[21], net1255[22], net1255[23]}), .sp12_h_r_02({net1256[0],
     net1256[1], net1256[2], net1256[3], net1256[4], net1256[5],
     net1256[6], net1256[7], net1256[8], net1256[9], net1256[10],
     net1256[11], net1256[12], net1256[13], net1256[14], net1256[15],
     net1256[16], net1256[17], net1256[18], net1256[19], net1256[20],
     net1256[21], net1256[22], net1256[23]}), .sp12_h_r_01({net1257[0],
     net1257[1], net1257[2], net1257[3], net1257[4], net1257[5],
     net1257[6], net1257[7], net1257[8], net1257[9], net1257[10],
     net1257[11], net1257[12], net1257[13], net1257[14], net1257[15],
     net1257[16], net1257[17], net1257[18], net1257[19], net1257[20],
     net1257[21], net1257[22], net1257[23]}),
     .glb_netwk_col(clk_tree_drv_br[7:0]), .sp4_v_b_01({net889[0],
     net889[1], net889[2], net889[3], net889[4], net889[5], net889[6],
     net889[7], net889[8], net889[9], net889[10], net889[11],
     net889[12], net889[13], net889[14], net889[15], net889[16],
     net889[17], net889[18], net889[19], net889[20], net889[21],
     net889[22], net889[23], net889[24], net889[25], net889[26],
     net889[27], net889[28], net889[29], net889[30], net889[31],
     net889[32], net889[33], net889[34], net889[35], net889[36],
     net889[37], net889[38], net889[39], net889[40], net889[41],
     net889[42], net889[43], net889[44], net889[45], net889[46],
     net889[47]}), .sp4_r_v_b_04({net1260[0], net1260[1], net1260[2],
     net1260[3], net1260[4], net1260[5], net1260[6], net1260[7],
     net1260[8], net1260[9], net1260[10], net1260[11], net1260[12],
     net1260[13], net1260[14], net1260[15], net1260[16], net1260[17],
     net1260[18], net1260[19], net1260[20], net1260[21], net1260[22],
     net1260[23], net1260[24], net1260[25], net1260[26], net1260[27],
     net1260[28], net1260[29], net1260[30], net1260[31], net1260[32],
     net1260[33], net1260[34], net1260[35], net1260[36], net1260[37],
     net1260[38], net1260[39], net1260[40], net1260[41], net1260[42],
     net1260[43], net1260[44], net1260[45], net1260[46], net1260[47]}),
     .sp4_r_v_b_03({net1261[0], net1261[1], net1261[2], net1261[3],
     net1261[4], net1261[5], net1261[6], net1261[7], net1261[8],
     net1261[9], net1261[10], net1261[11], net1261[12], net1261[13],
     net1261[14], net1261[15], net1261[16], net1261[17], net1261[18],
     net1261[19], net1261[20], net1261[21], net1261[22], net1261[23],
     net1261[24], net1261[25], net1261[26], net1261[27], net1261[28],
     net1261[29], net1261[30], net1261[31], net1261[32], net1261[33],
     net1261[34], net1261[35], net1261[36], net1261[37], net1261[38],
     net1261[39], net1261[40], net1261[41], net1261[42], net1261[43],
     net1261[44], net1261[45], net1261[46], net1261[47]}),
     .sp4_r_v_b_02({net1262[0], net1262[1], net1262[2], net1262[3],
     net1262[4], net1262[5], net1262[6], net1262[7], net1262[8],
     net1262[9], net1262[10], net1262[11], net1262[12], net1262[13],
     net1262[14], net1262[15], net1262[16], net1262[17], net1262[18],
     net1262[19], net1262[20], net1262[21], net1262[22], net1262[23],
     net1262[24], net1262[25], net1262[26], net1262[27], net1262[28],
     net1262[29], net1262[30], net1262[31], net1262[32], net1262[33],
     net1262[34], net1262[35], net1262[36], net1262[37], net1262[38],
     net1262[39], net1262[40], net1262[41], net1262[42], net1262[43],
     net1262[44], net1262[45], net1262[46], net1262[47]}),
     .sp4_r_v_b_01({net916[0], net916[1], net916[2], net916[3],
     net916[4], net916[5], net916[6], net916[7], net916[8], net916[9],
     net916[10], net916[11], net916[12], net916[13], net916[14],
     net916[15], net916[16], net916[17], net916[18], net916[19],
     net916[20], net916[21], net916[22], net916[23], net916[24],
     net916[25], net916[26], net916[27], net916[28], net916[29],
     net916[30], net916[31], net916[32], net916[33], net916[34],
     net916[35], net916[36], net916[37], net916[38], net916[39],
     net916[40], net916[41], net916[42], net916[43], net916[44],
     net916[45], net916[46], net916[47]}), .sp4_h_r_04({net1264[0],
     net1264[1], net1264[2], net1264[3], net1264[4], net1264[5],
     net1264[6], net1264[7], net1264[8], net1264[9], net1264[10],
     net1264[11], net1264[12], net1264[13], net1264[14], net1264[15],
     net1264[16], net1264[17], net1264[18], net1264[19], net1264[20],
     net1264[21], net1264[22], net1264[23], net1264[24], net1264[25],
     net1264[26], net1264[27], net1264[28], net1264[29], net1264[30],
     net1264[31], net1264[32], net1264[33], net1264[34], net1264[35],
     net1264[36], net1264[37], net1264[38], net1264[39], net1264[40],
     net1264[41], net1264[42], net1264[43], net1264[44], net1264[45],
     net1264[46], net1264[47]}), .sp4_h_r_03({net1265[0], net1265[1],
     net1265[2], net1265[3], net1265[4], net1265[5], net1265[6],
     net1265[7], net1265[8], net1265[9], net1265[10], net1265[11],
     net1265[12], net1265[13], net1265[14], net1265[15], net1265[16],
     net1265[17], net1265[18], net1265[19], net1265[20], net1265[21],
     net1265[22], net1265[23], net1265[24], net1265[25], net1265[26],
     net1265[27], net1265[28], net1265[29], net1265[30], net1265[31],
     net1265[32], net1265[33], net1265[34], net1265[35], net1265[36],
     net1265[37], net1265[38], net1265[39], net1265[40], net1265[41],
     net1265[42], net1265[43], net1265[44], net1265[45], net1265[46],
     net1265[47]}), .sp4_h_r_02({net1266[0], net1266[1], net1266[2],
     net1266[3], net1266[4], net1266[5], net1266[6], net1266[7],
     net1266[8], net1266[9], net1266[10], net1266[11], net1266[12],
     net1266[13], net1266[14], net1266[15], net1266[16], net1266[17],
     net1266[18], net1266[19], net1266[20], net1266[21], net1266[22],
     net1266[23], net1266[24], net1266[25], net1266[26], net1266[27],
     net1266[28], net1266[29], net1266[30], net1266[31], net1266[32],
     net1266[33], net1266[34], net1266[35], net1266[36], net1266[37],
     net1266[38], net1266[39], net1266[40], net1266[41], net1266[42],
     net1266[43], net1266[44], net1266[45], net1266[46], net1266[47]}),
     .sp4_h_r_01({net1267[0], net1267[1], net1267[2], net1267[3],
     net1267[4], net1267[5], net1267[6], net1267[7], net1267[8],
     net1267[9], net1267[10], net1267[11], net1267[12], net1267[13],
     net1267[14], net1267[15], net1267[16], net1267[17], net1267[18],
     net1267[19], net1267[20], net1267[21], net1267[22], net1267[23],
     net1267[24], net1267[25], net1267[26], net1267[27], net1267[28],
     net1267[29], net1267[30], net1267[31], net1267[32], net1267[33],
     net1267[34], net1267[35], net1267[36], net1267[37], net1267[38],
     net1267[39], net1267[40], net1267[41], net1267[42], net1267[43],
     net1267[44], net1267[45], net1267[46], net1267[47]}),
     .sp4_h_l_03({net1360[0], net1360[1], net1360[2], net1360[3],
     net1360[4], net1360[5], net1360[6], net1360[7], net1360[8],
     net1360[9], net1360[10], net1360[11], net1360[12], net1360[13],
     net1360[14], net1360[15], net1360[16], net1360[17], net1360[18],
     net1360[19], net1360[20], net1360[21], net1360[22], net1360[23],
     net1360[24], net1360[25], net1360[26], net1360[27], net1360[28],
     net1360[29], net1360[30], net1360[31], net1360[32], net1360[33],
     net1360[34], net1360[35], net1360[36], net1360[37], net1360[38],
     net1360[39], net1360[40], net1360[41], net1360[42], net1360[43],
     net1360[44], net1360[45], net1360[46], net1360[47]}),
     .sp4_h_l_02({net1361[0], net1361[1], net1361[2], net1361[3],
     net1361[4], net1361[5], net1361[6], net1361[7], net1361[8],
     net1361[9], net1361[10], net1361[11], net1361[12], net1361[13],
     net1361[14], net1361[15], net1361[16], net1361[17], net1361[18],
     net1361[19], net1361[20], net1361[21], net1361[22], net1361[23],
     net1361[24], net1361[25], net1361[26], net1361[27], net1361[28],
     net1361[29], net1361[30], net1361[31], net1361[32], net1361[33],
     net1361[34], net1361[35], net1361[36], net1361[37], net1361[38],
     net1361[39], net1361[40], net1361[41], net1361[42], net1361[43],
     net1361[44], net1361[45], net1361[46], net1361[47]}),
     .sp4_h_l_01({net1362[0], net1362[1], net1362[2], net1362[3],
     net1362[4], net1362[5], net1362[6], net1362[7], net1362[8],
     net1362[9], net1362[10], net1362[11], net1362[12], net1362[13],
     net1362[14], net1362[15], net1362[16], net1362[17], net1362[18],
     net1362[19], net1362[20], net1362[21], net1362[22], net1362[23],
     net1362[24], net1362[25], net1362[26], net1362[27], net1362[28],
     net1362[29], net1362[30], net1362[31], net1362[32], net1362[33],
     net1362[34], net1362[35], net1362[36], net1362[37], net1362[38],
     net1362[39], net1362[40], net1362[41], net1362[42], net1362[43],
     net1362[44], net1362[45], net1362[46], net1362[47]}),
     .bl(bl[107:54]), .bot_op_01({slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0], slf_op_08_00[3],
     slf_op_08_00[2], slf_op_08_00[1], slf_op_08_00[0]}),
     .sp12_h_l_01({net1352[0], net1352[1], net1352[2], net1352[3],
     net1352[4], net1352[5], net1352[6], net1352[7], net1352[8],
     net1352[9], net1352[10], net1352[11], net1352[12], net1352[13],
     net1352[14], net1352[15], net1352[16], net1352[17], net1352[18],
     net1352[19], net1352[20], net1352[21], net1352[22], net1352[23]}),
     .sp12_h_l_02({net1351[0], net1351[1], net1351[2], net1351[3],
     net1351[4], net1351[5], net1351[6], net1351[7], net1351[8],
     net1351[9], net1351[10], net1351[11], net1351[12], net1351[13],
     net1351[14], net1351[15], net1351[16], net1351[17], net1351[18],
     net1351[19], net1351[20], net1351[21], net1351[22], net1351[23]}),
     .sp12_h_l_03({net1350[0], net1350[1], net1350[2], net1350[3],
     net1350[4], net1350[5], net1350[6], net1350[7], net1350[8],
     net1350[9], net1350[10], net1350[11], net1350[12], net1350[13],
     net1350[14], net1350[15], net1350[16], net1350[17], net1350[18],
     net1350[19], net1350[20], net1350[21], net1350[22], net1350[23]}),
     .sp12_h_l_04({net1349[0], net1349[1], net1349[2], net1349[3],
     net1349[4], net1349[5], net1349[6], net1349[7], net1349[8],
     net1349[9], net1349[10], net1349[11], net1349[12], net1349[13],
     net1349[14], net1349[15], net1349[16], net1349[17], net1349[18],
     net1349[19], net1349[20], net1349[21], net1349[22], net1349[23]}),
     .sp4_v_b_04({net1355[0], net1355[1], net1355[2], net1355[3],
     net1355[4], net1355[5], net1355[6], net1355[7], net1355[8],
     net1355[9], net1355[10], net1355[11], net1355[12], net1355[13],
     net1355[14], net1355[15], net1355[16], net1355[17], net1355[18],
     net1355[19], net1355[20], net1355[21], net1355[22], net1355[23],
     net1355[24], net1355[25], net1355[26], net1355[27], net1355[28],
     net1355[29], net1355[30], net1355[31], net1355[32], net1355[33],
     net1355[34], net1355[35], net1355[36], net1355[37], net1355[38],
     net1355[39], net1355[40], net1355[41], net1355[42], net1355[43],
     net1355[44], net1355[45], net1355[46], net1355[47]}),
     .sp4_v_b_03({net1356[0], net1356[1], net1356[2], net1356[3],
     net1356[4], net1356[5], net1356[6], net1356[7], net1356[8],
     net1356[9], net1356[10], net1356[11], net1356[12], net1356[13],
     net1356[14], net1356[15], net1356[16], net1356[17], net1356[18],
     net1356[19], net1356[20], net1356[21], net1356[22], net1356[23],
     net1356[24], net1356[25], net1356[26], net1356[27], net1356[28],
     net1356[29], net1356[30], net1356[31], net1356[32], net1356[33],
     net1356[34], net1356[35], net1356[36], net1356[37], net1356[38],
     net1356[39], net1356[40], net1356[41], net1356[42], net1356[43],
     net1356[44], net1356[45], net1356[46], net1356[47]}),
     .sp4_v_b_02({net1357[0], net1357[1], net1357[2], net1357[3],
     net1357[4], net1357[5], net1357[6], net1357[7], net1357[8],
     net1357[9], net1357[10], net1357[11], net1357[12], net1357[13],
     net1357[14], net1357[15], net1357[16], net1357[17], net1357[18],
     net1357[19], net1357[20], net1357[21], net1357[22], net1357[23],
     net1357[24], net1357[25], net1357[26], net1357[27], net1357[28],
     net1357[29], net1357[30], net1357[31], net1357[32], net1357[33],
     net1357[34], net1357[35], net1357[36], net1357[37], net1357[38],
     net1357[39], net1357[40], net1357[41], net1357[42], net1357[43],
     net1357[44], net1357[45], net1357[46], net1357[47]}),
     .bnr_op_01({slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0], slf_op_09_00[3], slf_op_09_00[2],
     slf_op_09_00[1], slf_op_09_00[0]}), .sp4_h_l_05({net1383[0],
     net1383[1], net1383[2], net1383[3], net1383[4], net1383[5],
     net1383[6], net1383[7], net1383[8], net1383[9], net1383[10],
     net1383[11], net1383[12], net1383[13], net1383[14], net1383[15],
     net1383[16], net1383[17], net1383[18], net1383[19], net1383[20],
     net1383[21], net1383[22], net1383[23], net1383[24], net1383[25],
     net1383[26], net1383[27], net1383[28], net1383[29], net1383[30],
     net1383[31], net1383[32], net1383[33], net1383[34], net1383[35],
     net1383[36], net1383[37], net1383[38], net1383[39], net1383[40],
     net1383[41], net1383[42], net1383[43], net1383[44], net1383[45],
     net1383[46], net1383[47]}), .sp4_h_l_06({net1382[0], net1382[1],
     net1382[2], net1382[3], net1382[4], net1382[5], net1382[6],
     net1382[7], net1382[8], net1382[9], net1382[10], net1382[11],
     net1382[12], net1382[13], net1382[14], net1382[15], net1382[16],
     net1382[17], net1382[18], net1382[19], net1382[20], net1382[21],
     net1382[22], net1382[23], net1382[24], net1382[25], net1382[26],
     net1382[27], net1382[28], net1382[29], net1382[30], net1382[31],
     net1382[32], net1382[33], net1382[34], net1382[35], net1382[36],
     net1382[37], net1382[38], net1382[39], net1382[40], net1382[41],
     net1382[42], net1382[43], net1382[44], net1382[45], net1382[46],
     net1382[47]}), .sp4_h_l_07({net1381[0], net1381[1], net1381[2],
     net1381[3], net1381[4], net1381[5], net1381[6], net1381[7],
     net1381[8], net1381[9], net1381[10], net1381[11], net1381[12],
     net1381[13], net1381[14], net1381[15], net1381[16], net1381[17],
     net1381[18], net1381[19], net1381[20], net1381[21], net1381[22],
     net1381[23], net1381[24], net1381[25], net1381[26], net1381[27],
     net1381[28], net1381[29], net1381[30], net1381[31], net1381[32],
     net1381[33], net1381[34], net1381[35], net1381[36], net1381[37],
     net1381[38], net1381[39], net1381[40], net1381[41], net1381[42],
     net1381[43], net1381[44], net1381[45], net1381[46], net1381[47]}),
     .sp4_h_l_08({net1380[0], net1380[1], net1380[2], net1380[3],
     net1380[4], net1380[5], net1380[6], net1380[7], net1380[8],
     net1380[9], net1380[10], net1380[11], net1380[12], net1380[13],
     net1380[14], net1380[15], net1380[16], net1380[17], net1380[18],
     net1380[19], net1380[20], net1380[21], net1380[22], net1380[23],
     net1380[24], net1380[25], net1380[26], net1380[27], net1380[28],
     net1380[29], net1380[30], net1380[31], net1380[32], net1380[33],
     net1380[34], net1380[35], net1380[36], net1380[37], net1380[38],
     net1380[39], net1380[40], net1380[41], net1380[42], net1380[43],
     net1380[44], net1380[45], net1380[46], net1380[47]}),
     .sp4_h_r_08({net1285[0], net1285[1], net1285[2], net1285[3],
     net1285[4], net1285[5], net1285[6], net1285[7], net1285[8],
     net1285[9], net1285[10], net1285[11], net1285[12], net1285[13],
     net1285[14], net1285[15], net1285[16], net1285[17], net1285[18],
     net1285[19], net1285[20], net1285[21], net1285[22], net1285[23],
     net1285[24], net1285[25], net1285[26], net1285[27], net1285[28],
     net1285[29], net1285[30], net1285[31], net1285[32], net1285[33],
     net1285[34], net1285[35], net1285[36], net1285[37], net1285[38],
     net1285[39], net1285[40], net1285[41], net1285[42], net1285[43],
     net1285[44], net1285[45], net1285[46], net1285[47]}),
     .sp4_h_r_07({net1286[0], net1286[1], net1286[2], net1286[3],
     net1286[4], net1286[5], net1286[6], net1286[7], net1286[8],
     net1286[9], net1286[10], net1286[11], net1286[12], net1286[13],
     net1286[14], net1286[15], net1286[16], net1286[17], net1286[18],
     net1286[19], net1286[20], net1286[21], net1286[22], net1286[23],
     net1286[24], net1286[25], net1286[26], net1286[27], net1286[28],
     net1286[29], net1286[30], net1286[31], net1286[32], net1286[33],
     net1286[34], net1286[35], net1286[36], net1286[37], net1286[38],
     net1286[39], net1286[40], net1286[41], net1286[42], net1286[43],
     net1286[44], net1286[45], net1286[46], net1286[47]}),
     .sp4_h_r_06({net1287[0], net1287[1], net1287[2], net1287[3],
     net1287[4], net1287[5], net1287[6], net1287[7], net1287[8],
     net1287[9], net1287[10], net1287[11], net1287[12], net1287[13],
     net1287[14], net1287[15], net1287[16], net1287[17], net1287[18],
     net1287[19], net1287[20], net1287[21], net1287[22], net1287[23],
     net1287[24], net1287[25], net1287[26], net1287[27], net1287[28],
     net1287[29], net1287[30], net1287[31], net1287[32], net1287[33],
     net1287[34], net1287[35], net1287[36], net1287[37], net1287[38],
     net1287[39], net1287[40], net1287[41], net1287[42], net1287[43],
     net1287[44], net1287[45], net1287[46], net1287[47]}),
     .sp4_h_r_05({net1288[0], net1288[1], net1288[2], net1288[3],
     net1288[4], net1288[5], net1288[6], net1288[7], net1288[8],
     net1288[9], net1288[10], net1288[11], net1288[12], net1288[13],
     net1288[14], net1288[15], net1288[16], net1288[17], net1288[18],
     net1288[19], net1288[20], net1288[21], net1288[22], net1288[23],
     net1288[24], net1288[25], net1288[26], net1288[27], net1288[28],
     net1288[29], net1288[30], net1288[31], net1288[32], net1288[33],
     net1288[34], net1288[35], net1288[36], net1288[37], net1288[38],
     net1288[39], net1288[40], net1288[41], net1288[42], net1288[43],
     net1288[44], net1288[45], net1288[46], net1288[47]}),
     .slf_op_05({net1391[0], net1391[1], net1391[2], net1391[3],
     net1391[4], net1391[5], net1391[6], net1391[7]}),
     .slf_op_06({net1390[0], net1390[1], net1390[2], net1390[3],
     net1390[4], net1390[5], net1390[6], net1390[7]}),
     .slf_op_07({net1389[0], net1389[1], net1389[2], net1389[3],
     net1389[4], net1389[5], net1389[6], net1389[7]}),
     .slf_op_08(slf_op_08_08[7:0]), .rgt_op_08(slf_op_09_08[7:0]),
     .rgt_op_07({net1294[0], net1294[1], net1294[2], net1294[3],
     net1294[4], net1294[5], net1294[6], net1294[7]}),
     .rgt_op_06({net1295[0], net1295[1], net1295[2], net1295[3],
     net1295[4], net1295[5], net1295[6], net1295[7]}),
     .rgt_op_05({net1296[0], net1296[1], net1296[2], net1296[3],
     net1296[4], net1296[5], net1296[6], net1296[7]}),
     .lft_op_08(slf_op_07_08[7:0]), .lft_op_07(slf_op_07_07[7:0]),
     .lft_op_06(slf_op_07_06[7:0]), .lft_op_05(slf_op_07_05[7:0]),
     .sp12_h_l_08({net1402[0], net1402[1], net1402[2], net1402[3],
     net1402[4], net1402[5], net1402[6], net1402[7], net1402[8],
     net1402[9], net1402[10], net1402[11], net1402[12], net1402[13],
     net1402[14], net1402[15], net1402[16], net1402[17], net1402[18],
     net1402[19], net1402[20], net1402[21], net1402[22], net1402[23]}),
     .sp12_h_l_07({net1401[0], net1401[1], net1401[2], net1401[3],
     net1401[4], net1401[5], net1401[6], net1401[7], net1401[8],
     net1401[9], net1401[10], net1401[11], net1401[12], net1401[13],
     net1401[14], net1401[15], net1401[16], net1401[17], net1401[18],
     net1401[19], net1401[20], net1401[21], net1401[22], net1401[23]}),
     .sp12_h_l_06({net1400[0], net1400[1], net1400[2], net1400[3],
     net1400[4], net1400[5], net1400[6], net1400[7], net1400[8],
     net1400[9], net1400[10], net1400[11], net1400[12], net1400[13],
     net1400[14], net1400[15], net1400[16], net1400[17], net1400[18],
     net1400[19], net1400[20], net1400[21], net1400[22], net1400[23]}),
     .sp12_h_r_05({net1304[0], net1304[1], net1304[2], net1304[3],
     net1304[4], net1304[5], net1304[6], net1304[7], net1304[8],
     net1304[9], net1304[10], net1304[11], net1304[12], net1304[13],
     net1304[14], net1304[15], net1304[16], net1304[17], net1304[18],
     net1304[19], net1304[20], net1304[21], net1304[22], net1304[23]}),
     .sp12_h_r_06({net1305[0], net1305[1], net1305[2], net1305[3],
     net1305[4], net1305[5], net1305[6], net1305[7], net1305[8],
     net1305[9], net1305[10], net1305[11], net1305[12], net1305[13],
     net1305[14], net1305[15], net1305[16], net1305[17], net1305[18],
     net1305[19], net1305[20], net1305[21], net1305[22], net1305[23]}),
     .sp12_h_r_07({net1306[0], net1306[1], net1306[2], net1306[3],
     net1306[4], net1306[5], net1306[6], net1306[7], net1306[8],
     net1306[9], net1306[10], net1306[11], net1306[12], net1306[13],
     net1306[14], net1306[15], net1306[16], net1306[17], net1306[18],
     net1306[19], net1306[20], net1306[21], net1306[22], net1306[23]}),
     .sp12_h_r_08({net1307[0], net1307[1], net1307[2], net1307[3],
     net1307[4], net1307[5], net1307[6], net1307[7], net1307[8],
     net1307[9], net1307[10], net1307[11], net1307[12], net1307[13],
     net1307[14], net1307[15], net1307[16], net1307[17], net1307[18],
     net1307[19], net1307[20], net1307[21], net1307[22], net1307[23]}),
     .sp12_h_l_05({net1399[0], net1399[1], net1399[2], net1399[3],
     net1399[4], net1399[5], net1399[6], net1399[7], net1399[8],
     net1399[9], net1399[10], net1399[11], net1399[12], net1399[13],
     net1399[14], net1399[15], net1399[16], net1399[17], net1399[18],
     net1399[19], net1399[20], net1399[21], net1399[22], net1399[23]}),
     .sp4_r_v_b_05({net1309[0], net1309[1], net1309[2], net1309[3],
     net1309[4], net1309[5], net1309[6], net1309[7], net1309[8],
     net1309[9], net1309[10], net1309[11], net1309[12], net1309[13],
     net1309[14], net1309[15], net1309[16], net1309[17], net1309[18],
     net1309[19], net1309[20], net1309[21], net1309[22], net1309[23],
     net1309[24], net1309[25], net1309[26], net1309[27], net1309[28],
     net1309[29], net1309[30], net1309[31], net1309[32], net1309[33],
     net1309[34], net1309[35], net1309[36], net1309[37], net1309[38],
     net1309[39], net1309[40], net1309[41], net1309[42], net1309[43],
     net1309[44], net1309[45], net1309[46], net1309[47]}),
     .sp4_r_v_b_06({net1310[0], net1310[1], net1310[2], net1310[3],
     net1310[4], net1310[5], net1310[6], net1310[7], net1310[8],
     net1310[9], net1310[10], net1310[11], net1310[12], net1310[13],
     net1310[14], net1310[15], net1310[16], net1310[17], net1310[18],
     net1310[19], net1310[20], net1310[21], net1310[22], net1310[23],
     net1310[24], net1310[25], net1310[26], net1310[27], net1310[28],
     net1310[29], net1310[30], net1310[31], net1310[32], net1310[33],
     net1310[34], net1310[35], net1310[36], net1310[37], net1310[38],
     net1310[39], net1310[40], net1310[41], net1310[42], net1310[43],
     net1310[44], net1310[45], net1310[46], net1310[47]}),
     .sp4_r_v_b_07({net1311[0], net1311[1], net1311[2], net1311[3],
     net1311[4], net1311[5], net1311[6], net1311[7], net1311[8],
     net1311[9], net1311[10], net1311[11], net1311[12], net1311[13],
     net1311[14], net1311[15], net1311[16], net1311[17], net1311[18],
     net1311[19], net1311[20], net1311[21], net1311[22], net1311[23],
     net1311[24], net1311[25], net1311[26], net1311[27], net1311[28],
     net1311[29], net1311[30], net1311[31], net1311[32], net1311[33],
     net1311[34], net1311[35], net1311[36], net1311[37], net1311[38],
     net1311[39], net1311[40], net1311[41], net1311[42], net1311[43],
     net1311[44], net1311[45], net1311[46], net1311[47]}),
     .sp4_r_v_b_08({net1312[0], net1312[1], net1312[2], net1312[3],
     net1312[4], net1312[5], net1312[6], net1312[7], net1312[8],
     net1312[9], net1312[10], net1312[11], net1312[12], net1312[13],
     net1312[14], net1312[15], net1312[16], net1312[17], net1312[18],
     net1312[19], net1312[20], net1312[21], net1312[22], net1312[23],
     net1312[24], net1312[25], net1312[26], net1312[27], net1312[28],
     net1312[29], net1312[30], net1312[31], net1312[32], net1312[33],
     net1312[34], net1312[35], net1312[36], net1312[37], net1312[38],
     net1312[39], net1312[40], net1312[41], net1312[42], net1312[43],
     net1312[44], net1312[45], net1312[46], net1312[47]}),
     .sp4_v_b_08({net1407[0], net1407[1], net1407[2], net1407[3],
     net1407[4], net1407[5], net1407[6], net1407[7], net1407[8],
     net1407[9], net1407[10], net1407[11], net1407[12], net1407[13],
     net1407[14], net1407[15], net1407[16], net1407[17], net1407[18],
     net1407[19], net1407[20], net1407[21], net1407[22], net1407[23],
     net1407[24], net1407[25], net1407[26], net1407[27], net1407[28],
     net1407[29], net1407[30], net1407[31], net1407[32], net1407[33],
     net1407[34], net1407[35], net1407[36], net1407[37], net1407[38],
     net1407[39], net1407[40], net1407[41], net1407[42], net1407[43],
     net1407[44], net1407[45], net1407[46], net1407[47]}),
     .sp4_v_b_07({net1406[0], net1406[1], net1406[2], net1406[3],
     net1406[4], net1406[5], net1406[6], net1406[7], net1406[8],
     net1406[9], net1406[10], net1406[11], net1406[12], net1406[13],
     net1406[14], net1406[15], net1406[16], net1406[17], net1406[18],
     net1406[19], net1406[20], net1406[21], net1406[22], net1406[23],
     net1406[24], net1406[25], net1406[26], net1406[27], net1406[28],
     net1406[29], net1406[30], net1406[31], net1406[32], net1406[33],
     net1406[34], net1406[35], net1406[36], net1406[37], net1406[38],
     net1406[39], net1406[40], net1406[41], net1406[42], net1406[43],
     net1406[44], net1406[45], net1406[46], net1406[47]}),
     .sp4_v_b_06({net1405[0], net1405[1], net1405[2], net1405[3],
     net1405[4], net1405[5], net1405[6], net1405[7], net1405[8],
     net1405[9], net1405[10], net1405[11], net1405[12], net1405[13],
     net1405[14], net1405[15], net1405[16], net1405[17], net1405[18],
     net1405[19], net1405[20], net1405[21], net1405[22], net1405[23],
     net1405[24], net1405[25], net1405[26], net1405[27], net1405[28],
     net1405[29], net1405[30], net1405[31], net1405[32], net1405[33],
     net1405[34], net1405[35], net1405[36], net1405[37], net1405[38],
     net1405[39], net1405[40], net1405[41], net1405[42], net1405[43],
     net1405[44], net1405[45], net1405[46], net1405[47]}),
     .sp4_v_b_05({net1404[0], net1404[1], net1404[2], net1404[3],
     net1404[4], net1404[5], net1404[6], net1404[7], net1404[8],
     net1404[9], net1404[10], net1404[11], net1404[12], net1404[13],
     net1404[14], net1404[15], net1404[16], net1404[17], net1404[18],
     net1404[19], net1404[20], net1404[21], net1404[22], net1404[23],
     net1404[24], net1404[25], net1404[26], net1404[27], net1404[28],
     net1404[29], net1404[30], net1404[31], net1404[32], net1404[33],
     net1404[34], net1404[35], net1404[36], net1404[37], net1404[38],
     net1404[39], net1404[40], net1404[41], net1404[42], net1404[43],
     net1404[44], net1404[45], net1404[46], net1404[47]}),
     .pgate(pgate_r[143:16]), .reset_b(reset_b_r[143:16]),
     .wl(wl_r[143:16]), .sp12_v_t_08(sp12_v_t_08_08[23:0]),
     .tnr_op_08(tnr_op_08_08[7:0]), .top_op_08(top_op_08_08[7:0]),
     .tnl_op_08(tnl_op_08_08[7:0]), .sp4_v_t_08(sp4_v_t_08_08[47:0]),
     .lc_bot(tgnd_br_q), .op_vic(op_vic_08_08),
     .sp12_v_b_01({net901[0], net901[1], net901[2], net901[3],
     net901[4], net901[5], net901[6], net901[7], net901[8], net901[9],
     net901[10], net901[11], net901[12], net901[13], net901[14],
     net901[15], net901[16], net901[17], net901[18], net901[19],
     net901[20], net901[21], net901[22], net901[23]}));
lt_1x8_bot_ice1f I_lt_col_b07 ( .glb_netwk_bot({net939[0], net939[1],
     net939[2], net939[3], net939[4], net939[5], net939[6],
     net939[7]}), .rgt_op_03({net1330[0], net1330[1], net1330[2],
     net1330[3], net1330[4], net1330[5], net1330[6], net1330[7]}),
     .slf_op_02(slf_op_07_02[7:0]), .rgt_op_02({net1332[0], net1332[1],
     net1332[2], net1332[3], net1332[4], net1332[5], net1332[6],
     net1332[7]}), .rgt_op_01({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7]}),
     .purst(purst), .prog(prog), .lft_op_04(lft_op_07_04[7:0]),
     .lft_op_03(lft_op_07_03[7:0]), .lft_op_02(lft_op_07_02[7:0]),
     .lft_op_01(lft_op_07_01[7:0]), .rgt_op_04({net1340[0], net1340[1],
     net1340[2], net1340[3], net1340[4], net1340[5], net1340[6],
     net1340[7]}), .carry_in(tgnd_br_q), .bnl_op_01({bnl_op_07_01[3],
     bnl_op_07_01[2], bnl_op_07_01[1], bnl_op_07_01[0],
     bnl_op_07_01[3], bnl_op_07_01[2], bnl_op_07_01[1],
     bnl_op_07_01[0]}), .slf_op_04(slf_op_07_04[7:0]),
     .slf_op_03(slf_op_07_03[7:0]), .slf_op_01(slf_op_07_01[7:0]),
     .sp4_h_l_04(sp4_h_l_07_04[47:0]), .carry_out(carry_out_07_08),
     .vdd_cntl(vdd_cntl_r[143:16]), .sp12_h_r_04({net1349[0],
     net1349[1], net1349[2], net1349[3], net1349[4], net1349[5],
     net1349[6], net1349[7], net1349[8], net1349[9], net1349[10],
     net1349[11], net1349[12], net1349[13], net1349[14], net1349[15],
     net1349[16], net1349[17], net1349[18], net1349[19], net1349[20],
     net1349[21], net1349[22], net1349[23]}), .sp12_h_r_03({net1350[0],
     net1350[1], net1350[2], net1350[3], net1350[4], net1350[5],
     net1350[6], net1350[7], net1350[8], net1350[9], net1350[10],
     net1350[11], net1350[12], net1350[13], net1350[14], net1350[15],
     net1350[16], net1350[17], net1350[18], net1350[19], net1350[20],
     net1350[21], net1350[22], net1350[23]}), .sp12_h_r_02({net1351[0],
     net1351[1], net1351[2], net1351[3], net1351[4], net1351[5],
     net1351[6], net1351[7], net1351[8], net1351[9], net1351[10],
     net1351[11], net1351[12], net1351[13], net1351[14], net1351[15],
     net1351[16], net1351[17], net1351[18], net1351[19], net1351[20],
     net1351[21], net1351[22], net1351[23]}), .sp12_h_r_01({net1352[0],
     net1352[1], net1352[2], net1352[3], net1352[4], net1352[5],
     net1352[6], net1352[7], net1352[8], net1352[9], net1352[10],
     net1352[11], net1352[12], net1352[13], net1352[14], net1352[15],
     net1352[16], net1352[17], net1352[18], net1352[19], net1352[20],
     net1352[21], net1352[22], net1352[23]}),
     .glb_netwk_col(clk_tree_drv_br[7:0]),
     .sp4_v_b_01(sp4_v_b_07_01[47:0]), .sp4_r_v_b_04({net1355[0],
     net1355[1], net1355[2], net1355[3], net1355[4], net1355[5],
     net1355[6], net1355[7], net1355[8], net1355[9], net1355[10],
     net1355[11], net1355[12], net1355[13], net1355[14], net1355[15],
     net1355[16], net1355[17], net1355[18], net1355[19], net1355[20],
     net1355[21], net1355[22], net1355[23], net1355[24], net1355[25],
     net1355[26], net1355[27], net1355[28], net1355[29], net1355[30],
     net1355[31], net1355[32], net1355[33], net1355[34], net1355[35],
     net1355[36], net1355[37], net1355[38], net1355[39], net1355[40],
     net1355[41], net1355[42], net1355[43], net1355[44], net1355[45],
     net1355[46], net1355[47]}), .sp4_r_v_b_03({net1356[0], net1356[1],
     net1356[2], net1356[3], net1356[4], net1356[5], net1356[6],
     net1356[7], net1356[8], net1356[9], net1356[10], net1356[11],
     net1356[12], net1356[13], net1356[14], net1356[15], net1356[16],
     net1356[17], net1356[18], net1356[19], net1356[20], net1356[21],
     net1356[22], net1356[23], net1356[24], net1356[25], net1356[26],
     net1356[27], net1356[28], net1356[29], net1356[30], net1356[31],
     net1356[32], net1356[33], net1356[34], net1356[35], net1356[36],
     net1356[37], net1356[38], net1356[39], net1356[40], net1356[41],
     net1356[42], net1356[43], net1356[44], net1356[45], net1356[46],
     net1356[47]}), .sp4_r_v_b_02({net1357[0], net1357[1], net1357[2],
     net1357[3], net1357[4], net1357[5], net1357[6], net1357[7],
     net1357[8], net1357[9], net1357[10], net1357[11], net1357[12],
     net1357[13], net1357[14], net1357[15], net1357[16], net1357[17],
     net1357[18], net1357[19], net1357[20], net1357[21], net1357[22],
     net1357[23], net1357[24], net1357[25], net1357[26], net1357[27],
     net1357[28], net1357[29], net1357[30], net1357[31], net1357[32],
     net1357[33], net1357[34], net1357[35], net1357[36], net1357[37],
     net1357[38], net1357[39], net1357[40], net1357[41], net1357[42],
     net1357[43], net1357[44], net1357[45], net1357[46], net1357[47]}),
     .sp4_r_v_b_01({net889[0], net889[1], net889[2], net889[3],
     net889[4], net889[5], net889[6], net889[7], net889[8], net889[9],
     net889[10], net889[11], net889[12], net889[13], net889[14],
     net889[15], net889[16], net889[17], net889[18], net889[19],
     net889[20], net889[21], net889[22], net889[23], net889[24],
     net889[25], net889[26], net889[27], net889[28], net889[29],
     net889[30], net889[31], net889[32], net889[33], net889[34],
     net889[35], net889[36], net889[37], net889[38], net889[39],
     net889[40], net889[41], net889[42], net889[43], net889[44],
     net889[45], net889[46], net889[47]}), .sp4_h_r_04({net1359[0],
     net1359[1], net1359[2], net1359[3], net1359[4], net1359[5],
     net1359[6], net1359[7], net1359[8], net1359[9], net1359[10],
     net1359[11], net1359[12], net1359[13], net1359[14], net1359[15],
     net1359[16], net1359[17], net1359[18], net1359[19], net1359[20],
     net1359[21], net1359[22], net1359[23], net1359[24], net1359[25],
     net1359[26], net1359[27], net1359[28], net1359[29], net1359[30],
     net1359[31], net1359[32], net1359[33], net1359[34], net1359[35],
     net1359[36], net1359[37], net1359[38], net1359[39], net1359[40],
     net1359[41], net1359[42], net1359[43], net1359[44], net1359[45],
     net1359[46], net1359[47]}), .sp4_h_r_03({net1360[0], net1360[1],
     net1360[2], net1360[3], net1360[4], net1360[5], net1360[6],
     net1360[7], net1360[8], net1360[9], net1360[10], net1360[11],
     net1360[12], net1360[13], net1360[14], net1360[15], net1360[16],
     net1360[17], net1360[18], net1360[19], net1360[20], net1360[21],
     net1360[22], net1360[23], net1360[24], net1360[25], net1360[26],
     net1360[27], net1360[28], net1360[29], net1360[30], net1360[31],
     net1360[32], net1360[33], net1360[34], net1360[35], net1360[36],
     net1360[37], net1360[38], net1360[39], net1360[40], net1360[41],
     net1360[42], net1360[43], net1360[44], net1360[45], net1360[46],
     net1360[47]}), .sp4_h_r_02({net1361[0], net1361[1], net1361[2],
     net1361[3], net1361[4], net1361[5], net1361[6], net1361[7],
     net1361[8], net1361[9], net1361[10], net1361[11], net1361[12],
     net1361[13], net1361[14], net1361[15], net1361[16], net1361[17],
     net1361[18], net1361[19], net1361[20], net1361[21], net1361[22],
     net1361[23], net1361[24], net1361[25], net1361[26], net1361[27],
     net1361[28], net1361[29], net1361[30], net1361[31], net1361[32],
     net1361[33], net1361[34], net1361[35], net1361[36], net1361[37],
     net1361[38], net1361[39], net1361[40], net1361[41], net1361[42],
     net1361[43], net1361[44], net1361[45], net1361[46], net1361[47]}),
     .sp4_h_r_01({net1362[0], net1362[1], net1362[2], net1362[3],
     net1362[4], net1362[5], net1362[6], net1362[7], net1362[8],
     net1362[9], net1362[10], net1362[11], net1362[12], net1362[13],
     net1362[14], net1362[15], net1362[16], net1362[17], net1362[18],
     net1362[19], net1362[20], net1362[21], net1362[22], net1362[23],
     net1362[24], net1362[25], net1362[26], net1362[27], net1362[28],
     net1362[29], net1362[30], net1362[31], net1362[32], net1362[33],
     net1362[34], net1362[35], net1362[36], net1362[37], net1362[38],
     net1362[39], net1362[40], net1362[41], net1362[42], net1362[43],
     net1362[44], net1362[45], net1362[46], net1362[47]}),
     .sp4_h_l_03(sp4_h_l_07_03[47:0]),
     .sp4_h_l_02(sp4_h_l_07_02[47:0]),
     .sp4_h_l_01(sp4_h_l_07_01[47:0]), .bl(bl[53:0]),
     .bot_op_01({slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0], slf_op_07_00[3], slf_op_07_00[2],
     slf_op_07_00[1], slf_op_07_00[0]}),
     .sp12_h_l_01(sp12_h_l_07_01[23:0]),
     .sp12_h_l_02(sp12_h_l_07_02[23:0]),
     .sp12_h_l_03(sp12_h_l_07_03[23:0]),
     .sp12_h_l_04(sp12_h_l_07_04[23:0]),
     .sp4_v_b_04(sp4_v_b_07_04[47:0]),
     .sp4_v_b_03(sp4_v_b_07_03[47:0]),
     .sp4_v_b_02(sp4_v_b_07_02[47:0]), .bnr_op_01({slf_op_08_00[3],
     slf_op_08_00[2], slf_op_08_00[1], slf_op_08_00[0],
     slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0]}), .sp4_h_l_05(sp4_h_l_07_05[47:0]),
     .sp4_h_l_06(sp4_h_l_07_06[47:0]),
     .sp4_h_l_07(sp4_h_l_07_07[47:0]),
     .sp4_h_l_08(sp4_h_l_07_08[47:0]), .sp4_h_r_08({net1380[0],
     net1380[1], net1380[2], net1380[3], net1380[4], net1380[5],
     net1380[6], net1380[7], net1380[8], net1380[9], net1380[10],
     net1380[11], net1380[12], net1380[13], net1380[14], net1380[15],
     net1380[16], net1380[17], net1380[18], net1380[19], net1380[20],
     net1380[21], net1380[22], net1380[23], net1380[24], net1380[25],
     net1380[26], net1380[27], net1380[28], net1380[29], net1380[30],
     net1380[31], net1380[32], net1380[33], net1380[34], net1380[35],
     net1380[36], net1380[37], net1380[38], net1380[39], net1380[40],
     net1380[41], net1380[42], net1380[43], net1380[44], net1380[45],
     net1380[46], net1380[47]}), .sp4_h_r_07({net1381[0], net1381[1],
     net1381[2], net1381[3], net1381[4], net1381[5], net1381[6],
     net1381[7], net1381[8], net1381[9], net1381[10], net1381[11],
     net1381[12], net1381[13], net1381[14], net1381[15], net1381[16],
     net1381[17], net1381[18], net1381[19], net1381[20], net1381[21],
     net1381[22], net1381[23], net1381[24], net1381[25], net1381[26],
     net1381[27], net1381[28], net1381[29], net1381[30], net1381[31],
     net1381[32], net1381[33], net1381[34], net1381[35], net1381[36],
     net1381[37], net1381[38], net1381[39], net1381[40], net1381[41],
     net1381[42], net1381[43], net1381[44], net1381[45], net1381[46],
     net1381[47]}), .sp4_h_r_06({net1382[0], net1382[1], net1382[2],
     net1382[3], net1382[4], net1382[5], net1382[6], net1382[7],
     net1382[8], net1382[9], net1382[10], net1382[11], net1382[12],
     net1382[13], net1382[14], net1382[15], net1382[16], net1382[17],
     net1382[18], net1382[19], net1382[20], net1382[21], net1382[22],
     net1382[23], net1382[24], net1382[25], net1382[26], net1382[27],
     net1382[28], net1382[29], net1382[30], net1382[31], net1382[32],
     net1382[33], net1382[34], net1382[35], net1382[36], net1382[37],
     net1382[38], net1382[39], net1382[40], net1382[41], net1382[42],
     net1382[43], net1382[44], net1382[45], net1382[46], net1382[47]}),
     .sp4_h_r_05({net1383[0], net1383[1], net1383[2], net1383[3],
     net1383[4], net1383[5], net1383[6], net1383[7], net1383[8],
     net1383[9], net1383[10], net1383[11], net1383[12], net1383[13],
     net1383[14], net1383[15], net1383[16], net1383[17], net1383[18],
     net1383[19], net1383[20], net1383[21], net1383[22], net1383[23],
     net1383[24], net1383[25], net1383[26], net1383[27], net1383[28],
     net1383[29], net1383[30], net1383[31], net1383[32], net1383[33],
     net1383[34], net1383[35], net1383[36], net1383[37], net1383[38],
     net1383[39], net1383[40], net1383[41], net1383[42], net1383[43],
     net1383[44], net1383[45], net1383[46], net1383[47]}),
     .slf_op_05(slf_op_07_05[7:0]), .slf_op_06(slf_op_07_06[7:0]),
     .slf_op_07(slf_op_07_07[7:0]), .slf_op_08(slf_op_07_08[7:0]),
     .rgt_op_08(slf_op_08_08[7:0]), .rgt_op_07({net1389[0], net1389[1],
     net1389[2], net1389[3], net1389[4], net1389[5], net1389[6],
     net1389[7]}), .rgt_op_06({net1390[0], net1390[1], net1390[2],
     net1390[3], net1390[4], net1390[5], net1390[6], net1390[7]}),
     .rgt_op_05({net1391[0], net1391[1], net1391[2], net1391[3],
     net1391[4], net1391[5], net1391[6], net1391[7]}),
     .lft_op_08(lft_op_07_08[7:0]), .lft_op_07(lft_op_07_07[7:0]),
     .lft_op_06(lft_op_07_06[7:0]), .lft_op_05(lft_op_07_05[7:0]),
     .sp12_h_l_08(sp12_h_l_07_08[23:0]),
     .sp12_h_l_07(sp12_h_l_07_07[23:0]),
     .sp12_h_l_06(sp12_h_l_07_06[23:0]), .sp12_h_r_05({net1399[0],
     net1399[1], net1399[2], net1399[3], net1399[4], net1399[5],
     net1399[6], net1399[7], net1399[8], net1399[9], net1399[10],
     net1399[11], net1399[12], net1399[13], net1399[14], net1399[15],
     net1399[16], net1399[17], net1399[18], net1399[19], net1399[20],
     net1399[21], net1399[22], net1399[23]}), .sp12_h_r_06({net1400[0],
     net1400[1], net1400[2], net1400[3], net1400[4], net1400[5],
     net1400[6], net1400[7], net1400[8], net1400[9], net1400[10],
     net1400[11], net1400[12], net1400[13], net1400[14], net1400[15],
     net1400[16], net1400[17], net1400[18], net1400[19], net1400[20],
     net1400[21], net1400[22], net1400[23]}), .sp12_h_r_07({net1401[0],
     net1401[1], net1401[2], net1401[3], net1401[4], net1401[5],
     net1401[6], net1401[7], net1401[8], net1401[9], net1401[10],
     net1401[11], net1401[12], net1401[13], net1401[14], net1401[15],
     net1401[16], net1401[17], net1401[18], net1401[19], net1401[20],
     net1401[21], net1401[22], net1401[23]}), .sp12_h_r_08({net1402[0],
     net1402[1], net1402[2], net1402[3], net1402[4], net1402[5],
     net1402[6], net1402[7], net1402[8], net1402[9], net1402[10],
     net1402[11], net1402[12], net1402[13], net1402[14], net1402[15],
     net1402[16], net1402[17], net1402[18], net1402[19], net1402[20],
     net1402[21], net1402[22], net1402[23]}),
     .sp12_h_l_05(sp12_h_l_07_05[23:0]), .sp4_r_v_b_05({net1404[0],
     net1404[1], net1404[2], net1404[3], net1404[4], net1404[5],
     net1404[6], net1404[7], net1404[8], net1404[9], net1404[10],
     net1404[11], net1404[12], net1404[13], net1404[14], net1404[15],
     net1404[16], net1404[17], net1404[18], net1404[19], net1404[20],
     net1404[21], net1404[22], net1404[23], net1404[24], net1404[25],
     net1404[26], net1404[27], net1404[28], net1404[29], net1404[30],
     net1404[31], net1404[32], net1404[33], net1404[34], net1404[35],
     net1404[36], net1404[37], net1404[38], net1404[39], net1404[40],
     net1404[41], net1404[42], net1404[43], net1404[44], net1404[45],
     net1404[46], net1404[47]}), .sp4_r_v_b_06({net1405[0], net1405[1],
     net1405[2], net1405[3], net1405[4], net1405[5], net1405[6],
     net1405[7], net1405[8], net1405[9], net1405[10], net1405[11],
     net1405[12], net1405[13], net1405[14], net1405[15], net1405[16],
     net1405[17], net1405[18], net1405[19], net1405[20], net1405[21],
     net1405[22], net1405[23], net1405[24], net1405[25], net1405[26],
     net1405[27], net1405[28], net1405[29], net1405[30], net1405[31],
     net1405[32], net1405[33], net1405[34], net1405[35], net1405[36],
     net1405[37], net1405[38], net1405[39], net1405[40], net1405[41],
     net1405[42], net1405[43], net1405[44], net1405[45], net1405[46],
     net1405[47]}), .sp4_r_v_b_07({net1406[0], net1406[1], net1406[2],
     net1406[3], net1406[4], net1406[5], net1406[6], net1406[7],
     net1406[8], net1406[9], net1406[10], net1406[11], net1406[12],
     net1406[13], net1406[14], net1406[15], net1406[16], net1406[17],
     net1406[18], net1406[19], net1406[20], net1406[21], net1406[22],
     net1406[23], net1406[24], net1406[25], net1406[26], net1406[27],
     net1406[28], net1406[29], net1406[30], net1406[31], net1406[32],
     net1406[33], net1406[34], net1406[35], net1406[36], net1406[37],
     net1406[38], net1406[39], net1406[40], net1406[41], net1406[42],
     net1406[43], net1406[44], net1406[45], net1406[46], net1406[47]}),
     .sp4_r_v_b_08({net1407[0], net1407[1], net1407[2], net1407[3],
     net1407[4], net1407[5], net1407[6], net1407[7], net1407[8],
     net1407[9], net1407[10], net1407[11], net1407[12], net1407[13],
     net1407[14], net1407[15], net1407[16], net1407[17], net1407[18],
     net1407[19], net1407[20], net1407[21], net1407[22], net1407[23],
     net1407[24], net1407[25], net1407[26], net1407[27], net1407[28],
     net1407[29], net1407[30], net1407[31], net1407[32], net1407[33],
     net1407[34], net1407[35], net1407[36], net1407[37], net1407[38],
     net1407[39], net1407[40], net1407[41], net1407[42], net1407[43],
     net1407[44], net1407[45], net1407[46], net1407[47]}),
     .sp4_v_b_08(sp4_v_b_07_08[47:0]),
     .sp4_v_b_07(sp4_v_b_07_07[47:0]),
     .sp4_v_b_06(sp4_v_b_07_06[47:0]),
     .sp4_v_b_05(sp4_v_b_07_05[47:0]), .pgate(pgate_r[143:16]),
     .reset_b(reset_b_r[143:16]), .wl(wl_r[143:16]),
     .sp12_v_t_08(sp12_v_t_07_08[23:0]), .tnr_op_08(tnr_op_07_08[7:0]),
     .top_op_08(top_op_07_08[7:0]), .tnl_op_08(tnl_op_07_08[7:0]),
     .sp4_v_t_08(sp4_v_t_07_08[47:0]), .lc_bot(tgnd_br_q),
     .op_vic(op_vic_07_08), .sp12_v_b_01({net903[0], net903[1],
     net903[2], net903[3], net903[4], net903[5], net903[6], net903[7],
     net903[8], net903[9], net903[10], net903[11], net903[12],
     net903[13], net903[14], net903[15], net903[16], net903[17],
     net903[18], net903[19], net903[20], net903[21], net903[22],
     net903[23]}));
fabric_buf_ice8p I485 ( .f_in(net0731), .f_out(padin_13_08b));
fabric_buf_ice8p I481 ( .f_in(net807), .f_out(fabric_out_13_02));
fabric_buf_ice8p I453 ( .f_in(net1437), .f_out(fabric_out_07_00));
fabric_buf_ice8p I482 ( .f_in(net808), .f_out(fabric_out_13_01));
fabric_buf_ice8p I480 ( .f_in(net809), .f_out(fabric_out_13_08));
fabric_buf_ice8p I454 ( .f_in(padinlat_b_r[11]), .f_out(padin_07_00a));
fabric_buf_ice8p I452 ( .f_in(net912), .f_out(fabric_out_12_00));
clk_quad_buf_x8_ice8p I428 ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));
clk_quad_buf_x8_ice8p I427 ( .clko(clk_tree_drv_br[7:0]),
     .clki(clk_center[7:0]));

endmodule
// Library - ice1chip, Cell - io_lft_bot_1x8_ice1f, View - schematic
// LAST TIME SAVED: Apr 11 16:03:08 2011
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module io_lft_bot_1x8_ice1f ( cf_l, fabric_out_07, fabric_out_08,
     fo_dlyadj, fo_fb, fo_ref, padeb, pado, sdo, slf_op_01, slf_op_02,
     slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07, slf_op_08,
     tclk_o, SP4_h_l_01, SP4_h_l_02, SP4_h_l_03, SP4_h_l_04,
     SP4_h_l_05, SP4_h_l_06, SP4_h_l_07, SP4_h_l_08, SP12_h_l_01,
     SP12_h_l_02, SP12_h_l_03, SP12_h_l_04, SP12_h_l_05, SP12_h_l_06,
     SP12_h_l_07, SP12_h_l_08, bl, pgate, reset_b, sp4_v_b_00_01,
     sp4_v_t_08, vdd_cntl, wl, bnr_op_00_01, bs_en, ceb, glb_netwk_col,
     hiz_b, hold, jtag_rowtest_mode_rowu0_b, last_rsr, mode, padin,
     prog, r, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04, rgt_op_05,
     rgt_op_06, rgt_op_07, rgt_op_08, sdi, shift, tclk, tnr_op_08,
     update );
output  fabric_out_07, fabric_out_08, fo_fb, fo_ref, sdo, tclk_o;


input  bs_en, ceb, hiz_b, hold, jtag_rowtest_mode_rowu0_b, mode, prog,
     r, sdi, shift, tclk, update;

output [3:0]  slf_op_08;
output [3:0]  slf_op_07;
output [3:0]  slf_op_05;
output [3:0]  slf_op_04;
output [3:0]  slf_op_03;
output [3:0]  slf_op_02;
output [3:0]  slf_op_06;
output [2:0]  fo_dlyadj;
output [11:0]  padeb;
output [3:0]  slf_op_01;
output [11:0]  pado;
output [191:0]  cf_l;

inout [47:0]  SP4_h_l_05;
inout [47:0]  SP4_h_l_02;
inout [47:0]  SP4_h_l_01;
inout [17:0]  bl;
inout [15:0]  sp4_v_t_08;
inout [23:0]  SP12_h_l_04;
inout [23:0]  SP12_h_l_03;
inout [47:0]  SP4_h_l_07;
inout [47:0]  SP4_h_l_03;
inout [23:0]  SP12_h_l_02;
inout [23:0]  SP12_h_l_06;
inout [47:0]  SP4_h_l_06;
inout [47:0]  SP4_h_l_04;
inout [23:0]  SP12_h_l_07;
inout [127:0]  pgate;
inout [127:0]  vdd_cntl;
inout [127:0]  wl;
inout [127:0]  reset_b;
inout [23:0]  SP12_h_l_05;
inout [47:0]  SP4_h_l_08;
inout [23:0]  SP12_h_l_08;
inout [15:0]  sp4_v_b_00_01;
inout [23:0]  SP12_h_l_01;

input [7:0]  bnr_op_00_01;
input [7:0]  tnr_op_08;
input [7:0]  rgt_op_02;
input [7:0]  rgt_op_03;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_04;
input [0:0]  last_rsr;
input [11:0]  padin;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_08;
input [7:0]  rgt_op_07;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net1009;

wire  [1:0]  net1014;

wire  [1:0]  net1003;

wire  [7:0]  glb_netwk_t;

wire  [1:0]  net0539;

wire  [1:0]  net1001;

wire  [1:0]  net0540;

wire  [1:0]  net1005;

wire  [7:0]  net884;

wire  [1:0]  net1010;

wire  [15:0]  net937;

wire  [1:0]  net1002;

wire  [15:0]  net901;

wire  [7:0]  net1007;

wire  [15:0]  net829;

wire  [1:0]  net1013;

wire  [1:0]  net1012;

wire  [15:0]  net793;

wire  [7:0]  net704;

wire  [7:0]  net1008;

wire  [15:0]  net757;

wire  [1:0]  net755;

wire  [7:0]  net1017;

wire  [7:0]  colbuf_cntl_b;

wire  [7:0]  net1016;

wire  [15:0]  net973;

wire  [1:0]  net0538;

wire  [7:0]  colbuf_cntl_t;

wire  [15:0]  net865;

wire  [7:0]  glb_netwk_b;



fabric_buf_ice8p I_fabric_buf_8p_0015 ( .f_in(net0546),
     .f_out(fo_ref));
fabric_buf_ice8p I162 ( .f_in(net883), .f_out(fo_fb));
tckbufx32_ice8p I_tck_halfbankcenter ( .in(tclk), .out(tclk_o));
tielo4x I483 ( .tielo(tiegnd));
tiehi4x I482 ( .tiehi(tievdd));
io_col4_lft_ice8p_v2 I_io_00_08 ( .cbit_colcntl({net704[0], net704[1],
     net704[2], net704[3], net704[4], net704[5], net704[6],
     net704[7]}), .ceb(ceb), .sdo(net743), .sdi(sdi), .spiout({tiegnd,
     last_rsr[0]}), .cdone_in(jtag_rowtest_mode_rowu0_b),
     .spioeb({tievdd, tiegnd}), .mode(mode), .shift(shift),
     .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[11:10]), .pado(pado[11:10]),
     .padeb(padeb[11:10]), .sp4_v_t(sp4_v_t_08[15:0]),
     .sp4_h_l(SP4_h_l_08[47:0]), .sp12_h_l(SP12_h_l_08[23:0]),
     .prog(prog), .spi_ss_in_b({net1012[0], net1012[1]}),
     .tnl_op(tnr_op_08[7:0]), .lft_op(rgt_op_08[7:0]),
     .bnl_op(rgt_op_07[7:0]), .pgate(pgate[127:112]),
     .reset(reset_b[127:112]), .sp4_v_b({net757[0], net757[1],
     net757[2], net757[3], net757[4], net757[5], net757[6], net757[7],
     net757[8], net757[9], net757[10], net757[11], net757[12],
     net757[13], net757[14], net757[15]}), .wl(wl[127:112]),
     .cf(cf_l[191:168]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_08[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fabric_out_08));
io_col4_lft_ice8p_v2 I_io_00_07 ( .cbit_colcntl({net1016[0],
     net1016[1], net1016[2], net1016[3], net1016[4], net1016[5],
     net1016[6], net1016[7]}), .ceb(ceb), .sdo(net815), .sdi(net743),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin({net755[0],
     net755[1]}), .pado({net755[0], net755[1]}), .padeb({net1001[0],
     net1001[1]}), .sp4_v_t({net757[0], net757[1], net757[2],
     net757[3], net757[4], net757[5], net757[6], net757[7], net757[8],
     net757[9], net757[10], net757[11], net757[12], net757[13],
     net757[14], net757[15]}), .sp4_h_l(SP4_h_l_07[47:0]),
     .sp12_h_l(SP12_h_l_07[23:0]), .prog(prog),
     .spi_ss_in_b({net1013[0], net1013[1]}), .tnl_op(rgt_op_08[7:0]),
     .lft_op(rgt_op_07[7:0]), .bnl_op(rgt_op_06[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b({net829[0], net829[1], net829[2], net829[3], net829[4],
     net829[5], net829[6], net829[7], net829[8], net829[9], net829[10],
     net829[11], net829[12], net829[13], net829[14], net829[15]}),
     .wl(wl[111:96]), .cf(cf_l[167:144]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[111:96]), .slf_op(slf_op_07[3:0]),
     .glb_netwk(glb_netwk_t[7:0]), .hold(hold),
     .fabric_out(fabric_out_07));
io_col4_lft_ice8p_v2 I_io_00_05 ( .cbit_colcntl(colbuf_cntl_t[7:0]),
     .ceb(ceb), .sdo(net959), .sdi(net779), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[7:6]), .pado(pado[7:6]),
     .padeb(padeb[7:6]), .sp4_v_t({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7], net793[8],
     net793[9], net793[10], net793[11], net793[12], net793[13],
     net793[14], net793[15]}), .sp4_h_l(SP4_h_l_05[47:0]),
     .sp12_h_l(SP12_h_l_05[23:0]), .prog(prog),
     .spi_ss_in_b({net1003[0], net1003[1]}), .tnl_op(rgt_op_06[7:0]),
     .lft_op(rgt_op_05[7:0]), .bnl_op(rgt_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]), .sp4_v_b({net973[0],
     net973[1], net973[2], net973[3], net973[4], net973[5], net973[6],
     net973[7], net973[8], net973[9], net973[10], net973[11],
     net973[12], net973[13], net973[14], net973[15]}), .wl(wl[79:64]),
     .cf(cf_l[119:96]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[1]));
io_col4_lft_ice8p_v2 I_io_00_06 ( .cbit_colcntl({net1017[0],
     net1017[1], net1017[2], net1017[3], net1017[4], net1017[5],
     net1017[6], net1017[7]}), .ceb(ceb), .sdo(net779), .sdi(net815),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin(padin[9:8]),
     .pado(pado[9:8]), .padeb(padeb[9:8]), .sp4_v_t({net829[0],
     net829[1], net829[2], net829[3], net829[4], net829[5], net829[6],
     net829[7], net829[8], net829[9], net829[10], net829[11],
     net829[12], net829[13], net829[14], net829[15]}),
     .sp4_h_l(SP4_h_l_06[47:0]), .sp12_h_l(SP12_h_l_06[23:0]),
     .prog(prog), .spi_ss_in_b({net1010[0], net1010[1]}),
     .tnl_op(rgt_op_07[7:0]), .lft_op(rgt_op_06[7:0]),
     .bnl_op(rgt_op_05[7:0]), .pgate(pgate[95:80]),
     .reset(reset_b[95:80]), .sp4_v_b({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7], net793[8],
     net793[9], net793[10], net793[11], net793[12], net793[13],
     net793[14], net793[15]}), .wl(wl[95:80]), .cf(cf_l[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk_t[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[2]));
io_col4_lft_ice8p_v2 I_io_00_02 ( .cbit_colcntl({net1007[0],
     net1007[1], net1007[2], net1007[3], net1007[4], net1007[5],
     net1007[6], net1007[7]}), .ceb(ceb), .sdo(net887), .sdi(net851),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin(padin[1:0]),
     .pado(pado[1:0]), .padeb(padeb[1:0]), .sp4_v_t({net865[0],
     net865[1], net865[2], net865[3], net865[4], net865[5], net865[6],
     net865[7], net865[8], net865[9], net865[10], net865[11],
     net865[12], net865[13], net865[14], net865[15]}),
     .sp4_h_l(SP4_h_l_02[47:0]), .sp12_h_l(SP12_h_l_02[23:0]),
     .prog(prog), .spi_ss_in_b({net1014[0], net1014[1]}),
     .tnl_op(rgt_op_03[7:0]), .lft_op(rgt_op_02[7:0]),
     .bnl_op(rgt_op_01[7:0]), .pgate(pgate[31:16]),
     .reset(reset_b[31:16]), .sp4_v_b({net901[0], net901[1], net901[2],
     net901[3], net901[4], net901[5], net901[6], net901[7], net901[8],
     net901[9], net901[10], net901[11], net901[12], net901[13],
     net901[14], net901[15]}), .wl(wl[31:16]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net883));
io_col4_lft_ice8p_v2 I_io_00_01 ( .cbit_colcntl({net884[0], net884[1],
     net884[2], net884[3], net884[4], net884[5], net884[6],
     net884[7]}), .ceb(ceb), .sdo(sdo), .sdi(net887), .spiout({tiegnd,
     tiegnd}), .cdone_in(tievdd), .spioeb({tievdd, tievdd}),
     .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en),
     .tclk(tclk_o), .update(update), .padin({net0538[0], net0538[1]}),
     .pado({net0539[0], net0539[1]}), .padeb({net0540[0], net0540[1]}),
     .sp4_v_t({net901[0], net901[1], net901[2], net901[3], net901[4],
     net901[5], net901[6], net901[7], net901[8], net901[9], net901[10],
     net901[11], net901[12], net901[13], net901[14], net901[15]}),
     .sp4_h_l(SP4_h_l_01[47:0]), .sp12_h_l(SP12_h_l_01[23:0]),
     .prog(prog), .spi_ss_in_b({net1005[0], net1005[1]}),
     .tnl_op(rgt_op_02[7:0]), .lft_op(rgt_op_01[7:0]),
     .bnl_op(bnr_op_00_01[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(sp4_v_b_00_01[15:0]),
     .wl(wl[15:0]), .cf(cf_l[23:0]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk_b[7:0]), .hold(hold), .fabric_out(net0546));
io_col4_lft_ice8p_v2 I_io_00_03 ( .cbit_colcntl({net1008[0],
     net1008[1], net1008[2], net1008[3], net1008[4], net1008[5],
     net1008[6], net1008[7]}), .ceb(ceb), .sdo(net851), .sdi(net923),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode), .shift(shift), .hiz_b(hiz_b), .r(r),
     .bs_en(bs_en), .tclk(tclk_o), .update(update), .padin(padin[3:2]),
     .pado(pado[3:2]), .padeb(padeb[3:2]), .sp4_v_t({net937[0],
     net937[1], net937[2], net937[3], net937[4], net937[5], net937[6],
     net937[7], net937[8], net937[9], net937[10], net937[11],
     net937[12], net937[13], net937[14], net937[15]}),
     .sp4_h_l(SP4_h_l_03[47:0]), .sp12_h_l(SP12_h_l_03[23:0]),
     .prog(prog), .spi_ss_in_b({net1009[0], net1009[1]}),
     .tnl_op(rgt_op_04[7:0]), .lft_op(rgt_op_03[7:0]),
     .bnl_op(rgt_op_02[7:0]), .pgate(pgate[47:32]),
     .reset(reset_b[47:32]), .sp4_v_b({net865[0], net865[1], net865[2],
     net865[3], net865[4], net865[5], net865[6], net865[7], net865[8],
     net865[9], net865[10], net865[11], net865[12], net865[13],
     net865[14], net865[15]}), .wl(wl[47:32]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(net955));
io_col4_lft_ice8p_v2 I_io_00_04 ( .cbit_colcntl(colbuf_cntl_b[7:0]),
     .ceb(ceb), .sdo(net923), .sdi(net959), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode),
     .shift(shift), .hiz_b(hiz_b), .r(r), .bs_en(bs_en), .tclk(tclk_o),
     .update(update), .padin(padin[5:4]), .pado(pado[5:4]),
     .padeb(padeb[5:4]), .sp4_v_t({net973[0], net973[1], net973[2],
     net973[3], net973[4], net973[5], net973[6], net973[7], net973[8],
     net973[9], net973[10], net973[11], net973[12], net973[13],
     net973[14], net973[15]}), .sp4_h_l(SP4_h_l_04[47:0]),
     .sp12_h_l(SP12_h_l_04[23:0]), .prog(prog),
     .spi_ss_in_b({net1002[0], net1002[1]}), .tnl_op(rgt_op_05[7:0]),
     .lft_op(rgt_op_04[7:0]), .bnl_op(rgt_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]), .sp4_v_b({net937[0],
     net937[1], net937[2], net937[3], net937[4], net937[5], net937[6],
     net937[7], net937[8], net937[9], net937[10], net937[11],
     net937[12], net937[13], net937[14], net937[15]}), .wl(wl[63:48]),
     .cf(cf_l[95:72]), .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk_b[7:0]),
     .hold(hold), .fabric_out(fo_dlyadj[0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_bot (
     .colbuf_cntl(colbuf_cntl_b[7:0]), .col_clk(glb_netwk_b[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_colbuf12kx8_top (
     .colbuf_cntl(colbuf_cntl_t[7:0]), .col_clk(glb_netwk_t[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - ice1chip, Cell - io_bot_lft_1x6_ice1f, View - schematic
// LAST TIME SAVED: May  3 11:55:27 2011
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module io_bot_lft_1x6_ice1f ( bs_en_o, ceb_o, cf_bot_l[143:0],
     fabric_out_05_00, fabric_out_06_00, fo_bypass, fo_reset, fo_sck,
     fo_sdi, hiz_b_o, mode_o, padeb_b_l[10:0], padeb_b_l[12],
     pado_b_l[10:0], pado_b_l[12], r_o, sdo, shift_o,
     slf_op_01_00[3:0], slf_op_02_00[3:0], slf_op_03_00[3:0],
     slf_op_04_00[3:0], slf_op_05_00[3:0], slf_op_06_00[3:0], tclk_o,
     update_o, bl_01[53:0], bl_02[53:0], bl_03[41:0], bl_04[53:0],
     bl_05[53:0], bl_06[53:0], sp4_h_l_01_00[15:0],
     sp4_h_r_06_00[15:0], sp4_v_b_01_00[47:0], sp4_v_b_02_00[47:0],
     sp4_v_b_03_00[47:0], sp4_v_b_04_00[47:0], sp4_v_b_05_00[47:0],
     sp4_v_b_06_00[47:0], sp12_v_b_01_00[23:0], sp12_v_b_02_00[23:0],
     sp12_v_b_03_00[23:0], sp12_v_b_04_00[23:0], sp12_v_b_05_00[23:0],
     sp12_v_b_06_00[23:0], bnl_op_01_00[7:0], bs_en_i, ceb_i,
     glb_net_01[7:0], glb_net_02[7:0], glb_net_03[7:0],
     glb_net_04[7:0], glb_net_05[7:0], glb_net_06[7:0], hiz_b_i,
     hold_b_l, lft_op_01_00[7:0], lft_op_02_00[7:0], lft_op_03_00[7:0],
     lft_op_04_00[7:0], lft_op_05_00[7:0], lft_op_06_00[7:0], mode_i,
     padin_b_l[10:0], padin_b_l[12], pgate_l[15:0], prog, r_i,
     reset_l[15:0], sdi, shift_i, tclk_i, tnr_op_06_00[7:0], update_i,
     vdd_cntl_l[15:0], wl_l[15:0] );
output  bs_en_o, ceb_o, fabric_out_05_00, fabric_out_06_00, fo_bypass,
     fo_reset, fo_sck, fo_sdi, hiz_b_o, mode_o, r_o, sdo, shift_o,
     tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_02_00;
output [3:0]  slf_op_04_00;
output [3:0]  slf_op_06_00;
output [3:0]  slf_op_01_00;
output [12:0]  pado_b_l;
output [12:0]  padeb_b_l;
output [3:0]  slf_op_05_00;
output [143:0]  cf_bot_l;
output [3:0]  slf_op_03_00;

inout [47:0]  sp4_v_b_02_00;
inout [23:0]  sp12_v_b_02_00;
inout [23:0]  sp12_v_b_06_00;
inout [47:0]  sp4_v_b_03_00;
inout [23:0]  sp12_v_b_03_00;
inout [23:0]  sp12_v_b_01_00;
inout [47:0]  sp4_v_b_04_00;
inout [53:0]  bl_02;
inout [15:0]  sp4_h_l_01_00;
inout [47:0]  sp4_v_b_06_00;
inout [47:0]  sp4_v_b_01_00;
inout [41:0]  bl_03;
inout [23:0]  sp12_v_b_04_00;
inout [15:0]  sp4_h_r_06_00;
inout [53:0]  bl_04;
inout [47:0]  sp4_v_b_05_00;
inout [53:0]  bl_01;
inout [53:0]  bl_05;
inout [23:0]  sp12_v_b_05_00;
inout [53:0]  bl_06;

input [15:0]  pgate_l;
input [7:0]  lft_op_02_00;
input [7:0]  lft_op_06_00;
input [15:0]  wl_l;
input [7:0]  tnr_op_06_00;
input [7:0]  glb_net_01;
input [7:0]  lft_op_04_00;
input [7:0]  lft_op_03_00;
input [7:0]  bnl_op_01_00;
input [15:0]  reset_l;
input [7:0]  glb_net_05;
input [7:0]  glb_net_03;
input [7:0]  glb_net_06;
input [7:0]  lft_op_01_00;
input [12:0]  padin_b_l;
input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_04;
input [7:0]  glb_net_02;
input [7:0]  lft_op_05_00;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net519;

wire  [1:0]  net312;

wire  [1:0]  net520;

wire  [1:0]  net452;

wire  [1:0]  net487;

wire  [15:0]  net483;

wire  [15:0]  net308;

wire  [15:0]  net343;

wire  [15:0]  net413;

wire  [15:0]  net378;

wire  [1:0]  net382;



scan_buf_ice8p I_scanbuf_bl ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(update_o), .tclk_o(net284), .shift_o(shift_o),
     .sdo(net286), .r_o(r_o), .mode_o(mode_o), .hiz_b_o(hiz_b_o),
     .ceb_o(ceb_o), .bs_en_o(bs_en_o));
io_col4_bot_ice8p I_IO_02_00 ( .sdo(net292), .sdi(net362),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net378[0], net378[1], net378[2], net378[3],
     net378[4], net378[5], net378[6], net378[7], net378[8], net378[9],
     net378[10], net378[11], net378[12], net378[13], net378[14],
     net378[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_b_l[3:2]), .pado(pado_b_l[3:2]),
     .padeb(padeb_b_l[3:2]), .sp4_v_b({net308[0], net308[1], net308[2],
     net308[3], net308[4], net308[5], net308[6], net308[7], net308[8],
     net308[9], net308[10], net308[11], net308[12], net308[13],
     net308[14], net308[15]}), .sp4_h_l(sp4_v_b_02_00[47:0]),
     .sp12_h_l(sp12_v_b_02_00[23:0]), .prog(prog),
     .spi_ss_in_b({net312[0], net312[1]}), .tnl_op(lft_op_01_00[7:0]),
     .lft_op(lft_op_02_00[7:0]), .bnl_op(lft_op_03_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_02[5],
     bl_02[4], bl_02[37], bl_02[36], bl_02[35], bl_02[34], bl_02[33],
     bl_02[32], bl_02[14], bl_02[20], bl_02[19], bl_02[18], bl_02[17],
     bl_02[16], bl_02[27], bl_02[26], bl_02[25], bl_02[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[47:24]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_02_00[3:0]),
     .glb_netwk(glb_net_02[7:0]), .hold(hold_b_l),
     .fabric_out(fo_reset));
io_col4_bot_ice8p I_IO_03_00_bram ( .sdo(net327), .sdi(net292),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net308[0], net308[1], net308[2], net308[3],
     net308[4], net308[5], net308[6], net308[7], net308[8], net308[9],
     net308[10], net308[11], net308[12], net308[13], net308[14],
     net308[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_b_l[5:4]), .pado(pado_b_l[5:4]),
     .padeb(padeb_b_l[5:4]), .sp4_v_b({net343[0], net343[1], net343[2],
     net343[3], net343[4], net343[5], net343[6], net343[7], net343[8],
     net343[9], net343[10], net343[11], net343[12], net343[13],
     net343[14], net343[15]}), .sp4_h_l(sp4_v_b_03_00[47:0]),
     .sp12_h_l(sp12_v_b_03_00[23:0]), .prog(prog),
     .spi_ss_in_b({net519[0], net519[1]}), .tnl_op(lft_op_02_00[7:0]),
     .lft_op(lft_op_03_00[7:0]), .bnl_op(lft_op_04_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_03[5],
     bl_03[4], bl_03[37], bl_03[36], bl_03[35], bl_03[34], bl_03[33],
     bl_03[32], bl_03[14], bl_03[20], bl_03[19], bl_03[18], bl_03[17],
     bl_03[16], bl_03[27], bl_03[26], bl_03[25], bl_03[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[71:48]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_03_00[3:0]),
     .glb_netwk(glb_net_03[7:0]), .hold(hold_b_l),
     .fabric_out(fo_sck));
io_col4_bot_ice8p I_IO_01_00 ( .sdo(net362), .sdi(net286),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t(sp4_h_l_01_00[15:0]), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b_l[1:0]),
     .pado(pado_b_l[1:0]), .padeb(padeb_b_l[1:0]), .sp4_v_b({net378[0],
     net378[1], net378[2], net378[3], net378[4], net378[5], net378[6],
     net378[7], net378[8], net378[9], net378[10], net378[11],
     net378[12], net378[13], net378[14], net378[15]}),
     .sp4_h_l(sp4_v_b_01_00[47:0]), .sp12_h_l(sp12_v_b_01_00[23:0]),
     .prog(prog), .spi_ss_in_b({net382[0], net382[1]}),
     .tnl_op(bnl_op_01_00[7:0]), .lft_op(lft_op_01_00[7:0]),
     .bnl_op(lft_op_02_00[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .bl({bl_01[5], bl_01[4], bl_01[37],
     bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32], bl_01[14],
     bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16], bl_01[27],
     bl_01[26], bl_01[25], bl_01[23]}), .wl(wl_l[15:0]),
     .cf(cf_bot_l[23:0]), .ceb(ceb_o), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_00[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_b_l), .fabric_out(fo_bypass));
io_col4_bot_ice8p I_IO_05_00 ( .sdo(net397), .sdi(net467),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net483[0], net483[1], net483[2], net483[3],
     net483[4], net483[5], net483[6], net483[7], net483[8], net483[9],
     net483[10], net483[11], net483[12], net483[13], net483[14],
     net483[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_b_l[9:8]), .pado(pado_b_l[9:8]),
     .padeb(padeb_b_l[9:8]), .sp4_v_b({net413[0], net413[1], net413[2],
     net413[3], net413[4], net413[5], net413[6], net413[7], net413[8],
     net413[9], net413[10], net413[11], net413[12], net413[13],
     net413[14], net413[15]}), .sp4_h_l(sp4_v_b_05_00[47:0]),
     .sp12_h_l(sp12_v_b_05_00[23:0]), .prog(prog),
     .spi_ss_in_b({net520[0], net520[1]}), .tnl_op(lft_op_04_00[7:0]),
     .lft_op(lft_op_05_00[7:0]), .bnl_op(lft_op_06_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_05[5],
     bl_05[4], bl_05[37], bl_05[36], bl_05[35], bl_05[34], bl_05[33],
     bl_05[32], bl_05[14], bl_05[20], bl_05[19], bl_05[18], bl_05[17],
     bl_05[16], bl_05[27], bl_05[26], bl_05[25], bl_05[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[119:96]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_05_00[3:0]),
     .glb_netwk(glb_net_05[7:0]), .hold(hold_b_l),
     .fabric_out(fabric_out_05_00));
io_col4_bot_ice8p I_IO_06_00 ( .sdo(sdo), .sdi(net397),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net413[0], net413[1], net413[2], net413[3],
     net413[4], net413[5], net413[6], net413[7], net413[8], net413[9],
     net413[10], net413[11], net413[12], net413[13], net413[14],
     net413[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin({padin_b_l[10], padin_b_l[12]}), .pado({pado_b_l[10],
     pado_b_l[12]}), .padeb({padeb_b_l[10], padeb_b_l[12]}),
     .sp4_v_b(sp4_h_r_06_00[15:0]), .sp4_h_l(sp4_v_b_06_00[47:0]),
     .sp12_h_l(sp12_v_b_06_00[23:0]), .prog(prog),
     .spi_ss_in_b({net452[0], net452[1]}), .tnl_op(lft_op_05_00[7:0]),
     .lft_op(lft_op_06_00[7:0]), .bnl_op(tnr_op_06_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_06[5],
     bl_06[4], bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33],
     bl_06[32], bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17],
     bl_06[16], bl_06[27], bl_06[26], bl_06[25], bl_06[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[143:120]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_06_00[3:0]),
     .glb_netwk(glb_net_06[7:0]), .hold(hold_b_l),
     .fabric_out(fabric_out_06_00));
io_col4_bot_ice8p I_IO_04_00 ( .sdo(net467), .sdi(net327),
     .spiout({tielow, tielow}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .sp4_v_t({net343[0], net343[1], net343[2], net343[3],
     net343[4], net343[5], net343[6], net343[7], net343[8], net343[9],
     net343[10], net343[11], net343[12], net343[13], net343[14],
     net343[15]}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_b_l[7:6]), .pado(pado_b_l[7:6]),
     .padeb(padeb_b_l[7:6]), .sp4_v_b({net483[0], net483[1], net483[2],
     net483[3], net483[4], net483[5], net483[6], net483[7], net483[8],
     net483[9], net483[10], net483[11], net483[12], net483[13],
     net483[14], net483[15]}), .sp4_h_l(sp4_v_b_04_00[47:0]),
     .sp12_h_l(sp12_v_b_04_00[23:0]), .prog(prog),
     .spi_ss_in_b({net487[0], net487[1]}), .tnl_op(lft_op_03_00[7:0]),
     .lft_op(lft_op_04_00[7:0]), .bnl_op(lft_op_05_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .bl({bl_04[5],
     bl_04[4], bl_04[37], bl_04[36], bl_04[35], bl_04[34], bl_04[33],
     bl_04[32], bl_04[14], bl_04[20], bl_04[19], bl_04[18], bl_04[17],
     bl_04[16], bl_04[27], bl_04[26], bl_04[25], bl_04[23]}),
     .wl(wl_l[15:0]), .cf(cf_bot_l[95:72]), .ceb(ceb_o),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_04_00[3:0]),
     .glb_netwk(glb_net_04[7:0]), .hold(hold_b_l),
     .fabric_out(fo_sdi));
tckbufx32_ice8p I354 ( .in(net284), .out(tclk_o));
tiehi4x I482 ( .tiehi(tievdd));
tielo4x I483 ( .tielo(tielow));

endmodule
// Library - ice1chip, Cell - quad_bl_ice1, View - schematic
// LAST TIME SAVED: May  3 11:44:07 2011
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module quad_bl_ice1 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o[7:0],
     bm_sclk_o, bm_sclkrw_o[1:0], bm_sdi_o[1:0], bm_sdo_o[1:0],
     bm_sreb_o, bm_sweb_o[1:0], bm_wdummymux_en_o, bs_en_o,
     carry_out_01_08, carry_out_02_08, carry_out_04_08,
     carry_out_05_08, carry_out_06_08, ceb_o, cf_b_l[143:0],
     cf_l[191:0], fabric_out_00_07, fabric_out_00_08, fabric_out_05_00,
     fabric_out_06_00, fo_bypass, fo_dlyadj[2:0], fo_fb, fo_ref,
     fo_reset, fo_sck, fo_sdi, hiz_b_o, mode_o, op_vic_01_08,
     op_vic_02_08, op_vic_04_08, op_vic_05_08, op_vic_06_08,
     padeb_b_l[10:0], padeb_b_l[12], padeb_l_b[11:0], padin_00_08,
     padin_06_00, pado_b_l[10:0], pado_b_l[12], pado_l_b[11:0], r_o,
     sdo, shift_o, slf_op_00_08[3:0], slf_op_01_08[7:0],
     slf_op_02_08[7:0], slf_op_03_08[7:0], slf_op_04_08[7:0],
     slf_op_05_08[7:0], slf_op_06_00[3:0], slf_op_06_01[7:0],
     slf_op_06_02[7:0], slf_op_06_03[7:0], slf_op_06_04[7:0],
     slf_op_06_05[7:0], slf_op_06_06[7:0], slf_op_06_07[7:0],
     slf_op_06_08[7:0], tclk_o, update_o, bl[329:0], pgate_l[143:0],
     reset_b_l[143:0], sp4_h_r_06_00[15:0], sp4_h_r_06_01[47:0],
     sp4_h_r_06_02[47:0], sp4_h_r_06_03[47:0], sp4_h_r_06_04[47:0],
     sp4_h_r_06_05[47:0], sp4_h_r_06_06[47:0], sp4_h_r_06_07[47:0],
     sp4_h_r_06_08[47:0], sp4_r_v_b_06_01[47:0], sp4_r_v_b_06_02[47:0],
     sp4_r_v_b_06_03[47:0], sp4_r_v_b_06_04[47:0],
     sp4_r_v_b_06_05[47:0], sp4_r_v_b_06_06[47:0],
     sp4_r_v_b_06_07[47:0], sp4_r_v_b_06_08[47:0], sp4_v_t_00_08[15:0],
     sp4_v_t_01_08[47:0], sp4_v_t_02_08[47:0], sp4_v_t_03_08[47:0],
     sp4_v_t_04_08[47:0], sp4_v_t_05_08[47:0], sp4_v_t_06_08[47:0],
     sp12_h_r_06_01[23:0], sp12_h_r_06_02[23:0], sp12_h_r_06_03[23:0],
     sp12_h_r_06_04[23:0], sp12_h_r_06_05[23:0], sp12_h_r_06_06[23:0],
     sp12_h_r_06_07[23:0], sp12_h_r_06_08[23:0], sp12_v_t_01_08[23:0],
     sp12_v_t_02_08[23:0], sp12_v_t_03_08[23:0], sp12_v_t_04_08[23:0],
     sp12_v_t_05_08[23:0], sp12_v_t_06_08[23:0], vdd_cntl_l[143:0],
     wl_l[143:0], bm_aa_top[10:0], bm_ab_top[10:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i[1:0],
     bm_sdi_i[1:0], bm_sdo_i[1:0], bm_sreb_i, bm_sweb_i[1:0],
     bm_wdummymux_en_i, bnr_op_06_01[3:0], bs_en_i, ceb_i, glb_in[7:0],
     hiz_b_i, hold_b_l, hold_l_b, jtag_rowtest_mode_rowu0_b,
     last_rsr[0], mode_i, padin_b_l[10:0], padin_b_l[12],
     padin_l_b[11:0], pll_lock_out, prog, purst, r_i,
     rgt_op_06_01[7:0], rgt_op_06_02[7:0], rgt_op_06_03[7:0],
     rgt_op_06_04[7:0], rgt_op_06_05[7:0], rgt_op_06_06[7:0],
     rgt_op_06_07[7:0], rgt_op_06_08[7:0], sdi, shift_i, tclk_i,
     tnl_op_01_08[7:0], tnl_op_02_08[7:0], tnl_op_03_08[7:0],
     tnl_op_04_08[7:0], tnl_op_05_08[7:0], tnl_op_06_08[7:0],
     tnr_op_00_08[7:0], tnr_op_01_08[7:0], tnr_op_02_08[7:0],
     tnr_op_03_08[7:0], tnr_op_04_08[7:0], tnr_op_05_08[7:0],
     tnr_op_06_08[7:0], top_op_01_08[7:0], top_op_02_08[7:0],
     top_op_03_08[7:0], top_op_04_08[7:0], top_op_05_08[7:0],
     top_op_06_08[7:0], update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_08, carry_out_02_08,
     carry_out_04_08, carry_out_05_08, carry_out_06_08, ceb_o,
     fabric_out_00_07, fabric_out_00_08, fabric_out_05_00,
     fabric_out_06_00, fo_bypass, fo_fb, fo_ref, fo_reset, fo_sck,
     fo_sdi, hiz_b_o, mode_o, op_vic_01_08, op_vic_02_08, op_vic_04_08,
     op_vic_05_08, op_vic_06_08, padin_00_08, padin_06_00, r_o, sdo,
     shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, ceb_i, hiz_b_i, hold_b_l, hold_l_b,
     jtag_rowtest_mode_rowu0_b, mode_i, pll_lock_out, prog, purst, r_i,
     sdi, shift_i, tclk_i, update_i;

output [7:0]  slf_op_06_02;
output [7:0]  slf_op_06_08;
output [7:0]  slf_op_06_05;
output [11:0]  pado_l_b;
output [7:0]  slf_op_06_07;
output [191:0]  cf_l;
output [3:0]  slf_op_06_00;
output [3:0]  slf_op_00_08;
output [11:0]  padeb_l_b;
output [7:0]  slf_op_05_08;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_01_08;
output [12:0]  padeb_b_l;
output [12:0]  pado_b_l;
output [7:0]  slf_op_06_06;
output [7:0]  slf_op_03_08;
output [7:0]  slf_op_06_03;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_06_01;
output [7:0]  slf_op_04_08;
output [7:0]  slf_op_02_08;
output [1:0]  bm_sclkrw_o;
output [143:0]  cf_b_l;
output [7:0]  slf_op_06_04;
output [2:0]  fo_dlyadj;
output [1:0]  bm_sweb_o;

inout [47:0]  sp4_h_r_06_03;
inout [47:0]  sp4_v_t_06_08;
inout [47:0]  sp4_h_r_06_06;
inout [47:0]  sp4_v_t_03_08;
inout [23:0]  sp12_v_t_03_08;
inout [47:0]  sp4_v_t_05_08;
inout [23:0]  sp12_v_t_06_08;
inout [47:0]  sp4_r_v_b_06_01;
inout [47:0]  sp4_r_v_b_06_02;
inout [47:0]  sp4_r_v_b_06_05;
inout [47:0]  sp4_v_t_02_08;
inout [23:0]  sp12_h_r_06_02;
inout [23:0]  sp12_h_r_06_01;
inout [23:0]  sp12_h_r_06_07;
inout [143:0]  reset_b_l;
inout [15:0]  sp4_h_r_06_00;
inout [47:0]  sp4_h_r_06_05;
inout [47:0]  sp4_h_r_06_04;
inout [47:0]  sp4_v_t_04_08;
inout [47:0]  sp4_v_t_01_08;
inout [23:0]  sp12_h_r_06_03;
inout [15:0]  sp4_v_t_00_08;
inout [143:0]  vdd_cntl_l;
inout [47:0]  sp4_r_v_b_06_06;
inout [23:0]  sp12_h_r_06_05;
inout [47:0]  sp4_h_r_06_02;
inout [47:0]  sp4_r_v_b_06_08;
inout [23:0]  sp12_h_r_06_04;
inout [23:0]  sp12_h_r_06_08;
inout [23:0]  sp12_v_t_04_08;
inout [143:0]  pgate_l;
inout [23:0]  sp12_h_r_06_06;
inout [47:0]  sp4_h_r_06_01;
inout [329:0]  bl;
inout [47:0]  sp4_r_v_b_06_03;
inout [23:0]  sp12_v_t_01_08;
inout [23:0]  sp12_v_t_05_08;
inout [47:0]  sp4_r_v_b_06_04;
inout [23:0]  sp12_v_t_02_08;
inout [47:0]  sp4_h_r_06_08;
inout [47:0]  sp4_r_v_b_06_07;
inout [143:0]  wl_l;
inout [47:0]  sp4_h_r_06_07;

input [7:0]  top_op_04_08;
input [7:0]  rgt_op_06_04;
input [7:0]  top_op_03_08;
input [7:0]  tnr_op_05_08;
input [1:0]  bm_sdi_i;
input [7:0]  tnr_op_01_08;
input [7:0]  top_op_01_08;
input [7:0]  top_op_05_08;
input [7:0]  rgt_op_06_08;
input [7:0]  tnr_op_02_08;
input [7:0]  rgt_op_06_02;
input [7:0]  rgt_op_06_07;
input [1:0]  bm_sdo_i;
input [7:0]  top_op_02_08;
input [0:0]  last_rsr;
input [7:0]  rgt_op_06_03;
input [7:0]  tnl_op_02_08;
input [7:0]  tnl_op_01_08;
input [11:0]  padin_l_b;
input [10:0]  bm_ab_top;
input [7:0]  tnr_op_04_08;
input [7:0]  tnr_op_06_08;
input [12:0]  padin_b_l;
input [7:0]  tnl_op_04_08;
input [10:0]  bm_aa_top;
input [1:0]  bm_sweb_i;
input [7:0]  tnr_op_00_08;
input [7:0]  bm_sa_i;
input [7:0]  top_op_06_08;
input [3:0]  bnr_op_06_01;
input [7:0]  rgt_op_06_06;
input [7:0]  rgt_op_06_01;
input [7:0]  tnl_op_06_08;
input [1:0]  bm_sclkrw_i;
input [7:0]  tnl_op_05_08;
input [7:0]  tnl_op_03_08;
input [7:0]  tnr_op_03_08;
input [7:0]  glb_in;
input [7:0]  rgt_op_06_05;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [47:0]  net1315;

wire  [47:0]  net1261;

wire  [7:0]  net1408;

wire  [47:0]  net1128;

wire  [47:0]  net1289;

wire  [47:0]  net1325;

wire  [47:0]  net776;

wire  [47:0]  net751;

wire  [47:0]  net1291;

wire  [7:0]  net1344;

wire  [47:0]  net1125;

wire  [23:0]  net1144;

wire  [7:0]  net1268;

wire  [7:0]  net981;

wire  [23:0]  net1095;

wire  [23:0]  net1236;

wire  [23:0]  net1051;

wire  [47:0]  net1106;

wire  [23:0]  net813;

wire  [7:0]  net1040;

wire  [7:0]  net1355;

wire  [47:0]  net728;

wire  [7:0]  net1385;

wire  [10:10]  padinlat_b_l;

wire  [23:0]  net769;

wire  [23:0]  net770;

wire  [23:0]  net1212;

wire  [11:11]  padinlat_l_b;

wire  [47:0]  net1304;

wire  [3:0]  slf_op_00_01;

wire  [7:0]  net760;

wire  [7:0]  clk_center;

wire  [47:0]  net774;

wire  [47:0]  net1321;

wire  [10:0]  net1257;

wire  [3:0]  slf_op_02_00;

wire  [47:0]  net1290;

wire  [3:0]  slf_op_03_00;

wire  [3:0]  slf_op_01_00;

wire  [47:0]  net1260;

wire  [47:0]  net872;

wire  [47:0]  net868;

wire  [7:0]  net1388;

wire  [47:0]  net1402;

wire  [7:0]  net1328;

wire  [23:0]  net1003;

wire  [23:0]  net1145;

wire  [23:0]  net1050;

wire  [47:0]  net1440;

wire  [47:0]  net835;

wire  [47:0]  net730;

wire  [7:0]  net700;

wire  [7:0]  net1384;

wire  [47:0]  net1437;

wire  [47:0]  net1152;

wire  [47:0]  net1149;

wire  [3:0]  slf_op_00_06;

wire  [3:0]  slf_op_00_05;

wire  [3:0]  slf_op_00_07;

wire  [3:0]  slf_op_00_03;

wire  [23:0]  net1146;

wire  [3:0]  slf_op_00_02;

wire  [23:0]  net1404;

wire  [3:0]  slf_op_00_04;

wire  [7:0]  net1419;

wire  [47:0]  net1006;

wire  [7:0]  net1042;

wire  [3:0]  slf_op_05_00;

wire  [3:0]  slf_op_04_00;

wire  [23:0]  net719;

wire  [47:0]  net773;

wire  [47:0]  net1324;

wire  [23:0]  net1217;

wire  [47:0]  net845;

wire  [7:0]  net1383;

wire  [7:0]  net1041;

wire  [23:0]  net1342;

wire  [23:0]  net1413;

wire  [47:0]  net1032;

wire  [23:0]  net1096;

wire  [23:0]  net1097;

wire  [47:0]  net1287;

wire  [23:0]  net1147;

wire  [47:0]  net1436;

wire  [23:0]  net720;

wire  [7:0]  net1282;

wire  [47:0]  net1007;

wire  [23:0]  net771;

wire  [47:0]  net724;

wire  [23:0]  net1052;

wire  [23:0]  net815;

wire  [23:0]  net862;

wire  [47:0]  net844;

wire  [23:0]  net1345;

wire  [47:0]  net1151;

wire  [7:0]  net1410;

wire  [47:0]  net1414;

wire  [23:0]  net1407;

wire  [7:0]  net1269;

wire  [47:0]  net726;

wire  [23:0]  net1348;

wire  [47:0]  net846;

wire  [7:0]  net793;

wire  [7:0]  net708;

wire  [7:0]  net1409;

wire  [47:0]  net1105;

wire  [47:0]  net869;

wire  [47:0]  net1127;

wire  [7:0]  net1387;

wire  [47:0]  net1008;

wire  [7:0]  net1327;

wire  [47:0]  net1231;

wire  [23:0]  net812;

wire  [47:0]  net1228;

wire  [47:0]  net1411;

wire  [47:0]  net1013;

wire  [47:0]  net1031;

wire  [7:0]  net1265;

wire  [47:0]  net1227;

wire  [47:0]  net1323;

wire  [23:0]  net718;

wire  [47:0]  net843;

wire  [47:0]  net1058;

wire  [47:0]  net775;

wire  [23:0]  net768;

wire  [23:0]  net1341;

wire  [47:0]  net729;

wire  [47:0]  net867;

wire  [47:0]  net1101;

wire  [47:0]  net1056;

wire  [47:0]  net1104;

wire  [47:0]  net1055;

wire  [47:0]  net1150;

wire  [23:0]  net1214;

wire  [23:0]  net864;

wire  [23:0]  net865;

wire  [47:0]  net1100;

wire  [23:0]  net1350;

wire  [47:0]  net1011;

wire  [7:0]  net1266;

wire  [23:0]  net1001;

wire  [47:0]  net870;

wire  [7:0]  net795;

wire  [47:0]  net1288;

wire  [7:0]  net1329;

wire  [47:0]  net1435;

wire  [47:0]  net1286;

wire  [47:0]  net1010;

wire  [7:0]  net758;

wire  [47:0]  net752;

wire  [7:0]  net991;

wire  [7:0]  net803;

wire  [47:0]  net1012;

wire  [23:0]  net814;

wire  [7:0]  net853;

wire  [47:0]  net731;

wire  [7:0]  net698;

wire  [47:0]  net1126;

wire  [47:0]  net1412;

wire  [23:0]  net721;

wire  [23:0]  net1200;

wire  [47:0]  net824;

wire  [23:0]  net1340;

wire  [15:0]  net1311;

wire  [47:0]  net1326;

wire  [23:0]  net1216;

wire  [47:0]  net823;

wire  [7:0]  net1267;

wire  [23:0]  net1053;

wire  [47:0]  net1107;

wire  [47:0]  net1322;

wire  [23:0]  net1343;

wire  [23:0]  net1002;

wire  [23:0]  net1426;

wire  [7:0]  net759;

wire  [47:0]  net750;

wire  [7:0]  net1417;

wire  [7:0]  net983;

wire  [47:0]  net1406;

wire  [47:0]  net1430;

wire  [47:0]  net1102;

wire  [47:0]  net1242;

wire  [23:0]  net863;

wire  [47:0]  net819;

wire  [47:0]  net1057;

wire  [23:0]  net1000;

wire  [47:0]  net1220;

wire  [7:0]  net1386;

wire  [47:0]  net725;

wire  [47:0]  net825;

wire  [23:0]  net1390;

wire  [47:0]  net871;

wire  [47:0]  net818;

wire  [23:0]  net1373;

wire  [23:0]  net1094;

wire  [47:0]  net749;

wire  [7:0]  net852;

wire  [47:0]  net822;

wire  [47:0]  net1034;

wire  [47:0]  net1033;

wire  [47:0]  net820;

wire  [7:0]  net1264;

wire  [7:0]  net1330;

wire  [23:0]  net1244;

wire  [10:0]  net1256;

wire  [47:0]  net1259;

wire  [23:0]  net1245;

wire  [7:0]  net854;

wire  [7:0]  net1314;

wire  [47:0]  net1224;

wire  [23:0]  net1346;



bram1x4_ice1f I_bram_col_t03 ( .prog(prog), .glb_netwk_col({net1344[0],
     net1344[1], net1344[2], net1344[3], net1344[4], net1344[5],
     net1344[6], net1344[7]}), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .reset_b(reset_b_l[143:16]),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sreb_o(bm_sreb_o),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .lft_op_05({net854[0], net854[1],
     net854[2], net854[3], net854[4], net854[5], net854[6],
     net854[7]}), .bl(bl[167:126]), .sp4_h_l_06({net751[0], net751[1],
     net751[2], net751[3], net751[4], net751[5], net751[6], net751[7],
     net751[8], net751[9], net751[10], net751[11], net751[12],
     net751[13], net751[14], net751[15], net751[16], net751[17],
     net751[18], net751[19], net751[20], net751[21], net751[22],
     net751[23], net751[24], net751[25], net751[26], net751[27],
     net751[28], net751[29], net751[30], net751[31], net751[32],
     net751[33], net751[34], net751[35], net751[36], net751[37],
     net751[38], net751[39], net751[40], net751[41], net751[42],
     net751[43], net751[44], net751[45], net751[46], net751[47]}),
     .sp12_h_l_02({net720[0], net720[1], net720[2], net720[3],
     net720[4], net720[5], net720[6], net720[7], net720[8], net720[9],
     net720[10], net720[11], net720[12], net720[13], net720[14],
     net720[15], net720[16], net720[17], net720[18], net720[19],
     net720[20], net720[21], net720[22], net720[23]}),
     .lft_op_06({net853[0], net853[1], net853[2], net853[3], net853[4],
     net853[5], net853[6], net853[7]}), .sp12_h_l_03({net719[0],
     net719[1], net719[2], net719[3], net719[4], net719[5], net719[6],
     net719[7], net719[8], net719[9], net719[10], net719[11],
     net719[12], net719[13], net719[14], net719[15], net719[16],
     net719[17], net719[18], net719[19], net719[20], net719[21],
     net719[22], net719[23]}), .sp12_h_r_03({net1200[0], net1200[1],
     net1200[2], net1200[3], net1200[4], net1200[5], net1200[6],
     net1200[7], net1200[8], net1200[9], net1200[10], net1200[11],
     net1200[12], net1200[13], net1200[14], net1200[15], net1200[16],
     net1200[17], net1200[18], net1200[19], net1200[20], net1200[21],
     net1200[22], net1200[23]}), .sp12_h_l_01({net721[0], net721[1],
     net721[2], net721[3], net721[4], net721[5], net721[6], net721[7],
     net721[8], net721[9], net721[10], net721[11], net721[12],
     net721[13], net721[14], net721[15], net721[16], net721[17],
     net721[18], net721[19], net721[20], net721[21], net721[22],
     net721[23]}), .sp4_v_b_04({net724[0], net724[1], net724[2],
     net724[3], net724[4], net724[5], net724[6], net724[7], net724[8],
     net724[9], net724[10], net724[11], net724[12], net724[13],
     net724[14], net724[15], net724[16], net724[17], net724[18],
     net724[19], net724[20], net724[21], net724[22], net724[23],
     net724[24], net724[25], net724[26], net724[27], net724[28],
     net724[29], net724[30], net724[31], net724[32], net724[33],
     net724[34], net724[35], net724[36], net724[37], net724[38],
     net724[39], net724[40], net724[41], net724[42], net724[43],
     net724[44], net724[45], net724[46], net724[47]}),
     .sp4_v_b_05({net773[0], net773[1], net773[2], net773[3],
     net773[4], net773[5], net773[6], net773[7], net773[8], net773[9],
     net773[10], net773[11], net773[12], net773[13], net773[14],
     net773[15], net773[16], net773[17], net773[18], net773[19],
     net773[20], net773[21], net773[22], net773[23], net773[24],
     net773[25], net773[26], net773[27], net773[28], net773[29],
     net773[30], net773[31], net773[32], net773[33], net773[34],
     net773[35], net773[36], net773[37], net773[38], net773[39],
     net773[40], net773[41], net773[42], net773[43], net773[44],
     net773[45], net773[46], net773[47]}), .lft_op_07({net852[0],
     net852[1], net852[2], net852[3], net852[4], net852[5], net852[6],
     net852[7]}), .sp4_v_b_06({net774[0], net774[1], net774[2],
     net774[3], net774[4], net774[5], net774[6], net774[7], net774[8],
     net774[9], net774[10], net774[11], net774[12], net774[13],
     net774[14], net774[15], net774[16], net774[17], net774[18],
     net774[19], net774[20], net774[21], net774[22], net774[23],
     net774[24], net774[25], net774[26], net774[27], net774[28],
     net774[29], net774[30], net774[31], net774[32], net774[33],
     net774[34], net774[35], net774[36], net774[37], net774[38],
     net774[39], net774[40], net774[41], net774[42], net774[43],
     net774[44], net774[45], net774[46], net774[47]}),
     .sp4_v_b_08({net776[0], net776[1], net776[2], net776[3],
     net776[4], net776[5], net776[6], net776[7], net776[8], net776[9],
     net776[10], net776[11], net776[12], net776[13], net776[14],
     net776[15], net776[16], net776[17], net776[18], net776[19],
     net776[20], net776[21], net776[22], net776[23], net776[24],
     net776[25], net776[26], net776[27], net776[28], net776[29],
     net776[30], net776[31], net776[32], net776[33], net776[34],
     net776[35], net776[36], net776[37], net776[38], net776[39],
     net776[40], net776[41], net776[42], net776[43], net776[44],
     net776[45], net776[46], net776[47]}), .sp4_v_b_07({net775[0],
     net775[1], net775[2], net775[3], net775[4], net775[5], net775[6],
     net775[7], net775[8], net775[9], net775[10], net775[11],
     net775[12], net775[13], net775[14], net775[15], net775[16],
     net775[17], net775[18], net775[19], net775[20], net775[21],
     net775[22], net775[23], net775[24], net775[25], net775[26],
     net775[27], net775[28], net775[29], net775[30], net775[31],
     net775[32], net775[33], net775[34], net775[35], net775[36],
     net775[37], net775[38], net775[39], net775[40], net775[41],
     net775[42], net775[43], net775[44], net775[45], net775[46],
     net775[47]}), .lft_op_03({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7]}),
     .lft_op_01({net1419[0], net1419[1], net1419[2], net1419[3],
     net1419[4], net1419[5], net1419[6], net1419[7]}),
     .sp4_h_l_02({net730[0], net730[1], net730[2], net730[3],
     net730[4], net730[5], net730[6], net730[7], net730[8], net730[9],
     net730[10], net730[11], net730[12], net730[13], net730[14],
     net730[15], net730[16], net730[17], net730[18], net730[19],
     net730[20], net730[21], net730[22], net730[23], net730[24],
     net730[25], net730[26], net730[27], net730[28], net730[29],
     net730[30], net730[31], net730[32], net730[33], net730[34],
     net730[35], net730[36], net730[37], net730[38], net730[39],
     net730[40], net730[41], net730[42], net730[43], net730[44],
     net730[45], net730[46], net730[47]}), .sp12_h_l_06({net769[0],
     net769[1], net769[2], net769[3], net769[4], net769[5], net769[6],
     net769[7], net769[8], net769[9], net769[10], net769[11],
     net769[12], net769[13], net769[14], net769[15], net769[16],
     net769[17], net769[18], net769[19], net769[20], net769[21],
     net769[22], net769[23]}), .sp12_h_r_07({net1212[0], net1212[1],
     net1212[2], net1212[3], net1212[4], net1212[5], net1212[6],
     net1212[7], net1212[8], net1212[9], net1212[10], net1212[11],
     net1212[12], net1212[13], net1212[14], net1212[15], net1212[16],
     net1212[17], net1212[18], net1212[19], net1212[20], net1212[21],
     net1212[22], net1212[23]}), .sp12_h_l_05({net768[0], net768[1],
     net768[2], net768[3], net768[4], net768[5], net768[6], net768[7],
     net768[8], net768[9], net768[10], net768[11], net768[12],
     net768[13], net768[14], net768[15], net768[16], net768[17],
     net768[18], net768[19], net768[20], net768[21], net768[22],
     net768[23]}), .sp12_h_r_06({net1214[0], net1214[1], net1214[2],
     net1214[3], net1214[4], net1214[5], net1214[6], net1214[7],
     net1214[8], net1214[9], net1214[10], net1214[11], net1214[12],
     net1214[13], net1214[14], net1214[15], net1214[16], net1214[17],
     net1214[18], net1214[19], net1214[20], net1214[21], net1214[22],
     net1214[23]}), .sp12_h_l_04({net718[0], net718[1], net718[2],
     net718[3], net718[4], net718[5], net718[6], net718[7], net718[8],
     net718[9], net718[10], net718[11], net718[12], net718[13],
     net718[14], net718[15], net718[16], net718[17], net718[18],
     net718[19], net718[20], net718[21], net718[22], net718[23]}),
     .sp12_h_r_05({net1216[0], net1216[1], net1216[2], net1216[3],
     net1216[4], net1216[5], net1216[6], net1216[7], net1216[8],
     net1216[9], net1216[10], net1216[11], net1216[12], net1216[13],
     net1216[14], net1216[15], net1216[16], net1216[17], net1216[18],
     net1216[19], net1216[20], net1216[21], net1216[22], net1216[23]}),
     .sp12_h_r_08({net1217[0], net1217[1], net1217[2], net1217[3],
     net1217[4], net1217[5], net1217[6], net1217[7], net1217[8],
     net1217[9], net1217[10], net1217[11], net1217[12], net1217[13],
     net1217[14], net1217[15], net1217[16], net1217[17], net1217[18],
     net1217[19], net1217[20], net1217[21], net1217[22], net1217[23]}),
     .sp12_h_l_07({net770[0], net770[1], net770[2], net770[3],
     net770[4], net770[5], net770[6], net770[7], net770[8], net770[9],
     net770[10], net770[11], net770[12], net770[13], net770[14],
     net770[15], net770[16], net770[17], net770[18], net770[19],
     net770[20], net770[21], net770[22], net770[23]}),
     .sp12_h_l_08({net771[0], net771[1], net771[2], net771[3],
     net771[4], net771[5], net771[6], net771[7], net771[8], net771[9],
     net771[10], net771[11], net771[12], net771[13], net771[14],
     net771[15], net771[16], net771[17], net771[18], net771[19],
     net771[20], net771[21], net771[22], net771[23]}),
     .sp4_r_v_b_03({net1220[0], net1220[1], net1220[2], net1220[3],
     net1220[4], net1220[5], net1220[6], net1220[7], net1220[8],
     net1220[9], net1220[10], net1220[11], net1220[12], net1220[13],
     net1220[14], net1220[15], net1220[16], net1220[17], net1220[18],
     net1220[19], net1220[20], net1220[21], net1220[22], net1220[23],
     net1220[24], net1220[25], net1220[26], net1220[27], net1220[28],
     net1220[29], net1220[30], net1220[31], net1220[32], net1220[33],
     net1220[34], net1220[35], net1220[36], net1220[37], net1220[38],
     net1220[39], net1220[40], net1220[41], net1220[42], net1220[43],
     net1220[44], net1220[45], net1220[46], net1220[47]}),
     .vdd_cntl(vdd_cntl_l[143:16]), .pgate(pgate_l[143:16]),
     .bot_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .sp4_r_v_b_04({net1224[0],
     net1224[1], net1224[2], net1224[3], net1224[4], net1224[5],
     net1224[6], net1224[7], net1224[8], net1224[9], net1224[10],
     net1224[11], net1224[12], net1224[13], net1224[14], net1224[15],
     net1224[16], net1224[17], net1224[18], net1224[19], net1224[20],
     net1224[21], net1224[22], net1224[23], net1224[24], net1224[25],
     net1224[26], net1224[27], net1224[28], net1224[29], net1224[30],
     net1224[31], net1224[32], net1224[33], net1224[34], net1224[35],
     net1224[36], net1224[37], net1224[38], net1224[39], net1224[40],
     net1224[41], net1224[42], net1224[43], net1224[44], net1224[45],
     net1224[46], net1224[47]}), .sp4_v_b_01({net1412[0], net1412[1],
     net1412[2], net1412[3], net1412[4], net1412[5], net1412[6],
     net1412[7], net1412[8], net1412[9], net1412[10], net1412[11],
     net1412[12], net1412[13], net1412[14], net1412[15], net1412[16],
     net1412[17], net1412[18], net1412[19], net1412[20], net1412[21],
     net1412[22], net1412[23], net1412[24], net1412[25], net1412[26],
     net1412[27], net1412[28], net1412[29], net1412[30], net1412[31],
     net1412[32], net1412[33], net1412[34], net1412[35], net1412[36],
     net1412[37], net1412[38], net1412[39], net1412[40], net1412[41],
     net1412[42], net1412[43], net1412[44], net1412[45], net1412[46],
     net1412[47]}), .sp4_v_b_03({net725[0], net725[1], net725[2],
     net725[3], net725[4], net725[5], net725[6], net725[7], net725[8],
     net725[9], net725[10], net725[11], net725[12], net725[13],
     net725[14], net725[15], net725[16], net725[17], net725[18],
     net725[19], net725[20], net725[21], net725[22], net725[23],
     net725[24], net725[25], net725[26], net725[27], net725[28],
     net725[29], net725[30], net725[31], net725[32], net725[33],
     net725[34], net725[35], net725[36], net725[37], net725[38],
     net725[39], net725[40], net725[41], net725[42], net725[43],
     net725[44], net725[45], net725[46], net725[47]}),
     .sp4_h_r_08({net1227[0], net1227[1], net1227[2], net1227[3],
     net1227[4], net1227[5], net1227[6], net1227[7], net1227[8],
     net1227[9], net1227[10], net1227[11], net1227[12], net1227[13],
     net1227[14], net1227[15], net1227[16], net1227[17], net1227[18],
     net1227[19], net1227[20], net1227[21], net1227[22], net1227[23],
     net1227[24], net1227[25], net1227[26], net1227[27], net1227[28],
     net1227[29], net1227[30], net1227[31], net1227[32], net1227[33],
     net1227[34], net1227[35], net1227[36], net1227[37], net1227[38],
     net1227[39], net1227[40], net1227[41], net1227[42], net1227[43],
     net1227[44], net1227[45], net1227[46], net1227[47]}),
     .sp4_r_v_b_05({net1228[0], net1228[1], net1228[2], net1228[3],
     net1228[4], net1228[5], net1228[6], net1228[7], net1228[8],
     net1228[9], net1228[10], net1228[11], net1228[12], net1228[13],
     net1228[14], net1228[15], net1228[16], net1228[17], net1228[18],
     net1228[19], net1228[20], net1228[21], net1228[22], net1228[23],
     net1228[24], net1228[25], net1228[26], net1228[27], net1228[28],
     net1228[29], net1228[30], net1228[31], net1228[32], net1228[33],
     net1228[34], net1228[35], net1228[36], net1228[37], net1228[38],
     net1228[39], net1228[40], net1228[41], net1228[42], net1228[43],
     net1228[44], net1228[45], net1228[46], net1228[47]}),
     .sp4_v_b_02({net726[0], net726[1], net726[2], net726[3],
     net726[4], net726[5], net726[6], net726[7], net726[8], net726[9],
     net726[10], net726[11], net726[12], net726[13], net726[14],
     net726[15], net726[16], net726[17], net726[18], net726[19],
     net726[20], net726[21], net726[22], net726[23], net726[24],
     net726[25], net726[26], net726[27], net726[28], net726[29],
     net726[30], net726[31], net726[32], net726[33], net726[34],
     net726[35], net726[36], net726[37], net726[38], net726[39],
     net726[40], net726[41], net726[42], net726[43], net726[44],
     net726[45], net726[46], net726[47]}),
     .sp4_v_t_08(sp4_v_t_03_08[47:0]), .sp4_r_v_b_02({net1231[0],
     net1231[1], net1231[2], net1231[3], net1231[4], net1231[5],
     net1231[6], net1231[7], net1231[8], net1231[9], net1231[10],
     net1231[11], net1231[12], net1231[13], net1231[14], net1231[15],
     net1231[16], net1231[17], net1231[18], net1231[19], net1231[20],
     net1231[21], net1231[22], net1231[23], net1231[24], net1231[25],
     net1231[26], net1231[27], net1231[28], net1231[29], net1231[30],
     net1231[31], net1231[32], net1231[33], net1231[34], net1231[35],
     net1231[36], net1231[37], net1231[38], net1231[39], net1231[40],
     net1231[41], net1231[42], net1231[43], net1231[44], net1231[45],
     net1231[46], net1231[47]}), .bnr_op_01({slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0],
     slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0]}), .bm_sdi_o(bm_sdi_o[1:0]),
     .sp4_h_l_04({net728[0], net728[1], net728[2], net728[3],
     net728[4], net728[5], net728[6], net728[7], net728[8], net728[9],
     net728[10], net728[11], net728[12], net728[13], net728[14],
     net728[15], net728[16], net728[17], net728[18], net728[19],
     net728[20], net728[21], net728[22], net728[23], net728[24],
     net728[25], net728[26], net728[27], net728[28], net728[29],
     net728[30], net728[31], net728[32], net728[33], net728[34],
     net728[35], net728[36], net728[37], net728[38], net728[39],
     net728[40], net728[41], net728[42], net728[43], net728[44],
     net728[45], net728[46], net728[47]}),
     .lft_op_08(slf_op_02_08[7:0]), .sp12_h_r_01({net1236[0],
     net1236[1], net1236[2], net1236[3], net1236[4], net1236[5],
     net1236[6], net1236[7], net1236[8], net1236[9], net1236[10],
     net1236[11], net1236[12], net1236[13], net1236[14], net1236[15],
     net1236[16], net1236[17], net1236[18], net1236[19], net1236[20],
     net1236[21], net1236[22], net1236[23]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdo_o(bm_sdo_o[1:0]), .bm_sweb_o(bm_sweb_o[1:0]),
     .sp4_h_l_03({net729[0], net729[1], net729[2], net729[3],
     net729[4], net729[5], net729[6], net729[7], net729[8], net729[9],
     net729[10], net729[11], net729[12], net729[13], net729[14],
     net729[15], net729[16], net729[17], net729[18], net729[19],
     net729[20], net729[21], net729[22], net729[23], net729[24],
     net729[25], net729[26], net729[27], net729[28], net729[29],
     net729[30], net729[31], net729[32], net729[33], net729[34],
     net729[35], net729[36], net729[37], net729[38], net729[39],
     net729[40], net729[41], net729[42], net729[43], net729[44],
     net729[45], net729[46], net729[47]}), .sp4_h_l_01({net731[0],
     net731[1], net731[2], net731[3], net731[4], net731[5], net731[6],
     net731[7], net731[8], net731[9], net731[10], net731[11],
     net731[12], net731[13], net731[14], net731[15], net731[16],
     net731[17], net731[18], net731[19], net731[20], net731[21],
     net731[22], net731[23], net731[24], net731[25], net731[26],
     net731[27], net731[28], net731[29], net731[30], net731[31],
     net731[32], net731[33], net731[34], net731[35], net731[36],
     net731[37], net731[38], net731[39], net731[40], net731[41],
     net731[42], net731[43], net731[44], net731[45], net731[46],
     net731[47]}), .sp4_h_r_01({net1242[0], net1242[1], net1242[2],
     net1242[3], net1242[4], net1242[5], net1242[6], net1242[7],
     net1242[8], net1242[9], net1242[10], net1242[11], net1242[12],
     net1242[13], net1242[14], net1242[15], net1242[16], net1242[17],
     net1242[18], net1242[19], net1242[20], net1242[21], net1242[22],
     net1242[23], net1242[24], net1242[25], net1242[26], net1242[27],
     net1242[28], net1242[29], net1242[30], net1242[31], net1242[32],
     net1242[33], net1242[34], net1242[35], net1242[36], net1242[37],
     net1242[38], net1242[39], net1242[40], net1242[41], net1242[42],
     net1242[43], net1242[44], net1242[45], net1242[46], net1242[47]}),
     .tnr_op_08(tnr_op_03_08[7:0]), .sp12_h_r_02({net1244[0],
     net1244[1], net1244[2], net1244[3], net1244[4], net1244[5],
     net1244[6], net1244[7], net1244[8], net1244[9], net1244[10],
     net1244[11], net1244[12], net1244[13], net1244[14], net1244[15],
     net1244[16], net1244[17], net1244[18], net1244[19], net1244[20],
     net1244[21], net1244[22], net1244[23]}), .sp12_h_r_04({net1245[0],
     net1245[1], net1245[2], net1245[3], net1245[4], net1245[5],
     net1245[6], net1245[7], net1245[8], net1245[9], net1245[10],
     net1245[11], net1245[12], net1245[13], net1245[14], net1245[15],
     net1245[16], net1245[17], net1245[18], net1245[19], net1245[20],
     net1245[21], net1245[22], net1245[23]}),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .lft_op_02({net795[0], net795[1], net795[2], net795[3], net795[4],
     net795[5], net795[6], net795[7]}), .lft_op_04({net803[0],
     net803[1], net803[2], net803[3], net803[4], net803[5], net803[6],
     net803[7]}), .bm_sweb_i(bm_sweb_i[1:0]),
     .bnl_op_01({slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0], slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0]}),
     .sp12_v_t_08(sp12_v_t_03_08[23:0]), .wl(wl_l[143:16]),
     .tnl_op_08(tnl_op_03_08[7:0]), .top_op_08(top_op_03_08[7:0]),
     .bm_ab_2bot({net1256[0], net1256[1], net1256[2], net1256[3],
     net1256[4], net1256[5], net1256[6], net1256[7], net1256[8],
     net1256[9], net1256[10]}), .bm_aa_2bot({net1257[0], net1257[1],
     net1257[2], net1257[3], net1257[4], net1257[5], net1257[6],
     net1257[7], net1257[8], net1257[9], net1257[10]}),
     .sp12_v_b_01({net1413[0], net1413[1], net1413[2], net1413[3],
     net1413[4], net1413[5], net1413[6], net1413[7], net1413[8],
     net1413[9], net1413[10], net1413[11], net1413[12], net1413[13],
     net1413[14], net1413[15], net1413[16], net1413[17], net1413[18],
     net1413[19], net1413[20], net1413[21], net1413[22], net1413[23]}),
     .sp4_r_v_b_08({net1259[0], net1259[1], net1259[2], net1259[3],
     net1259[4], net1259[5], net1259[6], net1259[7], net1259[8],
     net1259[9], net1259[10], net1259[11], net1259[12], net1259[13],
     net1259[14], net1259[15], net1259[16], net1259[17], net1259[18],
     net1259[19], net1259[20], net1259[21], net1259[22], net1259[23],
     net1259[24], net1259[25], net1259[26], net1259[27], net1259[28],
     net1259[29], net1259[30], net1259[31], net1259[32], net1259[33],
     net1259[34], net1259[35], net1259[36], net1259[37], net1259[38],
     net1259[39], net1259[40], net1259[41], net1259[42], net1259[43],
     net1259[44], net1259[45], net1259[46], net1259[47]}),
     .sp4_r_v_b_07({net1260[0], net1260[1], net1260[2], net1260[3],
     net1260[4], net1260[5], net1260[6], net1260[7], net1260[8],
     net1260[9], net1260[10], net1260[11], net1260[12], net1260[13],
     net1260[14], net1260[15], net1260[16], net1260[17], net1260[18],
     net1260[19], net1260[20], net1260[21], net1260[22], net1260[23],
     net1260[24], net1260[25], net1260[26], net1260[27], net1260[28],
     net1260[29], net1260[30], net1260[31], net1260[32], net1260[33],
     net1260[34], net1260[35], net1260[36], net1260[37], net1260[38],
     net1260[39], net1260[40], net1260[41], net1260[42], net1260[43],
     net1260[44], net1260[45], net1260[46], net1260[47]}),
     .sp4_r_v_b_06({net1261[0], net1261[1], net1261[2], net1261[3],
     net1261[4], net1261[5], net1261[6], net1261[7], net1261[8],
     net1261[9], net1261[10], net1261[11], net1261[12], net1261[13],
     net1261[14], net1261[15], net1261[16], net1261[17], net1261[18],
     net1261[19], net1261[20], net1261[21], net1261[22], net1261[23],
     net1261[24], net1261[25], net1261[26], net1261[27], net1261[28],
     net1261[29], net1261[30], net1261[31], net1261[32], net1261[33],
     net1261[34], net1261[35], net1261[36], net1261[37], net1261[38],
     net1261[39], net1261[40], net1261[41], net1261[42], net1261[43],
     net1261[44], net1261[45], net1261[46], net1261[47]}),
     .sp4_r_v_b_01({net1414[0], net1414[1], net1414[2], net1414[3],
     net1414[4], net1414[5], net1414[6], net1414[7], net1414[8],
     net1414[9], net1414[10], net1414[11], net1414[12], net1414[13],
     net1414[14], net1414[15], net1414[16], net1414[17], net1414[18],
     net1414[19], net1414[20], net1414[21], net1414[22], net1414[23],
     net1414[24], net1414[25], net1414[26], net1414[27], net1414[28],
     net1414[29], net1414[30], net1414[31], net1414[32], net1414[33],
     net1414[34], net1414[35], net1414[36], net1414[37], net1414[38],
     net1414[39], net1414[40], net1414[41], net1414[42], net1414[43],
     net1414[44], net1414[45], net1414[46], net1414[47]}),
     .rgt_op_08(slf_op_04_08[7:0]), .rgt_op_07({net1264[0], net1264[1],
     net1264[2], net1264[3], net1264[4], net1264[5], net1264[6],
     net1264[7]}), .rgt_op_06({net1265[0], net1265[1], net1265[2],
     net1265[3], net1265[4], net1265[5], net1265[6], net1265[7]}),
     .rgt_op_05({net1266[0], net1266[1], net1266[2], net1266[3],
     net1266[4], net1266[5], net1266[6], net1266[7]}),
     .rgt_op_04({net1267[0], net1267[1], net1267[2], net1267[3],
     net1267[4], net1267[5], net1267[6], net1267[7]}),
     .rgt_op_03({net1268[0], net1268[1], net1268[2], net1268[3],
     net1268[4], net1268[5], net1268[6], net1268[7]}),
     .rgt_op_02({net1269[0], net1269[1], net1269[2], net1269[3],
     net1269[4], net1269[5], net1269[6], net1269[7]}),
     .rgt_op_01({net1408[0], net1408[1], net1408[2], net1408[3],
     net1408[4], net1408[5], net1408[6], net1408[7]}),
     .slf_op_02({net700[0], net700[1], net700[2], net700[3], net700[4],
     net700[5], net700[6], net700[7]}), .slf_op_01({net1410[0],
     net1410[1], net1410[2], net1410[3], net1410[4], net1410[5],
     net1410[6], net1410[7]}), .slf_op_03({net698[0], net698[1],
     net698[2], net698[3], net698[4], net698[5], net698[6],
     net698[7]}), .slf_op_04({net708[0], net708[1], net708[2],
     net708[3], net708[4], net708[5], net708[6], net708[7]}),
     .slf_op_05({net760[0], net760[1], net760[2], net760[3], net760[4],
     net760[5], net760[6], net760[7]}), .slf_op_06({net759[0],
     net759[1], net759[2], net759[3], net759[4], net759[5], net759[6],
     net759[7]}), .slf_op_07({net758[0], net758[1], net758[2],
     net758[3], net758[4], net758[5], net758[6], net758[7]}),
     .slf_op_08(slf_op_03_08[7:0]), .bm_ab_top(bm_ab_top[10:0]),
     .bm_aa_top(bm_aa_top[10:0]), .glb_netwk_bot({net1386[0],
     net1386[1], net1386[2], net1386[3], net1386[4], net1386[5],
     net1386[6], net1386[7]}), .glb_netwk_top({net1282[0], net1282[1],
     net1282[2], net1282[3], net1282[4], net1282[5], net1282[6],
     net1282[7]}), .sp4_h_l_08({net749[0], net749[1], net749[2],
     net749[3], net749[4], net749[5], net749[6], net749[7], net749[8],
     net749[9], net749[10], net749[11], net749[12], net749[13],
     net749[14], net749[15], net749[16], net749[17], net749[18],
     net749[19], net749[20], net749[21], net749[22], net749[23],
     net749[24], net749[25], net749[26], net749[27], net749[28],
     net749[29], net749[30], net749[31], net749[32], net749[33],
     net749[34], net749[35], net749[36], net749[37], net749[38],
     net749[39], net749[40], net749[41], net749[42], net749[43],
     net749[44], net749[45], net749[46], net749[47]}),
     .sp4_h_l_07({net750[0], net750[1], net750[2], net750[3],
     net750[4], net750[5], net750[6], net750[7], net750[8], net750[9],
     net750[10], net750[11], net750[12], net750[13], net750[14],
     net750[15], net750[16], net750[17], net750[18], net750[19],
     net750[20], net750[21], net750[22], net750[23], net750[24],
     net750[25], net750[26], net750[27], net750[28], net750[29],
     net750[30], net750[31], net750[32], net750[33], net750[34],
     net750[35], net750[36], net750[37], net750[38], net750[39],
     net750[40], net750[41], net750[42], net750[43], net750[44],
     net750[45], net750[46], net750[47]}), .sp4_h_l_05({net752[0],
     net752[1], net752[2], net752[3], net752[4], net752[5], net752[6],
     net752[7], net752[8], net752[9], net752[10], net752[11],
     net752[12], net752[13], net752[14], net752[15], net752[16],
     net752[17], net752[18], net752[19], net752[20], net752[21],
     net752[22], net752[23], net752[24], net752[25], net752[26],
     net752[27], net752[28], net752[29], net752[30], net752[31],
     net752[32], net752[33], net752[34], net752[35], net752[36],
     net752[37], net752[38], net752[39], net752[40], net752[41],
     net752[42], net752[43], net752[44], net752[45], net752[46],
     net752[47]}), .sp4_h_r_02({net1286[0], net1286[1], net1286[2],
     net1286[3], net1286[4], net1286[5], net1286[6], net1286[7],
     net1286[8], net1286[9], net1286[10], net1286[11], net1286[12],
     net1286[13], net1286[14], net1286[15], net1286[16], net1286[17],
     net1286[18], net1286[19], net1286[20], net1286[21], net1286[22],
     net1286[23], net1286[24], net1286[25], net1286[26], net1286[27],
     net1286[28], net1286[29], net1286[30], net1286[31], net1286[32],
     net1286[33], net1286[34], net1286[35], net1286[36], net1286[37],
     net1286[38], net1286[39], net1286[40], net1286[41], net1286[42],
     net1286[43], net1286[44], net1286[45], net1286[46], net1286[47]}),
     .sp4_h_r_03({net1287[0], net1287[1], net1287[2], net1287[3],
     net1287[4], net1287[5], net1287[6], net1287[7], net1287[8],
     net1287[9], net1287[10], net1287[11], net1287[12], net1287[13],
     net1287[14], net1287[15], net1287[16], net1287[17], net1287[18],
     net1287[19], net1287[20], net1287[21], net1287[22], net1287[23],
     net1287[24], net1287[25], net1287[26], net1287[27], net1287[28],
     net1287[29], net1287[30], net1287[31], net1287[32], net1287[33],
     net1287[34], net1287[35], net1287[36], net1287[37], net1287[38],
     net1287[39], net1287[40], net1287[41], net1287[42], net1287[43],
     net1287[44], net1287[45], net1287[46], net1287[47]}),
     .sp4_h_r_04({net1288[0], net1288[1], net1288[2], net1288[3],
     net1288[4], net1288[5], net1288[6], net1288[7], net1288[8],
     net1288[9], net1288[10], net1288[11], net1288[12], net1288[13],
     net1288[14], net1288[15], net1288[16], net1288[17], net1288[18],
     net1288[19], net1288[20], net1288[21], net1288[22], net1288[23],
     net1288[24], net1288[25], net1288[26], net1288[27], net1288[28],
     net1288[29], net1288[30], net1288[31], net1288[32], net1288[33],
     net1288[34], net1288[35], net1288[36], net1288[37], net1288[38],
     net1288[39], net1288[40], net1288[41], net1288[42], net1288[43],
     net1288[44], net1288[45], net1288[46], net1288[47]}),
     .sp4_h_r_05({net1289[0], net1289[1], net1289[2], net1289[3],
     net1289[4], net1289[5], net1289[6], net1289[7], net1289[8],
     net1289[9], net1289[10], net1289[11], net1289[12], net1289[13],
     net1289[14], net1289[15], net1289[16], net1289[17], net1289[18],
     net1289[19], net1289[20], net1289[21], net1289[22], net1289[23],
     net1289[24], net1289[25], net1289[26], net1289[27], net1289[28],
     net1289[29], net1289[30], net1289[31], net1289[32], net1289[33],
     net1289[34], net1289[35], net1289[36], net1289[37], net1289[38],
     net1289[39], net1289[40], net1289[41], net1289[42], net1289[43],
     net1289[44], net1289[45], net1289[46], net1289[47]}),
     .sp4_h_r_06({net1290[0], net1290[1], net1290[2], net1290[3],
     net1290[4], net1290[5], net1290[6], net1290[7], net1290[8],
     net1290[9], net1290[10], net1290[11], net1290[12], net1290[13],
     net1290[14], net1290[15], net1290[16], net1290[17], net1290[18],
     net1290[19], net1290[20], net1290[21], net1290[22], net1290[23],
     net1290[24], net1290[25], net1290[26], net1290[27], net1290[28],
     net1290[29], net1290[30], net1290[31], net1290[32], net1290[33],
     net1290[34], net1290[35], net1290[36], net1290[37], net1290[38],
     net1290[39], net1290[40], net1290[41], net1290[42], net1290[43],
     net1290[44], net1290[45], net1290[46], net1290[47]}),
     .sp4_h_r_07({net1291[0], net1291[1], net1291[2], net1291[3],
     net1291[4], net1291[5], net1291[6], net1291[7], net1291[8],
     net1291[9], net1291[10], net1291[11], net1291[12], net1291[13],
     net1291[14], net1291[15], net1291[16], net1291[17], net1291[18],
     net1291[19], net1291[20], net1291[21], net1291[22], net1291[23],
     net1291[24], net1291[25], net1291[26], net1291[27], net1291[28],
     net1291[29], net1291[30], net1291[31], net1291[32], net1291[33],
     net1291[34], net1291[35], net1291[36], net1291[37], net1291[38],
     net1291[39], net1291[40], net1291[41], net1291[42], net1291[43],
     net1291[44], net1291[45], net1291[46], net1291[47]}));
lt_1x8_bot_ice1f I_lt_col_t02 ( .rgt_op_03({net698[0], net698[1],
     net698[2], net698[3], net698[4], net698[5], net698[6],
     net698[7]}), .slf_op_02({net795[0], net795[1], net795[2],
     net795[3], net795[4], net795[5], net795[6], net795[7]}),
     .rgt_op_02({net700[0], net700[1], net700[2], net700[3], net700[4],
     net700[5], net700[6], net700[7]}), .rgt_op_01({net1410[0],
     net1410[1], net1410[2], net1410[3], net1410[4], net1410[5],
     net1410[6], net1410[7]}), .purst(purst), .prog(prog),
     .lft_op_04({net1355[0], net1355[1], net1355[2], net1355[3],
     net1355[4], net1355[5], net1355[6], net1355[7]}),
     .lft_op_03({net1330[0], net1330[1], net1330[2], net1330[3],
     net1330[4], net1330[5], net1330[6], net1330[7]}),
     .lft_op_02({net1314[0], net1314[1], net1314[2], net1314[3],
     net1314[4], net1314[5], net1314[6], net1314[7]}),
     .lft_op_01({net1417[0], net1417[1], net1417[2], net1417[3],
     net1417[4], net1417[5], net1417[6], net1417[7]}),
     .rgt_op_04({net708[0], net708[1], net708[2], net708[3], net708[4],
     net708[5], net708[6], net708[7]}), .glb_netwk_bot({net1387[0],
     net1387[1], net1387[2], net1387[3], net1387[4], net1387[5],
     net1387[6], net1387[7]}), .carry_in(tiegnd_bl),
     .bnl_op_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}), .slf_op_04({net803[0],
     net803[1], net803[2], net803[3], net803[4], net803[5], net803[6],
     net803[7]}), .slf_op_03({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7]}),
     .slf_op_01({net1419[0], net1419[1], net1419[2], net1419[3],
     net1419[4], net1419[5], net1419[6], net1419[7]}),
     .sp4_h_l_04({net822[0], net822[1], net822[2], net822[3],
     net822[4], net822[5], net822[6], net822[7], net822[8], net822[9],
     net822[10], net822[11], net822[12], net822[13], net822[14],
     net822[15], net822[16], net822[17], net822[18], net822[19],
     net822[20], net822[21], net822[22], net822[23], net822[24],
     net822[25], net822[26], net822[27], net822[28], net822[29],
     net822[30], net822[31], net822[32], net822[33], net822[34],
     net822[35], net822[36], net822[37], net822[38], net822[39],
     net822[40], net822[41], net822[42], net822[43], net822[44],
     net822[45], net822[46], net822[47]}), .carry_out(carry_out_02_08),
     .vdd_cntl(vdd_cntl_l[143:16]), .sp12_h_r_04({net718[0], net718[1],
     net718[2], net718[3], net718[4], net718[5], net718[6], net718[7],
     net718[8], net718[9], net718[10], net718[11], net718[12],
     net718[13], net718[14], net718[15], net718[16], net718[17],
     net718[18], net718[19], net718[20], net718[21], net718[22],
     net718[23]}), .sp12_h_r_03({net719[0], net719[1], net719[2],
     net719[3], net719[4], net719[5], net719[6], net719[7], net719[8],
     net719[9], net719[10], net719[11], net719[12], net719[13],
     net719[14], net719[15], net719[16], net719[17], net719[18],
     net719[19], net719[20], net719[21], net719[22], net719[23]}),
     .sp12_h_r_02({net720[0], net720[1], net720[2], net720[3],
     net720[4], net720[5], net720[6], net720[7], net720[8], net720[9],
     net720[10], net720[11], net720[12], net720[13], net720[14],
     net720[15], net720[16], net720[17], net720[18], net720[19],
     net720[20], net720[21], net720[22], net720[23]}),
     .sp12_h_r_01({net721[0], net721[1], net721[2], net721[3],
     net721[4], net721[5], net721[6], net721[7], net721[8], net721[9],
     net721[10], net721[11], net721[12], net721[13], net721[14],
     net721[15], net721[16], net721[17], net721[18], net721[19],
     net721[20], net721[21], net721[22], net721[23]}),
     .glb_netwk_col({net1344[0], net1344[1], net1344[2], net1344[3],
     net1344[4], net1344[5], net1344[6], net1344[7]}),
     .sp4_v_b_01({net1411[0], net1411[1], net1411[2], net1411[3],
     net1411[4], net1411[5], net1411[6], net1411[7], net1411[8],
     net1411[9], net1411[10], net1411[11], net1411[12], net1411[13],
     net1411[14], net1411[15], net1411[16], net1411[17], net1411[18],
     net1411[19], net1411[20], net1411[21], net1411[22], net1411[23],
     net1411[24], net1411[25], net1411[26], net1411[27], net1411[28],
     net1411[29], net1411[30], net1411[31], net1411[32], net1411[33],
     net1411[34], net1411[35], net1411[36], net1411[37], net1411[38],
     net1411[39], net1411[40], net1411[41], net1411[42], net1411[43],
     net1411[44], net1411[45], net1411[46], net1411[47]}),
     .sp4_r_v_b_04({net724[0], net724[1], net724[2], net724[3],
     net724[4], net724[5], net724[6], net724[7], net724[8], net724[9],
     net724[10], net724[11], net724[12], net724[13], net724[14],
     net724[15], net724[16], net724[17], net724[18], net724[19],
     net724[20], net724[21], net724[22], net724[23], net724[24],
     net724[25], net724[26], net724[27], net724[28], net724[29],
     net724[30], net724[31], net724[32], net724[33], net724[34],
     net724[35], net724[36], net724[37], net724[38], net724[39],
     net724[40], net724[41], net724[42], net724[43], net724[44],
     net724[45], net724[46], net724[47]}), .sp4_r_v_b_03({net725[0],
     net725[1], net725[2], net725[3], net725[4], net725[5], net725[6],
     net725[7], net725[8], net725[9], net725[10], net725[11],
     net725[12], net725[13], net725[14], net725[15], net725[16],
     net725[17], net725[18], net725[19], net725[20], net725[21],
     net725[22], net725[23], net725[24], net725[25], net725[26],
     net725[27], net725[28], net725[29], net725[30], net725[31],
     net725[32], net725[33], net725[34], net725[35], net725[36],
     net725[37], net725[38], net725[39], net725[40], net725[41],
     net725[42], net725[43], net725[44], net725[45], net725[46],
     net725[47]}), .sp4_r_v_b_02({net726[0], net726[1], net726[2],
     net726[3], net726[4], net726[5], net726[6], net726[7], net726[8],
     net726[9], net726[10], net726[11], net726[12], net726[13],
     net726[14], net726[15], net726[16], net726[17], net726[18],
     net726[19], net726[20], net726[21], net726[22], net726[23],
     net726[24], net726[25], net726[26], net726[27], net726[28],
     net726[29], net726[30], net726[31], net726[32], net726[33],
     net726[34], net726[35], net726[36], net726[37], net726[38],
     net726[39], net726[40], net726[41], net726[42], net726[43],
     net726[44], net726[45], net726[46], net726[47]}),
     .sp4_r_v_b_01({net1412[0], net1412[1], net1412[2], net1412[3],
     net1412[4], net1412[5], net1412[6], net1412[7], net1412[8],
     net1412[9], net1412[10], net1412[11], net1412[12], net1412[13],
     net1412[14], net1412[15], net1412[16], net1412[17], net1412[18],
     net1412[19], net1412[20], net1412[21], net1412[22], net1412[23],
     net1412[24], net1412[25], net1412[26], net1412[27], net1412[28],
     net1412[29], net1412[30], net1412[31], net1412[32], net1412[33],
     net1412[34], net1412[35], net1412[36], net1412[37], net1412[38],
     net1412[39], net1412[40], net1412[41], net1412[42], net1412[43],
     net1412[44], net1412[45], net1412[46], net1412[47]}),
     .sp4_h_r_04({net728[0], net728[1], net728[2], net728[3],
     net728[4], net728[5], net728[6], net728[7], net728[8], net728[9],
     net728[10], net728[11], net728[12], net728[13], net728[14],
     net728[15], net728[16], net728[17], net728[18], net728[19],
     net728[20], net728[21], net728[22], net728[23], net728[24],
     net728[25], net728[26], net728[27], net728[28], net728[29],
     net728[30], net728[31], net728[32], net728[33], net728[34],
     net728[35], net728[36], net728[37], net728[38], net728[39],
     net728[40], net728[41], net728[42], net728[43], net728[44],
     net728[45], net728[46], net728[47]}), .sp4_h_r_03({net729[0],
     net729[1], net729[2], net729[3], net729[4], net729[5], net729[6],
     net729[7], net729[8], net729[9], net729[10], net729[11],
     net729[12], net729[13], net729[14], net729[15], net729[16],
     net729[17], net729[18], net729[19], net729[20], net729[21],
     net729[22], net729[23], net729[24], net729[25], net729[26],
     net729[27], net729[28], net729[29], net729[30], net729[31],
     net729[32], net729[33], net729[34], net729[35], net729[36],
     net729[37], net729[38], net729[39], net729[40], net729[41],
     net729[42], net729[43], net729[44], net729[45], net729[46],
     net729[47]}), .sp4_h_r_02({net730[0], net730[1], net730[2],
     net730[3], net730[4], net730[5], net730[6], net730[7], net730[8],
     net730[9], net730[10], net730[11], net730[12], net730[13],
     net730[14], net730[15], net730[16], net730[17], net730[18],
     net730[19], net730[20], net730[21], net730[22], net730[23],
     net730[24], net730[25], net730[26], net730[27], net730[28],
     net730[29], net730[30], net730[31], net730[32], net730[33],
     net730[34], net730[35], net730[36], net730[37], net730[38],
     net730[39], net730[40], net730[41], net730[42], net730[43],
     net730[44], net730[45], net730[46], net730[47]}),
     .sp4_h_r_01({net731[0], net731[1], net731[2], net731[3],
     net731[4], net731[5], net731[6], net731[7], net731[8], net731[9],
     net731[10], net731[11], net731[12], net731[13], net731[14],
     net731[15], net731[16], net731[17], net731[18], net731[19],
     net731[20], net731[21], net731[22], net731[23], net731[24],
     net731[25], net731[26], net731[27], net731[28], net731[29],
     net731[30], net731[31], net731[32], net731[33], net731[34],
     net731[35], net731[36], net731[37], net731[38], net731[39],
     net731[40], net731[41], net731[42], net731[43], net731[44],
     net731[45], net731[46], net731[47]}), .sp4_h_l_03({net823[0],
     net823[1], net823[2], net823[3], net823[4], net823[5], net823[6],
     net823[7], net823[8], net823[9], net823[10], net823[11],
     net823[12], net823[13], net823[14], net823[15], net823[16],
     net823[17], net823[18], net823[19], net823[20], net823[21],
     net823[22], net823[23], net823[24], net823[25], net823[26],
     net823[27], net823[28], net823[29], net823[30], net823[31],
     net823[32], net823[33], net823[34], net823[35], net823[36],
     net823[37], net823[38], net823[39], net823[40], net823[41],
     net823[42], net823[43], net823[44], net823[45], net823[46],
     net823[47]}), .sp4_h_l_02({net824[0], net824[1], net824[2],
     net824[3], net824[4], net824[5], net824[6], net824[7], net824[8],
     net824[9], net824[10], net824[11], net824[12], net824[13],
     net824[14], net824[15], net824[16], net824[17], net824[18],
     net824[19], net824[20], net824[21], net824[22], net824[23],
     net824[24], net824[25], net824[26], net824[27], net824[28],
     net824[29], net824[30], net824[31], net824[32], net824[33],
     net824[34], net824[35], net824[36], net824[37], net824[38],
     net824[39], net824[40], net824[41], net824[42], net824[43],
     net824[44], net824[45], net824[46], net824[47]}),
     .sp4_h_l_01({net825[0], net825[1], net825[2], net825[3],
     net825[4], net825[5], net825[6], net825[7], net825[8], net825[9],
     net825[10], net825[11], net825[12], net825[13], net825[14],
     net825[15], net825[16], net825[17], net825[18], net825[19],
     net825[20], net825[21], net825[22], net825[23], net825[24],
     net825[25], net825[26], net825[27], net825[28], net825[29],
     net825[30], net825[31], net825[32], net825[33], net825[34],
     net825[35], net825[36], net825[37], net825[38], net825[39],
     net825[40], net825[41], net825[42], net825[43], net825[44],
     net825[45], net825[46], net825[47]}), .bl(bl[125:72]),
     .bot_op_01({slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0], slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0]}), .sp12_h_l_01({net815[0],
     net815[1], net815[2], net815[3], net815[4], net815[5], net815[6],
     net815[7], net815[8], net815[9], net815[10], net815[11],
     net815[12], net815[13], net815[14], net815[15], net815[16],
     net815[17], net815[18], net815[19], net815[20], net815[21],
     net815[22], net815[23]}), .sp12_h_l_02({net814[0], net814[1],
     net814[2], net814[3], net814[4], net814[5], net814[6], net814[7],
     net814[8], net814[9], net814[10], net814[11], net814[12],
     net814[13], net814[14], net814[15], net814[16], net814[17],
     net814[18], net814[19], net814[20], net814[21], net814[22],
     net814[23]}), .sp12_h_l_03({net813[0], net813[1], net813[2],
     net813[3], net813[4], net813[5], net813[6], net813[7], net813[8],
     net813[9], net813[10], net813[11], net813[12], net813[13],
     net813[14], net813[15], net813[16], net813[17], net813[18],
     net813[19], net813[20], net813[21], net813[22], net813[23]}),
     .sp12_h_l_04({net812[0], net812[1], net812[2], net812[3],
     net812[4], net812[5], net812[6], net812[7], net812[8], net812[9],
     net812[10], net812[11], net812[12], net812[13], net812[14],
     net812[15], net812[16], net812[17], net812[18], net812[19],
     net812[20], net812[21], net812[22], net812[23]}),
     .sp4_v_b_04({net818[0], net818[1], net818[2], net818[3],
     net818[4], net818[5], net818[6], net818[7], net818[8], net818[9],
     net818[10], net818[11], net818[12], net818[13], net818[14],
     net818[15], net818[16], net818[17], net818[18], net818[19],
     net818[20], net818[21], net818[22], net818[23], net818[24],
     net818[25], net818[26], net818[27], net818[28], net818[29],
     net818[30], net818[31], net818[32], net818[33], net818[34],
     net818[35], net818[36], net818[37], net818[38], net818[39],
     net818[40], net818[41], net818[42], net818[43], net818[44],
     net818[45], net818[46], net818[47]}), .sp4_v_b_03({net819[0],
     net819[1], net819[2], net819[3], net819[4], net819[5], net819[6],
     net819[7], net819[8], net819[9], net819[10], net819[11],
     net819[12], net819[13], net819[14], net819[15], net819[16],
     net819[17], net819[18], net819[19], net819[20], net819[21],
     net819[22], net819[23], net819[24], net819[25], net819[26],
     net819[27], net819[28], net819[29], net819[30], net819[31],
     net819[32], net819[33], net819[34], net819[35], net819[36],
     net819[37], net819[38], net819[39], net819[40], net819[41],
     net819[42], net819[43], net819[44], net819[45], net819[46],
     net819[47]}), .sp4_v_b_02({net820[0], net820[1], net820[2],
     net820[3], net820[4], net820[5], net820[6], net820[7], net820[8],
     net820[9], net820[10], net820[11], net820[12], net820[13],
     net820[14], net820[15], net820[16], net820[17], net820[18],
     net820[19], net820[20], net820[21], net820[22], net820[23],
     net820[24], net820[25], net820[26], net820[27], net820[28],
     net820[29], net820[30], net820[31], net820[32], net820[33],
     net820[34], net820[35], net820[36], net820[37], net820[38],
     net820[39], net820[40], net820[41], net820[42], net820[43],
     net820[44], net820[45], net820[46], net820[47]}),
     .bnr_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .sp4_h_l_05({net846[0],
     net846[1], net846[2], net846[3], net846[4], net846[5], net846[6],
     net846[7], net846[8], net846[9], net846[10], net846[11],
     net846[12], net846[13], net846[14], net846[15], net846[16],
     net846[17], net846[18], net846[19], net846[20], net846[21],
     net846[22], net846[23], net846[24], net846[25], net846[26],
     net846[27], net846[28], net846[29], net846[30], net846[31],
     net846[32], net846[33], net846[34], net846[35], net846[36],
     net846[37], net846[38], net846[39], net846[40], net846[41],
     net846[42], net846[43], net846[44], net846[45], net846[46],
     net846[47]}), .sp4_h_l_06({net845[0], net845[1], net845[2],
     net845[3], net845[4], net845[5], net845[6], net845[7], net845[8],
     net845[9], net845[10], net845[11], net845[12], net845[13],
     net845[14], net845[15], net845[16], net845[17], net845[18],
     net845[19], net845[20], net845[21], net845[22], net845[23],
     net845[24], net845[25], net845[26], net845[27], net845[28],
     net845[29], net845[30], net845[31], net845[32], net845[33],
     net845[34], net845[35], net845[36], net845[37], net845[38],
     net845[39], net845[40], net845[41], net845[42], net845[43],
     net845[44], net845[45], net845[46], net845[47]}),
     .sp4_h_l_07({net844[0], net844[1], net844[2], net844[3],
     net844[4], net844[5], net844[6], net844[7], net844[8], net844[9],
     net844[10], net844[11], net844[12], net844[13], net844[14],
     net844[15], net844[16], net844[17], net844[18], net844[19],
     net844[20], net844[21], net844[22], net844[23], net844[24],
     net844[25], net844[26], net844[27], net844[28], net844[29],
     net844[30], net844[31], net844[32], net844[33], net844[34],
     net844[35], net844[36], net844[37], net844[38], net844[39],
     net844[40], net844[41], net844[42], net844[43], net844[44],
     net844[45], net844[46], net844[47]}), .sp4_h_l_08({net843[0],
     net843[1], net843[2], net843[3], net843[4], net843[5], net843[6],
     net843[7], net843[8], net843[9], net843[10], net843[11],
     net843[12], net843[13], net843[14], net843[15], net843[16],
     net843[17], net843[18], net843[19], net843[20], net843[21],
     net843[22], net843[23], net843[24], net843[25], net843[26],
     net843[27], net843[28], net843[29], net843[30], net843[31],
     net843[32], net843[33], net843[34], net843[35], net843[36],
     net843[37], net843[38], net843[39], net843[40], net843[41],
     net843[42], net843[43], net843[44], net843[45], net843[46],
     net843[47]}), .sp4_h_r_08({net749[0], net749[1], net749[2],
     net749[3], net749[4], net749[5], net749[6], net749[7], net749[8],
     net749[9], net749[10], net749[11], net749[12], net749[13],
     net749[14], net749[15], net749[16], net749[17], net749[18],
     net749[19], net749[20], net749[21], net749[22], net749[23],
     net749[24], net749[25], net749[26], net749[27], net749[28],
     net749[29], net749[30], net749[31], net749[32], net749[33],
     net749[34], net749[35], net749[36], net749[37], net749[38],
     net749[39], net749[40], net749[41], net749[42], net749[43],
     net749[44], net749[45], net749[46], net749[47]}),
     .sp4_h_r_07({net750[0], net750[1], net750[2], net750[3],
     net750[4], net750[5], net750[6], net750[7], net750[8], net750[9],
     net750[10], net750[11], net750[12], net750[13], net750[14],
     net750[15], net750[16], net750[17], net750[18], net750[19],
     net750[20], net750[21], net750[22], net750[23], net750[24],
     net750[25], net750[26], net750[27], net750[28], net750[29],
     net750[30], net750[31], net750[32], net750[33], net750[34],
     net750[35], net750[36], net750[37], net750[38], net750[39],
     net750[40], net750[41], net750[42], net750[43], net750[44],
     net750[45], net750[46], net750[47]}), .sp4_h_r_06({net751[0],
     net751[1], net751[2], net751[3], net751[4], net751[5], net751[6],
     net751[7], net751[8], net751[9], net751[10], net751[11],
     net751[12], net751[13], net751[14], net751[15], net751[16],
     net751[17], net751[18], net751[19], net751[20], net751[21],
     net751[22], net751[23], net751[24], net751[25], net751[26],
     net751[27], net751[28], net751[29], net751[30], net751[31],
     net751[32], net751[33], net751[34], net751[35], net751[36],
     net751[37], net751[38], net751[39], net751[40], net751[41],
     net751[42], net751[43], net751[44], net751[45], net751[46],
     net751[47]}), .sp4_h_r_05({net752[0], net752[1], net752[2],
     net752[3], net752[4], net752[5], net752[6], net752[7], net752[8],
     net752[9], net752[10], net752[11], net752[12], net752[13],
     net752[14], net752[15], net752[16], net752[17], net752[18],
     net752[19], net752[20], net752[21], net752[22], net752[23],
     net752[24], net752[25], net752[26], net752[27], net752[28],
     net752[29], net752[30], net752[31], net752[32], net752[33],
     net752[34], net752[35], net752[36], net752[37], net752[38],
     net752[39], net752[40], net752[41], net752[42], net752[43],
     net752[44], net752[45], net752[46], net752[47]}),
     .slf_op_05({net854[0], net854[1], net854[2], net854[3], net854[4],
     net854[5], net854[6], net854[7]}), .slf_op_06({net853[0],
     net853[1], net853[2], net853[3], net853[4], net853[5], net853[6],
     net853[7]}), .slf_op_07({net852[0], net852[1], net852[2],
     net852[3], net852[4], net852[5], net852[6], net852[7]}),
     .slf_op_08(slf_op_02_08[7:0]), .rgt_op_08(slf_op_03_08[7:0]),
     .rgt_op_07({net758[0], net758[1], net758[2], net758[3], net758[4],
     net758[5], net758[6], net758[7]}), .rgt_op_06({net759[0],
     net759[1], net759[2], net759[3], net759[4], net759[5], net759[6],
     net759[7]}), .rgt_op_05({net760[0], net760[1], net760[2],
     net760[3], net760[4], net760[5], net760[6], net760[7]}),
     .lft_op_08(slf_op_01_08[7:0]), .lft_op_07({net1327[0], net1327[1],
     net1327[2], net1327[3], net1327[4], net1327[5], net1327[6],
     net1327[7]}), .lft_op_06({net1328[0], net1328[1], net1328[2],
     net1328[3], net1328[4], net1328[5], net1328[6], net1328[7]}),
     .lft_op_05({net1329[0], net1329[1], net1329[2], net1329[3],
     net1329[4], net1329[5], net1329[6], net1329[7]}),
     .sp12_h_l_08({net865[0], net865[1], net865[2], net865[3],
     net865[4], net865[5], net865[6], net865[7], net865[8], net865[9],
     net865[10], net865[11], net865[12], net865[13], net865[14],
     net865[15], net865[16], net865[17], net865[18], net865[19],
     net865[20], net865[21], net865[22], net865[23]}),
     .sp12_h_l_07({net864[0], net864[1], net864[2], net864[3],
     net864[4], net864[5], net864[6], net864[7], net864[8], net864[9],
     net864[10], net864[11], net864[12], net864[13], net864[14],
     net864[15], net864[16], net864[17], net864[18], net864[19],
     net864[20], net864[21], net864[22], net864[23]}),
     .sp12_h_l_06({net863[0], net863[1], net863[2], net863[3],
     net863[4], net863[5], net863[6], net863[7], net863[8], net863[9],
     net863[10], net863[11], net863[12], net863[13], net863[14],
     net863[15], net863[16], net863[17], net863[18], net863[19],
     net863[20], net863[21], net863[22], net863[23]}),
     .sp12_h_r_05({net768[0], net768[1], net768[2], net768[3],
     net768[4], net768[5], net768[6], net768[7], net768[8], net768[9],
     net768[10], net768[11], net768[12], net768[13], net768[14],
     net768[15], net768[16], net768[17], net768[18], net768[19],
     net768[20], net768[21], net768[22], net768[23]}),
     .sp12_h_r_06({net769[0], net769[1], net769[2], net769[3],
     net769[4], net769[5], net769[6], net769[7], net769[8], net769[9],
     net769[10], net769[11], net769[12], net769[13], net769[14],
     net769[15], net769[16], net769[17], net769[18], net769[19],
     net769[20], net769[21], net769[22], net769[23]}),
     .sp12_h_r_07({net770[0], net770[1], net770[2], net770[3],
     net770[4], net770[5], net770[6], net770[7], net770[8], net770[9],
     net770[10], net770[11], net770[12], net770[13], net770[14],
     net770[15], net770[16], net770[17], net770[18], net770[19],
     net770[20], net770[21], net770[22], net770[23]}),
     .sp12_h_r_08({net771[0], net771[1], net771[2], net771[3],
     net771[4], net771[5], net771[6], net771[7], net771[8], net771[9],
     net771[10], net771[11], net771[12], net771[13], net771[14],
     net771[15], net771[16], net771[17], net771[18], net771[19],
     net771[20], net771[21], net771[22], net771[23]}),
     .sp12_h_l_05({net862[0], net862[1], net862[2], net862[3],
     net862[4], net862[5], net862[6], net862[7], net862[8], net862[9],
     net862[10], net862[11], net862[12], net862[13], net862[14],
     net862[15], net862[16], net862[17], net862[18], net862[19],
     net862[20], net862[21], net862[22], net862[23]}),
     .sp4_r_v_b_05({net773[0], net773[1], net773[2], net773[3],
     net773[4], net773[5], net773[6], net773[7], net773[8], net773[9],
     net773[10], net773[11], net773[12], net773[13], net773[14],
     net773[15], net773[16], net773[17], net773[18], net773[19],
     net773[20], net773[21], net773[22], net773[23], net773[24],
     net773[25], net773[26], net773[27], net773[28], net773[29],
     net773[30], net773[31], net773[32], net773[33], net773[34],
     net773[35], net773[36], net773[37], net773[38], net773[39],
     net773[40], net773[41], net773[42], net773[43], net773[44],
     net773[45], net773[46], net773[47]}), .sp4_r_v_b_06({net774[0],
     net774[1], net774[2], net774[3], net774[4], net774[5], net774[6],
     net774[7], net774[8], net774[9], net774[10], net774[11],
     net774[12], net774[13], net774[14], net774[15], net774[16],
     net774[17], net774[18], net774[19], net774[20], net774[21],
     net774[22], net774[23], net774[24], net774[25], net774[26],
     net774[27], net774[28], net774[29], net774[30], net774[31],
     net774[32], net774[33], net774[34], net774[35], net774[36],
     net774[37], net774[38], net774[39], net774[40], net774[41],
     net774[42], net774[43], net774[44], net774[45], net774[46],
     net774[47]}), .sp4_r_v_b_07({net775[0], net775[1], net775[2],
     net775[3], net775[4], net775[5], net775[6], net775[7], net775[8],
     net775[9], net775[10], net775[11], net775[12], net775[13],
     net775[14], net775[15], net775[16], net775[17], net775[18],
     net775[19], net775[20], net775[21], net775[22], net775[23],
     net775[24], net775[25], net775[26], net775[27], net775[28],
     net775[29], net775[30], net775[31], net775[32], net775[33],
     net775[34], net775[35], net775[36], net775[37], net775[38],
     net775[39], net775[40], net775[41], net775[42], net775[43],
     net775[44], net775[45], net775[46], net775[47]}),
     .sp4_r_v_b_08({net776[0], net776[1], net776[2], net776[3],
     net776[4], net776[5], net776[6], net776[7], net776[8], net776[9],
     net776[10], net776[11], net776[12], net776[13], net776[14],
     net776[15], net776[16], net776[17], net776[18], net776[19],
     net776[20], net776[21], net776[22], net776[23], net776[24],
     net776[25], net776[26], net776[27], net776[28], net776[29],
     net776[30], net776[31], net776[32], net776[33], net776[34],
     net776[35], net776[36], net776[37], net776[38], net776[39],
     net776[40], net776[41], net776[42], net776[43], net776[44],
     net776[45], net776[46], net776[47]}), .sp4_v_b_08({net870[0],
     net870[1], net870[2], net870[3], net870[4], net870[5], net870[6],
     net870[7], net870[8], net870[9], net870[10], net870[11],
     net870[12], net870[13], net870[14], net870[15], net870[16],
     net870[17], net870[18], net870[19], net870[20], net870[21],
     net870[22], net870[23], net870[24], net870[25], net870[26],
     net870[27], net870[28], net870[29], net870[30], net870[31],
     net870[32], net870[33], net870[34], net870[35], net870[36],
     net870[37], net870[38], net870[39], net870[40], net870[41],
     net870[42], net870[43], net870[44], net870[45], net870[46],
     net870[47]}), .sp4_v_b_07({net869[0], net869[1], net869[2],
     net869[3], net869[4], net869[5], net869[6], net869[7], net869[8],
     net869[9], net869[10], net869[11], net869[12], net869[13],
     net869[14], net869[15], net869[16], net869[17], net869[18],
     net869[19], net869[20], net869[21], net869[22], net869[23],
     net869[24], net869[25], net869[26], net869[27], net869[28],
     net869[29], net869[30], net869[31], net869[32], net869[33],
     net869[34], net869[35], net869[36], net869[37], net869[38],
     net869[39], net869[40], net869[41], net869[42], net869[43],
     net869[44], net869[45], net869[46], net869[47]}),
     .sp4_v_b_06({net868[0], net868[1], net868[2], net868[3],
     net868[4], net868[5], net868[6], net868[7], net868[8], net868[9],
     net868[10], net868[11], net868[12], net868[13], net868[14],
     net868[15], net868[16], net868[17], net868[18], net868[19],
     net868[20], net868[21], net868[22], net868[23], net868[24],
     net868[25], net868[26], net868[27], net868[28], net868[29],
     net868[30], net868[31], net868[32], net868[33], net868[34],
     net868[35], net868[36], net868[37], net868[38], net868[39],
     net868[40], net868[41], net868[42], net868[43], net868[44],
     net868[45], net868[46], net868[47]}), .sp4_v_b_05({net867[0],
     net867[1], net867[2], net867[3], net867[4], net867[5], net867[6],
     net867[7], net867[8], net867[9], net867[10], net867[11],
     net867[12], net867[13], net867[14], net867[15], net867[16],
     net867[17], net867[18], net867[19], net867[20], net867[21],
     net867[22], net867[23], net867[24], net867[25], net867[26],
     net867[27], net867[28], net867[29], net867[30], net867[31],
     net867[32], net867[33], net867[34], net867[35], net867[36],
     net867[37], net867[38], net867[39], net867[40], net867[41],
     net867[42], net867[43], net867[44], net867[45], net867[46],
     net867[47]}), .pgate(pgate_l[143:16]),
     .reset_b(reset_b_l[143:16]), .wl(wl_l[143:16]),
     .top_op_08(top_op_02_08[7:0]), .tnr_op_08(tnr_op_02_08[7:0]),
     .tnl_op_08(tnl_op_02_08[7:0]), .sp12_v_t_08(sp12_v_t_02_08[23:0]),
     .sp4_v_t_08(sp4_v_t_02_08[47:0]), .lc_bot(tiegnd_bl),
     .op_vic(op_vic_02_08), .sp12_v_b_01({net1390[0], net1390[1],
     net1390[2], net1390[3], net1390[4], net1390[5], net1390[6],
     net1390[7], net1390[8], net1390[9], net1390[10], net1390[11],
     net1390[12], net1390[13], net1390[14], net1390[15], net1390[16],
     net1390[17], net1390[18], net1390[19], net1390[20], net1390[21],
     net1390[22], net1390[23]}));
lt_1x8_bot_ice1f I_lt_col_t01 ( .glb_netwk_bot({net1388[0], net1388[1],
     net1388[2], net1388[3], net1388[4], net1388[5], net1388[6],
     net1388[7]}), .rgt_op_03({net793[0], net793[1], net793[2],
     net793[3], net793[4], net793[5], net793[6], net793[7]}),
     .slf_op_02({net1314[0], net1314[1], net1314[2], net1314[3],
     net1314[4], net1314[5], net1314[6], net1314[7]}),
     .rgt_op_02({net795[0], net795[1], net795[2], net795[3], net795[4],
     net795[5], net795[6], net795[7]}), .rgt_op_01({net1419[0],
     net1419[1], net1419[2], net1419[3], net1419[4], net1419[5],
     net1419[6], net1419[7]}), .purst(purst), .prog(prog),
     .lft_op_04({slf_op_00_04[3], slf_op_00_04[2], slf_op_00_04[1],
     slf_op_00_04[0], slf_op_00_04[3], slf_op_00_04[2],
     slf_op_00_04[1], slf_op_00_04[0]}), .lft_op_03({slf_op_00_03[3],
     slf_op_00_03[2], slf_op_00_03[1], slf_op_00_03[0],
     slf_op_00_03[3], slf_op_00_03[2], slf_op_00_03[1],
     slf_op_00_03[0]}), .lft_op_02({slf_op_00_02[3], slf_op_00_02[2],
     slf_op_00_02[1], slf_op_00_02[0], slf_op_00_02[3],
     slf_op_00_02[2], slf_op_00_02[1], slf_op_00_02[0]}),
     .lft_op_01({slf_op_00_01[3], slf_op_00_01[2], slf_op_00_01[1],
     slf_op_00_01[0], slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0]}), .rgt_op_04({net803[0],
     net803[1], net803[2], net803[3], net803[4], net803[5], net803[6],
     net803[7]}), .carry_in(tiegnd_bl), .bnl_op_01({pll_lock_out,
     pll_lock_out, pll_lock_out, pll_lock_out, pll_lock_out,
     pll_lock_out, pll_lock_out, pll_lock_out}),
     .slf_op_04({net1355[0], net1355[1], net1355[2], net1355[3],
     net1355[4], net1355[5], net1355[6], net1355[7]}),
     .slf_op_03({net1330[0], net1330[1], net1330[2], net1330[3],
     net1330[4], net1330[5], net1330[6], net1330[7]}),
     .slf_op_01({net1417[0], net1417[1], net1417[2], net1417[3],
     net1417[4], net1417[5], net1417[6], net1417[7]}),
     .sp4_h_l_04({net1324[0], net1324[1], net1324[2], net1324[3],
     net1324[4], net1324[5], net1324[6], net1324[7], net1324[8],
     net1324[9], net1324[10], net1324[11], net1324[12], net1324[13],
     net1324[14], net1324[15], net1324[16], net1324[17], net1324[18],
     net1324[19], net1324[20], net1324[21], net1324[22], net1324[23],
     net1324[24], net1324[25], net1324[26], net1324[27], net1324[28],
     net1324[29], net1324[30], net1324[31], net1324[32], net1324[33],
     net1324[34], net1324[35], net1324[36], net1324[37], net1324[38],
     net1324[39], net1324[40], net1324[41], net1324[42], net1324[43],
     net1324[44], net1324[45], net1324[46], net1324[47]}),
     .carry_out(carry_out_01_08), .vdd_cntl(vdd_cntl_l[143:16]),
     .sp12_h_r_04({net812[0], net812[1], net812[2], net812[3],
     net812[4], net812[5], net812[6], net812[7], net812[8], net812[9],
     net812[10], net812[11], net812[12], net812[13], net812[14],
     net812[15], net812[16], net812[17], net812[18], net812[19],
     net812[20], net812[21], net812[22], net812[23]}),
     .sp12_h_r_03({net813[0], net813[1], net813[2], net813[3],
     net813[4], net813[5], net813[6], net813[7], net813[8], net813[9],
     net813[10], net813[11], net813[12], net813[13], net813[14],
     net813[15], net813[16], net813[17], net813[18], net813[19],
     net813[20], net813[21], net813[22], net813[23]}),
     .sp12_h_r_02({net814[0], net814[1], net814[2], net814[3],
     net814[4], net814[5], net814[6], net814[7], net814[8], net814[9],
     net814[10], net814[11], net814[12], net814[13], net814[14],
     net814[15], net814[16], net814[17], net814[18], net814[19],
     net814[20], net814[21], net814[22], net814[23]}),
     .sp12_h_r_01({net815[0], net815[1], net815[2], net815[3],
     net815[4], net815[5], net815[6], net815[7], net815[8], net815[9],
     net815[10], net815[11], net815[12], net815[13], net815[14],
     net815[15], net815[16], net815[17], net815[18], net815[19],
     net815[20], net815[21], net815[22], net815[23]}),
     .glb_netwk_col({net1344[0], net1344[1], net1344[2], net1344[3],
     net1344[4], net1344[5], net1344[6], net1344[7]}),
     .sp4_v_b_01({net1437[0], net1437[1], net1437[2], net1437[3],
     net1437[4], net1437[5], net1437[6], net1437[7], net1437[8],
     net1437[9], net1437[10], net1437[11], net1437[12], net1437[13],
     net1437[14], net1437[15], net1437[16], net1437[17], net1437[18],
     net1437[19], net1437[20], net1437[21], net1437[22], net1437[23],
     net1437[24], net1437[25], net1437[26], net1437[27], net1437[28],
     net1437[29], net1437[30], net1437[31], net1437[32], net1437[33],
     net1437[34], net1437[35], net1437[36], net1437[37], net1437[38],
     net1437[39], net1437[40], net1437[41], net1437[42], net1437[43],
     net1437[44], net1437[45], net1437[46], net1437[47]}),
     .sp4_r_v_b_04({net818[0], net818[1], net818[2], net818[3],
     net818[4], net818[5], net818[6], net818[7], net818[8], net818[9],
     net818[10], net818[11], net818[12], net818[13], net818[14],
     net818[15], net818[16], net818[17], net818[18], net818[19],
     net818[20], net818[21], net818[22], net818[23], net818[24],
     net818[25], net818[26], net818[27], net818[28], net818[29],
     net818[30], net818[31], net818[32], net818[33], net818[34],
     net818[35], net818[36], net818[37], net818[38], net818[39],
     net818[40], net818[41], net818[42], net818[43], net818[44],
     net818[45], net818[46], net818[47]}), .sp4_r_v_b_03({net819[0],
     net819[1], net819[2], net819[3], net819[4], net819[5], net819[6],
     net819[7], net819[8], net819[9], net819[10], net819[11],
     net819[12], net819[13], net819[14], net819[15], net819[16],
     net819[17], net819[18], net819[19], net819[20], net819[21],
     net819[22], net819[23], net819[24], net819[25], net819[26],
     net819[27], net819[28], net819[29], net819[30], net819[31],
     net819[32], net819[33], net819[34], net819[35], net819[36],
     net819[37], net819[38], net819[39], net819[40], net819[41],
     net819[42], net819[43], net819[44], net819[45], net819[46],
     net819[47]}), .sp4_r_v_b_02({net820[0], net820[1], net820[2],
     net820[3], net820[4], net820[5], net820[6], net820[7], net820[8],
     net820[9], net820[10], net820[11], net820[12], net820[13],
     net820[14], net820[15], net820[16], net820[17], net820[18],
     net820[19], net820[20], net820[21], net820[22], net820[23],
     net820[24], net820[25], net820[26], net820[27], net820[28],
     net820[29], net820[30], net820[31], net820[32], net820[33],
     net820[34], net820[35], net820[36], net820[37], net820[38],
     net820[39], net820[40], net820[41], net820[42], net820[43],
     net820[44], net820[45], net820[46], net820[47]}),
     .sp4_r_v_b_01({net1411[0], net1411[1], net1411[2], net1411[3],
     net1411[4], net1411[5], net1411[6], net1411[7], net1411[8],
     net1411[9], net1411[10], net1411[11], net1411[12], net1411[13],
     net1411[14], net1411[15], net1411[16], net1411[17], net1411[18],
     net1411[19], net1411[20], net1411[21], net1411[22], net1411[23],
     net1411[24], net1411[25], net1411[26], net1411[27], net1411[28],
     net1411[29], net1411[30], net1411[31], net1411[32], net1411[33],
     net1411[34], net1411[35], net1411[36], net1411[37], net1411[38],
     net1411[39], net1411[40], net1411[41], net1411[42], net1411[43],
     net1411[44], net1411[45], net1411[46], net1411[47]}),
     .sp4_h_r_04({net822[0], net822[1], net822[2], net822[3],
     net822[4], net822[5], net822[6], net822[7], net822[8], net822[9],
     net822[10], net822[11], net822[12], net822[13], net822[14],
     net822[15], net822[16], net822[17], net822[18], net822[19],
     net822[20], net822[21], net822[22], net822[23], net822[24],
     net822[25], net822[26], net822[27], net822[28], net822[29],
     net822[30], net822[31], net822[32], net822[33], net822[34],
     net822[35], net822[36], net822[37], net822[38], net822[39],
     net822[40], net822[41], net822[42], net822[43], net822[44],
     net822[45], net822[46], net822[47]}), .sp4_h_r_03({net823[0],
     net823[1], net823[2], net823[3], net823[4], net823[5], net823[6],
     net823[7], net823[8], net823[9], net823[10], net823[11],
     net823[12], net823[13], net823[14], net823[15], net823[16],
     net823[17], net823[18], net823[19], net823[20], net823[21],
     net823[22], net823[23], net823[24], net823[25], net823[26],
     net823[27], net823[28], net823[29], net823[30], net823[31],
     net823[32], net823[33], net823[34], net823[35], net823[36],
     net823[37], net823[38], net823[39], net823[40], net823[41],
     net823[42], net823[43], net823[44], net823[45], net823[46],
     net823[47]}), .sp4_h_r_02({net824[0], net824[1], net824[2],
     net824[3], net824[4], net824[5], net824[6], net824[7], net824[8],
     net824[9], net824[10], net824[11], net824[12], net824[13],
     net824[14], net824[15], net824[16], net824[17], net824[18],
     net824[19], net824[20], net824[21], net824[22], net824[23],
     net824[24], net824[25], net824[26], net824[27], net824[28],
     net824[29], net824[30], net824[31], net824[32], net824[33],
     net824[34], net824[35], net824[36], net824[37], net824[38],
     net824[39], net824[40], net824[41], net824[42], net824[43],
     net824[44], net824[45], net824[46], net824[47]}),
     .sp4_h_r_01({net825[0], net825[1], net825[2], net825[3],
     net825[4], net825[5], net825[6], net825[7], net825[8], net825[9],
     net825[10], net825[11], net825[12], net825[13], net825[14],
     net825[15], net825[16], net825[17], net825[18], net825[19],
     net825[20], net825[21], net825[22], net825[23], net825[24],
     net825[25], net825[26], net825[27], net825[28], net825[29],
     net825[30], net825[31], net825[32], net825[33], net825[34],
     net825[35], net825[36], net825[37], net825[38], net825[39],
     net825[40], net825[41], net825[42], net825[43], net825[44],
     net825[45], net825[46], net825[47]}), .sp4_h_l_03({net1323[0],
     net1323[1], net1323[2], net1323[3], net1323[4], net1323[5],
     net1323[6], net1323[7], net1323[8], net1323[9], net1323[10],
     net1323[11], net1323[12], net1323[13], net1323[14], net1323[15],
     net1323[16], net1323[17], net1323[18], net1323[19], net1323[20],
     net1323[21], net1323[22], net1323[23], net1323[24], net1323[25],
     net1323[26], net1323[27], net1323[28], net1323[29], net1323[30],
     net1323[31], net1323[32], net1323[33], net1323[34], net1323[35],
     net1323[36], net1323[37], net1323[38], net1323[39], net1323[40],
     net1323[41], net1323[42], net1323[43], net1323[44], net1323[45],
     net1323[46], net1323[47]}), .sp4_h_l_02({net1325[0], net1325[1],
     net1325[2], net1325[3], net1325[4], net1325[5], net1325[6],
     net1325[7], net1325[8], net1325[9], net1325[10], net1325[11],
     net1325[12], net1325[13], net1325[14], net1325[15], net1325[16],
     net1325[17], net1325[18], net1325[19], net1325[20], net1325[21],
     net1325[22], net1325[23], net1325[24], net1325[25], net1325[26],
     net1325[27], net1325[28], net1325[29], net1325[30], net1325[31],
     net1325[32], net1325[33], net1325[34], net1325[35], net1325[36],
     net1325[37], net1325[38], net1325[39], net1325[40], net1325[41],
     net1325[42], net1325[43], net1325[44], net1325[45], net1325[46],
     net1325[47]}), .sp4_h_l_01({net1326[0], net1326[1], net1326[2],
     net1326[3], net1326[4], net1326[5], net1326[6], net1326[7],
     net1326[8], net1326[9], net1326[10], net1326[11], net1326[12],
     net1326[13], net1326[14], net1326[15], net1326[16], net1326[17],
     net1326[18], net1326[19], net1326[20], net1326[21], net1326[22],
     net1326[23], net1326[24], net1326[25], net1326[26], net1326[27],
     net1326[28], net1326[29], net1326[30], net1326[31], net1326[32],
     net1326[33], net1326[34], net1326[35], net1326[36], net1326[37],
     net1326[38], net1326[39], net1326[40], net1326[41], net1326[42],
     net1326[43], net1326[44], net1326[45], net1326[46], net1326[47]}),
     .bl(bl[71:18]), .bot_op_01({slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0], slf_op_01_00[3],
     slf_op_01_00[2], slf_op_01_00[1], slf_op_01_00[0]}),
     .sp12_h_l_01({net1346[0], net1346[1], net1346[2], net1346[3],
     net1346[4], net1346[5], net1346[6], net1346[7], net1346[8],
     net1346[9], net1346[10], net1346[11], net1346[12], net1346[13],
     net1346[14], net1346[15], net1346[16], net1346[17], net1346[18],
     net1346[19], net1346[20], net1346[21], net1346[22], net1346[23]}),
     .sp12_h_l_02({net1340[0], net1340[1], net1340[2], net1340[3],
     net1340[4], net1340[5], net1340[6], net1340[7], net1340[8],
     net1340[9], net1340[10], net1340[11], net1340[12], net1340[13],
     net1340[14], net1340[15], net1340[16], net1340[17], net1340[18],
     net1340[19], net1340[20], net1340[21], net1340[22], net1340[23]}),
     .sp12_h_l_03({net1348[0], net1348[1], net1348[2], net1348[3],
     net1348[4], net1348[5], net1348[6], net1348[7], net1348[8],
     net1348[9], net1348[10], net1348[11], net1348[12], net1348[13],
     net1348[14], net1348[15], net1348[16], net1348[17], net1348[18],
     net1348[19], net1348[20], net1348[21], net1348[22], net1348[23]}),
     .sp12_h_l_04({net1341[0], net1341[1], net1341[2], net1341[3],
     net1341[4], net1341[5], net1341[6], net1341[7], net1341[8],
     net1341[9], net1341[10], net1341[11], net1341[12], net1341[13],
     net1341[14], net1341[15], net1341[16], net1341[17], net1341[18],
     net1341[19], net1341[20], net1341[21], net1341[22], net1341[23]}),
     .sp4_v_b_04({net835[0], net835[1], net835[2], net835[3],
     net835[4], net835[5], net835[6], net835[7], net835[8], net835[9],
     net835[10], net835[11], net835[12], net835[13], net835[14],
     net835[15], net835[16], net835[17], net835[18], net835[19],
     net835[20], net835[21], net835[22], net835[23], net835[24],
     net835[25], net835[26], net835[27], net835[28], net835[29],
     net835[30], net835[31], net835[32], net835[33], net835[34],
     net835[35], net835[36], net835[37], net835[38], net835[39],
     net835[40], net835[41], net835[42], net835[43], net835[44],
     net835[45], net835[46], net835[47]}), .sp4_v_b_03({net1440[0],
     net1440[1], net1440[2], net1440[3], net1440[4], net1440[5],
     net1440[6], net1440[7], net1440[8], net1440[9], net1440[10],
     net1440[11], net1440[12], net1440[13], net1440[14], net1440[15],
     net1440[16], net1440[17], net1440[18], net1440[19], net1440[20],
     net1440[21], net1440[22], net1440[23], net1440[24], net1440[25],
     net1440[26], net1440[27], net1440[28], net1440[29], net1440[30],
     net1440[31], net1440[32], net1440[33], net1440[34], net1440[35],
     net1440[36], net1440[37], net1440[38], net1440[39], net1440[40],
     net1440[41], net1440[42], net1440[43], net1440[44], net1440[45],
     net1440[46], net1440[47]}), .sp4_v_b_02({net1435[0], net1435[1],
     net1435[2], net1435[3], net1435[4], net1435[5], net1435[6],
     net1435[7], net1435[8], net1435[9], net1435[10], net1435[11],
     net1435[12], net1435[13], net1435[14], net1435[15], net1435[16],
     net1435[17], net1435[18], net1435[19], net1435[20], net1435[21],
     net1435[22], net1435[23], net1435[24], net1435[25], net1435[26],
     net1435[27], net1435[28], net1435[29], net1435[30], net1435[31],
     net1435[32], net1435[33], net1435[34], net1435[35], net1435[36],
     net1435[37], net1435[38], net1435[39], net1435[40], net1435[41],
     net1435[42], net1435[43], net1435[44], net1435[45], net1435[46],
     net1435[47]}), .bnr_op_01({slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0], slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0]}),
     .sp4_h_l_05({net1304[0], net1304[1], net1304[2], net1304[3],
     net1304[4], net1304[5], net1304[6], net1304[7], net1304[8],
     net1304[9], net1304[10], net1304[11], net1304[12], net1304[13],
     net1304[14], net1304[15], net1304[16], net1304[17], net1304[18],
     net1304[19], net1304[20], net1304[21], net1304[22], net1304[23],
     net1304[24], net1304[25], net1304[26], net1304[27], net1304[28],
     net1304[29], net1304[30], net1304[31], net1304[32], net1304[33],
     net1304[34], net1304[35], net1304[36], net1304[37], net1304[38],
     net1304[39], net1304[40], net1304[41], net1304[42], net1304[43],
     net1304[44], net1304[45], net1304[46], net1304[47]}),
     .sp4_h_l_06({net1315[0], net1315[1], net1315[2], net1315[3],
     net1315[4], net1315[5], net1315[6], net1315[7], net1315[8],
     net1315[9], net1315[10], net1315[11], net1315[12], net1315[13],
     net1315[14], net1315[15], net1315[16], net1315[17], net1315[18],
     net1315[19], net1315[20], net1315[21], net1315[22], net1315[23],
     net1315[24], net1315[25], net1315[26], net1315[27], net1315[28],
     net1315[29], net1315[30], net1315[31], net1315[32], net1315[33],
     net1315[34], net1315[35], net1315[36], net1315[37], net1315[38],
     net1315[39], net1315[40], net1315[41], net1315[42], net1315[43],
     net1315[44], net1315[45], net1315[46], net1315[47]}),
     .sp4_h_l_07({net1322[0], net1322[1], net1322[2], net1322[3],
     net1322[4], net1322[5], net1322[6], net1322[7], net1322[8],
     net1322[9], net1322[10], net1322[11], net1322[12], net1322[13],
     net1322[14], net1322[15], net1322[16], net1322[17], net1322[18],
     net1322[19], net1322[20], net1322[21], net1322[22], net1322[23],
     net1322[24], net1322[25], net1322[26], net1322[27], net1322[28],
     net1322[29], net1322[30], net1322[31], net1322[32], net1322[33],
     net1322[34], net1322[35], net1322[36], net1322[37], net1322[38],
     net1322[39], net1322[40], net1322[41], net1322[42], net1322[43],
     net1322[44], net1322[45], net1322[46], net1322[47]}),
     .sp4_h_l_08({net1321[0], net1321[1], net1321[2], net1321[3],
     net1321[4], net1321[5], net1321[6], net1321[7], net1321[8],
     net1321[9], net1321[10], net1321[11], net1321[12], net1321[13],
     net1321[14], net1321[15], net1321[16], net1321[17], net1321[18],
     net1321[19], net1321[20], net1321[21], net1321[22], net1321[23],
     net1321[24], net1321[25], net1321[26], net1321[27], net1321[28],
     net1321[29], net1321[30], net1321[31], net1321[32], net1321[33],
     net1321[34], net1321[35], net1321[36], net1321[37], net1321[38],
     net1321[39], net1321[40], net1321[41], net1321[42], net1321[43],
     net1321[44], net1321[45], net1321[46], net1321[47]}),
     .sp4_h_r_08({net843[0], net843[1], net843[2], net843[3],
     net843[4], net843[5], net843[6], net843[7], net843[8], net843[9],
     net843[10], net843[11], net843[12], net843[13], net843[14],
     net843[15], net843[16], net843[17], net843[18], net843[19],
     net843[20], net843[21], net843[22], net843[23], net843[24],
     net843[25], net843[26], net843[27], net843[28], net843[29],
     net843[30], net843[31], net843[32], net843[33], net843[34],
     net843[35], net843[36], net843[37], net843[38], net843[39],
     net843[40], net843[41], net843[42], net843[43], net843[44],
     net843[45], net843[46], net843[47]}), .sp4_h_r_07({net844[0],
     net844[1], net844[2], net844[3], net844[4], net844[5], net844[6],
     net844[7], net844[8], net844[9], net844[10], net844[11],
     net844[12], net844[13], net844[14], net844[15], net844[16],
     net844[17], net844[18], net844[19], net844[20], net844[21],
     net844[22], net844[23], net844[24], net844[25], net844[26],
     net844[27], net844[28], net844[29], net844[30], net844[31],
     net844[32], net844[33], net844[34], net844[35], net844[36],
     net844[37], net844[38], net844[39], net844[40], net844[41],
     net844[42], net844[43], net844[44], net844[45], net844[46],
     net844[47]}), .sp4_h_r_06({net845[0], net845[1], net845[2],
     net845[3], net845[4], net845[5], net845[6], net845[7], net845[8],
     net845[9], net845[10], net845[11], net845[12], net845[13],
     net845[14], net845[15], net845[16], net845[17], net845[18],
     net845[19], net845[20], net845[21], net845[22], net845[23],
     net845[24], net845[25], net845[26], net845[27], net845[28],
     net845[29], net845[30], net845[31], net845[32], net845[33],
     net845[34], net845[35], net845[36], net845[37], net845[38],
     net845[39], net845[40], net845[41], net845[42], net845[43],
     net845[44], net845[45], net845[46], net845[47]}),
     .sp4_h_r_05({net846[0], net846[1], net846[2], net846[3],
     net846[4], net846[5], net846[6], net846[7], net846[8], net846[9],
     net846[10], net846[11], net846[12], net846[13], net846[14],
     net846[15], net846[16], net846[17], net846[18], net846[19],
     net846[20], net846[21], net846[22], net846[23], net846[24],
     net846[25], net846[26], net846[27], net846[28], net846[29],
     net846[30], net846[31], net846[32], net846[33], net846[34],
     net846[35], net846[36], net846[37], net846[38], net846[39],
     net846[40], net846[41], net846[42], net846[43], net846[44],
     net846[45], net846[46], net846[47]}), .slf_op_05({net1329[0],
     net1329[1], net1329[2], net1329[3], net1329[4], net1329[5],
     net1329[6], net1329[7]}), .slf_op_06({net1328[0], net1328[1],
     net1328[2], net1328[3], net1328[4], net1328[5], net1328[6],
     net1328[7]}), .slf_op_07({net1327[0], net1327[1], net1327[2],
     net1327[3], net1327[4], net1327[5], net1327[6], net1327[7]}),
     .slf_op_08(slf_op_01_08[7:0]), .rgt_op_08(slf_op_02_08[7:0]),
     .rgt_op_07({net852[0], net852[1], net852[2], net852[3], net852[4],
     net852[5], net852[6], net852[7]}), .rgt_op_06({net853[0],
     net853[1], net853[2], net853[3], net853[4], net853[5], net853[6],
     net853[7]}), .rgt_op_05({net854[0], net854[1], net854[2],
     net854[3], net854[4], net854[5], net854[6], net854[7]}),
     .lft_op_08({slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0], slf_op_00_08[3], slf_op_00_08[2],
     slf_op_00_08[1], slf_op_00_08[0]}), .lft_op_07({slf_op_00_07[3],
     slf_op_00_07[2], slf_op_00_07[1], slf_op_00_07[0],
     slf_op_00_07[3], slf_op_00_07[2], slf_op_00_07[1],
     slf_op_00_07[0]}), .lft_op_06({slf_op_00_06[3], slf_op_00_06[2],
     slf_op_00_06[1], slf_op_00_06[0], slf_op_00_06[3],
     slf_op_00_06[2], slf_op_00_06[1], slf_op_00_06[0]}),
     .lft_op_05({slf_op_00_05[3], slf_op_00_05[2], slf_op_00_05[1],
     slf_op_00_05[0], slf_op_00_05[3], slf_op_00_05[2],
     slf_op_00_05[1], slf_op_00_05[0]}), .sp12_h_l_08({net1342[0],
     net1342[1], net1342[2], net1342[3], net1342[4], net1342[5],
     net1342[6], net1342[7], net1342[8], net1342[9], net1342[10],
     net1342[11], net1342[12], net1342[13], net1342[14], net1342[15],
     net1342[16], net1342[17], net1342[18], net1342[19], net1342[20],
     net1342[21], net1342[22], net1342[23]}), .sp12_h_l_07({net1350[0],
     net1350[1], net1350[2], net1350[3], net1350[4], net1350[5],
     net1350[6], net1350[7], net1350[8], net1350[9], net1350[10],
     net1350[11], net1350[12], net1350[13], net1350[14], net1350[15],
     net1350[16], net1350[17], net1350[18], net1350[19], net1350[20],
     net1350[21], net1350[22], net1350[23]}), .sp12_h_l_06({net1343[0],
     net1343[1], net1343[2], net1343[3], net1343[4], net1343[5],
     net1343[6], net1343[7], net1343[8], net1343[9], net1343[10],
     net1343[11], net1343[12], net1343[13], net1343[14], net1343[15],
     net1343[16], net1343[17], net1343[18], net1343[19], net1343[20],
     net1343[21], net1343[22], net1343[23]}), .sp12_h_r_05({net862[0],
     net862[1], net862[2], net862[3], net862[4], net862[5], net862[6],
     net862[7], net862[8], net862[9], net862[10], net862[11],
     net862[12], net862[13], net862[14], net862[15], net862[16],
     net862[17], net862[18], net862[19], net862[20], net862[21],
     net862[22], net862[23]}), .sp12_h_r_06({net863[0], net863[1],
     net863[2], net863[3], net863[4], net863[5], net863[6], net863[7],
     net863[8], net863[9], net863[10], net863[11], net863[12],
     net863[13], net863[14], net863[15], net863[16], net863[17],
     net863[18], net863[19], net863[20], net863[21], net863[22],
     net863[23]}), .sp12_h_r_07({net864[0], net864[1], net864[2],
     net864[3], net864[4], net864[5], net864[6], net864[7], net864[8],
     net864[9], net864[10], net864[11], net864[12], net864[13],
     net864[14], net864[15], net864[16], net864[17], net864[18],
     net864[19], net864[20], net864[21], net864[22], net864[23]}),
     .sp12_h_r_08({net865[0], net865[1], net865[2], net865[3],
     net865[4], net865[5], net865[6], net865[7], net865[8], net865[9],
     net865[10], net865[11], net865[12], net865[13], net865[14],
     net865[15], net865[16], net865[17], net865[18], net865[19],
     net865[20], net865[21], net865[22], net865[23]}),
     .sp12_h_l_05({net1345[0], net1345[1], net1345[2], net1345[3],
     net1345[4], net1345[5], net1345[6], net1345[7], net1345[8],
     net1345[9], net1345[10], net1345[11], net1345[12], net1345[13],
     net1345[14], net1345[15], net1345[16], net1345[17], net1345[18],
     net1345[19], net1345[20], net1345[21], net1345[22], net1345[23]}),
     .sp4_r_v_b_05({net867[0], net867[1], net867[2], net867[3],
     net867[4], net867[5], net867[6], net867[7], net867[8], net867[9],
     net867[10], net867[11], net867[12], net867[13], net867[14],
     net867[15], net867[16], net867[17], net867[18], net867[19],
     net867[20], net867[21], net867[22], net867[23], net867[24],
     net867[25], net867[26], net867[27], net867[28], net867[29],
     net867[30], net867[31], net867[32], net867[33], net867[34],
     net867[35], net867[36], net867[37], net867[38], net867[39],
     net867[40], net867[41], net867[42], net867[43], net867[44],
     net867[45], net867[46], net867[47]}), .sp4_r_v_b_06({net868[0],
     net868[1], net868[2], net868[3], net868[4], net868[5], net868[6],
     net868[7], net868[8], net868[9], net868[10], net868[11],
     net868[12], net868[13], net868[14], net868[15], net868[16],
     net868[17], net868[18], net868[19], net868[20], net868[21],
     net868[22], net868[23], net868[24], net868[25], net868[26],
     net868[27], net868[28], net868[29], net868[30], net868[31],
     net868[32], net868[33], net868[34], net868[35], net868[36],
     net868[37], net868[38], net868[39], net868[40], net868[41],
     net868[42], net868[43], net868[44], net868[45], net868[46],
     net868[47]}), .sp4_r_v_b_07({net869[0], net869[1], net869[2],
     net869[3], net869[4], net869[5], net869[6], net869[7], net869[8],
     net869[9], net869[10], net869[11], net869[12], net869[13],
     net869[14], net869[15], net869[16], net869[17], net869[18],
     net869[19], net869[20], net869[21], net869[22], net869[23],
     net869[24], net869[25], net869[26], net869[27], net869[28],
     net869[29], net869[30], net869[31], net869[32], net869[33],
     net869[34], net869[35], net869[36], net869[37], net869[38],
     net869[39], net869[40], net869[41], net869[42], net869[43],
     net869[44], net869[45], net869[46], net869[47]}),
     .sp4_r_v_b_08({net870[0], net870[1], net870[2], net870[3],
     net870[4], net870[5], net870[6], net870[7], net870[8], net870[9],
     net870[10], net870[11], net870[12], net870[13], net870[14],
     net870[15], net870[16], net870[17], net870[18], net870[19],
     net870[20], net870[21], net870[22], net870[23], net870[24],
     net870[25], net870[26], net870[27], net870[28], net870[29],
     net870[30], net870[31], net870[32], net870[33], net870[34],
     net870[35], net870[36], net870[37], net870[38], net870[39],
     net870[40], net870[41], net870[42], net870[43], net870[44],
     net870[45], net870[46], net870[47]}), .sp4_v_b_08({net871[0],
     net871[1], net871[2], net871[3], net871[4], net871[5], net871[6],
     net871[7], net871[8], net871[9], net871[10], net871[11],
     net871[12], net871[13], net871[14], net871[15], net871[16],
     net871[17], net871[18], net871[19], net871[20], net871[21],
     net871[22], net871[23], net871[24], net871[25], net871[26],
     net871[27], net871[28], net871[29], net871[30], net871[31],
     net871[32], net871[33], net871[34], net871[35], net871[36],
     net871[37], net871[38], net871[39], net871[40], net871[41],
     net871[42], net871[43], net871[44], net871[45], net871[46],
     net871[47]}), .sp4_v_b_07({net872[0], net872[1], net872[2],
     net872[3], net872[4], net872[5], net872[6], net872[7], net872[8],
     net872[9], net872[10], net872[11], net872[12], net872[13],
     net872[14], net872[15], net872[16], net872[17], net872[18],
     net872[19], net872[20], net872[21], net872[22], net872[23],
     net872[24], net872[25], net872[26], net872[27], net872[28],
     net872[29], net872[30], net872[31], net872[32], net872[33],
     net872[34], net872[35], net872[36], net872[37], net872[38],
     net872[39], net872[40], net872[41], net872[42], net872[43],
     net872[44], net872[45], net872[46], net872[47]}),
     .sp4_v_b_06({net1430[0], net1430[1], net1430[2], net1430[3],
     net1430[4], net1430[5], net1430[6], net1430[7], net1430[8],
     net1430[9], net1430[10], net1430[11], net1430[12], net1430[13],
     net1430[14], net1430[15], net1430[16], net1430[17], net1430[18],
     net1430[19], net1430[20], net1430[21], net1430[22], net1430[23],
     net1430[24], net1430[25], net1430[26], net1430[27], net1430[28],
     net1430[29], net1430[30], net1430[31], net1430[32], net1430[33],
     net1430[34], net1430[35], net1430[36], net1430[37], net1430[38],
     net1430[39], net1430[40], net1430[41], net1430[42], net1430[43],
     net1430[44], net1430[45], net1430[46], net1430[47]}),
     .sp4_v_b_05({net1436[0], net1436[1], net1436[2], net1436[3],
     net1436[4], net1436[5], net1436[6], net1436[7], net1436[8],
     net1436[9], net1436[10], net1436[11], net1436[12], net1436[13],
     net1436[14], net1436[15], net1436[16], net1436[17], net1436[18],
     net1436[19], net1436[20], net1436[21], net1436[22], net1436[23],
     net1436[24], net1436[25], net1436[26], net1436[27], net1436[28],
     net1436[29], net1436[30], net1436[31], net1436[32], net1436[33],
     net1436[34], net1436[35], net1436[36], net1436[37], net1436[38],
     net1436[39], net1436[40], net1436[41], net1436[42], net1436[43],
     net1436[44], net1436[45], net1436[46], net1436[47]}),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .wl(wl_l[143:16]), .sp12_v_t_08(sp12_v_t_01_08[23:0]),
     .tnr_op_08(tnr_op_01_08[7:0]), .top_op_08(top_op_01_08[7:0]),
     .tnl_op_08(tnl_op_01_08[7:0]), .sp4_v_t_08(sp4_v_t_01_08[47:0]),
     .lc_bot(tiegnd_bl), .op_vic(op_vic_01_08),
     .sp12_v_b_01({net1373[0], net1373[1], net1373[2], net1373[3],
     net1373[4], net1373[5], net1373[6], net1373[7], net1373[8],
     net1373[9], net1373[10], net1373[11], net1373[12], net1373[13],
     net1373[14], net1373[15], net1373[16], net1373[17], net1373[18],
     net1373[19], net1373[20], net1373[21], net1373[22],
     net1373[23]}));
lt_1x8_bot_ice1f I_lt_col_t06 ( .glb_netwk_bot({net1383[0], net1383[1],
     net1383[2], net1383[3], net1383[4], net1383[5], net1383[6],
     net1383[7]}), .rgt_op_03(rgt_op_06_03[7:0]),
     .slf_op_02(slf_op_06_02[7:0]), .rgt_op_02(rgt_op_06_02[7:0]),
     .rgt_op_01(rgt_op_06_01[7:0]), .purst(purst), .prog(prog),
     .lft_op_04({net991[0], net991[1], net991[2], net991[3], net991[4],
     net991[5], net991[6], net991[7]}), .lft_op_03({net981[0],
     net981[1], net981[2], net981[3], net981[4], net981[5], net981[6],
     net981[7]}), .lft_op_02({net983[0], net983[1], net983[2],
     net983[3], net983[4], net983[5], net983[6], net983[7]}),
     .lft_op_01({net1409[0], net1409[1], net1409[2], net1409[3],
     net1409[4], net1409[5], net1409[6], net1409[7]}),
     .rgt_op_04(rgt_op_06_04[7:0]), .carry_in(tiegnd_bl),
     .bnl_op_01({slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0], slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0]}), .slf_op_04(slf_op_06_04[7:0]),
     .slf_op_03(slf_op_06_03[7:0]), .slf_op_01(slf_op_06_01[7:0]),
     .sp4_h_l_04({net1104[0], net1104[1], net1104[2], net1104[3],
     net1104[4], net1104[5], net1104[6], net1104[7], net1104[8],
     net1104[9], net1104[10], net1104[11], net1104[12], net1104[13],
     net1104[14], net1104[15], net1104[16], net1104[17], net1104[18],
     net1104[19], net1104[20], net1104[21], net1104[22], net1104[23],
     net1104[24], net1104[25], net1104[26], net1104[27], net1104[28],
     net1104[29], net1104[30], net1104[31], net1104[32], net1104[33],
     net1104[34], net1104[35], net1104[36], net1104[37], net1104[38],
     net1104[39], net1104[40], net1104[41], net1104[42], net1104[43],
     net1104[44], net1104[45], net1104[46], net1104[47]}),
     .carry_out(carry_out_06_08), .vdd_cntl(vdd_cntl_l[143:16]),
     .sp12_h_r_04(sp12_h_r_06_04[23:0]),
     .sp12_h_r_03(sp12_h_r_06_03[23:0]),
     .sp12_h_r_02(sp12_h_r_06_02[23:0]),
     .sp12_h_r_01(sp12_h_r_06_01[23:0]), .glb_netwk_col({net1344[0],
     net1344[1], net1344[2], net1344[3], net1344[4], net1344[5],
     net1344[6], net1344[7]}), .sp4_v_b_01({net1406[0], net1406[1],
     net1406[2], net1406[3], net1406[4], net1406[5], net1406[6],
     net1406[7], net1406[8], net1406[9], net1406[10], net1406[11],
     net1406[12], net1406[13], net1406[14], net1406[15], net1406[16],
     net1406[17], net1406[18], net1406[19], net1406[20], net1406[21],
     net1406[22], net1406[23], net1406[24], net1406[25], net1406[26],
     net1406[27], net1406[28], net1406[29], net1406[30], net1406[31],
     net1406[32], net1406[33], net1406[34], net1406[35], net1406[36],
     net1406[37], net1406[38], net1406[39], net1406[40], net1406[41],
     net1406[42], net1406[43], net1406[44], net1406[45], net1406[46],
     net1406[47]}), .sp4_r_v_b_04(sp4_r_v_b_06_04[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_06_03[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_06_02[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_06_01[47:0]),
     .sp4_h_r_04(sp4_h_r_06_04[47:0]),
     .sp4_h_r_03(sp4_h_r_06_03[47:0]),
     .sp4_h_r_02(sp4_h_r_06_02[47:0]),
     .sp4_h_r_01(sp4_h_r_06_01[47:0]), .sp4_h_l_03({net1105[0],
     net1105[1], net1105[2], net1105[3], net1105[4], net1105[5],
     net1105[6], net1105[7], net1105[8], net1105[9], net1105[10],
     net1105[11], net1105[12], net1105[13], net1105[14], net1105[15],
     net1105[16], net1105[17], net1105[18], net1105[19], net1105[20],
     net1105[21], net1105[22], net1105[23], net1105[24], net1105[25],
     net1105[26], net1105[27], net1105[28], net1105[29], net1105[30],
     net1105[31], net1105[32], net1105[33], net1105[34], net1105[35],
     net1105[36], net1105[37], net1105[38], net1105[39], net1105[40],
     net1105[41], net1105[42], net1105[43], net1105[44], net1105[45],
     net1105[46], net1105[47]}), .sp4_h_l_02({net1106[0], net1106[1],
     net1106[2], net1106[3], net1106[4], net1106[5], net1106[6],
     net1106[7], net1106[8], net1106[9], net1106[10], net1106[11],
     net1106[12], net1106[13], net1106[14], net1106[15], net1106[16],
     net1106[17], net1106[18], net1106[19], net1106[20], net1106[21],
     net1106[22], net1106[23], net1106[24], net1106[25], net1106[26],
     net1106[27], net1106[28], net1106[29], net1106[30], net1106[31],
     net1106[32], net1106[33], net1106[34], net1106[35], net1106[36],
     net1106[37], net1106[38], net1106[39], net1106[40], net1106[41],
     net1106[42], net1106[43], net1106[44], net1106[45], net1106[46],
     net1106[47]}), .sp4_h_l_01({net1107[0], net1107[1], net1107[2],
     net1107[3], net1107[4], net1107[5], net1107[6], net1107[7],
     net1107[8], net1107[9], net1107[10], net1107[11], net1107[12],
     net1107[13], net1107[14], net1107[15], net1107[16], net1107[17],
     net1107[18], net1107[19], net1107[20], net1107[21], net1107[22],
     net1107[23], net1107[24], net1107[25], net1107[26], net1107[27],
     net1107[28], net1107[29], net1107[30], net1107[31], net1107[32],
     net1107[33], net1107[34], net1107[35], net1107[36], net1107[37],
     net1107[38], net1107[39], net1107[40], net1107[41], net1107[42],
     net1107[43], net1107[44], net1107[45], net1107[46], net1107[47]}),
     .bl(bl[329:276]), .bot_op_01({slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0], slf_op_06_00[3],
     slf_op_06_00[2], slf_op_06_00[1], slf_op_06_00[0]}),
     .sp12_h_l_01({net1097[0], net1097[1], net1097[2], net1097[3],
     net1097[4], net1097[5], net1097[6], net1097[7], net1097[8],
     net1097[9], net1097[10], net1097[11], net1097[12], net1097[13],
     net1097[14], net1097[15], net1097[16], net1097[17], net1097[18],
     net1097[19], net1097[20], net1097[21], net1097[22], net1097[23]}),
     .sp12_h_l_02({net1096[0], net1096[1], net1096[2], net1096[3],
     net1096[4], net1096[5], net1096[6], net1096[7], net1096[8],
     net1096[9], net1096[10], net1096[11], net1096[12], net1096[13],
     net1096[14], net1096[15], net1096[16], net1096[17], net1096[18],
     net1096[19], net1096[20], net1096[21], net1096[22], net1096[23]}),
     .sp12_h_l_03({net1095[0], net1095[1], net1095[2], net1095[3],
     net1095[4], net1095[5], net1095[6], net1095[7], net1095[8],
     net1095[9], net1095[10], net1095[11], net1095[12], net1095[13],
     net1095[14], net1095[15], net1095[16], net1095[17], net1095[18],
     net1095[19], net1095[20], net1095[21], net1095[22], net1095[23]}),
     .sp12_h_l_04({net1094[0], net1094[1], net1094[2], net1094[3],
     net1094[4], net1094[5], net1094[6], net1094[7], net1094[8],
     net1094[9], net1094[10], net1094[11], net1094[12], net1094[13],
     net1094[14], net1094[15], net1094[16], net1094[17], net1094[18],
     net1094[19], net1094[20], net1094[21], net1094[22], net1094[23]}),
     .sp4_v_b_04({net1100[0], net1100[1], net1100[2], net1100[3],
     net1100[4], net1100[5], net1100[6], net1100[7], net1100[8],
     net1100[9], net1100[10], net1100[11], net1100[12], net1100[13],
     net1100[14], net1100[15], net1100[16], net1100[17], net1100[18],
     net1100[19], net1100[20], net1100[21], net1100[22], net1100[23],
     net1100[24], net1100[25], net1100[26], net1100[27], net1100[28],
     net1100[29], net1100[30], net1100[31], net1100[32], net1100[33],
     net1100[34], net1100[35], net1100[36], net1100[37], net1100[38],
     net1100[39], net1100[40], net1100[41], net1100[42], net1100[43],
     net1100[44], net1100[45], net1100[46], net1100[47]}),
     .sp4_v_b_03({net1101[0], net1101[1], net1101[2], net1101[3],
     net1101[4], net1101[5], net1101[6], net1101[7], net1101[8],
     net1101[9], net1101[10], net1101[11], net1101[12], net1101[13],
     net1101[14], net1101[15], net1101[16], net1101[17], net1101[18],
     net1101[19], net1101[20], net1101[21], net1101[22], net1101[23],
     net1101[24], net1101[25], net1101[26], net1101[27], net1101[28],
     net1101[29], net1101[30], net1101[31], net1101[32], net1101[33],
     net1101[34], net1101[35], net1101[36], net1101[37], net1101[38],
     net1101[39], net1101[40], net1101[41], net1101[42], net1101[43],
     net1101[44], net1101[45], net1101[46], net1101[47]}),
     .sp4_v_b_02({net1102[0], net1102[1], net1102[2], net1102[3],
     net1102[4], net1102[5], net1102[6], net1102[7], net1102[8],
     net1102[9], net1102[10], net1102[11], net1102[12], net1102[13],
     net1102[14], net1102[15], net1102[16], net1102[17], net1102[18],
     net1102[19], net1102[20], net1102[21], net1102[22], net1102[23],
     net1102[24], net1102[25], net1102[26], net1102[27], net1102[28],
     net1102[29], net1102[30], net1102[31], net1102[32], net1102[33],
     net1102[34], net1102[35], net1102[36], net1102[37], net1102[38],
     net1102[39], net1102[40], net1102[41], net1102[42], net1102[43],
     net1102[44], net1102[45], net1102[46], net1102[47]}),
     .bnr_op_01({bnr_op_06_01[3], bnr_op_06_01[2], bnr_op_06_01[1],
     bnr_op_06_01[0], bnr_op_06_01[3], bnr_op_06_01[2],
     bnr_op_06_01[1], bnr_op_06_01[0]}), .sp4_h_l_05({net1128[0],
     net1128[1], net1128[2], net1128[3], net1128[4], net1128[5],
     net1128[6], net1128[7], net1128[8], net1128[9], net1128[10],
     net1128[11], net1128[12], net1128[13], net1128[14], net1128[15],
     net1128[16], net1128[17], net1128[18], net1128[19], net1128[20],
     net1128[21], net1128[22], net1128[23], net1128[24], net1128[25],
     net1128[26], net1128[27], net1128[28], net1128[29], net1128[30],
     net1128[31], net1128[32], net1128[33], net1128[34], net1128[35],
     net1128[36], net1128[37], net1128[38], net1128[39], net1128[40],
     net1128[41], net1128[42], net1128[43], net1128[44], net1128[45],
     net1128[46], net1128[47]}), .sp4_h_l_06({net1127[0], net1127[1],
     net1127[2], net1127[3], net1127[4], net1127[5], net1127[6],
     net1127[7], net1127[8], net1127[9], net1127[10], net1127[11],
     net1127[12], net1127[13], net1127[14], net1127[15], net1127[16],
     net1127[17], net1127[18], net1127[19], net1127[20], net1127[21],
     net1127[22], net1127[23], net1127[24], net1127[25], net1127[26],
     net1127[27], net1127[28], net1127[29], net1127[30], net1127[31],
     net1127[32], net1127[33], net1127[34], net1127[35], net1127[36],
     net1127[37], net1127[38], net1127[39], net1127[40], net1127[41],
     net1127[42], net1127[43], net1127[44], net1127[45], net1127[46],
     net1127[47]}), .sp4_h_l_07({net1126[0], net1126[1], net1126[2],
     net1126[3], net1126[4], net1126[5], net1126[6], net1126[7],
     net1126[8], net1126[9], net1126[10], net1126[11], net1126[12],
     net1126[13], net1126[14], net1126[15], net1126[16], net1126[17],
     net1126[18], net1126[19], net1126[20], net1126[21], net1126[22],
     net1126[23], net1126[24], net1126[25], net1126[26], net1126[27],
     net1126[28], net1126[29], net1126[30], net1126[31], net1126[32],
     net1126[33], net1126[34], net1126[35], net1126[36], net1126[37],
     net1126[38], net1126[39], net1126[40], net1126[41], net1126[42],
     net1126[43], net1126[44], net1126[45], net1126[46], net1126[47]}),
     .sp4_h_l_08({net1125[0], net1125[1], net1125[2], net1125[3],
     net1125[4], net1125[5], net1125[6], net1125[7], net1125[8],
     net1125[9], net1125[10], net1125[11], net1125[12], net1125[13],
     net1125[14], net1125[15], net1125[16], net1125[17], net1125[18],
     net1125[19], net1125[20], net1125[21], net1125[22], net1125[23],
     net1125[24], net1125[25], net1125[26], net1125[27], net1125[28],
     net1125[29], net1125[30], net1125[31], net1125[32], net1125[33],
     net1125[34], net1125[35], net1125[36], net1125[37], net1125[38],
     net1125[39], net1125[40], net1125[41], net1125[42], net1125[43],
     net1125[44], net1125[45], net1125[46], net1125[47]}),
     .sp4_h_r_08(sp4_h_r_06_08[47:0]),
     .sp4_h_r_07(sp4_h_r_06_07[47:0]),
     .sp4_h_r_06(sp4_h_r_06_06[47:0]),
     .sp4_h_r_05(sp4_h_r_06_05[47:0]), .slf_op_05(slf_op_06_05[7:0]),
     .slf_op_06(slf_op_06_06[7:0]), .slf_op_07(slf_op_06_07[7:0]),
     .slf_op_08(slf_op_06_08[7:0]), .rgt_op_08(rgt_op_06_08[7:0]),
     .rgt_op_07(rgt_op_06_07[7:0]), .rgt_op_06(rgt_op_06_06[7:0]),
     .rgt_op_05(rgt_op_06_05[7:0]), .lft_op_08(slf_op_05_08[7:0]),
     .lft_op_07({net1040[0], net1040[1], net1040[2], net1040[3],
     net1040[4], net1040[5], net1040[6], net1040[7]}),
     .lft_op_06({net1041[0], net1041[1], net1041[2], net1041[3],
     net1041[4], net1041[5], net1041[6], net1041[7]}),
     .lft_op_05({net1042[0], net1042[1], net1042[2], net1042[3],
     net1042[4], net1042[5], net1042[6], net1042[7]}),
     .sp12_h_l_08({net1147[0], net1147[1], net1147[2], net1147[3],
     net1147[4], net1147[5], net1147[6], net1147[7], net1147[8],
     net1147[9], net1147[10], net1147[11], net1147[12], net1147[13],
     net1147[14], net1147[15], net1147[16], net1147[17], net1147[18],
     net1147[19], net1147[20], net1147[21], net1147[22], net1147[23]}),
     .sp12_h_l_07({net1146[0], net1146[1], net1146[2], net1146[3],
     net1146[4], net1146[5], net1146[6], net1146[7], net1146[8],
     net1146[9], net1146[10], net1146[11], net1146[12], net1146[13],
     net1146[14], net1146[15], net1146[16], net1146[17], net1146[18],
     net1146[19], net1146[20], net1146[21], net1146[22], net1146[23]}),
     .sp12_h_l_06({net1145[0], net1145[1], net1145[2], net1145[3],
     net1145[4], net1145[5], net1145[6], net1145[7], net1145[8],
     net1145[9], net1145[10], net1145[11], net1145[12], net1145[13],
     net1145[14], net1145[15], net1145[16], net1145[17], net1145[18],
     net1145[19], net1145[20], net1145[21], net1145[22], net1145[23]}),
     .sp12_h_r_05(sp12_h_r_06_05[23:0]),
     .sp12_h_r_06(sp12_h_r_06_06[23:0]),
     .sp12_h_r_07(sp12_h_r_06_07[23:0]),
     .sp12_h_r_08(sp12_h_r_06_08[23:0]), .sp12_h_l_05({net1144[0],
     net1144[1], net1144[2], net1144[3], net1144[4], net1144[5],
     net1144[6], net1144[7], net1144[8], net1144[9], net1144[10],
     net1144[11], net1144[12], net1144[13], net1144[14], net1144[15],
     net1144[16], net1144[17], net1144[18], net1144[19], net1144[20],
     net1144[21], net1144[22], net1144[23]}),
     .sp4_r_v_b_05(sp4_r_v_b_06_05[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_06_06[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_06_07[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_06_08[47:0]), .sp4_v_b_08({net1152[0],
     net1152[1], net1152[2], net1152[3], net1152[4], net1152[5],
     net1152[6], net1152[7], net1152[8], net1152[9], net1152[10],
     net1152[11], net1152[12], net1152[13], net1152[14], net1152[15],
     net1152[16], net1152[17], net1152[18], net1152[19], net1152[20],
     net1152[21], net1152[22], net1152[23], net1152[24], net1152[25],
     net1152[26], net1152[27], net1152[28], net1152[29], net1152[30],
     net1152[31], net1152[32], net1152[33], net1152[34], net1152[35],
     net1152[36], net1152[37], net1152[38], net1152[39], net1152[40],
     net1152[41], net1152[42], net1152[43], net1152[44], net1152[45],
     net1152[46], net1152[47]}), .sp4_v_b_07({net1151[0], net1151[1],
     net1151[2], net1151[3], net1151[4], net1151[5], net1151[6],
     net1151[7], net1151[8], net1151[9], net1151[10], net1151[11],
     net1151[12], net1151[13], net1151[14], net1151[15], net1151[16],
     net1151[17], net1151[18], net1151[19], net1151[20], net1151[21],
     net1151[22], net1151[23], net1151[24], net1151[25], net1151[26],
     net1151[27], net1151[28], net1151[29], net1151[30], net1151[31],
     net1151[32], net1151[33], net1151[34], net1151[35], net1151[36],
     net1151[37], net1151[38], net1151[39], net1151[40], net1151[41],
     net1151[42], net1151[43], net1151[44], net1151[45], net1151[46],
     net1151[47]}), .sp4_v_b_06({net1150[0], net1150[1], net1150[2],
     net1150[3], net1150[4], net1150[5], net1150[6], net1150[7],
     net1150[8], net1150[9], net1150[10], net1150[11], net1150[12],
     net1150[13], net1150[14], net1150[15], net1150[16], net1150[17],
     net1150[18], net1150[19], net1150[20], net1150[21], net1150[22],
     net1150[23], net1150[24], net1150[25], net1150[26], net1150[27],
     net1150[28], net1150[29], net1150[30], net1150[31], net1150[32],
     net1150[33], net1150[34], net1150[35], net1150[36], net1150[37],
     net1150[38], net1150[39], net1150[40], net1150[41], net1150[42],
     net1150[43], net1150[44], net1150[45], net1150[46], net1150[47]}),
     .sp4_v_b_05({net1149[0], net1149[1], net1149[2], net1149[3],
     net1149[4], net1149[5], net1149[6], net1149[7], net1149[8],
     net1149[9], net1149[10], net1149[11], net1149[12], net1149[13],
     net1149[14], net1149[15], net1149[16], net1149[17], net1149[18],
     net1149[19], net1149[20], net1149[21], net1149[22], net1149[23],
     net1149[24], net1149[25], net1149[26], net1149[27], net1149[28],
     net1149[29], net1149[30], net1149[31], net1149[32], net1149[33],
     net1149[34], net1149[35], net1149[36], net1149[37], net1149[38],
     net1149[39], net1149[40], net1149[41], net1149[42], net1149[43],
     net1149[44], net1149[45], net1149[46], net1149[47]}),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .wl(wl_l[143:16]), .sp12_v_t_08(sp12_v_t_06_08[23:0]),
     .tnr_op_08(tnr_op_06_08[7:0]), .top_op_08(top_op_06_08[7:0]),
     .tnl_op_08(tnl_op_06_08[7:0]), .sp4_v_t_08(sp4_v_t_06_08[47:0]),
     .lc_bot(tiegnd_bl), .op_vic(op_vic_06_08),
     .sp12_v_b_01({net1407[0], net1407[1], net1407[2], net1407[3],
     net1407[4], net1407[5], net1407[6], net1407[7], net1407[8],
     net1407[9], net1407[10], net1407[11], net1407[12], net1407[13],
     net1407[14], net1407[15], net1407[16], net1407[17], net1407[18],
     net1407[19], net1407[20], net1407[21], net1407[22],
     net1407[23]}));
lt_1x8_bot_ice1f I_lt_col_t04 ( .glb_netwk_bot({net1385[0], net1385[1],
     net1385[2], net1385[3], net1385[4], net1385[5], net1385[6],
     net1385[7]}), .rgt_op_03({net981[0], net981[1], net981[2],
     net981[3], net981[4], net981[5], net981[6], net981[7]}),
     .slf_op_02({net1269[0], net1269[1], net1269[2], net1269[3],
     net1269[4], net1269[5], net1269[6], net1269[7]}),
     .rgt_op_02({net983[0], net983[1], net983[2], net983[3], net983[4],
     net983[5], net983[6], net983[7]}), .rgt_op_01({net1409[0],
     net1409[1], net1409[2], net1409[3], net1409[4], net1409[5],
     net1409[6], net1409[7]}), .purst(purst), .prog(prog),
     .lft_op_04({net708[0], net708[1], net708[2], net708[3], net708[4],
     net708[5], net708[6], net708[7]}), .lft_op_03({net698[0],
     net698[1], net698[2], net698[3], net698[4], net698[5], net698[6],
     net698[7]}), .lft_op_02({net700[0], net700[1], net700[2],
     net700[3], net700[4], net700[5], net700[6], net700[7]}),
     .lft_op_01({net1410[0], net1410[1], net1410[2], net1410[3],
     net1410[4], net1410[5], net1410[6], net1410[7]}),
     .rgt_op_04({net991[0], net991[1], net991[2], net991[3], net991[4],
     net991[5], net991[6], net991[7]}), .carry_in(tiegnd_bl),
     .bnl_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .slf_op_04({net1267[0],
     net1267[1], net1267[2], net1267[3], net1267[4], net1267[5],
     net1267[6], net1267[7]}), .slf_op_03({net1268[0], net1268[1],
     net1268[2], net1268[3], net1268[4], net1268[5], net1268[6],
     net1268[7]}), .slf_op_01({net1408[0], net1408[1], net1408[2],
     net1408[3], net1408[4], net1408[5], net1408[6], net1408[7]}),
     .sp4_h_l_04({net1288[0], net1288[1], net1288[2], net1288[3],
     net1288[4], net1288[5], net1288[6], net1288[7], net1288[8],
     net1288[9], net1288[10], net1288[11], net1288[12], net1288[13],
     net1288[14], net1288[15], net1288[16], net1288[17], net1288[18],
     net1288[19], net1288[20], net1288[21], net1288[22], net1288[23],
     net1288[24], net1288[25], net1288[26], net1288[27], net1288[28],
     net1288[29], net1288[30], net1288[31], net1288[32], net1288[33],
     net1288[34], net1288[35], net1288[36], net1288[37], net1288[38],
     net1288[39], net1288[40], net1288[41], net1288[42], net1288[43],
     net1288[44], net1288[45], net1288[46], net1288[47]}),
     .carry_out(carry_out_04_08), .vdd_cntl(vdd_cntl_l[143:16]),
     .sp12_h_r_04({net1000[0], net1000[1], net1000[2], net1000[3],
     net1000[4], net1000[5], net1000[6], net1000[7], net1000[8],
     net1000[9], net1000[10], net1000[11], net1000[12], net1000[13],
     net1000[14], net1000[15], net1000[16], net1000[17], net1000[18],
     net1000[19], net1000[20], net1000[21], net1000[22], net1000[23]}),
     .sp12_h_r_03({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7], net1001[8],
     net1001[9], net1001[10], net1001[11], net1001[12], net1001[13],
     net1001[14], net1001[15], net1001[16], net1001[17], net1001[18],
     net1001[19], net1001[20], net1001[21], net1001[22], net1001[23]}),
     .sp12_h_r_02({net1002[0], net1002[1], net1002[2], net1002[3],
     net1002[4], net1002[5], net1002[6], net1002[7], net1002[8],
     net1002[9], net1002[10], net1002[11], net1002[12], net1002[13],
     net1002[14], net1002[15], net1002[16], net1002[17], net1002[18],
     net1002[19], net1002[20], net1002[21], net1002[22], net1002[23]}),
     .sp12_h_r_01({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7], net1003[8],
     net1003[9], net1003[10], net1003[11], net1003[12], net1003[13],
     net1003[14], net1003[15], net1003[16], net1003[17], net1003[18],
     net1003[19], net1003[20], net1003[21], net1003[22], net1003[23]}),
     .glb_netwk_col({net1344[0], net1344[1], net1344[2], net1344[3],
     net1344[4], net1344[5], net1344[6], net1344[7]}),
     .sp4_v_b_01({net1414[0], net1414[1], net1414[2], net1414[3],
     net1414[4], net1414[5], net1414[6], net1414[7], net1414[8],
     net1414[9], net1414[10], net1414[11], net1414[12], net1414[13],
     net1414[14], net1414[15], net1414[16], net1414[17], net1414[18],
     net1414[19], net1414[20], net1414[21], net1414[22], net1414[23],
     net1414[24], net1414[25], net1414[26], net1414[27], net1414[28],
     net1414[29], net1414[30], net1414[31], net1414[32], net1414[33],
     net1414[34], net1414[35], net1414[36], net1414[37], net1414[38],
     net1414[39], net1414[40], net1414[41], net1414[42], net1414[43],
     net1414[44], net1414[45], net1414[46], net1414[47]}),
     .sp4_r_v_b_04({net1006[0], net1006[1], net1006[2], net1006[3],
     net1006[4], net1006[5], net1006[6], net1006[7], net1006[8],
     net1006[9], net1006[10], net1006[11], net1006[12], net1006[13],
     net1006[14], net1006[15], net1006[16], net1006[17], net1006[18],
     net1006[19], net1006[20], net1006[21], net1006[22], net1006[23],
     net1006[24], net1006[25], net1006[26], net1006[27], net1006[28],
     net1006[29], net1006[30], net1006[31], net1006[32], net1006[33],
     net1006[34], net1006[35], net1006[36], net1006[37], net1006[38],
     net1006[39], net1006[40], net1006[41], net1006[42], net1006[43],
     net1006[44], net1006[45], net1006[46], net1006[47]}),
     .sp4_r_v_b_03({net1007[0], net1007[1], net1007[2], net1007[3],
     net1007[4], net1007[5], net1007[6], net1007[7], net1007[8],
     net1007[9], net1007[10], net1007[11], net1007[12], net1007[13],
     net1007[14], net1007[15], net1007[16], net1007[17], net1007[18],
     net1007[19], net1007[20], net1007[21], net1007[22], net1007[23],
     net1007[24], net1007[25], net1007[26], net1007[27], net1007[28],
     net1007[29], net1007[30], net1007[31], net1007[32], net1007[33],
     net1007[34], net1007[35], net1007[36], net1007[37], net1007[38],
     net1007[39], net1007[40], net1007[41], net1007[42], net1007[43],
     net1007[44], net1007[45], net1007[46], net1007[47]}),
     .sp4_r_v_b_02({net1008[0], net1008[1], net1008[2], net1008[3],
     net1008[4], net1008[5], net1008[6], net1008[7], net1008[8],
     net1008[9], net1008[10], net1008[11], net1008[12], net1008[13],
     net1008[14], net1008[15], net1008[16], net1008[17], net1008[18],
     net1008[19], net1008[20], net1008[21], net1008[22], net1008[23],
     net1008[24], net1008[25], net1008[26], net1008[27], net1008[28],
     net1008[29], net1008[30], net1008[31], net1008[32], net1008[33],
     net1008[34], net1008[35], net1008[36], net1008[37], net1008[38],
     net1008[39], net1008[40], net1008[41], net1008[42], net1008[43],
     net1008[44], net1008[45], net1008[46], net1008[47]}),
     .sp4_r_v_b_01({net1402[0], net1402[1], net1402[2], net1402[3],
     net1402[4], net1402[5], net1402[6], net1402[7], net1402[8],
     net1402[9], net1402[10], net1402[11], net1402[12], net1402[13],
     net1402[14], net1402[15], net1402[16], net1402[17], net1402[18],
     net1402[19], net1402[20], net1402[21], net1402[22], net1402[23],
     net1402[24], net1402[25], net1402[26], net1402[27], net1402[28],
     net1402[29], net1402[30], net1402[31], net1402[32], net1402[33],
     net1402[34], net1402[35], net1402[36], net1402[37], net1402[38],
     net1402[39], net1402[40], net1402[41], net1402[42], net1402[43],
     net1402[44], net1402[45], net1402[46], net1402[47]}),
     .sp4_h_r_04({net1010[0], net1010[1], net1010[2], net1010[3],
     net1010[4], net1010[5], net1010[6], net1010[7], net1010[8],
     net1010[9], net1010[10], net1010[11], net1010[12], net1010[13],
     net1010[14], net1010[15], net1010[16], net1010[17], net1010[18],
     net1010[19], net1010[20], net1010[21], net1010[22], net1010[23],
     net1010[24], net1010[25], net1010[26], net1010[27], net1010[28],
     net1010[29], net1010[30], net1010[31], net1010[32], net1010[33],
     net1010[34], net1010[35], net1010[36], net1010[37], net1010[38],
     net1010[39], net1010[40], net1010[41], net1010[42], net1010[43],
     net1010[44], net1010[45], net1010[46], net1010[47]}),
     .sp4_h_r_03({net1011[0], net1011[1], net1011[2], net1011[3],
     net1011[4], net1011[5], net1011[6], net1011[7], net1011[8],
     net1011[9], net1011[10], net1011[11], net1011[12], net1011[13],
     net1011[14], net1011[15], net1011[16], net1011[17], net1011[18],
     net1011[19], net1011[20], net1011[21], net1011[22], net1011[23],
     net1011[24], net1011[25], net1011[26], net1011[27], net1011[28],
     net1011[29], net1011[30], net1011[31], net1011[32], net1011[33],
     net1011[34], net1011[35], net1011[36], net1011[37], net1011[38],
     net1011[39], net1011[40], net1011[41], net1011[42], net1011[43],
     net1011[44], net1011[45], net1011[46], net1011[47]}),
     .sp4_h_r_02({net1012[0], net1012[1], net1012[2], net1012[3],
     net1012[4], net1012[5], net1012[6], net1012[7], net1012[8],
     net1012[9], net1012[10], net1012[11], net1012[12], net1012[13],
     net1012[14], net1012[15], net1012[16], net1012[17], net1012[18],
     net1012[19], net1012[20], net1012[21], net1012[22], net1012[23],
     net1012[24], net1012[25], net1012[26], net1012[27], net1012[28],
     net1012[29], net1012[30], net1012[31], net1012[32], net1012[33],
     net1012[34], net1012[35], net1012[36], net1012[37], net1012[38],
     net1012[39], net1012[40], net1012[41], net1012[42], net1012[43],
     net1012[44], net1012[45], net1012[46], net1012[47]}),
     .sp4_h_r_01({net1013[0], net1013[1], net1013[2], net1013[3],
     net1013[4], net1013[5], net1013[6], net1013[7], net1013[8],
     net1013[9], net1013[10], net1013[11], net1013[12], net1013[13],
     net1013[14], net1013[15], net1013[16], net1013[17], net1013[18],
     net1013[19], net1013[20], net1013[21], net1013[22], net1013[23],
     net1013[24], net1013[25], net1013[26], net1013[27], net1013[28],
     net1013[29], net1013[30], net1013[31], net1013[32], net1013[33],
     net1013[34], net1013[35], net1013[36], net1013[37], net1013[38],
     net1013[39], net1013[40], net1013[41], net1013[42], net1013[43],
     net1013[44], net1013[45], net1013[46], net1013[47]}),
     .sp4_h_l_03({net1287[0], net1287[1], net1287[2], net1287[3],
     net1287[4], net1287[5], net1287[6], net1287[7], net1287[8],
     net1287[9], net1287[10], net1287[11], net1287[12], net1287[13],
     net1287[14], net1287[15], net1287[16], net1287[17], net1287[18],
     net1287[19], net1287[20], net1287[21], net1287[22], net1287[23],
     net1287[24], net1287[25], net1287[26], net1287[27], net1287[28],
     net1287[29], net1287[30], net1287[31], net1287[32], net1287[33],
     net1287[34], net1287[35], net1287[36], net1287[37], net1287[38],
     net1287[39], net1287[40], net1287[41], net1287[42], net1287[43],
     net1287[44], net1287[45], net1287[46], net1287[47]}),
     .sp4_h_l_02({net1286[0], net1286[1], net1286[2], net1286[3],
     net1286[4], net1286[5], net1286[6], net1286[7], net1286[8],
     net1286[9], net1286[10], net1286[11], net1286[12], net1286[13],
     net1286[14], net1286[15], net1286[16], net1286[17], net1286[18],
     net1286[19], net1286[20], net1286[21], net1286[22], net1286[23],
     net1286[24], net1286[25], net1286[26], net1286[27], net1286[28],
     net1286[29], net1286[30], net1286[31], net1286[32], net1286[33],
     net1286[34], net1286[35], net1286[36], net1286[37], net1286[38],
     net1286[39], net1286[40], net1286[41], net1286[42], net1286[43],
     net1286[44], net1286[45], net1286[46], net1286[47]}),
     .sp4_h_l_01({net1242[0], net1242[1], net1242[2], net1242[3],
     net1242[4], net1242[5], net1242[6], net1242[7], net1242[8],
     net1242[9], net1242[10], net1242[11], net1242[12], net1242[13],
     net1242[14], net1242[15], net1242[16], net1242[17], net1242[18],
     net1242[19], net1242[20], net1242[21], net1242[22], net1242[23],
     net1242[24], net1242[25], net1242[26], net1242[27], net1242[28],
     net1242[29], net1242[30], net1242[31], net1242[32], net1242[33],
     net1242[34], net1242[35], net1242[36], net1242[37], net1242[38],
     net1242[39], net1242[40], net1242[41], net1242[42], net1242[43],
     net1242[44], net1242[45], net1242[46], net1242[47]}),
     .bl(bl[221:168]), .bot_op_01({slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0], slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0]}),
     .sp12_h_l_01({net1236[0], net1236[1], net1236[2], net1236[3],
     net1236[4], net1236[5], net1236[6], net1236[7], net1236[8],
     net1236[9], net1236[10], net1236[11], net1236[12], net1236[13],
     net1236[14], net1236[15], net1236[16], net1236[17], net1236[18],
     net1236[19], net1236[20], net1236[21], net1236[22], net1236[23]}),
     .sp12_h_l_02({net1244[0], net1244[1], net1244[2], net1244[3],
     net1244[4], net1244[5], net1244[6], net1244[7], net1244[8],
     net1244[9], net1244[10], net1244[11], net1244[12], net1244[13],
     net1244[14], net1244[15], net1244[16], net1244[17], net1244[18],
     net1244[19], net1244[20], net1244[21], net1244[22], net1244[23]}),
     .sp12_h_l_03({net1200[0], net1200[1], net1200[2], net1200[3],
     net1200[4], net1200[5], net1200[6], net1200[7], net1200[8],
     net1200[9], net1200[10], net1200[11], net1200[12], net1200[13],
     net1200[14], net1200[15], net1200[16], net1200[17], net1200[18],
     net1200[19], net1200[20], net1200[21], net1200[22], net1200[23]}),
     .sp12_h_l_04({net1245[0], net1245[1], net1245[2], net1245[3],
     net1245[4], net1245[5], net1245[6], net1245[7], net1245[8],
     net1245[9], net1245[10], net1245[11], net1245[12], net1245[13],
     net1245[14], net1245[15], net1245[16], net1245[17], net1245[18],
     net1245[19], net1245[20], net1245[21], net1245[22], net1245[23]}),
     .sp4_v_b_04({net1224[0], net1224[1], net1224[2], net1224[3],
     net1224[4], net1224[5], net1224[6], net1224[7], net1224[8],
     net1224[9], net1224[10], net1224[11], net1224[12], net1224[13],
     net1224[14], net1224[15], net1224[16], net1224[17], net1224[18],
     net1224[19], net1224[20], net1224[21], net1224[22], net1224[23],
     net1224[24], net1224[25], net1224[26], net1224[27], net1224[28],
     net1224[29], net1224[30], net1224[31], net1224[32], net1224[33],
     net1224[34], net1224[35], net1224[36], net1224[37], net1224[38],
     net1224[39], net1224[40], net1224[41], net1224[42], net1224[43],
     net1224[44], net1224[45], net1224[46], net1224[47]}),
     .sp4_v_b_03({net1220[0], net1220[1], net1220[2], net1220[3],
     net1220[4], net1220[5], net1220[6], net1220[7], net1220[8],
     net1220[9], net1220[10], net1220[11], net1220[12], net1220[13],
     net1220[14], net1220[15], net1220[16], net1220[17], net1220[18],
     net1220[19], net1220[20], net1220[21], net1220[22], net1220[23],
     net1220[24], net1220[25], net1220[26], net1220[27], net1220[28],
     net1220[29], net1220[30], net1220[31], net1220[32], net1220[33],
     net1220[34], net1220[35], net1220[36], net1220[37], net1220[38],
     net1220[39], net1220[40], net1220[41], net1220[42], net1220[43],
     net1220[44], net1220[45], net1220[46], net1220[47]}),
     .sp4_v_b_02({net1231[0], net1231[1], net1231[2], net1231[3],
     net1231[4], net1231[5], net1231[6], net1231[7], net1231[8],
     net1231[9], net1231[10], net1231[11], net1231[12], net1231[13],
     net1231[14], net1231[15], net1231[16], net1231[17], net1231[18],
     net1231[19], net1231[20], net1231[21], net1231[22], net1231[23],
     net1231[24], net1231[25], net1231[26], net1231[27], net1231[28],
     net1231[29], net1231[30], net1231[31], net1231[32], net1231[33],
     net1231[34], net1231[35], net1231[36], net1231[37], net1231[38],
     net1231[39], net1231[40], net1231[41], net1231[42], net1231[43],
     net1231[44], net1231[45], net1231[46], net1231[47]}),
     .bnr_op_01({slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0], slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0]}), .sp4_h_l_05({net1289[0],
     net1289[1], net1289[2], net1289[3], net1289[4], net1289[5],
     net1289[6], net1289[7], net1289[8], net1289[9], net1289[10],
     net1289[11], net1289[12], net1289[13], net1289[14], net1289[15],
     net1289[16], net1289[17], net1289[18], net1289[19], net1289[20],
     net1289[21], net1289[22], net1289[23], net1289[24], net1289[25],
     net1289[26], net1289[27], net1289[28], net1289[29], net1289[30],
     net1289[31], net1289[32], net1289[33], net1289[34], net1289[35],
     net1289[36], net1289[37], net1289[38], net1289[39], net1289[40],
     net1289[41], net1289[42], net1289[43], net1289[44], net1289[45],
     net1289[46], net1289[47]}), .sp4_h_l_06({net1290[0], net1290[1],
     net1290[2], net1290[3], net1290[4], net1290[5], net1290[6],
     net1290[7], net1290[8], net1290[9], net1290[10], net1290[11],
     net1290[12], net1290[13], net1290[14], net1290[15], net1290[16],
     net1290[17], net1290[18], net1290[19], net1290[20], net1290[21],
     net1290[22], net1290[23], net1290[24], net1290[25], net1290[26],
     net1290[27], net1290[28], net1290[29], net1290[30], net1290[31],
     net1290[32], net1290[33], net1290[34], net1290[35], net1290[36],
     net1290[37], net1290[38], net1290[39], net1290[40], net1290[41],
     net1290[42], net1290[43], net1290[44], net1290[45], net1290[46],
     net1290[47]}), .sp4_h_l_07({net1291[0], net1291[1], net1291[2],
     net1291[3], net1291[4], net1291[5], net1291[6], net1291[7],
     net1291[8], net1291[9], net1291[10], net1291[11], net1291[12],
     net1291[13], net1291[14], net1291[15], net1291[16], net1291[17],
     net1291[18], net1291[19], net1291[20], net1291[21], net1291[22],
     net1291[23], net1291[24], net1291[25], net1291[26], net1291[27],
     net1291[28], net1291[29], net1291[30], net1291[31], net1291[32],
     net1291[33], net1291[34], net1291[35], net1291[36], net1291[37],
     net1291[38], net1291[39], net1291[40], net1291[41], net1291[42],
     net1291[43], net1291[44], net1291[45], net1291[46], net1291[47]}),
     .sp4_h_l_08({net1227[0], net1227[1], net1227[2], net1227[3],
     net1227[4], net1227[5], net1227[6], net1227[7], net1227[8],
     net1227[9], net1227[10], net1227[11], net1227[12], net1227[13],
     net1227[14], net1227[15], net1227[16], net1227[17], net1227[18],
     net1227[19], net1227[20], net1227[21], net1227[22], net1227[23],
     net1227[24], net1227[25], net1227[26], net1227[27], net1227[28],
     net1227[29], net1227[30], net1227[31], net1227[32], net1227[33],
     net1227[34], net1227[35], net1227[36], net1227[37], net1227[38],
     net1227[39], net1227[40], net1227[41], net1227[42], net1227[43],
     net1227[44], net1227[45], net1227[46], net1227[47]}),
     .sp4_h_r_08({net1031[0], net1031[1], net1031[2], net1031[3],
     net1031[4], net1031[5], net1031[6], net1031[7], net1031[8],
     net1031[9], net1031[10], net1031[11], net1031[12], net1031[13],
     net1031[14], net1031[15], net1031[16], net1031[17], net1031[18],
     net1031[19], net1031[20], net1031[21], net1031[22], net1031[23],
     net1031[24], net1031[25], net1031[26], net1031[27], net1031[28],
     net1031[29], net1031[30], net1031[31], net1031[32], net1031[33],
     net1031[34], net1031[35], net1031[36], net1031[37], net1031[38],
     net1031[39], net1031[40], net1031[41], net1031[42], net1031[43],
     net1031[44], net1031[45], net1031[46], net1031[47]}),
     .sp4_h_r_07({net1032[0], net1032[1], net1032[2], net1032[3],
     net1032[4], net1032[5], net1032[6], net1032[7], net1032[8],
     net1032[9], net1032[10], net1032[11], net1032[12], net1032[13],
     net1032[14], net1032[15], net1032[16], net1032[17], net1032[18],
     net1032[19], net1032[20], net1032[21], net1032[22], net1032[23],
     net1032[24], net1032[25], net1032[26], net1032[27], net1032[28],
     net1032[29], net1032[30], net1032[31], net1032[32], net1032[33],
     net1032[34], net1032[35], net1032[36], net1032[37], net1032[38],
     net1032[39], net1032[40], net1032[41], net1032[42], net1032[43],
     net1032[44], net1032[45], net1032[46], net1032[47]}),
     .sp4_h_r_06({net1033[0], net1033[1], net1033[2], net1033[3],
     net1033[4], net1033[5], net1033[6], net1033[7], net1033[8],
     net1033[9], net1033[10], net1033[11], net1033[12], net1033[13],
     net1033[14], net1033[15], net1033[16], net1033[17], net1033[18],
     net1033[19], net1033[20], net1033[21], net1033[22], net1033[23],
     net1033[24], net1033[25], net1033[26], net1033[27], net1033[28],
     net1033[29], net1033[30], net1033[31], net1033[32], net1033[33],
     net1033[34], net1033[35], net1033[36], net1033[37], net1033[38],
     net1033[39], net1033[40], net1033[41], net1033[42], net1033[43],
     net1033[44], net1033[45], net1033[46], net1033[47]}),
     .sp4_h_r_05({net1034[0], net1034[1], net1034[2], net1034[3],
     net1034[4], net1034[5], net1034[6], net1034[7], net1034[8],
     net1034[9], net1034[10], net1034[11], net1034[12], net1034[13],
     net1034[14], net1034[15], net1034[16], net1034[17], net1034[18],
     net1034[19], net1034[20], net1034[21], net1034[22], net1034[23],
     net1034[24], net1034[25], net1034[26], net1034[27], net1034[28],
     net1034[29], net1034[30], net1034[31], net1034[32], net1034[33],
     net1034[34], net1034[35], net1034[36], net1034[37], net1034[38],
     net1034[39], net1034[40], net1034[41], net1034[42], net1034[43],
     net1034[44], net1034[45], net1034[46], net1034[47]}),
     .slf_op_05({net1266[0], net1266[1], net1266[2], net1266[3],
     net1266[4], net1266[5], net1266[6], net1266[7]}),
     .slf_op_06({net1265[0], net1265[1], net1265[2], net1265[3],
     net1265[4], net1265[5], net1265[6], net1265[7]}),
     .slf_op_07({net1264[0], net1264[1], net1264[2], net1264[3],
     net1264[4], net1264[5], net1264[6], net1264[7]}),
     .slf_op_08(slf_op_04_08[7:0]), .rgt_op_08(slf_op_05_08[7:0]),
     .rgt_op_07({net1040[0], net1040[1], net1040[2], net1040[3],
     net1040[4], net1040[5], net1040[6], net1040[7]}),
     .rgt_op_06({net1041[0], net1041[1], net1041[2], net1041[3],
     net1041[4], net1041[5], net1041[6], net1041[7]}),
     .rgt_op_05({net1042[0], net1042[1], net1042[2], net1042[3],
     net1042[4], net1042[5], net1042[6], net1042[7]}),
     .lft_op_08(slf_op_03_08[7:0]), .lft_op_07({net758[0], net758[1],
     net758[2], net758[3], net758[4], net758[5], net758[6],
     net758[7]}), .lft_op_06({net759[0], net759[1], net759[2],
     net759[3], net759[4], net759[5], net759[6], net759[7]}),
     .lft_op_05({net760[0], net760[1], net760[2], net760[3], net760[4],
     net760[5], net760[6], net760[7]}), .sp12_h_l_08({net1217[0],
     net1217[1], net1217[2], net1217[3], net1217[4], net1217[5],
     net1217[6], net1217[7], net1217[8], net1217[9], net1217[10],
     net1217[11], net1217[12], net1217[13], net1217[14], net1217[15],
     net1217[16], net1217[17], net1217[18], net1217[19], net1217[20],
     net1217[21], net1217[22], net1217[23]}), .sp12_h_l_07({net1212[0],
     net1212[1], net1212[2], net1212[3], net1212[4], net1212[5],
     net1212[6], net1212[7], net1212[8], net1212[9], net1212[10],
     net1212[11], net1212[12], net1212[13], net1212[14], net1212[15],
     net1212[16], net1212[17], net1212[18], net1212[19], net1212[20],
     net1212[21], net1212[22], net1212[23]}), .sp12_h_l_06({net1214[0],
     net1214[1], net1214[2], net1214[3], net1214[4], net1214[5],
     net1214[6], net1214[7], net1214[8], net1214[9], net1214[10],
     net1214[11], net1214[12], net1214[13], net1214[14], net1214[15],
     net1214[16], net1214[17], net1214[18], net1214[19], net1214[20],
     net1214[21], net1214[22], net1214[23]}), .sp12_h_r_05({net1050[0],
     net1050[1], net1050[2], net1050[3], net1050[4], net1050[5],
     net1050[6], net1050[7], net1050[8], net1050[9], net1050[10],
     net1050[11], net1050[12], net1050[13], net1050[14], net1050[15],
     net1050[16], net1050[17], net1050[18], net1050[19], net1050[20],
     net1050[21], net1050[22], net1050[23]}), .sp12_h_r_06({net1051[0],
     net1051[1], net1051[2], net1051[3], net1051[4], net1051[5],
     net1051[6], net1051[7], net1051[8], net1051[9], net1051[10],
     net1051[11], net1051[12], net1051[13], net1051[14], net1051[15],
     net1051[16], net1051[17], net1051[18], net1051[19], net1051[20],
     net1051[21], net1051[22], net1051[23]}), .sp12_h_r_07({net1052[0],
     net1052[1], net1052[2], net1052[3], net1052[4], net1052[5],
     net1052[6], net1052[7], net1052[8], net1052[9], net1052[10],
     net1052[11], net1052[12], net1052[13], net1052[14], net1052[15],
     net1052[16], net1052[17], net1052[18], net1052[19], net1052[20],
     net1052[21], net1052[22], net1052[23]}), .sp12_h_r_08({net1053[0],
     net1053[1], net1053[2], net1053[3], net1053[4], net1053[5],
     net1053[6], net1053[7], net1053[8], net1053[9], net1053[10],
     net1053[11], net1053[12], net1053[13], net1053[14], net1053[15],
     net1053[16], net1053[17], net1053[18], net1053[19], net1053[20],
     net1053[21], net1053[22], net1053[23]}), .sp12_h_l_05({net1216[0],
     net1216[1], net1216[2], net1216[3], net1216[4], net1216[5],
     net1216[6], net1216[7], net1216[8], net1216[9], net1216[10],
     net1216[11], net1216[12], net1216[13], net1216[14], net1216[15],
     net1216[16], net1216[17], net1216[18], net1216[19], net1216[20],
     net1216[21], net1216[22], net1216[23]}),
     .sp4_r_v_b_05({net1055[0], net1055[1], net1055[2], net1055[3],
     net1055[4], net1055[5], net1055[6], net1055[7], net1055[8],
     net1055[9], net1055[10], net1055[11], net1055[12], net1055[13],
     net1055[14], net1055[15], net1055[16], net1055[17], net1055[18],
     net1055[19], net1055[20], net1055[21], net1055[22], net1055[23],
     net1055[24], net1055[25], net1055[26], net1055[27], net1055[28],
     net1055[29], net1055[30], net1055[31], net1055[32], net1055[33],
     net1055[34], net1055[35], net1055[36], net1055[37], net1055[38],
     net1055[39], net1055[40], net1055[41], net1055[42], net1055[43],
     net1055[44], net1055[45], net1055[46], net1055[47]}),
     .sp4_r_v_b_06({net1056[0], net1056[1], net1056[2], net1056[3],
     net1056[4], net1056[5], net1056[6], net1056[7], net1056[8],
     net1056[9], net1056[10], net1056[11], net1056[12], net1056[13],
     net1056[14], net1056[15], net1056[16], net1056[17], net1056[18],
     net1056[19], net1056[20], net1056[21], net1056[22], net1056[23],
     net1056[24], net1056[25], net1056[26], net1056[27], net1056[28],
     net1056[29], net1056[30], net1056[31], net1056[32], net1056[33],
     net1056[34], net1056[35], net1056[36], net1056[37], net1056[38],
     net1056[39], net1056[40], net1056[41], net1056[42], net1056[43],
     net1056[44], net1056[45], net1056[46], net1056[47]}),
     .sp4_r_v_b_07({net1057[0], net1057[1], net1057[2], net1057[3],
     net1057[4], net1057[5], net1057[6], net1057[7], net1057[8],
     net1057[9], net1057[10], net1057[11], net1057[12], net1057[13],
     net1057[14], net1057[15], net1057[16], net1057[17], net1057[18],
     net1057[19], net1057[20], net1057[21], net1057[22], net1057[23],
     net1057[24], net1057[25], net1057[26], net1057[27], net1057[28],
     net1057[29], net1057[30], net1057[31], net1057[32], net1057[33],
     net1057[34], net1057[35], net1057[36], net1057[37], net1057[38],
     net1057[39], net1057[40], net1057[41], net1057[42], net1057[43],
     net1057[44], net1057[45], net1057[46], net1057[47]}),
     .sp4_r_v_b_08({net1058[0], net1058[1], net1058[2], net1058[3],
     net1058[4], net1058[5], net1058[6], net1058[7], net1058[8],
     net1058[9], net1058[10], net1058[11], net1058[12], net1058[13],
     net1058[14], net1058[15], net1058[16], net1058[17], net1058[18],
     net1058[19], net1058[20], net1058[21], net1058[22], net1058[23],
     net1058[24], net1058[25], net1058[26], net1058[27], net1058[28],
     net1058[29], net1058[30], net1058[31], net1058[32], net1058[33],
     net1058[34], net1058[35], net1058[36], net1058[37], net1058[38],
     net1058[39], net1058[40], net1058[41], net1058[42], net1058[43],
     net1058[44], net1058[45], net1058[46], net1058[47]}),
     .sp4_v_b_08({net1259[0], net1259[1], net1259[2], net1259[3],
     net1259[4], net1259[5], net1259[6], net1259[7], net1259[8],
     net1259[9], net1259[10], net1259[11], net1259[12], net1259[13],
     net1259[14], net1259[15], net1259[16], net1259[17], net1259[18],
     net1259[19], net1259[20], net1259[21], net1259[22], net1259[23],
     net1259[24], net1259[25], net1259[26], net1259[27], net1259[28],
     net1259[29], net1259[30], net1259[31], net1259[32], net1259[33],
     net1259[34], net1259[35], net1259[36], net1259[37], net1259[38],
     net1259[39], net1259[40], net1259[41], net1259[42], net1259[43],
     net1259[44], net1259[45], net1259[46], net1259[47]}),
     .sp4_v_b_07({net1260[0], net1260[1], net1260[2], net1260[3],
     net1260[4], net1260[5], net1260[6], net1260[7], net1260[8],
     net1260[9], net1260[10], net1260[11], net1260[12], net1260[13],
     net1260[14], net1260[15], net1260[16], net1260[17], net1260[18],
     net1260[19], net1260[20], net1260[21], net1260[22], net1260[23],
     net1260[24], net1260[25], net1260[26], net1260[27], net1260[28],
     net1260[29], net1260[30], net1260[31], net1260[32], net1260[33],
     net1260[34], net1260[35], net1260[36], net1260[37], net1260[38],
     net1260[39], net1260[40], net1260[41], net1260[42], net1260[43],
     net1260[44], net1260[45], net1260[46], net1260[47]}),
     .sp4_v_b_06({net1261[0], net1261[1], net1261[2], net1261[3],
     net1261[4], net1261[5], net1261[6], net1261[7], net1261[8],
     net1261[9], net1261[10], net1261[11], net1261[12], net1261[13],
     net1261[14], net1261[15], net1261[16], net1261[17], net1261[18],
     net1261[19], net1261[20], net1261[21], net1261[22], net1261[23],
     net1261[24], net1261[25], net1261[26], net1261[27], net1261[28],
     net1261[29], net1261[30], net1261[31], net1261[32], net1261[33],
     net1261[34], net1261[35], net1261[36], net1261[37], net1261[38],
     net1261[39], net1261[40], net1261[41], net1261[42], net1261[43],
     net1261[44], net1261[45], net1261[46], net1261[47]}),
     .sp4_v_b_05({net1228[0], net1228[1], net1228[2], net1228[3],
     net1228[4], net1228[5], net1228[6], net1228[7], net1228[8],
     net1228[9], net1228[10], net1228[11], net1228[12], net1228[13],
     net1228[14], net1228[15], net1228[16], net1228[17], net1228[18],
     net1228[19], net1228[20], net1228[21], net1228[22], net1228[23],
     net1228[24], net1228[25], net1228[26], net1228[27], net1228[28],
     net1228[29], net1228[30], net1228[31], net1228[32], net1228[33],
     net1228[34], net1228[35], net1228[36], net1228[37], net1228[38],
     net1228[39], net1228[40], net1228[41], net1228[42], net1228[43],
     net1228[44], net1228[45], net1228[46], net1228[47]}),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .wl(wl_l[143:16]), .sp12_v_t_08(sp12_v_t_04_08[23:0]),
     .tnr_op_08(tnr_op_04_08[7:0]), .top_op_08(top_op_04_08[7:0]),
     .tnl_op_08(tnl_op_04_08[7:0]), .sp4_v_t_08(sp4_v_t_04_08[47:0]),
     .lc_bot(tiegnd_bl), .op_vic(op_vic_04_08),
     .sp12_v_b_01({net1404[0], net1404[1], net1404[2], net1404[3],
     net1404[4], net1404[5], net1404[6], net1404[7], net1404[8],
     net1404[9], net1404[10], net1404[11], net1404[12], net1404[13],
     net1404[14], net1404[15], net1404[16], net1404[17], net1404[18],
     net1404[19], net1404[20], net1404[21], net1404[22],
     net1404[23]}));
lt_1x8_bot_ice1f I_lt_col_t05 ( .glb_netwk_bot({net1384[0], net1384[1],
     net1384[2], net1384[3], net1384[4], net1384[5], net1384[6],
     net1384[7]}), .rgt_op_03(slf_op_06_03[7:0]),
     .slf_op_02({net983[0], net983[1], net983[2], net983[3], net983[4],
     net983[5], net983[6], net983[7]}), .rgt_op_02(slf_op_06_02[7:0]),
     .rgt_op_01(slf_op_06_01[7:0]), .purst(purst), .prog(prog),
     .lft_op_04({net1267[0], net1267[1], net1267[2], net1267[3],
     net1267[4], net1267[5], net1267[6], net1267[7]}),
     .lft_op_03({net1268[0], net1268[1], net1268[2], net1268[3],
     net1268[4], net1268[5], net1268[6], net1268[7]}),
     .lft_op_02({net1269[0], net1269[1], net1269[2], net1269[3],
     net1269[4], net1269[5], net1269[6], net1269[7]}),
     .lft_op_01({net1408[0], net1408[1], net1408[2], net1408[3],
     net1408[4], net1408[5], net1408[6], net1408[7]}),
     .rgt_op_04(slf_op_06_04[7:0]), .carry_in(tiegnd_bl),
     .bnl_op_01({slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0], slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0]}), .slf_op_04({net991[0],
     net991[1], net991[2], net991[3], net991[4], net991[5], net991[6],
     net991[7]}), .slf_op_03({net981[0], net981[1], net981[2],
     net981[3], net981[4], net981[5], net981[6], net981[7]}),
     .slf_op_01({net1409[0], net1409[1], net1409[2], net1409[3],
     net1409[4], net1409[5], net1409[6], net1409[7]}),
     .sp4_h_l_04({net1010[0], net1010[1], net1010[2], net1010[3],
     net1010[4], net1010[5], net1010[6], net1010[7], net1010[8],
     net1010[9], net1010[10], net1010[11], net1010[12], net1010[13],
     net1010[14], net1010[15], net1010[16], net1010[17], net1010[18],
     net1010[19], net1010[20], net1010[21], net1010[22], net1010[23],
     net1010[24], net1010[25], net1010[26], net1010[27], net1010[28],
     net1010[29], net1010[30], net1010[31], net1010[32], net1010[33],
     net1010[34], net1010[35], net1010[36], net1010[37], net1010[38],
     net1010[39], net1010[40], net1010[41], net1010[42], net1010[43],
     net1010[44], net1010[45], net1010[46], net1010[47]}),
     .carry_out(carry_out_05_08), .vdd_cntl(vdd_cntl_l[143:16]),
     .sp12_h_r_04({net1094[0], net1094[1], net1094[2], net1094[3],
     net1094[4], net1094[5], net1094[6], net1094[7], net1094[8],
     net1094[9], net1094[10], net1094[11], net1094[12], net1094[13],
     net1094[14], net1094[15], net1094[16], net1094[17], net1094[18],
     net1094[19], net1094[20], net1094[21], net1094[22], net1094[23]}),
     .sp12_h_r_03({net1095[0], net1095[1], net1095[2], net1095[3],
     net1095[4], net1095[5], net1095[6], net1095[7], net1095[8],
     net1095[9], net1095[10], net1095[11], net1095[12], net1095[13],
     net1095[14], net1095[15], net1095[16], net1095[17], net1095[18],
     net1095[19], net1095[20], net1095[21], net1095[22], net1095[23]}),
     .sp12_h_r_02({net1096[0], net1096[1], net1096[2], net1096[3],
     net1096[4], net1096[5], net1096[6], net1096[7], net1096[8],
     net1096[9], net1096[10], net1096[11], net1096[12], net1096[13],
     net1096[14], net1096[15], net1096[16], net1096[17], net1096[18],
     net1096[19], net1096[20], net1096[21], net1096[22], net1096[23]}),
     .sp12_h_r_01({net1097[0], net1097[1], net1097[2], net1097[3],
     net1097[4], net1097[5], net1097[6], net1097[7], net1097[8],
     net1097[9], net1097[10], net1097[11], net1097[12], net1097[13],
     net1097[14], net1097[15], net1097[16], net1097[17], net1097[18],
     net1097[19], net1097[20], net1097[21], net1097[22], net1097[23]}),
     .glb_netwk_col({net1344[0], net1344[1], net1344[2], net1344[3],
     net1344[4], net1344[5], net1344[6], net1344[7]}),
     .sp4_v_b_01({net1402[0], net1402[1], net1402[2], net1402[3],
     net1402[4], net1402[5], net1402[6], net1402[7], net1402[8],
     net1402[9], net1402[10], net1402[11], net1402[12], net1402[13],
     net1402[14], net1402[15], net1402[16], net1402[17], net1402[18],
     net1402[19], net1402[20], net1402[21], net1402[22], net1402[23],
     net1402[24], net1402[25], net1402[26], net1402[27], net1402[28],
     net1402[29], net1402[30], net1402[31], net1402[32], net1402[33],
     net1402[34], net1402[35], net1402[36], net1402[37], net1402[38],
     net1402[39], net1402[40], net1402[41], net1402[42], net1402[43],
     net1402[44], net1402[45], net1402[46], net1402[47]}),
     .sp4_r_v_b_04({net1100[0], net1100[1], net1100[2], net1100[3],
     net1100[4], net1100[5], net1100[6], net1100[7], net1100[8],
     net1100[9], net1100[10], net1100[11], net1100[12], net1100[13],
     net1100[14], net1100[15], net1100[16], net1100[17], net1100[18],
     net1100[19], net1100[20], net1100[21], net1100[22], net1100[23],
     net1100[24], net1100[25], net1100[26], net1100[27], net1100[28],
     net1100[29], net1100[30], net1100[31], net1100[32], net1100[33],
     net1100[34], net1100[35], net1100[36], net1100[37], net1100[38],
     net1100[39], net1100[40], net1100[41], net1100[42], net1100[43],
     net1100[44], net1100[45], net1100[46], net1100[47]}),
     .sp4_r_v_b_03({net1101[0], net1101[1], net1101[2], net1101[3],
     net1101[4], net1101[5], net1101[6], net1101[7], net1101[8],
     net1101[9], net1101[10], net1101[11], net1101[12], net1101[13],
     net1101[14], net1101[15], net1101[16], net1101[17], net1101[18],
     net1101[19], net1101[20], net1101[21], net1101[22], net1101[23],
     net1101[24], net1101[25], net1101[26], net1101[27], net1101[28],
     net1101[29], net1101[30], net1101[31], net1101[32], net1101[33],
     net1101[34], net1101[35], net1101[36], net1101[37], net1101[38],
     net1101[39], net1101[40], net1101[41], net1101[42], net1101[43],
     net1101[44], net1101[45], net1101[46], net1101[47]}),
     .sp4_r_v_b_02({net1102[0], net1102[1], net1102[2], net1102[3],
     net1102[4], net1102[5], net1102[6], net1102[7], net1102[8],
     net1102[9], net1102[10], net1102[11], net1102[12], net1102[13],
     net1102[14], net1102[15], net1102[16], net1102[17], net1102[18],
     net1102[19], net1102[20], net1102[21], net1102[22], net1102[23],
     net1102[24], net1102[25], net1102[26], net1102[27], net1102[28],
     net1102[29], net1102[30], net1102[31], net1102[32], net1102[33],
     net1102[34], net1102[35], net1102[36], net1102[37], net1102[38],
     net1102[39], net1102[40], net1102[41], net1102[42], net1102[43],
     net1102[44], net1102[45], net1102[46], net1102[47]}),
     .sp4_r_v_b_01({net1406[0], net1406[1], net1406[2], net1406[3],
     net1406[4], net1406[5], net1406[6], net1406[7], net1406[8],
     net1406[9], net1406[10], net1406[11], net1406[12], net1406[13],
     net1406[14], net1406[15], net1406[16], net1406[17], net1406[18],
     net1406[19], net1406[20], net1406[21], net1406[22], net1406[23],
     net1406[24], net1406[25], net1406[26], net1406[27], net1406[28],
     net1406[29], net1406[30], net1406[31], net1406[32], net1406[33],
     net1406[34], net1406[35], net1406[36], net1406[37], net1406[38],
     net1406[39], net1406[40], net1406[41], net1406[42], net1406[43],
     net1406[44], net1406[45], net1406[46], net1406[47]}),
     .sp4_h_r_04({net1104[0], net1104[1], net1104[2], net1104[3],
     net1104[4], net1104[5], net1104[6], net1104[7], net1104[8],
     net1104[9], net1104[10], net1104[11], net1104[12], net1104[13],
     net1104[14], net1104[15], net1104[16], net1104[17], net1104[18],
     net1104[19], net1104[20], net1104[21], net1104[22], net1104[23],
     net1104[24], net1104[25], net1104[26], net1104[27], net1104[28],
     net1104[29], net1104[30], net1104[31], net1104[32], net1104[33],
     net1104[34], net1104[35], net1104[36], net1104[37], net1104[38],
     net1104[39], net1104[40], net1104[41], net1104[42], net1104[43],
     net1104[44], net1104[45], net1104[46], net1104[47]}),
     .sp4_h_r_03({net1105[0], net1105[1], net1105[2], net1105[3],
     net1105[4], net1105[5], net1105[6], net1105[7], net1105[8],
     net1105[9], net1105[10], net1105[11], net1105[12], net1105[13],
     net1105[14], net1105[15], net1105[16], net1105[17], net1105[18],
     net1105[19], net1105[20], net1105[21], net1105[22], net1105[23],
     net1105[24], net1105[25], net1105[26], net1105[27], net1105[28],
     net1105[29], net1105[30], net1105[31], net1105[32], net1105[33],
     net1105[34], net1105[35], net1105[36], net1105[37], net1105[38],
     net1105[39], net1105[40], net1105[41], net1105[42], net1105[43],
     net1105[44], net1105[45], net1105[46], net1105[47]}),
     .sp4_h_r_02({net1106[0], net1106[1], net1106[2], net1106[3],
     net1106[4], net1106[5], net1106[6], net1106[7], net1106[8],
     net1106[9], net1106[10], net1106[11], net1106[12], net1106[13],
     net1106[14], net1106[15], net1106[16], net1106[17], net1106[18],
     net1106[19], net1106[20], net1106[21], net1106[22], net1106[23],
     net1106[24], net1106[25], net1106[26], net1106[27], net1106[28],
     net1106[29], net1106[30], net1106[31], net1106[32], net1106[33],
     net1106[34], net1106[35], net1106[36], net1106[37], net1106[38],
     net1106[39], net1106[40], net1106[41], net1106[42], net1106[43],
     net1106[44], net1106[45], net1106[46], net1106[47]}),
     .sp4_h_r_01({net1107[0], net1107[1], net1107[2], net1107[3],
     net1107[4], net1107[5], net1107[6], net1107[7], net1107[8],
     net1107[9], net1107[10], net1107[11], net1107[12], net1107[13],
     net1107[14], net1107[15], net1107[16], net1107[17], net1107[18],
     net1107[19], net1107[20], net1107[21], net1107[22], net1107[23],
     net1107[24], net1107[25], net1107[26], net1107[27], net1107[28],
     net1107[29], net1107[30], net1107[31], net1107[32], net1107[33],
     net1107[34], net1107[35], net1107[36], net1107[37], net1107[38],
     net1107[39], net1107[40], net1107[41], net1107[42], net1107[43],
     net1107[44], net1107[45], net1107[46], net1107[47]}),
     .sp4_h_l_03({net1011[0], net1011[1], net1011[2], net1011[3],
     net1011[4], net1011[5], net1011[6], net1011[7], net1011[8],
     net1011[9], net1011[10], net1011[11], net1011[12], net1011[13],
     net1011[14], net1011[15], net1011[16], net1011[17], net1011[18],
     net1011[19], net1011[20], net1011[21], net1011[22], net1011[23],
     net1011[24], net1011[25], net1011[26], net1011[27], net1011[28],
     net1011[29], net1011[30], net1011[31], net1011[32], net1011[33],
     net1011[34], net1011[35], net1011[36], net1011[37], net1011[38],
     net1011[39], net1011[40], net1011[41], net1011[42], net1011[43],
     net1011[44], net1011[45], net1011[46], net1011[47]}),
     .sp4_h_l_02({net1012[0], net1012[1], net1012[2], net1012[3],
     net1012[4], net1012[5], net1012[6], net1012[7], net1012[8],
     net1012[9], net1012[10], net1012[11], net1012[12], net1012[13],
     net1012[14], net1012[15], net1012[16], net1012[17], net1012[18],
     net1012[19], net1012[20], net1012[21], net1012[22], net1012[23],
     net1012[24], net1012[25], net1012[26], net1012[27], net1012[28],
     net1012[29], net1012[30], net1012[31], net1012[32], net1012[33],
     net1012[34], net1012[35], net1012[36], net1012[37], net1012[38],
     net1012[39], net1012[40], net1012[41], net1012[42], net1012[43],
     net1012[44], net1012[45], net1012[46], net1012[47]}),
     .sp4_h_l_01({net1013[0], net1013[1], net1013[2], net1013[3],
     net1013[4], net1013[5], net1013[6], net1013[7], net1013[8],
     net1013[9], net1013[10], net1013[11], net1013[12], net1013[13],
     net1013[14], net1013[15], net1013[16], net1013[17], net1013[18],
     net1013[19], net1013[20], net1013[21], net1013[22], net1013[23],
     net1013[24], net1013[25], net1013[26], net1013[27], net1013[28],
     net1013[29], net1013[30], net1013[31], net1013[32], net1013[33],
     net1013[34], net1013[35], net1013[36], net1013[37], net1013[38],
     net1013[39], net1013[40], net1013[41], net1013[42], net1013[43],
     net1013[44], net1013[45], net1013[46], net1013[47]}),
     .bl(bl[275:222]), .bot_op_01({slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0], slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0]}),
     .sp12_h_l_01({net1003[0], net1003[1], net1003[2], net1003[3],
     net1003[4], net1003[5], net1003[6], net1003[7], net1003[8],
     net1003[9], net1003[10], net1003[11], net1003[12], net1003[13],
     net1003[14], net1003[15], net1003[16], net1003[17], net1003[18],
     net1003[19], net1003[20], net1003[21], net1003[22], net1003[23]}),
     .sp12_h_l_02({net1002[0], net1002[1], net1002[2], net1002[3],
     net1002[4], net1002[5], net1002[6], net1002[7], net1002[8],
     net1002[9], net1002[10], net1002[11], net1002[12], net1002[13],
     net1002[14], net1002[15], net1002[16], net1002[17], net1002[18],
     net1002[19], net1002[20], net1002[21], net1002[22], net1002[23]}),
     .sp12_h_l_03({net1001[0], net1001[1], net1001[2], net1001[3],
     net1001[4], net1001[5], net1001[6], net1001[7], net1001[8],
     net1001[9], net1001[10], net1001[11], net1001[12], net1001[13],
     net1001[14], net1001[15], net1001[16], net1001[17], net1001[18],
     net1001[19], net1001[20], net1001[21], net1001[22], net1001[23]}),
     .sp12_h_l_04({net1000[0], net1000[1], net1000[2], net1000[3],
     net1000[4], net1000[5], net1000[6], net1000[7], net1000[8],
     net1000[9], net1000[10], net1000[11], net1000[12], net1000[13],
     net1000[14], net1000[15], net1000[16], net1000[17], net1000[18],
     net1000[19], net1000[20], net1000[21], net1000[22], net1000[23]}),
     .sp4_v_b_04({net1006[0], net1006[1], net1006[2], net1006[3],
     net1006[4], net1006[5], net1006[6], net1006[7], net1006[8],
     net1006[9], net1006[10], net1006[11], net1006[12], net1006[13],
     net1006[14], net1006[15], net1006[16], net1006[17], net1006[18],
     net1006[19], net1006[20], net1006[21], net1006[22], net1006[23],
     net1006[24], net1006[25], net1006[26], net1006[27], net1006[28],
     net1006[29], net1006[30], net1006[31], net1006[32], net1006[33],
     net1006[34], net1006[35], net1006[36], net1006[37], net1006[38],
     net1006[39], net1006[40], net1006[41], net1006[42], net1006[43],
     net1006[44], net1006[45], net1006[46], net1006[47]}),
     .sp4_v_b_03({net1007[0], net1007[1], net1007[2], net1007[3],
     net1007[4], net1007[5], net1007[6], net1007[7], net1007[8],
     net1007[9], net1007[10], net1007[11], net1007[12], net1007[13],
     net1007[14], net1007[15], net1007[16], net1007[17], net1007[18],
     net1007[19], net1007[20], net1007[21], net1007[22], net1007[23],
     net1007[24], net1007[25], net1007[26], net1007[27], net1007[28],
     net1007[29], net1007[30], net1007[31], net1007[32], net1007[33],
     net1007[34], net1007[35], net1007[36], net1007[37], net1007[38],
     net1007[39], net1007[40], net1007[41], net1007[42], net1007[43],
     net1007[44], net1007[45], net1007[46], net1007[47]}),
     .sp4_v_b_02({net1008[0], net1008[1], net1008[2], net1008[3],
     net1008[4], net1008[5], net1008[6], net1008[7], net1008[8],
     net1008[9], net1008[10], net1008[11], net1008[12], net1008[13],
     net1008[14], net1008[15], net1008[16], net1008[17], net1008[18],
     net1008[19], net1008[20], net1008[21], net1008[22], net1008[23],
     net1008[24], net1008[25], net1008[26], net1008[27], net1008[28],
     net1008[29], net1008[30], net1008[31], net1008[32], net1008[33],
     net1008[34], net1008[35], net1008[36], net1008[37], net1008[38],
     net1008[39], net1008[40], net1008[41], net1008[42], net1008[43],
     net1008[44], net1008[45], net1008[46], net1008[47]}),
     .bnr_op_01({slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0], slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0]}), .sp4_h_l_05({net1034[0],
     net1034[1], net1034[2], net1034[3], net1034[4], net1034[5],
     net1034[6], net1034[7], net1034[8], net1034[9], net1034[10],
     net1034[11], net1034[12], net1034[13], net1034[14], net1034[15],
     net1034[16], net1034[17], net1034[18], net1034[19], net1034[20],
     net1034[21], net1034[22], net1034[23], net1034[24], net1034[25],
     net1034[26], net1034[27], net1034[28], net1034[29], net1034[30],
     net1034[31], net1034[32], net1034[33], net1034[34], net1034[35],
     net1034[36], net1034[37], net1034[38], net1034[39], net1034[40],
     net1034[41], net1034[42], net1034[43], net1034[44], net1034[45],
     net1034[46], net1034[47]}), .sp4_h_l_06({net1033[0], net1033[1],
     net1033[2], net1033[3], net1033[4], net1033[5], net1033[6],
     net1033[7], net1033[8], net1033[9], net1033[10], net1033[11],
     net1033[12], net1033[13], net1033[14], net1033[15], net1033[16],
     net1033[17], net1033[18], net1033[19], net1033[20], net1033[21],
     net1033[22], net1033[23], net1033[24], net1033[25], net1033[26],
     net1033[27], net1033[28], net1033[29], net1033[30], net1033[31],
     net1033[32], net1033[33], net1033[34], net1033[35], net1033[36],
     net1033[37], net1033[38], net1033[39], net1033[40], net1033[41],
     net1033[42], net1033[43], net1033[44], net1033[45], net1033[46],
     net1033[47]}), .sp4_h_l_07({net1032[0], net1032[1], net1032[2],
     net1032[3], net1032[4], net1032[5], net1032[6], net1032[7],
     net1032[8], net1032[9], net1032[10], net1032[11], net1032[12],
     net1032[13], net1032[14], net1032[15], net1032[16], net1032[17],
     net1032[18], net1032[19], net1032[20], net1032[21], net1032[22],
     net1032[23], net1032[24], net1032[25], net1032[26], net1032[27],
     net1032[28], net1032[29], net1032[30], net1032[31], net1032[32],
     net1032[33], net1032[34], net1032[35], net1032[36], net1032[37],
     net1032[38], net1032[39], net1032[40], net1032[41], net1032[42],
     net1032[43], net1032[44], net1032[45], net1032[46], net1032[47]}),
     .sp4_h_l_08({net1031[0], net1031[1], net1031[2], net1031[3],
     net1031[4], net1031[5], net1031[6], net1031[7], net1031[8],
     net1031[9], net1031[10], net1031[11], net1031[12], net1031[13],
     net1031[14], net1031[15], net1031[16], net1031[17], net1031[18],
     net1031[19], net1031[20], net1031[21], net1031[22], net1031[23],
     net1031[24], net1031[25], net1031[26], net1031[27], net1031[28],
     net1031[29], net1031[30], net1031[31], net1031[32], net1031[33],
     net1031[34], net1031[35], net1031[36], net1031[37], net1031[38],
     net1031[39], net1031[40], net1031[41], net1031[42], net1031[43],
     net1031[44], net1031[45], net1031[46], net1031[47]}),
     .sp4_h_r_08({net1125[0], net1125[1], net1125[2], net1125[3],
     net1125[4], net1125[5], net1125[6], net1125[7], net1125[8],
     net1125[9], net1125[10], net1125[11], net1125[12], net1125[13],
     net1125[14], net1125[15], net1125[16], net1125[17], net1125[18],
     net1125[19], net1125[20], net1125[21], net1125[22], net1125[23],
     net1125[24], net1125[25], net1125[26], net1125[27], net1125[28],
     net1125[29], net1125[30], net1125[31], net1125[32], net1125[33],
     net1125[34], net1125[35], net1125[36], net1125[37], net1125[38],
     net1125[39], net1125[40], net1125[41], net1125[42], net1125[43],
     net1125[44], net1125[45], net1125[46], net1125[47]}),
     .sp4_h_r_07({net1126[0], net1126[1], net1126[2], net1126[3],
     net1126[4], net1126[5], net1126[6], net1126[7], net1126[8],
     net1126[9], net1126[10], net1126[11], net1126[12], net1126[13],
     net1126[14], net1126[15], net1126[16], net1126[17], net1126[18],
     net1126[19], net1126[20], net1126[21], net1126[22], net1126[23],
     net1126[24], net1126[25], net1126[26], net1126[27], net1126[28],
     net1126[29], net1126[30], net1126[31], net1126[32], net1126[33],
     net1126[34], net1126[35], net1126[36], net1126[37], net1126[38],
     net1126[39], net1126[40], net1126[41], net1126[42], net1126[43],
     net1126[44], net1126[45], net1126[46], net1126[47]}),
     .sp4_h_r_06({net1127[0], net1127[1], net1127[2], net1127[3],
     net1127[4], net1127[5], net1127[6], net1127[7], net1127[8],
     net1127[9], net1127[10], net1127[11], net1127[12], net1127[13],
     net1127[14], net1127[15], net1127[16], net1127[17], net1127[18],
     net1127[19], net1127[20], net1127[21], net1127[22], net1127[23],
     net1127[24], net1127[25], net1127[26], net1127[27], net1127[28],
     net1127[29], net1127[30], net1127[31], net1127[32], net1127[33],
     net1127[34], net1127[35], net1127[36], net1127[37], net1127[38],
     net1127[39], net1127[40], net1127[41], net1127[42], net1127[43],
     net1127[44], net1127[45], net1127[46], net1127[47]}),
     .sp4_h_r_05({net1128[0], net1128[1], net1128[2], net1128[3],
     net1128[4], net1128[5], net1128[6], net1128[7], net1128[8],
     net1128[9], net1128[10], net1128[11], net1128[12], net1128[13],
     net1128[14], net1128[15], net1128[16], net1128[17], net1128[18],
     net1128[19], net1128[20], net1128[21], net1128[22], net1128[23],
     net1128[24], net1128[25], net1128[26], net1128[27], net1128[28],
     net1128[29], net1128[30], net1128[31], net1128[32], net1128[33],
     net1128[34], net1128[35], net1128[36], net1128[37], net1128[38],
     net1128[39], net1128[40], net1128[41], net1128[42], net1128[43],
     net1128[44], net1128[45], net1128[46], net1128[47]}),
     .slf_op_05({net1042[0], net1042[1], net1042[2], net1042[3],
     net1042[4], net1042[5], net1042[6], net1042[7]}),
     .slf_op_06({net1041[0], net1041[1], net1041[2], net1041[3],
     net1041[4], net1041[5], net1041[6], net1041[7]}),
     .slf_op_07({net1040[0], net1040[1], net1040[2], net1040[3],
     net1040[4], net1040[5], net1040[6], net1040[7]}),
     .slf_op_08(slf_op_05_08[7:0]), .rgt_op_08(slf_op_06_08[7:0]),
     .rgt_op_07(slf_op_06_07[7:0]), .rgt_op_06(slf_op_06_06[7:0]),
     .rgt_op_05(slf_op_06_05[7:0]), .lft_op_08(slf_op_04_08[7:0]),
     .lft_op_07({net1264[0], net1264[1], net1264[2], net1264[3],
     net1264[4], net1264[5], net1264[6], net1264[7]}),
     .lft_op_06({net1265[0], net1265[1], net1265[2], net1265[3],
     net1265[4], net1265[5], net1265[6], net1265[7]}),
     .lft_op_05({net1266[0], net1266[1], net1266[2], net1266[3],
     net1266[4], net1266[5], net1266[6], net1266[7]}),
     .sp12_h_l_08({net1053[0], net1053[1], net1053[2], net1053[3],
     net1053[4], net1053[5], net1053[6], net1053[7], net1053[8],
     net1053[9], net1053[10], net1053[11], net1053[12], net1053[13],
     net1053[14], net1053[15], net1053[16], net1053[17], net1053[18],
     net1053[19], net1053[20], net1053[21], net1053[22], net1053[23]}),
     .sp12_h_l_07({net1052[0], net1052[1], net1052[2], net1052[3],
     net1052[4], net1052[5], net1052[6], net1052[7], net1052[8],
     net1052[9], net1052[10], net1052[11], net1052[12], net1052[13],
     net1052[14], net1052[15], net1052[16], net1052[17], net1052[18],
     net1052[19], net1052[20], net1052[21], net1052[22], net1052[23]}),
     .sp12_h_l_06({net1051[0], net1051[1], net1051[2], net1051[3],
     net1051[4], net1051[5], net1051[6], net1051[7], net1051[8],
     net1051[9], net1051[10], net1051[11], net1051[12], net1051[13],
     net1051[14], net1051[15], net1051[16], net1051[17], net1051[18],
     net1051[19], net1051[20], net1051[21], net1051[22], net1051[23]}),
     .sp12_h_r_05({net1144[0], net1144[1], net1144[2], net1144[3],
     net1144[4], net1144[5], net1144[6], net1144[7], net1144[8],
     net1144[9], net1144[10], net1144[11], net1144[12], net1144[13],
     net1144[14], net1144[15], net1144[16], net1144[17], net1144[18],
     net1144[19], net1144[20], net1144[21], net1144[22], net1144[23]}),
     .sp12_h_r_06({net1145[0], net1145[1], net1145[2], net1145[3],
     net1145[4], net1145[5], net1145[6], net1145[7], net1145[8],
     net1145[9], net1145[10], net1145[11], net1145[12], net1145[13],
     net1145[14], net1145[15], net1145[16], net1145[17], net1145[18],
     net1145[19], net1145[20], net1145[21], net1145[22], net1145[23]}),
     .sp12_h_r_07({net1146[0], net1146[1], net1146[2], net1146[3],
     net1146[4], net1146[5], net1146[6], net1146[7], net1146[8],
     net1146[9], net1146[10], net1146[11], net1146[12], net1146[13],
     net1146[14], net1146[15], net1146[16], net1146[17], net1146[18],
     net1146[19], net1146[20], net1146[21], net1146[22], net1146[23]}),
     .sp12_h_r_08({net1147[0], net1147[1], net1147[2], net1147[3],
     net1147[4], net1147[5], net1147[6], net1147[7], net1147[8],
     net1147[9], net1147[10], net1147[11], net1147[12], net1147[13],
     net1147[14], net1147[15], net1147[16], net1147[17], net1147[18],
     net1147[19], net1147[20], net1147[21], net1147[22], net1147[23]}),
     .sp12_h_l_05({net1050[0], net1050[1], net1050[2], net1050[3],
     net1050[4], net1050[5], net1050[6], net1050[7], net1050[8],
     net1050[9], net1050[10], net1050[11], net1050[12], net1050[13],
     net1050[14], net1050[15], net1050[16], net1050[17], net1050[18],
     net1050[19], net1050[20], net1050[21], net1050[22], net1050[23]}),
     .sp4_r_v_b_05({net1149[0], net1149[1], net1149[2], net1149[3],
     net1149[4], net1149[5], net1149[6], net1149[7], net1149[8],
     net1149[9], net1149[10], net1149[11], net1149[12], net1149[13],
     net1149[14], net1149[15], net1149[16], net1149[17], net1149[18],
     net1149[19], net1149[20], net1149[21], net1149[22], net1149[23],
     net1149[24], net1149[25], net1149[26], net1149[27], net1149[28],
     net1149[29], net1149[30], net1149[31], net1149[32], net1149[33],
     net1149[34], net1149[35], net1149[36], net1149[37], net1149[38],
     net1149[39], net1149[40], net1149[41], net1149[42], net1149[43],
     net1149[44], net1149[45], net1149[46], net1149[47]}),
     .sp4_r_v_b_06({net1150[0], net1150[1], net1150[2], net1150[3],
     net1150[4], net1150[5], net1150[6], net1150[7], net1150[8],
     net1150[9], net1150[10], net1150[11], net1150[12], net1150[13],
     net1150[14], net1150[15], net1150[16], net1150[17], net1150[18],
     net1150[19], net1150[20], net1150[21], net1150[22], net1150[23],
     net1150[24], net1150[25], net1150[26], net1150[27], net1150[28],
     net1150[29], net1150[30], net1150[31], net1150[32], net1150[33],
     net1150[34], net1150[35], net1150[36], net1150[37], net1150[38],
     net1150[39], net1150[40], net1150[41], net1150[42], net1150[43],
     net1150[44], net1150[45], net1150[46], net1150[47]}),
     .sp4_r_v_b_07({net1151[0], net1151[1], net1151[2], net1151[3],
     net1151[4], net1151[5], net1151[6], net1151[7], net1151[8],
     net1151[9], net1151[10], net1151[11], net1151[12], net1151[13],
     net1151[14], net1151[15], net1151[16], net1151[17], net1151[18],
     net1151[19], net1151[20], net1151[21], net1151[22], net1151[23],
     net1151[24], net1151[25], net1151[26], net1151[27], net1151[28],
     net1151[29], net1151[30], net1151[31], net1151[32], net1151[33],
     net1151[34], net1151[35], net1151[36], net1151[37], net1151[38],
     net1151[39], net1151[40], net1151[41], net1151[42], net1151[43],
     net1151[44], net1151[45], net1151[46], net1151[47]}),
     .sp4_r_v_b_08({net1152[0], net1152[1], net1152[2], net1152[3],
     net1152[4], net1152[5], net1152[6], net1152[7], net1152[8],
     net1152[9], net1152[10], net1152[11], net1152[12], net1152[13],
     net1152[14], net1152[15], net1152[16], net1152[17], net1152[18],
     net1152[19], net1152[20], net1152[21], net1152[22], net1152[23],
     net1152[24], net1152[25], net1152[26], net1152[27], net1152[28],
     net1152[29], net1152[30], net1152[31], net1152[32], net1152[33],
     net1152[34], net1152[35], net1152[36], net1152[37], net1152[38],
     net1152[39], net1152[40], net1152[41], net1152[42], net1152[43],
     net1152[44], net1152[45], net1152[46], net1152[47]}),
     .sp4_v_b_08({net1058[0], net1058[1], net1058[2], net1058[3],
     net1058[4], net1058[5], net1058[6], net1058[7], net1058[8],
     net1058[9], net1058[10], net1058[11], net1058[12], net1058[13],
     net1058[14], net1058[15], net1058[16], net1058[17], net1058[18],
     net1058[19], net1058[20], net1058[21], net1058[22], net1058[23],
     net1058[24], net1058[25], net1058[26], net1058[27], net1058[28],
     net1058[29], net1058[30], net1058[31], net1058[32], net1058[33],
     net1058[34], net1058[35], net1058[36], net1058[37], net1058[38],
     net1058[39], net1058[40], net1058[41], net1058[42], net1058[43],
     net1058[44], net1058[45], net1058[46], net1058[47]}),
     .sp4_v_b_07({net1057[0], net1057[1], net1057[2], net1057[3],
     net1057[4], net1057[5], net1057[6], net1057[7], net1057[8],
     net1057[9], net1057[10], net1057[11], net1057[12], net1057[13],
     net1057[14], net1057[15], net1057[16], net1057[17], net1057[18],
     net1057[19], net1057[20], net1057[21], net1057[22], net1057[23],
     net1057[24], net1057[25], net1057[26], net1057[27], net1057[28],
     net1057[29], net1057[30], net1057[31], net1057[32], net1057[33],
     net1057[34], net1057[35], net1057[36], net1057[37], net1057[38],
     net1057[39], net1057[40], net1057[41], net1057[42], net1057[43],
     net1057[44], net1057[45], net1057[46], net1057[47]}),
     .sp4_v_b_06({net1056[0], net1056[1], net1056[2], net1056[3],
     net1056[4], net1056[5], net1056[6], net1056[7], net1056[8],
     net1056[9], net1056[10], net1056[11], net1056[12], net1056[13],
     net1056[14], net1056[15], net1056[16], net1056[17], net1056[18],
     net1056[19], net1056[20], net1056[21], net1056[22], net1056[23],
     net1056[24], net1056[25], net1056[26], net1056[27], net1056[28],
     net1056[29], net1056[30], net1056[31], net1056[32], net1056[33],
     net1056[34], net1056[35], net1056[36], net1056[37], net1056[38],
     net1056[39], net1056[40], net1056[41], net1056[42], net1056[43],
     net1056[44], net1056[45], net1056[46], net1056[47]}),
     .sp4_v_b_05({net1055[0], net1055[1], net1055[2], net1055[3],
     net1055[4], net1055[5], net1055[6], net1055[7], net1055[8],
     net1055[9], net1055[10], net1055[11], net1055[12], net1055[13],
     net1055[14], net1055[15], net1055[16], net1055[17], net1055[18],
     net1055[19], net1055[20], net1055[21], net1055[22], net1055[23],
     net1055[24], net1055[25], net1055[26], net1055[27], net1055[28],
     net1055[29], net1055[30], net1055[31], net1055[32], net1055[33],
     net1055[34], net1055[35], net1055[36], net1055[37], net1055[38],
     net1055[39], net1055[40], net1055[41], net1055[42], net1055[43],
     net1055[44], net1055[45], net1055[46], net1055[47]}),
     .pgate(pgate_l[143:16]), .reset_b(reset_b_l[143:16]),
     .wl(wl_l[143:16]), .sp12_v_t_08(sp12_v_t_05_08[23:0]),
     .tnr_op_08(tnr_op_05_08[7:0]), .top_op_08(top_op_05_08[7:0]),
     .tnl_op_08(tnl_op_05_08[7:0]), .sp4_v_t_08(sp4_v_t_05_08[47:0]),
     .lc_bot(tiegnd_bl), .op_vic(op_vic_05_08),
     .sp12_v_b_01({net1426[0], net1426[1], net1426[2], net1426[3],
     net1426[4], net1426[5], net1426[6], net1426[7], net1426[8],
     net1426[9], net1426[10], net1426[11], net1426[12], net1426[13],
     net1426[14], net1426[15], net1426[16], net1426[17], net1426[18],
     net1426[19], net1426[20], net1426[21], net1426[22],
     net1426[23]}));
clk_quad_buf_x8_ice8p I_clktree_quad_drv_tl ( .clko(clk_center[7:0]),
     .clki(glb_in[7:0]));
clk_quad_buf_x8_ice8p I_clk_qtl_center ( .clko({net1344[0], net1344[1],
     net1344[2], net1344[3], net1344[4], net1344[5], net1344[6],
     net1344[7]}), .clki(clk_center[7:0]));
tielo I450 ( .tielo(tiegnd_bl));
pinlatbuf12p I_pinlatbuf12p_b ( .pad_in(padin_b_l[10]),
     .icegate(hold_l_b), .cbit(cf_b_l[135]), .cout(padinlat_b_l[10]),
     .prog(prog));
io_lft_bot_1x8_ice1f I_io_bot_00 ( .padeb(padeb_l_b[11:0]),
     .pado(pado_l_b[11:0]), .padin(padin_l_b[11:0]), .fo_fb(fo_fb),
     .fo_dlyadj(fo_dlyadj[2:0]), .fo_ref(fo_ref), .shift(net1295),
     .bs_en(net1296), .mode(net1297), .sdi(net1298), .hiz_b(net1299),
     .prog(prog), .hold(hold_l_b), .update(net1302), .r(net1303),
     .SP4_h_l_05({net1304[0], net1304[1], net1304[2], net1304[3],
     net1304[4], net1304[5], net1304[6], net1304[7], net1304[8],
     net1304[9], net1304[10], net1304[11], net1304[12], net1304[13],
     net1304[14], net1304[15], net1304[16], net1304[17], net1304[18],
     net1304[19], net1304[20], net1304[21], net1304[22], net1304[23],
     net1304[24], net1304[25], net1304[26], net1304[27], net1304[28],
     net1304[29], net1304[30], net1304[31], net1304[32], net1304[33],
     net1304[34], net1304[35], net1304[36], net1304[37], net1304[38],
     net1304[39], net1304[40], net1304[41], net1304[42], net1304[43],
     net1304[44], net1304[45], net1304[46], net1304[47]}),
     .slf_op_05(slf_op_00_05[3:0]), .slf_op_01(slf_op_00_01[3:0]),
     .slf_op_06(slf_op_00_06[3:0]), .slf_op_02(slf_op_00_02[3:0]),
     .sdo(net1309), .bl({bl[0], bl[1], bl[2], bl[3], bl[4], bl[5],
     bl[6], bl[7], bl[8], bl[9], bl[10], bl[11], bl[12], bl[13],
     bl[14], bl[15], bl[16], bl[17]}), .sp4_v_b_00_01({net1311[0],
     net1311[1], net1311[2], net1311[3], net1311[4], net1311[5],
     net1311[6], net1311[7], net1311[8], net1311[9], net1311[10],
     net1311[11], net1311[12], net1311[13], net1311[14], net1311[15]}),
     .tclk(net1312), .reset_b(reset_b_l[143:16]),
     .rgt_op_02({net1314[0], net1314[1], net1314[2], net1314[3],
     net1314[4], net1314[5], net1314[6], net1314[7]}),
     .SP4_h_l_06({net1315[0], net1315[1], net1315[2], net1315[3],
     net1315[4], net1315[5], net1315[6], net1315[7], net1315[8],
     net1315[9], net1315[10], net1315[11], net1315[12], net1315[13],
     net1315[14], net1315[15], net1315[16], net1315[17], net1315[18],
     net1315[19], net1315[20], net1315[21], net1315[22], net1315[23],
     net1315[24], net1315[25], net1315[26], net1315[27], net1315[28],
     net1315[29], net1315[30], net1315[31], net1315[32], net1315[33],
     net1315[34], net1315[35], net1315[36], net1315[37], net1315[38],
     net1315[39], net1315[40], net1315[41], net1315[42], net1315[43],
     net1315[44], net1315[45], net1315[46], net1315[47]}),
     .sp4_v_t_08(sp4_v_t_00_08[15:0]), .slf_op_04(slf_op_00_04[3:0]),
     .slf_op_03(slf_op_00_03[3:0]), .slf_op_07(slf_op_00_07[3:0]),
     .slf_op_08(slf_op_00_08[3:0]), .SP4_h_l_08({net1321[0],
     net1321[1], net1321[2], net1321[3], net1321[4], net1321[5],
     net1321[6], net1321[7], net1321[8], net1321[9], net1321[10],
     net1321[11], net1321[12], net1321[13], net1321[14], net1321[15],
     net1321[16], net1321[17], net1321[18], net1321[19], net1321[20],
     net1321[21], net1321[22], net1321[23], net1321[24], net1321[25],
     net1321[26], net1321[27], net1321[28], net1321[29], net1321[30],
     net1321[31], net1321[32], net1321[33], net1321[34], net1321[35],
     net1321[36], net1321[37], net1321[38], net1321[39], net1321[40],
     net1321[41], net1321[42], net1321[43], net1321[44], net1321[45],
     net1321[46], net1321[47]}), .SP4_h_l_07({net1322[0], net1322[1],
     net1322[2], net1322[3], net1322[4], net1322[5], net1322[6],
     net1322[7], net1322[8], net1322[9], net1322[10], net1322[11],
     net1322[12], net1322[13], net1322[14], net1322[15], net1322[16],
     net1322[17], net1322[18], net1322[19], net1322[20], net1322[21],
     net1322[22], net1322[23], net1322[24], net1322[25], net1322[26],
     net1322[27], net1322[28], net1322[29], net1322[30], net1322[31],
     net1322[32], net1322[33], net1322[34], net1322[35], net1322[36],
     net1322[37], net1322[38], net1322[39], net1322[40], net1322[41],
     net1322[42], net1322[43], net1322[44], net1322[45], net1322[46],
     net1322[47]}), .SP4_h_l_03({net1323[0], net1323[1], net1323[2],
     net1323[3], net1323[4], net1323[5], net1323[6], net1323[7],
     net1323[8], net1323[9], net1323[10], net1323[11], net1323[12],
     net1323[13], net1323[14], net1323[15], net1323[16], net1323[17],
     net1323[18], net1323[19], net1323[20], net1323[21], net1323[22],
     net1323[23], net1323[24], net1323[25], net1323[26], net1323[27],
     net1323[28], net1323[29], net1323[30], net1323[31], net1323[32],
     net1323[33], net1323[34], net1323[35], net1323[36], net1323[37],
     net1323[38], net1323[39], net1323[40], net1323[41], net1323[42],
     net1323[43], net1323[44], net1323[45], net1323[46], net1323[47]}),
     .SP4_h_l_04({net1324[0], net1324[1], net1324[2], net1324[3],
     net1324[4], net1324[5], net1324[6], net1324[7], net1324[8],
     net1324[9], net1324[10], net1324[11], net1324[12], net1324[13],
     net1324[14], net1324[15], net1324[16], net1324[17], net1324[18],
     net1324[19], net1324[20], net1324[21], net1324[22], net1324[23],
     net1324[24], net1324[25], net1324[26], net1324[27], net1324[28],
     net1324[29], net1324[30], net1324[31], net1324[32], net1324[33],
     net1324[34], net1324[35], net1324[36], net1324[37], net1324[38],
     net1324[39], net1324[40], net1324[41], net1324[42], net1324[43],
     net1324[44], net1324[45], net1324[46], net1324[47]}),
     .SP4_h_l_02({net1325[0], net1325[1], net1325[2], net1325[3],
     net1325[4], net1325[5], net1325[6], net1325[7], net1325[8],
     net1325[9], net1325[10], net1325[11], net1325[12], net1325[13],
     net1325[14], net1325[15], net1325[16], net1325[17], net1325[18],
     net1325[19], net1325[20], net1325[21], net1325[22], net1325[23],
     net1325[24], net1325[25], net1325[26], net1325[27], net1325[28],
     net1325[29], net1325[30], net1325[31], net1325[32], net1325[33],
     net1325[34], net1325[35], net1325[36], net1325[37], net1325[38],
     net1325[39], net1325[40], net1325[41], net1325[42], net1325[43],
     net1325[44], net1325[45], net1325[46], net1325[47]}),
     .SP4_h_l_01({net1326[0], net1326[1], net1326[2], net1326[3],
     net1326[4], net1326[5], net1326[6], net1326[7], net1326[8],
     net1326[9], net1326[10], net1326[11], net1326[12], net1326[13],
     net1326[14], net1326[15], net1326[16], net1326[17], net1326[18],
     net1326[19], net1326[20], net1326[21], net1326[22], net1326[23],
     net1326[24], net1326[25], net1326[26], net1326[27], net1326[28],
     net1326[29], net1326[30], net1326[31], net1326[32], net1326[33],
     net1326[34], net1326[35], net1326[36], net1326[37], net1326[38],
     net1326[39], net1326[40], net1326[41], net1326[42], net1326[43],
     net1326[44], net1326[45], net1326[46], net1326[47]}),
     .rgt_op_07({net1327[0], net1327[1], net1327[2], net1327[3],
     net1327[4], net1327[5], net1327[6], net1327[7]}),
     .rgt_op_06({net1328[0], net1328[1], net1328[2], net1328[3],
     net1328[4], net1328[5], net1328[6], net1328[7]}),
     .rgt_op_05({net1329[0], net1329[1], net1329[2], net1329[3],
     net1329[4], net1329[5], net1329[6], net1329[7]}),
     .rgt_op_03({net1330[0], net1330[1], net1330[2], net1330[3],
     net1330[4], net1330[5], net1330[6], net1330[7]}),
     .rgt_op_01({net1417[0], net1417[1], net1417[2], net1417[3],
     net1417[4], net1417[5], net1417[6], net1417[7]}),
     .rgt_op_08(slf_op_01_08[7:0]), .pgate(pgate_l[143:16]),
     .vdd_cntl(vdd_cntl_l[143:16]), .cf_l(cf_l[191:0]),
     .wl(wl_l[143:16]),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .tclk_o(net1338), .ceb(net1339), .SP12_h_l_02({net1340[0],
     net1340[1], net1340[2], net1340[3], net1340[4], net1340[5],
     net1340[6], net1340[7], net1340[8], net1340[9], net1340[10],
     net1340[11], net1340[12], net1340[13], net1340[14], net1340[15],
     net1340[16], net1340[17], net1340[18], net1340[19], net1340[20],
     net1340[21], net1340[22], net1340[23]}), .SP12_h_l_04({net1341[0],
     net1341[1], net1341[2], net1341[3], net1341[4], net1341[5],
     net1341[6], net1341[7], net1341[8], net1341[9], net1341[10],
     net1341[11], net1341[12], net1341[13], net1341[14], net1341[15],
     net1341[16], net1341[17], net1341[18], net1341[19], net1341[20],
     net1341[21], net1341[22], net1341[23]}), .SP12_h_l_08({net1342[0],
     net1342[1], net1342[2], net1342[3], net1342[4], net1342[5],
     net1342[6], net1342[7], net1342[8], net1342[9], net1342[10],
     net1342[11], net1342[12], net1342[13], net1342[14], net1342[15],
     net1342[16], net1342[17], net1342[18], net1342[19], net1342[20],
     net1342[21], net1342[22], net1342[23]}), .SP12_h_l_06({net1343[0],
     net1343[1], net1343[2], net1343[3], net1343[4], net1343[5],
     net1343[6], net1343[7], net1343[8], net1343[9], net1343[10],
     net1343[11], net1343[12], net1343[13], net1343[14], net1343[15],
     net1343[16], net1343[17], net1343[18], net1343[19], net1343[20],
     net1343[21], net1343[22], net1343[23]}),
     .glb_netwk_col({net1344[0], net1344[1], net1344[2], net1344[3],
     net1344[4], net1344[5], net1344[6], net1344[7]}),
     .SP12_h_l_05({net1345[0], net1345[1], net1345[2], net1345[3],
     net1345[4], net1345[5], net1345[6], net1345[7], net1345[8],
     net1345[9], net1345[10], net1345[11], net1345[12], net1345[13],
     net1345[14], net1345[15], net1345[16], net1345[17], net1345[18],
     net1345[19], net1345[20], net1345[21], net1345[22], net1345[23]}),
     .SP12_h_l_01({net1346[0], net1346[1], net1346[2], net1346[3],
     net1346[4], net1346[5], net1346[6], net1346[7], net1346[8],
     net1346[9], net1346[10], net1346[11], net1346[12], net1346[13],
     net1346[14], net1346[15], net1346[16], net1346[17], net1346[18],
     net1346[19], net1346[20], net1346[21], net1346[22], net1346[23]}),
     .fabric_out_07(fo_00_07), .SP12_h_l_03({net1348[0], net1348[1],
     net1348[2], net1348[3], net1348[4], net1348[5], net1348[6],
     net1348[7], net1348[8], net1348[9], net1348[10], net1348[11],
     net1348[12], net1348[13], net1348[14], net1348[15], net1348[16],
     net1348[17], net1348[18], net1348[19], net1348[20], net1348[21],
     net1348[22], net1348[23]}), .fabric_out_08(fo_00_08),
     .SP12_h_l_07({net1350[0], net1350[1], net1350[2], net1350[3],
     net1350[4], net1350[5], net1350[6], net1350[7], net1350[8],
     net1350[9], net1350[10], net1350[11], net1350[12], net1350[13],
     net1350[14], net1350[15], net1350[16], net1350[17], net1350[18],
     net1350[19], net1350[20], net1350[21], net1350[22], net1350[23]}),
     .last_rsr(last_rsr[0]), .rgt_op_04({net1355[0], net1355[1],
     net1355[2], net1355[3], net1355[4], net1355[5], net1355[6],
     net1355[7]}), .bnr_op_00_01({slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0], slf_op_01_00[3],
     slf_op_01_00[2], slf_op_01_00[1], slf_op_01_00[0]}),
     .tnr_op_08(tnr_op_00_08[7:0]));
io_bot_lft_1x6_ice1f test ( bs_en_o, ceb_o, cf_b_l[143:0], net1461,
     net1459, fo_bypass, fo_reset, fo_sck, fo_sdi, hiz_b_o, mode_o,
     padeb_b_l[10:0], padeb_b_l[12], pado_b_l[10:0], pado_b_l[12], r_o,
     sdo, shift_o, slf_op_01_00[3:0], slf_op_02_00[3:0],
     slf_op_03_00[3:0], slf_op_04_00[3:0], slf_op_05_00[3:0],
     slf_op_06_00[3:0], tclk_o, update_o, bl[71:18], bl[125:72],
     bl[167:126], bl[221:168], bl[275:222], bl[329:276], {net1311[0],
     net1311[1], net1311[2], net1311[3], net1311[4], net1311[5],
     net1311[6], net1311[7], net1311[8], net1311[9], net1311[10],
     net1311[11], net1311[12], net1311[13], net1311[14], net1311[15]},
     sp4_h_r_06_00[15:0], {net1437[0], net1437[1], net1437[2],
     net1437[3], net1437[4], net1437[5], net1437[6], net1437[7],
     net1437[8], net1437[9], net1437[10], net1437[11], net1437[12],
     net1437[13], net1437[14], net1437[15], net1437[16], net1437[17],
     net1437[18], net1437[19], net1437[20], net1437[21], net1437[22],
     net1437[23], net1437[24], net1437[25], net1437[26], net1437[27],
     net1437[28], net1437[29], net1437[30], net1437[31], net1437[32],
     net1437[33], net1437[34], net1437[35], net1437[36], net1437[37],
     net1437[38], net1437[39], net1437[40], net1437[41], net1437[42],
     net1437[43], net1437[44], net1437[45], net1437[46], net1437[47]},
     {net1411[0], net1411[1], net1411[2], net1411[3], net1411[4],
     net1411[5], net1411[6], net1411[7], net1411[8], net1411[9],
     net1411[10], net1411[11], net1411[12], net1411[13], net1411[14],
     net1411[15], net1411[16], net1411[17], net1411[18], net1411[19],
     net1411[20], net1411[21], net1411[22], net1411[23], net1411[24],
     net1411[25], net1411[26], net1411[27], net1411[28], net1411[29],
     net1411[30], net1411[31], net1411[32], net1411[33], net1411[34],
     net1411[35], net1411[36], net1411[37], net1411[38], net1411[39],
     net1411[40], net1411[41], net1411[42], net1411[43], net1411[44],
     net1411[45], net1411[46], net1411[47]}, {net1412[0], net1412[1],
     net1412[2], net1412[3], net1412[4], net1412[5], net1412[6],
     net1412[7], net1412[8], net1412[9], net1412[10], net1412[11],
     net1412[12], net1412[13], net1412[14], net1412[15], net1412[16],
     net1412[17], net1412[18], net1412[19], net1412[20], net1412[21],
     net1412[22], net1412[23], net1412[24], net1412[25], net1412[26],
     net1412[27], net1412[28], net1412[29], net1412[30], net1412[31],
     net1412[32], net1412[33], net1412[34], net1412[35], net1412[36],
     net1412[37], net1412[38], net1412[39], net1412[40], net1412[41],
     net1412[42], net1412[43], net1412[44], net1412[45], net1412[46],
     net1412[47]}, {net1414[0], net1414[1], net1414[2], net1414[3],
     net1414[4], net1414[5], net1414[6], net1414[7], net1414[8],
     net1414[9], net1414[10], net1414[11], net1414[12], net1414[13],
     net1414[14], net1414[15], net1414[16], net1414[17], net1414[18],
     net1414[19], net1414[20], net1414[21], net1414[22], net1414[23],
     net1414[24], net1414[25], net1414[26], net1414[27], net1414[28],
     net1414[29], net1414[30], net1414[31], net1414[32], net1414[33],
     net1414[34], net1414[35], net1414[36], net1414[37], net1414[38],
     net1414[39], net1414[40], net1414[41], net1414[42], net1414[43],
     net1414[44], net1414[45], net1414[46], net1414[47]}, {net1402[0],
     net1402[1], net1402[2], net1402[3], net1402[4], net1402[5],
     net1402[6], net1402[7], net1402[8], net1402[9], net1402[10],
     net1402[11], net1402[12], net1402[13], net1402[14], net1402[15],
     net1402[16], net1402[17], net1402[18], net1402[19], net1402[20],
     net1402[21], net1402[22], net1402[23], net1402[24], net1402[25],
     net1402[26], net1402[27], net1402[28], net1402[29], net1402[30],
     net1402[31], net1402[32], net1402[33], net1402[34], net1402[35],
     net1402[36], net1402[37], net1402[38], net1402[39], net1402[40],
     net1402[41], net1402[42], net1402[43], net1402[44], net1402[45],
     net1402[46], net1402[47]}, {net1406[0], net1406[1], net1406[2],
     net1406[3], net1406[4], net1406[5], net1406[6], net1406[7],
     net1406[8], net1406[9], net1406[10], net1406[11], net1406[12],
     net1406[13], net1406[14], net1406[15], net1406[16], net1406[17],
     net1406[18], net1406[19], net1406[20], net1406[21], net1406[22],
     net1406[23], net1406[24], net1406[25], net1406[26], net1406[27],
     net1406[28], net1406[29], net1406[30], net1406[31], net1406[32],
     net1406[33], net1406[34], net1406[35], net1406[36], net1406[37],
     net1406[38], net1406[39], net1406[40], net1406[41], net1406[42],
     net1406[43], net1406[44], net1406[45], net1406[46], net1406[47]},
     {net1373[0], net1373[1], net1373[2], net1373[3], net1373[4],
     net1373[5], net1373[6], net1373[7], net1373[8], net1373[9],
     net1373[10], net1373[11], net1373[12], net1373[13], net1373[14],
     net1373[15], net1373[16], net1373[17], net1373[18], net1373[19],
     net1373[20], net1373[21], net1373[22], net1373[23]}, {net1390[0],
     net1390[1], net1390[2], net1390[3], net1390[4], net1390[5],
     net1390[6], net1390[7], net1390[8], net1390[9], net1390[10],
     net1390[11], net1390[12], net1390[13], net1390[14], net1390[15],
     net1390[16], net1390[17], net1390[18], net1390[19], net1390[20],
     net1390[21], net1390[22], net1390[23]}, {net1413[0], net1413[1],
     net1413[2], net1413[3], net1413[4], net1413[5], net1413[6],
     net1413[7], net1413[8], net1413[9], net1413[10], net1413[11],
     net1413[12], net1413[13], net1413[14], net1413[15], net1413[16],
     net1413[17], net1413[18], net1413[19], net1413[20], net1413[21],
     net1413[22], net1413[23]}, {net1404[0], net1404[1], net1404[2],
     net1404[3], net1404[4], net1404[5], net1404[6], net1404[7],
     net1404[8], net1404[9], net1404[10], net1404[11], net1404[12],
     net1404[13], net1404[14], net1404[15], net1404[16], net1404[17],
     net1404[18], net1404[19], net1404[20], net1404[21], net1404[22],
     net1404[23]}, {net1426[0], net1426[1], net1426[2], net1426[3],
     net1426[4], net1426[5], net1426[6], net1426[7], net1426[8],
     net1426[9], net1426[10], net1426[11], net1426[12], net1426[13],
     net1426[14], net1426[15], net1426[16], net1426[17], net1426[18],
     net1426[19], net1426[20], net1426[21], net1426[22], net1426[23]},
     {net1407[0], net1407[1], net1407[2], net1407[3], net1407[4],
     net1407[5], net1407[6], net1407[7], net1407[8], net1407[9],
     net1407[10], net1407[11], net1407[12], net1407[13], net1407[14],
     net1407[15], net1407[16], net1407[17], net1407[18], net1407[19],
     net1407[20], net1407[21], net1407[22], net1407[23]},
     {slf_op_00_01[3], slf_op_00_01[2], slf_op_00_01[1],
     slf_op_00_01[0], slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0]}, net1296, net1339, {net1388[0],
     net1388[1], net1388[2], net1388[3], net1388[4], net1388[5],
     net1388[6], net1388[7]}, {net1387[0], net1387[1], net1387[2],
     net1387[3], net1387[4], net1387[5], net1387[6], net1387[7]},
     {net1386[0], net1386[1], net1386[2], net1386[3], net1386[4],
     net1386[5], net1386[6], net1386[7]}, {net1385[0], net1385[1],
     net1385[2], net1385[3], net1385[4], net1385[5], net1385[6],
     net1385[7]}, {net1384[0], net1384[1], net1384[2], net1384[3],
     net1384[4], net1384[5], net1384[6], net1384[7]}, {net1383[0],
     net1383[1], net1383[2], net1383[3], net1383[4], net1383[5],
     net1383[6], net1383[7]}, net1299, hold_b_l, {net1417[0],
     net1417[1], net1417[2], net1417[3], net1417[4], net1417[5],
     net1417[6], net1417[7]}, {net1419[0], net1419[1], net1419[2],
     net1419[3], net1419[4], net1419[5], net1419[6], net1419[7]},
     {net1410[0], net1410[1], net1410[2], net1410[3], net1410[4],
     net1410[5], net1410[6], net1410[7]}, {net1408[0], net1408[1],
     net1408[2], net1408[3], net1408[4], net1408[5], net1408[6],
     net1408[7]}, {net1409[0], net1409[1], net1409[2], net1409[3],
     net1409[4], net1409[5], net1409[6], net1409[7]},
     slf_op_06_01[7:0], net1297, padin_b_l[10:0], padin_b_l[12],
     {pgate_l[1], pgate_l[0], pgate_l[2], pgate_l[3], pgate_l[5],
     pgate_l[4], pgate_l[6], pgate_l[7], pgate_l[9], pgate_l[8],
     pgate_l[10], pgate_l[11], pgate_l[13], pgate_l[12], pgate_l[14],
     pgate_l[15]}, prog, net1303, {reset_b_l[1], reset_b_l[0],
     reset_b_l[2], reset_b_l[3], reset_b_l[5], reset_b_l[4],
     reset_b_l[6], reset_b_l[7], reset_b_l[9], reset_b_l[8],
     reset_b_l[10], reset_b_l[11], reset_b_l[13], reset_b_l[12],
     reset_b_l[14], reset_b_l[15]}, net1309, net1295, net1338,
     rgt_op_06_01[7:0], net1302, {vdd_cntl_l[1], vdd_cntl_l[0],
     vdd_cntl_l[2], vdd_cntl_l[3], vdd_cntl_l[5], vdd_cntl_l[4],
     vdd_cntl_l[6], vdd_cntl_l[7], vdd_cntl_l[9], vdd_cntl_l[8],
     vdd_cntl_l[10], vdd_cntl_l[11], vdd_cntl_l[13], vdd_cntl_l[12],
     vdd_cntl_l[14], vdd_cntl_l[15]}, {wl_l[1], wl_l[0], wl_l[2],
     wl_l[3], wl_l[5], wl_l[4], wl_l[6], wl_l[7], wl_l[9], wl_l[8],
     wl_l[10], wl_l[11], wl_l[13], wl_l[12], wl_l[14], wl_l[15]});
scan_buf_ice8p I_scanbuf_8p_ml ( .update_i(update_i), .tclk_i(tclk_i),
     .shift_i(shift_i), .sdi(sdi), .r_i(r_i), .mode_i(mode_i),
     .hiz_b_i(hiz_b_i), .ceb_i(ceb_i), .bs_en_i(bs_en_i),
     .update_o(net1302), .tclk_o(net1312), .shift_o(net1295),
     .sdo(net1298), .r_o(net1303), .mode_o(net1297), .hiz_b_o(net1299),
     .ceb_o(net1339), .bs_en_o(net1296));
fabric_buf_ice8p I785 ( .f_in(net1459), .f_out(fabric_out_06_00));
fabric_buf_ice8p I786 ( .f_in(net1461), .f_out(fabric_out_05_00));
fabric_buf_ice8p I_fabric_buf_8p_0016 ( .f_in(fo_00_08),
     .f_out(fabric_out_00_08));
fabric_buf_ice8p I_fabric_buf_8p_0015 ( .f_in(fo_00_07),
     .f_out(fabric_out_00_07));
fabric_buf_ice8p I_fabric_buf8p_25 ( .f_in(padinlat_l_b[11]),
     .f_out(padin_00_08));
fabric_buf_ice8p I784 ( .f_in(padinlat_b_l[10]), .f_out(padin_06_00));
pinlatbuf12p_1 I_pinlatbuf12p ( .pad_in(padin_l_b[11]),
     .icegate(hold_l_b), .cbit(cf_l[183]), .cout(padinlat_l_b[11]),
     .prog(prog));

endmodule
// Library - leafcell, Cell - bram_bufferx2e, View - schematic
// LAST TIME SAVED: May 13 10:18:51 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module bram_bufferx2e ( out, en, in );
output  out;

input  en, in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I391 ( .A(net7), .Y(out));
nand2 I193 ( .A(en), .Y(net7), .B(in));

endmodule
// Library - leafcell, Cell - bram_bank_logic_bot, View - schematic
// LAST TIME SAVED: Jul  8 10:16:10 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module bram_bank_logic_bot ( bm_sclkrw_o, bm_sdo_o, bm_sweb_o,
     bm_banksel_i, bm_sclk_i, bm_sclkrw_i, bm_sdo_i, bm_sweb_i );

input  bm_sclk_i, bm_sclkrw_i, bm_sweb_i;

output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sclkrw_o;

input [1:0]  bm_banksel_i;
input [1:0]  bm_sdo_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net26;

wire  [1:0]  net25;



ml_dff I52_1_ ( .R(net020), .D(bm_sdo_i[1]), .CLK(bm_sclk_i),
     .QN(net25[0]), .Q(net26[1]));
ml_dff I52_0_ ( .R(net020), .D(bm_sdo_i[0]), .CLK(bm_sclk_i),
     .QN(net25[1]), .Q(net26[0]));
bram_bufferx16_2inv I51_1_ ( .in(net26[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I51_0_ ( .in(net26[0]), .out(bm_sdo_o[0]));
bram_bufferx2e I54_1_ ( .in(bm_sweb_i), .en(bm_banksel_i[1]),
     .out(bm_sweb_o[1]));
bram_bufferx2e I54_0_ ( .in(bm_sweb_i), .en(bm_banksel_i[0]),
     .out(bm_sweb_o[0]));
bram_bufferx2e I48_1_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[1]),
     .out(bm_sclkrw_o[1]));
bram_bufferx2e I48_0_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[0]),
     .out(bm_sclkrw_o[0]));
tielo I55 ( .tielo(net020));

endmodule
// Library - leafcell, Cell - bram_icg, View - schematic
// LAST TIME SAVED: Oct 22 11:07:43 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module bram_icg ( clkout, clk, en );
output  clkout;

input  clk, en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I391 ( .A(net014), .Y(clkout));
inv I6 ( .A(net023), .Y(net027));
inv I4 ( .A(cn), .Y(c));
inv I3 ( .A(clk), .Y(cn));
nand2 I193 ( .A(net027), .Y(net014), .B(c));
inv_tri_2 I7 ( .Tb(cn), .T(c), .A(net027), .Y(net023));
inv_tri_2 I5 ( .Tb(c), .T(cn), .A(en), .Y(net023));

endmodule
// Library - leafcell, Cell - bram_hbuffer_dff_2xbank, View - schematic
// LAST TIME SAVED: Oct 22 09:16:56 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module bram_hbuffer_dff_2xbank ( bm_banksel_o, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclkrw_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [3:0]  bm_sdi_o;
output [3:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [3:0]  bm_banksel_o;
output [1:0]  bm_sclk_o;

input [3:0]  bm_sdi_i;
input [7:0]  bm_sa_i;
input [3:0]  bm_sdo_i;
input [3:0]  bm_banksel_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net103;

wire  [3:0]  net102;



ml_dff I48_3_ ( .R(net057), .D(bm_sdo_i[3]), .CLK(bm_sclk_i),
     .QN(net102[0]), .Q(net103[0]));
ml_dff I48_2_ ( .R(net057), .D(bm_sdo_i[2]), .CLK(bm_sclk_i),
     .QN(net102[1]), .Q(net103[1]));
ml_dff I48_1_ ( .R(net057), .D(bm_sdo_i[1]), .CLK(bm_sclk_i),
     .QN(net102[2]), .Q(net103[2]));
ml_dff I48_0_ ( .R(net057), .D(bm_sdo_i[0]), .CLK(bm_sclk_i),
     .QN(net102[3]), .Q(net103[3]));
nor2 I20 ( .A(bm_banksel_i[2]), .B(bm_banksel_i[3]), .Y(net67));
nor2 I49 ( .A(bm_banksel_i[0]), .B(bm_banksel_i[1]), .Y(net70));
inv I21 ( .A(net67), .Y(net72));
inv I17 ( .A(net70), .Y(net74));
tielo I23 ( .tielo(net057));
bram_icg I47 ( .en(net74), .clk(bm_sclk_i), .clkout(net61));
bram_icg I19 ( .en(net72), .clk(bm_sclk_i), .clkout(net64));
bram_bufferx16_2inv I16_3_ ( .in(net103[0]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I16_2_ ( .in(net103[1]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I16_1_ ( .in(net103[2]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I16_0_ ( .in(net103[3]), .out(bm_sdo_o[0]));
bram_bufferx4 I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx4 I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx4 I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx4 I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx4 I22 ( .in(net64), .out(bm_sclk_o[1]));
bram_bufferx4 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx4 I13_3_ ( .in(bm_banksel_i[3]), .out(bm_banksel_o[3]));
bram_bufferx4 I13_2_ ( .in(bm_banksel_i[2]), .out(bm_banksel_o[2]));
bram_bufferx4 I13_1_ ( .in(bm_banksel_i[1]), .out(bm_banksel_o[1]));
bram_bufferx4 I13_0_ ( .in(bm_banksel_i[0]), .out(bm_banksel_o[0]));
bram_bufferx4 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx4 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx4 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx4 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx4 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx4 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx4 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx4 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx4 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx4 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx4 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx4 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx4 I18 ( .in(net61), .out(bm_sclk_o[0]));
bram_bufferx4 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_hbuffer_1xbank, View - schematic
// LAST TIME SAVED: Jun 11 17:38:23 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module bram_hbuffer_1xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [1:0]  bm_banksel_o;
output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;

input [1:0]  bm_sdi_i;
input [1:0]  bm_sdo_i;
input [1:0]  bm_banksel_i;
input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - ice1chip, Cell - quad_x4_ice1, View - schematic
// LAST TIME SAVED: May  3 11:40:33 2011
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module quad_x4_ice1 ( bm_sdo_o[3:0], cf_b[287:0], cf_l[383:0],
     cf_r[383:0], cf_t[287:0], fabric_out_05_00_bicegate,
     fabric_out_06_00, fabric_out_07_00, fabric_out_12_00_wb,
     fabric_out_13_01, fabric_out_13_02, fo_bypass, fo_dlyadj[7:0],
     fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, padeb_b[23:0],
     padeb_l[23:0], padeb_r[24:0], padeb_t[23:0], pado_b[23:0],
     pado_l[23:0], pado_r[24:0], pado_t[23:0], sdo_pad,
     spi_ss_in_bbank[4:0], tck_pad, tdi_pad, tms_pad, bl_bot[663:0],
     bl_top[663:0], bm_banksel_i[3:0], bm_init_i, bm_rcapmux_en_i,
     bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i, bm_sdi_i[3:0], bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb, end_of_startup,
     gclk_l2clktv[1:0], gclk_r2clktv[1:0], hiz_b,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[0],
     last_rsr[1], last_rsr[2], last_rsr[3], md_spi_b, mode,
     mux_jtag_sel_b, padin_b[23:0], padin_l[23:0], padin_r[24:0],
     padin_t[23:0], pgate_l[287:0], pgate_r[287:0], pll_lock_out,
     pll_sdo, prog, purst, r, reset_b_l[287:0], reset_b_r[287:0],
     sdi_pad, sdo_enable, shift, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk, totdopad, trstb_pad, update, vdd_cntl_l[287:0],
     vdd_cntl_r[287:0], wl_l[287:0], wl_r[287:0] );
output  fabric_out_05_00_bicegate, fabric_out_06_00, fabric_out_07_00,
     fabric_out_12_00_wb, fabric_out_13_01, fabric_out_13_02,
     fo_bypass, fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, sdo_pad,
     tck_pad, tdi_pad, tms_pad;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb, end_of_startup, hiz_b,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode, mux_jtag_sel_b, pll_lock_out, pll_sdo, prog, purst, r,
     sdi_pad, sdo_enable, shift, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, tclk, totdopad, trstb_pad, update;

output [4:0]  spi_ss_in_bbank;
output [3:0]  bm_sdo_o;
output [23:0]  pado_l;
output [23:0]  padeb_l;
output [383:0]  cf_l;
output [23:0]  pado_t;
output [383:0]  cf_r;
output [24:0]  padeb_r;
output [23:0]  padeb_b;
output [23:0]  padeb_t;
output [287:0]  cf_t;
output [287:0]  cf_b;
output [7:0]  fo_dlyadj;
output [23:0]  pado_b;
output [24:0]  pado_r;

inout [663:0]  bl_bot;
inout [663:0]  bl_top;

input [3:0]  bm_sdi_i;
input [7:0]  bm_sa_i;
input [1:0]  gclk_r2clktv;
input [3:0]  bm_banksel_i;
input [287:0]  pgate_l;
input [23:0]  padin_l;
input [287:0]  pgate_r;
input [287:0]  vdd_cntl_r;
input [287:0]  reset_b_r;
input [287:0]  wl_r;
input [1:0]  gclk_l2clktv;
input [23:0]  padin_b;
input [3:0]  last_rsr;
input [287:0]  reset_b_l;
input [23:0]  padin_t;
input [24:0]  padin_r;
input [287:0]  wl_l;
input [287:0]  vdd_cntl_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  slf_op_07_13;

wire  [7:0]  slf_op_07_14;

wire  [23:0]  net1208;

wire  [23:0]  net983;

wire  [47:0]  net816;

wire  [3:0]  slf_op_06_17;

wire  [23:0]  net984;

wire  [23:0]  net1171;

wire  [23:0]  net1209;

wire  [7:0]  net995;

wire  [15:0]  net818;

wire  [23:0]  net1103;

wire  [7:0]  slf_op_07_11;

wire  [23:0]  net777;

wire  [7:0]  slf_op_01_09;

wire  [47:0]  net1225;

wire  [23:0]  net772;

wire  [47:0]  net1220;

wire  [23:0]  net771;

wire  [23:0]  net1198;

wire  [7:0]  slf_op_12_09;

wire  [10:0]  net1046;

wire  [1:0]  net1147;

wire  [7:0]  slf_op_08_09;

wire  [47:0]  net811;

wire  [47:0]  net1165;

wire  [47:0]  net1213;

wire  [47:0]  net849;

wire  [7:0]  slf_op_09_09;

wire  [7:0]  slf_op_07_08;

wire  [47:0]  net1218;

wire  [47:0]  net1001;

wire  [7:0]  net1190;

wire  [7:0]  slf_op_07_05;

wire  [47:0]  net1215;

wire  [23:0]  net985;

wire  [47:0]  net1224;

wire  [7:0]  slf_op_06_08;

wire  [23:0]  net1231;

wire  [47:0]  net1219;

wire  [23:0]  net986;

wire  [7:0]  slf_op_06_05;

wire  [47:0]  net1227;

wire  [23:0]  net1205;

wire  [7:0]  slf_op_06_06;

wire  [47:0]  net1115;

wire  [7:0]  slf_op_07_16;

wire  [7:0]  net1149;

wire  [47:0]  net1223;

wire  [7:0]  slf_op_04_08;

wire  [7:0]  slf_op_01_08;

wire  [47:0]  net921;

wire  [47:0]  net1212;

wire  [23:0]  net1222;

wire  [1:0]  bm_sweb_b2_o;

wire  [47:0]  net1242;

wire  [47:0]  net1228;

wire  [3:0]  slf_op_07_00;

wire  [47:0]  net998;

wire  [47:0]  net812;

wire  [1:0]  net1275;

wire  [1:0]  bm_sdo_b1_o;

wire  [23:0]  net773;

wire  [23:0]  net1206;

wire  [47:0]  net819;

wire  [7:0]  slf_op_07_15;

wire  [23:0]  net1170;

wire  [7:0]  slf_op_08_08;

wire  [7:0]  slf_op_07_12;

wire  [7:0]  slf_op_02_08;

wire  [23:0]  net1207;

wire  [7:0]  slf_op_06_11;

wire  [7:0]  slf_op_07_06;

wire  [47:0]  net820;

wire  [7:0]  slf_op_07_07;

wire  [7:0]  slf_op_04_09;

wire  [23:0]  net776;

wire  [47:0]  net1200;

wire  [7:0]  slf_op_02_09;

wire  [7:0]  slf_op_06_07;

wire  [7:0]  slf_op_06_03;

wire  [7:0]  slf_op_06_02;

wire  [7:0]  slf_op_07_01;

wire  [1:0]  net1146;

wire  [7:0]  slf_op_11_08;

wire  [7:0]  slf_op_07_03;

wire  [1:0]  bm_bank10_banksel_o;

wire  [7:0]  bm_bank30_sa_o;

wire  [7:0]  slf_op_03_09;

wire  [47:0]  net824;

wire  [47:0]  net1000;

wire  [23:0]  net774;

wire  [10:0]  net1232;

wire  [1:0]  net952;

wire  [7:0]  slf_op_05_08;

wire  [3:0]  slf_op_07_17;

wire  [47:0]  net814;

wire  [10:0]  net1071;

wire  [47:0]  net1221;

wire  [23:0]  net1195;

wire  [47:0]  net1241;

wire  [47:0]  net815;

wire  [7:0]  slf_op_06_14;

wire  [7:0]  slf_op_06_01;

wire  [7:0]  slf_op_05_09;

wire  [47:0]  net1217;

wire  [47:0]  net822;

wire  [7:0]  slf_op_06_16;

wire  [7:0]  slf_op_06_10;

wire  [7:0]  slf_op_03_08;

wire  [7:0]  slf_op_10_09;

wire  [47:0]  net848;

wire  [1:0]  bm_sdo_b0_o;

wire  [15:0]  net1250;

wire  [3:0]  slf_op_13_09;

wire  [47:0]  net810;

wire  [7:0]  gclk;

wire  [7:0]  slf_op_06_12;

wire  [1:0]  bm_sdo_b3_o;

wire  [47:0]  net813;

wire  [3:0]  slf_op_06_00;

wire  [1:0]  bm_sclkrw_b0_o;

wire  [1:0]  bm_bank30_sclk_o;

wire  [7:0]  slf_op_07_10;

wire  [47:0]  net1216;

wire  [1:0]  bm_sweb_b0_o;

wire  [3:0]  slf_op_00_08;

wire  [23:0]  net1197;

wire  [7:0]  slf_op_09_08;

wire  [1:0]  bm_sdi_b0_o;

wire  [7:0]  slf_op_12_08;

wire  [47:0]  net967;

wire  [7:0]  slf_op_06_15;

wire  [47:0]  net1214;

wire  [23:0]  net982;

wire  [7:0]  slf_op_06_04;

wire  [47:0]  net823;

wire  [23:0]  net775;

wire  [1:0]  bm_sclkrw_b2_o;

wire  [23:0]  net770;

wire  [47:0]  net1226;

wire  [1:0]  bm_sdi_b2_o;

wire  [47:0]  net999;

wire  [7:0]  slf_op_07_04;

wire  [3:0]  bm_bank30_sdi_o;

wire  [23:0]  net1196;

wire  [7:0]  slf_op_11_09;

wire  [7:0]  slf_op_07_02;

wire  [7:0]  slf_op_06_13;

wire  [47:0]  net821;

wire  [47:0]  net1199;

wire  [7:0]  slf_op_07_09;

wire  [3:0]  bm_bank30_sdo_i;

wire  [23:0]  net981;

wire  [15:0]  net911;

wire  [7:0]  slf_op_06_09;

wire  [1:0]  net1143;

wire  [3:0]  slf_op_00_09;

wire  [1:0]  net948;

wire  [10:0]  net1138;

wire  [7:0]  slf_op_10_08;

wire  [3:0]  bm_bank30_banksel_o;

wire  [15:0]  net1154;

wire  [3:0]  slf_op_13_08;

wire  [1:0]  bm_sdo_b2_o;



ice1f_cram_row142col4 I64 ( .vdd_cntl_l(vdd_cntl_l[287:146]),
     .bl(bl_top[333:330]), .vdd_cntl_r(vdd_cntl_r[287:146]),
     .reset_r(reset_b_r[287:146]), .pgate_r(pgate_r[287:146]),
     .reset_l(reset_b_l[287:146]), .pgate_l(pgate_l[287:146]),
     .wl_r(wl_r[287:146]), .wl_l(wl_l[287:146]));
ice1f_cram_row142col4 I65 ( .vdd_cntl_l(vdd_cntl_l[141:0]),
     .bl(bl_bot[333:330]), .vdd_cntl_r(vdd_cntl_r[141:0]),
     .reset_r(reset_b_r[141:0]), .pgate_r(pgate_r[141:0]),
     .reset_l(reset_b_l[141:0]), .pgate_l(pgate_l[141:0]),
     .wl_r(wl_r[141:0]), .wl_l(wl_l[141:0]));
bram_sdo_reg I_bm_sdo_reg_b0 ( .do(bm_sdo_b0_o_0), .di(bm_sdo_b0_o[0]),
     .clk(bm_sck_b0_i), .tielo(net1262));
bram_sdo_reg I_bm_sdo_reg_b2 ( .do(bm_sdo_b2_o_0), .di(bm_sdo_b2_o[0]),
     .clk(bm_bank30_sclk_o[1]), .tielo(net1256));
bram_sdo_reg I_bm_sdo_reg_b3 ( .do(bm_sdo_b3_o_0), .di(bm_sdo_b3_o[0]),
     .clk(bm_sck_b2_o), .tielo(tielo_4bram3));
bram_sdo_reg I_bm_sdo_reg_b1 ( .do(bm_sdo_b1_o_0), .di(bm_sdo_b1_o[0]),
     .clk(bm_sck_b0_o), .tielo(tielo_4bram1));
clk_mux2to1_ice8p I_glb_ck_tree_top5432 ( .bl(bl_top[333:330]),
     .gnet(gclk[5:2]), .reset_r(reset_b_r[145:144]),
     .min0({padin_0717a_ck, fabric_out_13_09}), .min1({gclk_r2clktv[0],
     fabric_out_00_09}), .min2({padin_0009a_ck, fabric_out_06_17}),
     .min3({padin_1309a_ck, gclk_l2clktv[1]}),
     .pgate_l(pgate_l[145:144]), .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[145:144]), .reset_l(reset_b_l[145:144]),
     .wl_l(wl_l[145:144]), .wl_r(wl_r[145:144]),
     .pgate_r(pgate_r[145:144]), .vdd_cntl_r(vdd_cntl_r[145:144]));
clk_mux2to1_ice8p I_glb_ck_tree_bot7610 ( .bl(bl_bot[333:330]),
     .gnet({gclk[7], gclk[6], gclk[1], gclk[0]}),
     .reset_r(reset_b_r[143:142]), .min0({padin_1308b_ck,
     gclk_r2clktv[1]}), .min1({padin_0008b_ck, fabric_out_07_17}),
     .min2({gclk_l2clktv[0], fabric_out_00_08}), .min3({padin_0617b_ck,
     fabric_out_13_08}), .pgate_l(pgate_l[143:142]), .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[143:142]), .reset_l(reset_b_l[143:142]),
     .wl_l(wl_l[143:142]), .wl_r(wl_r[143:142]),
     .pgate_r(pgate_r[143:142]), .vdd_cntl_r(vdd_cntl_r[143:142]));
quad_tr_ice1 i_tr_quad ( .update_i(net957), .sp4_h_l_07_17({net818[0],
     net818[1], net818[2], net818[3], net818[4], net818[5], net818[6],
     net818[7], net818[8], net818[9], net818[10], net818[11],
     net818[12], net818[13], net818[14], net818[15]}),
     .lc_bot_07_09(n_inter_07), .bm_sdi_i({tielo_4bram3,
     bm_sdi_b2_o[1]}), .lc_bot_09_09(n_inter_09), .tclk_i(tclkio_mr),
     .shift_i(net969), .sdi(sdio_mr), .r_i(net971), .purst(purst),
     .prog(prog), .mode_i(net974), .slf_op_07_16(slf_op_07_16[7:0]),
     .slf_op_07_15(slf_op_07_15[7:0]),
     .slf_op_07_14(slf_op_07_14[7:0]),
     .slf_op_07_13(slf_op_07_13[7:0]),
     .slf_op_07_12(slf_op_07_12[7:0]),
     .slf_op_07_11(slf_op_07_11[7:0]),
     .slf_op_07_10(slf_op_07_10[7:0]),
     .slf_op_07_09(slf_op_07_09[7:0]),
     .hold_t_r(fabric_out_08_17_ticegate),
     .hold_r_t(fabric_out_13_10_ricegate), .hiz_b_i(net975),
     .glb_in(gclk[7:0]), .ceb_i(net980),
     .carry_in_12_09(carry_io_12_0809),
     .carry_in_11_09(carry_io_11_0809),
     .carry_in_09_09(carry_io_09_0809),
     .carry_in_08_09(carry_io_08_0809), .bs_en_i(net987),
     .sp4_v_b_12_09({net999[0], net999[1], net999[2], net999[3],
     net999[4], net999[5], net999[6], net999[7], net999[8], net999[9],
     net999[10], net999[11], net999[12], net999[13], net999[14],
     net999[15], net999[16], net999[17], net999[18], net999[19],
     net999[20], net999[21], net999[22], net999[23], net999[24],
     net999[25], net999[26], net999[27], net999[28], net999[29],
     net999[30], net999[31], net999[32], net999[33], net999[34],
     net999[35], net999[36], net999[37], net999[38], net999[39],
     net999[40], net999[41], net999[42], net999[43], net999[44],
     net999[45], net999[46], net999[47]}), .sp4_v_b_11_09({net1000[0],
     net1000[1], net1000[2], net1000[3], net1000[4], net1000[5],
     net1000[6], net1000[7], net1000[8], net1000[9], net1000[10],
     net1000[11], net1000[12], net1000[13], net1000[14], net1000[15],
     net1000[16], net1000[17], net1000[18], net1000[19], net1000[20],
     net1000[21], net1000[22], net1000[23], net1000[24], net1000[25],
     net1000[26], net1000[27], net1000[28], net1000[29], net1000[30],
     net1000[31], net1000[32], net1000[33], net1000[34], net1000[35],
     net1000[36], net1000[37], net1000[38], net1000[39], net1000[40],
     net1000[41], net1000[42], net1000[43], net1000[44], net1000[45],
     net1000[46], net1000[47]}), .sp4_v_b_10_09({net1001[0],
     net1001[1], net1001[2], net1001[3], net1001[4], net1001[5],
     net1001[6], net1001[7], net1001[8], net1001[9], net1001[10],
     net1001[11], net1001[12], net1001[13], net1001[14], net1001[15],
     net1001[16], net1001[17], net1001[18], net1001[19], net1001[20],
     net1001[21], net1001[22], net1001[23], net1001[24], net1001[25],
     net1001[26], net1001[27], net1001[28], net1001[29], net1001[30],
     net1001[31], net1001[32], net1001[33], net1001[34], net1001[35],
     net1001[36], net1001[37], net1001[38], net1001[39], net1001[40],
     net1001[41], net1001[42], net1001[43], net1001[44], net1001[45],
     net1001[46], net1001[47]}), .sp4_v_b_09_09({net998[0], net998[1],
     net998[2], net998[3], net998[4], net998[5], net998[6], net998[7],
     net998[8], net998[9], net998[10], net998[11], net998[12],
     net998[13], net998[14], net998[15], net998[16], net998[17],
     net998[18], net998[19], net998[20], net998[21], net998[22],
     net998[23], net998[24], net998[25], net998[26], net998[27],
     net998[28], net998[29], net998[30], net998[31], net998[32],
     net998[33], net998[34], net998[35], net998[36], net998[37],
     net998[38], net998[39], net998[40], net998[41], net998[42],
     net998[43], net998[44], net998[45], net998[46], net998[47]}),
     .sp4_v_b_08_09({net967[0], net967[1], net967[2], net967[3],
     net967[4], net967[5], net967[6], net967[7], net967[8], net967[9],
     net967[10], net967[11], net967[12], net967[13], net967[14],
     net967[15], net967[16], net967[17], net967[18], net967[19],
     net967[20], net967[21], net967[22], net967[23], net967[24],
     net967[25], net967[26], net967[27], net967[28], net967[29],
     net967[30], net967[31], net967[32], net967[33], net967[34],
     net967[35], net967[36], net967[37], net967[38], net967[39],
     net967[40], net967[41], net967[42], net967[43], net967[44],
     net967[45], net967[46], net967[47]}),
     .bnl_op_12_09(slf_op_11_08[7:0]),
     .bnl_op_11_09(slf_op_10_08[7:0]),
     .bnl_op_10_09(slf_op_09_08[7:0]),
     .bnl_op_09_09(slf_op_08_08[7:0]),
     .slf_op_08_09(slf_op_08_09[7:0]),
     .bot_op_12_09(slf_op_12_08[7:0]),
     .bot_op_11_09(slf_op_11_08[7:0]),
     .bot_op_10_09(slf_op_10_08[7:0]),
     .bot_op_09_09(slf_op_09_08[7:0]),
     .bot_op_08_09(slf_op_08_08[7:0]),
     .bot_op_07_09(slf_op_07_08[7:0]), .update_o(net863),
     .tclk_o(tclkio_mt), .bm_wdummymux_en_i(net988),
     .lft_op_07_09(slf_op_06_09[7:0]),
     .carry_in_07_09(carry_io_07_0809),
     .lft_op_07_16(slf_op_06_16[7:0]),
     .slf_op_13_09(slf_op_13_09[3:0]),
     .fabric_out_13_10(fabric_out_13_10_ricegate),
     .slf_op_12_09(slf_op_12_09[7:0]),
     .slf_op_11_09(slf_op_11_09[7:0]),
     .slf_op_10_09(slf_op_10_09[7:0]),
     .slf_op_09_09(slf_op_09_09[7:0]),
     .slf_op_07_17(slf_op_07_17[3:0]), .sp12_h_l_07_16({net770[0],
     net770[1], net770[2], net770[3], net770[4], net770[5], net770[6],
     net770[7], net770[8], net770[9], net770[10], net770[11],
     net770[12], net770[13], net770[14], net770[15], net770[16],
     net770[17], net770[18], net770[19], net770[20], net770[21],
     net770[22], net770[23]}), .sp12_h_l_07_15({net771[0], net771[1],
     net771[2], net771[3], net771[4], net771[5], net771[6], net771[7],
     net771[8], net771[9], net771[10], net771[11], net771[12],
     net771[13], net771[14], net771[15], net771[16], net771[17],
     net771[18], net771[19], net771[20], net771[21], net771[22],
     net771[23]}), .sp12_h_l_07_14({net772[0], net772[1], net772[2],
     net772[3], net772[4], net772[5], net772[6], net772[7], net772[8],
     net772[9], net772[10], net772[11], net772[12], net772[13],
     net772[14], net772[15], net772[16], net772[17], net772[18],
     net772[19], net772[20], net772[21], net772[22], net772[23]}),
     .sp12_h_l_07_13({net773[0], net773[1], net773[2], net773[3],
     net773[4], net773[5], net773[6], net773[7], net773[8], net773[9],
     net773[10], net773[11], net773[12], net773[13], net773[14],
     net773[15], net773[16], net773[17], net773[18], net773[19],
     net773[20], net773[21], net773[22], net773[23]}),
     .sp12_h_l_07_12({net774[0], net774[1], net774[2], net774[3],
     net774[4], net774[5], net774[6], net774[7], net774[8], net774[9],
     net774[10], net774[11], net774[12], net774[13], net774[14],
     net774[15], net774[16], net774[17], net774[18], net774[19],
     net774[20], net774[21], net774[22], net774[23]}),
     .sp12_h_l_07_11({net775[0], net775[1], net775[2], net775[3],
     net775[4], net775[5], net775[6], net775[7], net775[8], net775[9],
     net775[10], net775[11], net775[12], net775[13], net775[14],
     net775[15], net775[16], net775[17], net775[18], net775[19],
     net775[20], net775[21], net775[22], net775[23]}),
     .sp12_h_l_07_10({net776[0], net776[1], net776[2], net776[3],
     net776[4], net776[5], net776[6], net776[7], net776[8], net776[9],
     net776[10], net776[11], net776[12], net776[13], net776[14],
     net776[15], net776[16], net776[17], net776[18], net776[19],
     net776[20], net776[21], net776[22], net776[23]}),
     .sp12_v_b_07_09({net986[0], net986[1], net986[2], net986[3],
     net986[4], net986[5], net986[6], net986[7], net986[8], net986[9],
     net986[10], net986[11], net986[12], net986[13], net986[14],
     net986[15], net986[16], net986[17], net986[18], net986[19],
     net986[20], net986[21], net986[22], net986[23]}),
     .shift_o(net866), .sdo(sdio_mt), .r_o(net876),
     .padin_13_09a(padin_1309a_ck),
     .fabric_out_07_17(fabric_out_07_17),
     .padin_07_17a(padin_0717a_ck), .mode_o(net880), .hiz_b_o(net883),
     .cf_r(cf_r[383:192]), .ceb_o(net858), .bs_en_o(net888),
     .bnr_op_12_09({slf_op_13_08[3], slf_op_13_08[2], slf_op_13_08[1],
     slf_op_13_08[0], slf_op_13_08[3], slf_op_13_08[2],
     slf_op_13_08[1], slf_op_13_08[0]}),
     .bnr_op_11_09(slf_op_12_08[7:0]),
     .bnr_op_10_09(slf_op_11_08[7:0]),
     .bnr_op_09_09(slf_op_10_08[7:0]),
     .bnr_op_08_09(slf_op_09_08[7:0]),
     .bnr_op_07_09(slf_op_08_08[7:0]), .sp4_v_b_07_16({net810[0],
     net810[1], net810[2], net810[3], net810[4], net810[5], net810[6],
     net810[7], net810[8], net810[9], net810[10], net810[11],
     net810[12], net810[13], net810[14], net810[15], net810[16],
     net810[17], net810[18], net810[19], net810[20], net810[21],
     net810[22], net810[23], net810[24], net810[25], net810[26],
     net810[27], net810[28], net810[29], net810[30], net810[31],
     net810[32], net810[33], net810[34], net810[35], net810[36],
     net810[37], net810[38], net810[39], net810[40], net810[41],
     net810[42], net810[43], net810[44], net810[45], net810[46],
     net810[47]}), .sp4_v_b_07_15({net811[0], net811[1], net811[2],
     net811[3], net811[4], net811[5], net811[6], net811[7], net811[8],
     net811[9], net811[10], net811[11], net811[12], net811[13],
     net811[14], net811[15], net811[16], net811[17], net811[18],
     net811[19], net811[20], net811[21], net811[22], net811[23],
     net811[24], net811[25], net811[26], net811[27], net811[28],
     net811[29], net811[30], net811[31], net811[32], net811[33],
     net811[34], net811[35], net811[36], net811[37], net811[38],
     net811[39], net811[40], net811[41], net811[42], net811[43],
     net811[44], net811[45], net811[46], net811[47]}),
     .sp4_v_b_07_14({net812[0], net812[1], net812[2], net812[3],
     net812[4], net812[5], net812[6], net812[7], net812[8], net812[9],
     net812[10], net812[11], net812[12], net812[13], net812[14],
     net812[15], net812[16], net812[17], net812[18], net812[19],
     net812[20], net812[21], net812[22], net812[23], net812[24],
     net812[25], net812[26], net812[27], net812[28], net812[29],
     net812[30], net812[31], net812[32], net812[33], net812[34],
     net812[35], net812[36], net812[37], net812[38], net812[39],
     net812[40], net812[41], net812[42], net812[43], net812[44],
     net812[45], net812[46], net812[47]}), .sp4_v_b_07_13({net813[0],
     net813[1], net813[2], net813[3], net813[4], net813[5], net813[6],
     net813[7], net813[8], net813[9], net813[10], net813[11],
     net813[12], net813[13], net813[14], net813[15], net813[16],
     net813[17], net813[18], net813[19], net813[20], net813[21],
     net813[22], net813[23], net813[24], net813[25], net813[26],
     net813[27], net813[28], net813[29], net813[30], net813[31],
     net813[32], net813[33], net813[34], net813[35], net813[36],
     net813[37], net813[38], net813[39], net813[40], net813[41],
     net813[42], net813[43], net813[44], net813[45], net813[46],
     net813[47]}), .sp4_v_b_07_12({net814[0], net814[1], net814[2],
     net814[3], net814[4], net814[5], net814[6], net814[7], net814[8],
     net814[9], net814[10], net814[11], net814[12], net814[13],
     net814[14], net814[15], net814[16], net814[17], net814[18],
     net814[19], net814[20], net814[21], net814[22], net814[23],
     net814[24], net814[25], net814[26], net814[27], net814[28],
     net814[29], net814[30], net814[31], net814[32], net814[33],
     net814[34], net814[35], net814[36], net814[37], net814[38],
     net814[39], net814[40], net814[41], net814[42], net814[43],
     net814[44], net814[45], net814[46], net814[47]}),
     .sp4_v_b_07_11({net815[0], net815[1], net815[2], net815[3],
     net815[4], net815[5], net815[6], net815[7], net815[8], net815[9],
     net815[10], net815[11], net815[12], net815[13], net815[14],
     net815[15], net815[16], net815[17], net815[18], net815[19],
     net815[20], net815[21], net815[22], net815[23], net815[24],
     net815[25], net815[26], net815[27], net815[28], net815[29],
     net815[30], net815[31], net815[32], net815[33], net815[34],
     net815[35], net815[36], net815[37], net815[38], net815[39],
     net815[40], net815[41], net815[42], net815[43], net815[44],
     net815[45], net815[46], net815[47]}), .sp4_v_b_07_10({net816[0],
     net816[1], net816[2], net816[3], net816[4], net816[5], net816[6],
     net816[7], net816[8], net816[9], net816[10], net816[11],
     net816[12], net816[13], net816[14], net816[15], net816[16],
     net816[17], net816[18], net816[19], net816[20], net816[21],
     net816[22], net816[23], net816[24], net816[25], net816[26],
     net816[27], net816[28], net816[29], net816[30], net816[31],
     net816[32], net816[33], net816[34], net816[35], net816[36],
     net816[37], net816[38], net816[39], net816[40], net816[41],
     net816[42], net816[43], net816[44], net816[45], net816[46],
     net816[47]}), .sp4_v_b_07_09({net921[0], net921[1], net921[2],
     net921[3], net921[4], net921[5], net921[6], net921[7], net921[8],
     net921[9], net921[10], net921[11], net921[12], net921[13],
     net921[14], net921[15], net921[16], net921[17], net921[18],
     net921[19], net921[20], net921[21], net921[22], net921[23],
     net921[24], net921[25], net921[26], net921[27], net921[28],
     net921[29], net921[30], net921[31], net921[32], net921[33],
     net921[34], net921[35], net921[36], net921[37], net921[38],
     net921[39], net921[40], net921[41], net921[42], net921[43],
     net921[44], net921[45], net921[46], net921[47]}),
     .sp12_v_b_12_09({net981[0], net981[1], net981[2], net981[3],
     net981[4], net981[5], net981[6], net981[7], net981[8], net981[9],
     net981[10], net981[11], net981[12], net981[13], net981[14],
     net981[15], net981[16], net981[17], net981[18], net981[19],
     net981[20], net981[21], net981[22], net981[23]}),
     .sp12_v_b_11_09({net982[0], net982[1], net982[2], net982[3],
     net982[4], net982[5], net982[6], net982[7], net982[8], net982[9],
     net982[10], net982[11], net982[12], net982[13], net982[14],
     net982[15], net982[16], net982[17], net982[18], net982[19],
     net982[20], net982[21], net982[22], net982[23]}),
     .sp12_v_b_10_09({net983[0], net983[1], net983[2], net983[3],
     net983[4], net983[5], net983[6], net983[7], net983[8], net983[9],
     net983[10], net983[11], net983[12], net983[13], net983[14],
     net983[15], net983[16], net983[17], net983[18], net983[19],
     net983[20], net983[21], net983[22], net983[23]}),
     .sp12_v_b_09_09({net984[0], net984[1], net984[2], net984[3],
     net984[4], net984[5], net984[6], net984[7], net984[8], net984[9],
     net984[10], net984[11], net984[12], net984[13], net984[14],
     net984[15], net984[16], net984[17], net984[18], net984[19],
     net984[20], net984[21], net984[22], net984[23]}),
     .sp12_v_b_08_09({net985[0], net985[1], net985[2], net985[3],
     net985[4], net985[5], net985[6], net985[7], net985[8], net985[9],
     net985[10], net985[11], net985[12], net985[13], net985[14],
     net985[15], net985[16], net985[17], net985[18], net985[19],
     net985[20], net985[21], net985[22], net985[23]}),
     .fabric_out_13_09(fabric_out_13_09), .pado_t_r(pado_t[23:12]),
     .sp4_h_l_07_16({net819[0], net819[1], net819[2], net819[3],
     net819[4], net819[5], net819[6], net819[7], net819[8], net819[9],
     net819[10], net819[11], net819[12], net819[13], net819[14],
     net819[15], net819[16], net819[17], net819[18], net819[19],
     net819[20], net819[21], net819[22], net819[23], net819[24],
     net819[25], net819[26], net819[27], net819[28], net819[29],
     net819[30], net819[31], net819[32], net819[33], net819[34],
     net819[35], net819[36], net819[37], net819[38], net819[39],
     net819[40], net819[41], net819[42], net819[43], net819[44],
     net819[45], net819[46], net819[47]}), .sp4_h_l_07_15({net820[0],
     net820[1], net820[2], net820[3], net820[4], net820[5], net820[6],
     net820[7], net820[8], net820[9], net820[10], net820[11],
     net820[12], net820[13], net820[14], net820[15], net820[16],
     net820[17], net820[18], net820[19], net820[20], net820[21],
     net820[22], net820[23], net820[24], net820[25], net820[26],
     net820[27], net820[28], net820[29], net820[30], net820[31],
     net820[32], net820[33], net820[34], net820[35], net820[36],
     net820[37], net820[38], net820[39], net820[40], net820[41],
     net820[42], net820[43], net820[44], net820[45], net820[46],
     net820[47]}), .sp4_h_l_07_14({net821[0], net821[1], net821[2],
     net821[3], net821[4], net821[5], net821[6], net821[7], net821[8],
     net821[9], net821[10], net821[11], net821[12], net821[13],
     net821[14], net821[15], net821[16], net821[17], net821[18],
     net821[19], net821[20], net821[21], net821[22], net821[23],
     net821[24], net821[25], net821[26], net821[27], net821[28],
     net821[29], net821[30], net821[31], net821[32], net821[33],
     net821[34], net821[35], net821[36], net821[37], net821[38],
     net821[39], net821[40], net821[41], net821[42], net821[43],
     net821[44], net821[45], net821[46], net821[47]}),
     .sp4_h_l_07_13({net822[0], net822[1], net822[2], net822[3],
     net822[4], net822[5], net822[6], net822[7], net822[8], net822[9],
     net822[10], net822[11], net822[12], net822[13], net822[14],
     net822[15], net822[16], net822[17], net822[18], net822[19],
     net822[20], net822[21], net822[22], net822[23], net822[24],
     net822[25], net822[26], net822[27], net822[28], net822[29],
     net822[30], net822[31], net822[32], net822[33], net822[34],
     net822[35], net822[36], net822[37], net822[38], net822[39],
     net822[40], net822[41], net822[42], net822[43], net822[44],
     net822[45], net822[46], net822[47]}), .sp4_h_l_07_12({net823[0],
     net823[1], net823[2], net823[3], net823[4], net823[5], net823[6],
     net823[7], net823[8], net823[9], net823[10], net823[11],
     net823[12], net823[13], net823[14], net823[15], net823[16],
     net823[17], net823[18], net823[19], net823[20], net823[21],
     net823[22], net823[23], net823[24], net823[25], net823[26],
     net823[27], net823[28], net823[29], net823[30], net823[31],
     net823[32], net823[33], net823[34], net823[35], net823[36],
     net823[37], net823[38], net823[39], net823[40], net823[41],
     net823[42], net823[43], net823[44], net823[45], net823[46],
     net823[47]}), .sp4_h_l_07_11({net824[0], net824[1], net824[2],
     net824[3], net824[4], net824[5], net824[6], net824[7], net824[8],
     net824[9], net824[10], net824[11], net824[12], net824[13],
     net824[14], net824[15], net824[16], net824[17], net824[18],
     net824[19], net824[20], net824[21], net824[22], net824[23],
     net824[24], net824[25], net824[26], net824[27], net824[28],
     net824[29], net824[30], net824[31], net824[32], net824[33],
     net824[34], net824[35], net824[36], net824[37], net824[38],
     net824[39], net824[40], net824[41], net824[42], net824[43],
     net824[44], net824[45], net824[46], net824[47]}),
     .sp4_h_l_07_10({net849[0], net849[1], net849[2], net849[3],
     net849[4], net849[5], net849[6], net849[7], net849[8], net849[9],
     net849[10], net849[11], net849[12], net849[13], net849[14],
     net849[15], net849[16], net849[17], net849[18], net849[19],
     net849[20], net849[21], net849[22], net849[23], net849[24],
     net849[25], net849[26], net849[27], net849[28], net849[29],
     net849[30], net849[31], net849[32], net849[33], net849[34],
     net849[35], net849[36], net849[37], net849[38], net849[39],
     net849[40], net849[41], net849[42], net849[43], net849[44],
     net849[45], net849[46], net849[47]}),
     .bnl_op_08_09(slf_op_07_08[7:0]),
     .bnl_op_13_09(slf_op_12_08[7:0]),
     .lft_op_07_15(slf_op_06_15[7:0]),
     .lft_op_07_14(slf_op_06_14[7:0]),
     .lft_op_07_13(slf_op_06_13[7:0]),
     .lft_op_07_12(slf_op_06_12[7:0]),
     .lft_op_07_11(slf_op_06_11[7:0]),
     .lft_op_07_10(slf_op_06_10[7:0]),
     .vdd_cntl_r(vdd_cntl_r[287:144]), .wl_r(wl_r[287:144]),
     .reset_b_r(reset_b_r[287:144]), .pado_r(pado_r[24:13]),
     .padeb_r(padeb_r[24:13]), .padin_r(padin_r[24:13]),
     .bnl_op_07_09(slf_op_06_08[7:0]), .sp4_h_l_07_09({net848[0],
     net848[1], net848[2], net848[3], net848[4], net848[5], net848[6],
     net848[7], net848[8], net848[9], net848[10], net848[11],
     net848[12], net848[13], net848[14], net848[15], net848[16],
     net848[17], net848[18], net848[19], net848[20], net848[21],
     net848[22], net848[23], net848[24], net848[25], net848[26],
     net848[27], net848[28], net848[29], net848[30], net848[31],
     net848[32], net848[33], net848[34], net848[35], net848[36],
     net848[37], net848[38], net848[39], net848[40], net848[41],
     net848[42], net848[43], net848[44], net848[45], net848[46],
     net848[47]}), .sp12_h_l_07_09({net777[0], net777[1], net777[2],
     net777[3], net777[4], net777[5], net777[6], net777[7], net777[8],
     net777[9], net777[10], net777[11], net777[12], net777[13],
     net777[14], net777[15], net777[16], net777[17], net777[18],
     net777[19], net777[20], net777[21], net777[22], net777[23]}),
     .lc_bot_11_09(n_inter_11), .lc_bot_12_09(n_inter_12),
     .sp4_h_r_13_09({net911[0], net911[1], net911[2], net911[3],
     net911[4], net911[5], net911[6], net911[7], net911[8], net911[9],
     net911[10], net911[11], net911[12], net911[13], net911[14],
     net911[15]}), .bl(bl_top[663:334]), .pgate_r(pgate_r[287:144]),
     .cf_t(cf_t[287:144]), .lc_bot_08_09(n_inter_08),
     .bm_aa_2bot({net1071[0], net1071[1], net1071[2], net1071[3],
     net1071[4], net1071[5], net1071[6], net1071[7], net1071[8],
     net1071[9], net1071[10]}), .bm_ab_2bot({net1046[0], net1046[1],
     net1046[2], net1046[3], net1046[4], net1046[5], net1046[6],
     net1046[7], net1046[8], net1046[9], net1046[10]}),
     .bm_init_i(net997), .bm_rcapmux_en_i(net996), .bm_sa_i({net995[0],
     net995[1], net995[2], net995[3], net995[4], net995[5], net995[6],
     net995[7]}), .bm_sclk_i(bm_sck_b2_o), .bm_sclkrw_i({tielo_4bram3,
     bm_sclkrw_b2_o[1]}), .bm_sdo_o(bm_sdo_b3_o[1:0]),
     .padin_t_r(padin_t[23:12]), .bm_sreb_i(net990),
     .bm_sweb_i({tielo_4bram3, bm_sweb_b2_o[1]}),
     .padeb_t_r(padeb_t[23:12]),
     .fabric_out_08_17(fabric_out_08_17_ticegate),
     .tnl_op_07_16(slf_op_06_17[3:0]));
quad_tl_ice1 i_tl_quad ( .padin_l_t(padin_l[23:12]),
     .pado_l_t(pado_l[23:12]), .padeb_l_t(padeb_l[23:12]),
     .fo_dlyadj(fo_dlyadj[7:3]), .padin_06_17b(padin_0617b_ck),
     .padin_00_09a(padin_0009a_ck), .padeb_t_l(padeb_t[11:0]),
     .mode_o(net1135), .hiz_b_o(net1136),
     .fabric_out_06_17(fabric_out_06_17),
     .fabric_out_00_09(fabric_out_00_09), .cf_t(cf_t[143:0]),
     .cf_l(cf_l[383:192]), .ceb_o(net1139), .bs_en_o(net1140),
     .bm_sdi_i({tielo_4bram1, bm_sdi_b0_o[1]}),
     .bm_sdo_o(bm_sdo_b1_o[1:0]), .sp12_v_b_02_09({net1171[0],
     net1171[1], net1171[2], net1171[3], net1171[4], net1171[5],
     net1171[6], net1171[7], net1171[8], net1171[9], net1171[10],
     net1171[11], net1171[12], net1171[13], net1171[14], net1171[15],
     net1171[16], net1171[17], net1171[18], net1171[19], net1171[20],
     net1171[21], net1171[22], net1171[23]}),
     .sp12_v_b_01_09({net1103[0], net1103[1], net1103[2], net1103[3],
     net1103[4], net1103[5], net1103[6], net1103[7], net1103[8],
     net1103[9], net1103[10], net1103[11], net1103[12], net1103[13],
     net1103[14], net1103[15], net1103[16], net1103[17], net1103[18],
     net1103[19], net1103[20], net1103[21], net1103[22], net1103[23]}),
     .sp12_h_r_06_16({net770[0], net770[1], net770[2], net770[3],
     net770[4], net770[5], net770[6], net770[7], net770[8], net770[9],
     net770[10], net770[11], net770[12], net770[13], net770[14],
     net770[15], net770[16], net770[17], net770[18], net770[19],
     net770[20], net770[21], net770[22], net770[23]}),
     .sp12_h_r_06_15({net771[0], net771[1], net771[2], net771[3],
     net771[4], net771[5], net771[6], net771[7], net771[8], net771[9],
     net771[10], net771[11], net771[12], net771[13], net771[14],
     net771[15], net771[16], net771[17], net771[18], net771[19],
     net771[20], net771[21], net771[22], net771[23]}),
     .sp12_h_r_06_14({net772[0], net772[1], net772[2], net772[3],
     net772[4], net772[5], net772[6], net772[7], net772[8], net772[9],
     net772[10], net772[11], net772[12], net772[13], net772[14],
     net772[15], net772[16], net772[17], net772[18], net772[19],
     net772[20], net772[21], net772[22], net772[23]}),
     .sp12_h_r_06_13({net773[0], net773[1], net773[2], net773[3],
     net773[4], net773[5], net773[6], net773[7], net773[8], net773[9],
     net773[10], net773[11], net773[12], net773[13], net773[14],
     net773[15], net773[16], net773[17], net773[18], net773[19],
     net773[20], net773[21], net773[22], net773[23]}),
     .sp12_h_r_06_12({net774[0], net774[1], net774[2], net774[3],
     net774[4], net774[5], net774[6], net774[7], net774[8], net774[9],
     net774[10], net774[11], net774[12], net774[13], net774[14],
     net774[15], net774[16], net774[17], net774[18], net774[19],
     net774[20], net774[21], net774[22], net774[23]}),
     .sp12_h_r_06_11({net775[0], net775[1], net775[2], net775[3],
     net775[4], net775[5], net775[6], net775[7], net775[8], net775[9],
     net775[10], net775[11], net775[12], net775[13], net775[14],
     net775[15], net775[16], net775[17], net775[18], net775[19],
     net775[20], net775[21], net775[22], net775[23]}),
     .sp12_h_r_06_10({net776[0], net776[1], net776[2], net776[3],
     net776[4], net776[5], net776[6], net776[7], net776[8], net776[9],
     net776[10], net776[11], net776[12], net776[13], net776[14],
     net776[15], net776[16], net776[17], net776[18], net776[19],
     net776[20], net776[21], net776[22], net776[23]}),
     .sp12_h_r_06_09({net777[0], net777[1], net777[2], net777[3],
     net777[4], net777[5], net777[6], net777[7], net777[8], net777[9],
     net777[10], net777[11], net777[12], net777[13], net777[14],
     net777[15], net777[16], net777[17], net777[18], net777[19],
     net777[20], net777[21], net777[22], net777[23]}),
     .vdd_cntl_l(vdd_cntl_l[287:144]), .sp12_v_b_05_09({net1170[0],
     net1170[1], net1170[2], net1170[3], net1170[4], net1170[5],
     net1170[6], net1170[7], net1170[8], net1170[9], net1170[10],
     net1170[11], net1170[12], net1170[13], net1170[14], net1170[15],
     net1170[16], net1170[17], net1170[18], net1170[19], net1170[20],
     net1170[21], net1170[22], net1170[23]}),
     .slf_op_06_17(slf_op_06_17[3:0]), .tclk_o(tclkio_ml),
     .update_o(net1102), .wl_l(wl_l[287:144]),
     .slf_op_06_16(slf_op_06_16[7:0]),
     .slf_op_06_15(slf_op_06_15[7:0]),
     .slf_op_06_14(slf_op_06_14[7:0]),
     .slf_op_06_13(slf_op_06_13[7:0]),
     .slf_op_06_12(slf_op_06_12[7:0]),
     .slf_op_06_11(slf_op_06_11[7:0]), .bm_wdummymux_en_i(net1183),
     .bm_sreb_i(net1185), .bm_sweb_i({tielo_4bram1, bm_sweb_b0_o[1]}),
     .sp12_v_b_03_09({net1231[0], net1231[1], net1231[2], net1231[3],
     net1231[4], net1231[5], net1231[6], net1231[7], net1231[8],
     net1231[9], net1231[10], net1231[11], net1231[12], net1231[13],
     net1231[14], net1231[15], net1231[16], net1231[17], net1231[18],
     net1231[19], net1231[20], net1231[21], net1231[22], net1231[23]}),
     .shift_o(net1124), .sdo(sdio_ml), .r_o(net1132),
     .pado_t_l(pado_t[11:0]), .sp12_v_b_04_09({net1196[0], net1196[1],
     net1196[2], net1196[3], net1196[4], net1196[5], net1196[6],
     net1196[7], net1196[8], net1196[9], net1196[10], net1196[11],
     net1196[12], net1196[13], net1196[14], net1196[15], net1196[16],
     net1196[17], net1196[18], net1196[19], net1196[20], net1196[21],
     net1196[22], net1196[23]}), .sp12_v_b_06_09({net1195[0],
     net1195[1], net1195[2], net1195[3], net1195[4], net1195[5],
     net1195[6], net1195[7], net1195[8], net1195[9], net1195[10],
     net1195[11], net1195[12], net1195[13], net1195[14], net1195[15],
     net1195[16], net1195[17], net1195[18], net1195[19], net1195[20],
     net1195[21], net1195[22], net1195[23]}),
     .sp4_v_b_06_09({net1212[0], net1212[1], net1212[2], net1212[3],
     net1212[4], net1212[5], net1212[6], net1212[7], net1212[8],
     net1212[9], net1212[10], net1212[11], net1212[12], net1212[13],
     net1212[14], net1212[15], net1212[16], net1212[17], net1212[18],
     net1212[19], net1212[20], net1212[21], net1212[22], net1212[23],
     net1212[24], net1212[25], net1212[26], net1212[27], net1212[28],
     net1212[29], net1212[30], net1212[31], net1212[32], net1212[33],
     net1212[34], net1212[35], net1212[36], net1212[37], net1212[38],
     net1212[39], net1212[40], net1212[41], net1212[42], net1212[43],
     net1212[44], net1212[45], net1212[46], net1212[47]}),
     .slf_op_06_10(slf_op_06_10[7:0]), .sp4_v_b_05_09({net1213[0],
     net1213[1], net1213[2], net1213[3], net1213[4], net1213[5],
     net1213[6], net1213[7], net1213[8], net1213[9], net1213[10],
     net1213[11], net1213[12], net1213[13], net1213[14], net1213[15],
     net1213[16], net1213[17], net1213[18], net1213[19], net1213[20],
     net1213[21], net1213[22], net1213[23], net1213[24], net1213[25],
     net1213[26], net1213[27], net1213[28], net1213[29], net1213[30],
     net1213[31], net1213[32], net1213[33], net1213[34], net1213[35],
     net1213[36], net1213[37], net1213[38], net1213[39], net1213[40],
     net1213[41], net1213[42], net1213[43], net1213[44], net1213[45],
     net1213[46], net1213[47]}), .sp4_v_b_04_09({net1214[0],
     net1214[1], net1214[2], net1214[3], net1214[4], net1214[5],
     net1214[6], net1214[7], net1214[8], net1214[9], net1214[10],
     net1214[11], net1214[12], net1214[13], net1214[14], net1214[15],
     net1214[16], net1214[17], net1214[18], net1214[19], net1214[20],
     net1214[21], net1214[22], net1214[23], net1214[24], net1214[25],
     net1214[26], net1214[27], net1214[28], net1214[29], net1214[30],
     net1214[31], net1214[32], net1214[33], net1214[34], net1214[35],
     net1214[36], net1214[37], net1214[38], net1214[39], net1214[40],
     net1214[41], net1214[42], net1214[43], net1214[44], net1214[45],
     net1214[46], net1214[47]}), .bnl_op_04_09(slf_op_03_08[7:0]),
     .bnl_op_05_09(slf_op_04_08[7:0]), .lc_bot_05_09(n_inter_05),
     .sp4_v_b_02_09({net1216[0], net1216[1], net1216[2], net1216[3],
     net1216[4], net1216[5], net1216[6], net1216[7], net1216[8],
     net1216[9], net1216[10], net1216[11], net1216[12], net1216[13],
     net1216[14], net1216[15], net1216[16], net1216[17], net1216[18],
     net1216[19], net1216[20], net1216[21], net1216[22], net1216[23],
     net1216[24], net1216[25], net1216[26], net1216[27], net1216[28],
     net1216[29], net1216[30], net1216[31], net1216[32], net1216[33],
     net1216[34], net1216[35], net1216[36], net1216[37], net1216[38],
     net1216[39], net1216[40], net1216[41], net1216[42], net1216[43],
     net1216[44], net1216[45], net1216[46], net1216[47]}),
     .sp4_v_b_01_09({net1115[0], net1115[1], net1115[2], net1115[3],
     net1115[4], net1115[5], net1115[6], net1115[7], net1115[8],
     net1115[9], net1115[10], net1115[11], net1115[12], net1115[13],
     net1115[14], net1115[15], net1115[16], net1115[17], net1115[18],
     net1115[19], net1115[20], net1115[21], net1115[22], net1115[23],
     net1115[24], net1115[25], net1115[26], net1115[27], net1115[28],
     net1115[29], net1115[30], net1115[31], net1115[32], net1115[33],
     net1115[34], net1115[35], net1115[36], net1115[37], net1115[38],
     net1115[39], net1115[40], net1115[41], net1115[42], net1115[43],
     net1115[44], net1115[45], net1115[46], net1115[47]}),
     .sp4_v_b_00_09({net1250[0], net1250[1], net1250[2], net1250[3],
     net1250[4], net1250[5], net1250[6], net1250[7], net1250[8],
     net1250[9], net1250[10], net1250[11], net1250[12], net1250[13],
     net1250[14], net1250[15]}), .sp4_r_v_b_06_16({net810[0],
     net810[1], net810[2], net810[3], net810[4], net810[5], net810[6],
     net810[7], net810[8], net810[9], net810[10], net810[11],
     net810[12], net810[13], net810[14], net810[15], net810[16],
     net810[17], net810[18], net810[19], net810[20], net810[21],
     net810[22], net810[23], net810[24], net810[25], net810[26],
     net810[27], net810[28], net810[29], net810[30], net810[31],
     net810[32], net810[33], net810[34], net810[35], net810[36],
     net810[37], net810[38], net810[39], net810[40], net810[41],
     net810[42], net810[43], net810[44], net810[45], net810[46],
     net810[47]}), .sp4_r_v_b_06_15({net811[0], net811[1], net811[2],
     net811[3], net811[4], net811[5], net811[6], net811[7], net811[8],
     net811[9], net811[10], net811[11], net811[12], net811[13],
     net811[14], net811[15], net811[16], net811[17], net811[18],
     net811[19], net811[20], net811[21], net811[22], net811[23],
     net811[24], net811[25], net811[26], net811[27], net811[28],
     net811[29], net811[30], net811[31], net811[32], net811[33],
     net811[34], net811[35], net811[36], net811[37], net811[38],
     net811[39], net811[40], net811[41], net811[42], net811[43],
     net811[44], net811[45], net811[46], net811[47]}),
     .sp4_r_v_b_06_14({net812[0], net812[1], net812[2], net812[3],
     net812[4], net812[5], net812[6], net812[7], net812[8], net812[9],
     net812[10], net812[11], net812[12], net812[13], net812[14],
     net812[15], net812[16], net812[17], net812[18], net812[19],
     net812[20], net812[21], net812[22], net812[23], net812[24],
     net812[25], net812[26], net812[27], net812[28], net812[29],
     net812[30], net812[31], net812[32], net812[33], net812[34],
     net812[35], net812[36], net812[37], net812[38], net812[39],
     net812[40], net812[41], net812[42], net812[43], net812[44],
     net812[45], net812[46], net812[47]}), .sp4_r_v_b_06_13({net813[0],
     net813[1], net813[2], net813[3], net813[4], net813[5], net813[6],
     net813[7], net813[8], net813[9], net813[10], net813[11],
     net813[12], net813[13], net813[14], net813[15], net813[16],
     net813[17], net813[18], net813[19], net813[20], net813[21],
     net813[22], net813[23], net813[24], net813[25], net813[26],
     net813[27], net813[28], net813[29], net813[30], net813[31],
     net813[32], net813[33], net813[34], net813[35], net813[36],
     net813[37], net813[38], net813[39], net813[40], net813[41],
     net813[42], net813[43], net813[44], net813[45], net813[46],
     net813[47]}), .sp4_r_v_b_06_12({net814[0], net814[1], net814[2],
     net814[3], net814[4], net814[5], net814[6], net814[7], net814[8],
     net814[9], net814[10], net814[11], net814[12], net814[13],
     net814[14], net814[15], net814[16], net814[17], net814[18],
     net814[19], net814[20], net814[21], net814[22], net814[23],
     net814[24], net814[25], net814[26], net814[27], net814[28],
     net814[29], net814[30], net814[31], net814[32], net814[33],
     net814[34], net814[35], net814[36], net814[37], net814[38],
     net814[39], net814[40], net814[41], net814[42], net814[43],
     net814[44], net814[45], net814[46], net814[47]}),
     .sp4_r_v_b_06_11({net815[0], net815[1], net815[2], net815[3],
     net815[4], net815[5], net815[6], net815[7], net815[8], net815[9],
     net815[10], net815[11], net815[12], net815[13], net815[14],
     net815[15], net815[16], net815[17], net815[18], net815[19],
     net815[20], net815[21], net815[22], net815[23], net815[24],
     net815[25], net815[26], net815[27], net815[28], net815[29],
     net815[30], net815[31], net815[32], net815[33], net815[34],
     net815[35], net815[36], net815[37], net815[38], net815[39],
     net815[40], net815[41], net815[42], net815[43], net815[44],
     net815[45], net815[46], net815[47]}), .sp4_r_v_b_06_10({net816[0],
     net816[1], net816[2], net816[3], net816[4], net816[5], net816[6],
     net816[7], net816[8], net816[9], net816[10], net816[11],
     net816[12], net816[13], net816[14], net816[15], net816[16],
     net816[17], net816[18], net816[19], net816[20], net816[21],
     net816[22], net816[23], net816[24], net816[25], net816[26],
     net816[27], net816[28], net816[29], net816[30], net816[31],
     net816[32], net816[33], net816[34], net816[35], net816[36],
     net816[37], net816[38], net816[39], net816[40], net816[41],
     net816[42], net816[43], net816[44], net816[45], net816[46],
     net816[47]}), .sp4_r_v_b_06_09({net921[0], net921[1], net921[2],
     net921[3], net921[4], net921[5], net921[6], net921[7], net921[8],
     net921[9], net921[10], net921[11], net921[12], net921[13],
     net921[14], net921[15], net921[16], net921[17], net921[18],
     net921[19], net921[20], net921[21], net921[22], net921[23],
     net921[24], net921[25], net921[26], net921[27], net921[28],
     net921[29], net921[30], net921[31], net921[32], net921[33],
     net921[34], net921[35], net921[36], net921[37], net921[38],
     net921[39], net921[40], net921[41], net921[42], net921[43],
     net921[44], net921[45], net921[46], net921[47]}),
     .sp4_h_r_06_17({net818[0], net818[1], net818[2], net818[3],
     net818[4], net818[5], net818[6], net818[7], net818[8], net818[9],
     net818[10], net818[11], net818[12], net818[13], net818[14],
     net818[15]}), .sp4_h_r_06_16({net819[0], net819[1], net819[2],
     net819[3], net819[4], net819[5], net819[6], net819[7], net819[8],
     net819[9], net819[10], net819[11], net819[12], net819[13],
     net819[14], net819[15], net819[16], net819[17], net819[18],
     net819[19], net819[20], net819[21], net819[22], net819[23],
     net819[24], net819[25], net819[26], net819[27], net819[28],
     net819[29], net819[30], net819[31], net819[32], net819[33],
     net819[34], net819[35], net819[36], net819[37], net819[38],
     net819[39], net819[40], net819[41], net819[42], net819[43],
     net819[44], net819[45], net819[46], net819[47]}),
     .sp4_h_r_06_15({net820[0], net820[1], net820[2], net820[3],
     net820[4], net820[5], net820[6], net820[7], net820[8], net820[9],
     net820[10], net820[11], net820[12], net820[13], net820[14],
     net820[15], net820[16], net820[17], net820[18], net820[19],
     net820[20], net820[21], net820[22], net820[23], net820[24],
     net820[25], net820[26], net820[27], net820[28], net820[29],
     net820[30], net820[31], net820[32], net820[33], net820[34],
     net820[35], net820[36], net820[37], net820[38], net820[39],
     net820[40], net820[41], net820[42], net820[43], net820[44],
     net820[45], net820[46], net820[47]}), .sp4_h_r_06_14({net821[0],
     net821[1], net821[2], net821[3], net821[4], net821[5], net821[6],
     net821[7], net821[8], net821[9], net821[10], net821[11],
     net821[12], net821[13], net821[14], net821[15], net821[16],
     net821[17], net821[18], net821[19], net821[20], net821[21],
     net821[22], net821[23], net821[24], net821[25], net821[26],
     net821[27], net821[28], net821[29], net821[30], net821[31],
     net821[32], net821[33], net821[34], net821[35], net821[36],
     net821[37], net821[38], net821[39], net821[40], net821[41],
     net821[42], net821[43], net821[44], net821[45], net821[46],
     net821[47]}), .sp4_h_r_06_13({net822[0], net822[1], net822[2],
     net822[3], net822[4], net822[5], net822[6], net822[7], net822[8],
     net822[9], net822[10], net822[11], net822[12], net822[13],
     net822[14], net822[15], net822[16], net822[17], net822[18],
     net822[19], net822[20], net822[21], net822[22], net822[23],
     net822[24], net822[25], net822[26], net822[27], net822[28],
     net822[29], net822[30], net822[31], net822[32], net822[33],
     net822[34], net822[35], net822[36], net822[37], net822[38],
     net822[39], net822[40], net822[41], net822[42], net822[43],
     net822[44], net822[45], net822[46], net822[47]}),
     .sp4_h_r_06_12({net823[0], net823[1], net823[2], net823[3],
     net823[4], net823[5], net823[6], net823[7], net823[8], net823[9],
     net823[10], net823[11], net823[12], net823[13], net823[14],
     net823[15], net823[16], net823[17], net823[18], net823[19],
     net823[20], net823[21], net823[22], net823[23], net823[24],
     net823[25], net823[26], net823[27], net823[28], net823[29],
     net823[30], net823[31], net823[32], net823[33], net823[34],
     net823[35], net823[36], net823[37], net823[38], net823[39],
     net823[40], net823[41], net823[42], net823[43], net823[44],
     net823[45], net823[46], net823[47]}), .sp4_h_r_06_11({net824[0],
     net824[1], net824[2], net824[3], net824[4], net824[5], net824[6],
     net824[7], net824[8], net824[9], net824[10], net824[11],
     net824[12], net824[13], net824[14], net824[15], net824[16],
     net824[17], net824[18], net824[19], net824[20], net824[21],
     net824[22], net824[23], net824[24], net824[25], net824[26],
     net824[27], net824[28], net824[29], net824[30], net824[31],
     net824[32], net824[33], net824[34], net824[35], net824[36],
     net824[37], net824[38], net824[39], net824[40], net824[41],
     net824[42], net824[43], net824[44], net824[45], net824[46],
     net824[47]}), .bnl_op_03_09(slf_op_02_08[7:0]),
     .bnl_op_02_09(slf_op_01_08[7:0]), .bnl_op_01_09({slf_op_00_08[3],
     slf_op_00_08[2], slf_op_00_08[1], slf_op_00_08[0],
     slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0]}), .slf_op_00_09(slf_op_00_09[3:0]),
     .slf_op_06_09(slf_op_06_09[7:0]),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .lc_bot_01_09(n_inter_01), .lc_bot_02_09(n_inter_02),
     .lc_bot_04_09(n_inter_04), .bnl_op_06_09(slf_op_05_08[7:0]),
     .bnr_op_00_09(slf_op_01_08[7:0]),
     .bnr_op_01_09(slf_op_02_08[7:0]),
     .bnr_op_02_09(slf_op_03_08[7:0]),
     .bnr_op_03_09(slf_op_04_08[7:0]), .last_rsr(last_rsr[1]),
     .slf_op_05_09(slf_op_05_09[7:0]),
     .slf_op_04_09(slf_op_04_09[7:0]),
     .slf_op_03_09(slf_op_03_09[7:0]),
     .slf_op_02_09(slf_op_02_09[7:0]),
     .slf_op_01_09(slf_op_01_09[7:0]), .bl(bl_top[329:0]),
     .pgate_l(pgate_l[287:144]), .reset_b_l(reset_b_l[287:144]),
     .sp4_h_r_06_09({net848[0], net848[1], net848[2], net848[3],
     net848[4], net848[5], net848[6], net848[7], net848[8], net848[9],
     net848[10], net848[11], net848[12], net848[13], net848[14],
     net848[15], net848[16], net848[17], net848[18], net848[19],
     net848[20], net848[21], net848[22], net848[23], net848[24],
     net848[25], net848[26], net848[27], net848[28], net848[29],
     net848[30], net848[31], net848[32], net848[33], net848[34],
     net848[35], net848[36], net848[37], net848[38], net848[39],
     net848[40], net848[41], net848[42], net848[43], net848[44],
     net848[45], net848[46], net848[47]}), .sp4_h_r_06_10({net849[0],
     net849[1], net849[2], net849[3], net849[4], net849[5], net849[6],
     net849[7], net849[8], net849[9], net849[10], net849[11],
     net849[12], net849[13], net849[14], net849[15], net849[16],
     net849[17], net849[18], net849[19], net849[20], net849[21],
     net849[22], net849[23], net849[24], net849[25], net849[26],
     net849[27], net849[28], net849[29], net849[30], net849[31],
     net849[32], net849[33], net849[34], net849[35], net849[36],
     net849[37], net849[38], net849[39], net849[40], net849[41],
     net849[42], net849[43], net849[44], net849[45], net849[46],
     net849[47]}), .bnr_op_04_09(slf_op_05_08[7:0]),
     .bnr_op_05_09(slf_op_06_08[7:0]),
     .bnr_op_06_09(slf_op_07_08[7:0]),
     .bot_op_01_09(slf_op_01_08[7:0]),
     .carry_in_05_09(carry_io_05_0809),
     .carry_in_02_09(carry_io_02_0809),
     .carry_in_04_09(carry_io_04_0809),
     .carry_in_06_09(carry_io_06_0809), .ceb_i(net858),
     .bot_op_05_09(slf_op_05_08[7:0]),
     .bot_op_02_09(slf_op_02_08[7:0]),
     .bot_op_03_09(slf_op_03_08[7:0]),
     .bot_op_04_09(slf_op_04_08[7:0]), .update_i(net863),
     .tnr_op_06_16(slf_op_07_17[3:0]), .tclk_i(tclkio_mt),
     .shift_i(net866), .sdi(sdio_mt), .rgt_op_06_16(slf_op_07_16[7:0]),
     .rgt_op_06_15(slf_op_07_15[7:0]),
     .rgt_op_06_14(slf_op_07_14[7:0]),
     .rgt_op_06_13(slf_op_07_13[7:0]),
     .rgt_op_06_12(slf_op_07_12[7:0]),
     .rgt_op_06_11(slf_op_07_11[7:0]),
     .rgt_op_06_10(slf_op_07_10[7:0]),
     .rgt_op_06_09(slf_op_07_09[7:0]), .r_i(net876), .purst(purst),
     .prog(prog), .padin_t_l(padin_t[11:0]), .mode_i(net880),
     .hold_t_l(fabric_out_08_17_ticegate),
     .hold_l_t(fabric_out_00_07_licegate), .hiz_b_i(net883),
     .glb_in(gclk[7:0]), .lc_bot_06_09(n_inter_06),
     .sp4_v_b_03_09({net1215[0], net1215[1], net1215[2], net1215[3],
     net1215[4], net1215[5], net1215[6], net1215[7], net1215[8],
     net1215[9], net1215[10], net1215[11], net1215[12], net1215[13],
     net1215[14], net1215[15], net1215[16], net1215[17], net1215[18],
     net1215[19], net1215[20], net1215[21], net1215[22], net1215[23],
     net1215[24], net1215[25], net1215[26], net1215[27], net1215[28],
     net1215[29], net1215[30], net1215[31], net1215[32], net1215[33],
     net1215[34], net1215[35], net1215[36], net1215[37], net1215[38],
     net1215[39], net1215[40], net1215[41], net1215[42], net1215[43],
     net1215[44], net1215[45], net1215[46], net1215[47]}),
     .carry_in_01_09(carry_io_01_0809), .bs_en_i(net888),
     .bot_op_06_09(slf_op_06_08[7:0]), .bm_ab_2bot({net1232[0],
     net1232[1], net1232[2], net1232[3], net1232[4], net1232[5],
     net1232[6], net1232[7], net1232[8], net1232[9], net1232[10]}),
     .bm_aa_2bot({net1138[0], net1138[1], net1138[2], net1138[3],
     net1138[4], net1138[5], net1138[6], net1138[7], net1138[8],
     net1138[9], net1138[10]}), .bm_init_i(net1192),
     .bm_rcapmux_en_i(net1191), .bm_sa_i({net1190[0], net1190[1],
     net1190[2], net1190[3], net1190[4], net1190[5], net1190[6],
     net1190[7]}), .bm_sclk_i(bm_sck_b0_o), .bm_sclkrw_i({tielo_4bram1,
     bm_sclkrw_b0_o[1]}));
quad_br_ice1 i_br_quad ( net997, net996, {net995[0], net995[1],
     net995[2], net995[3], net995[4], net995[5], net995[6], net995[7]},
     bm_sck_b2_o, bm_sclkrw_b2_o[1:0], bm_sdi_b2_o[1:0],
     bm_sdo_b2_o[1:0], net990, bm_sweb_b2_o[1:0], net988, net987,
     carry_io_07_0809, carry_io_08_0809, carry_io_09_0809,
     carry_io_11_0809, carry_io_12_0809, net980, cf_b[287:144],
     cf_r[191:0], fabric_out_07_00, fabric_out_12_00_wb,
     fabric_out_13_01, fabric_out_13_02, fabric_out_13_08, net975,
     net974, n_inter_07, n_inter_08, n_inter_09, n_inter_11,
     n_inter_12, padeb_b[11], padeb_b[23:13], padeb_r[12:0],
     padin_0700a_ck, padin_1308b_ck, pado_b[11], pado_b[23:13],
     pado_r[12:0], net971, sdio_mr, sdo_pad, net969, slf_op_07_00[3:0],
     slf_op_07_01[7:0], slf_op_07_02[7:0], slf_op_07_03[7:0],
     slf_op_07_04[7:0], slf_op_07_05[7:0], slf_op_07_06[7:0],
     slf_op_07_07[7:0], slf_op_07_08[7:0], slf_op_08_08[7:0],
     slf_op_09_08[7:0], slf_op_10_08[7:0], slf_op_11_08[7:0],
     slf_op_12_08[7:0], slf_op_13_08[3:0], spi_ss_in_bbank[4:0],
     tck_pad, tclkio_mr, tdi_pad, tms_pad, net957, bl_bot[663:334],
     pgate_r[143:0], reset_b_r[143:0], {net1154[0], net1154[1],
     net1154[2], net1154[3], net1154[4], net1154[5], net1154[6],
     net1154[7], net1154[8], net1154[9], net1154[10], net1154[11],
     net1154[12], net1154[13], net1154[14], net1154[15]}, {net1227[0],
     net1227[1], net1227[2], net1227[3], net1227[4], net1227[5],
     net1227[6], net1227[7], net1227[8], net1227[9], net1227[10],
     net1227[11], net1227[12], net1227[13], net1227[14], net1227[15],
     net1227[16], net1227[17], net1227[18], net1227[19], net1227[20],
     net1227[21], net1227[22], net1227[23], net1227[24], net1227[25],
     net1227[26], net1227[27], net1227[28], net1227[29], net1227[30],
     net1227[31], net1227[32], net1227[33], net1227[34], net1227[35],
     net1227[36], net1227[37], net1227[38], net1227[39], net1227[40],
     net1227[41], net1227[42], net1227[43], net1227[44], net1227[45],
     net1227[46], net1227[47]}, {net1226[0], net1226[1], net1226[2],
     net1226[3], net1226[4], net1226[5], net1226[6], net1226[7],
     net1226[8], net1226[9], net1226[10], net1226[11], net1226[12],
     net1226[13], net1226[14], net1226[15], net1226[16], net1226[17],
     net1226[18], net1226[19], net1226[20], net1226[21], net1226[22],
     net1226[23], net1226[24], net1226[25], net1226[26], net1226[27],
     net1226[28], net1226[29], net1226[30], net1226[31], net1226[32],
     net1226[33], net1226[34], net1226[35], net1226[36], net1226[37],
     net1226[38], net1226[39], net1226[40], net1226[41], net1226[42],
     net1226[43], net1226[44], net1226[45], net1226[46], net1226[47]},
     {net1225[0], net1225[1], net1225[2], net1225[3], net1225[4],
     net1225[5], net1225[6], net1225[7], net1225[8], net1225[9],
     net1225[10], net1225[11], net1225[12], net1225[13], net1225[14],
     net1225[15], net1225[16], net1225[17], net1225[18], net1225[19],
     net1225[20], net1225[21], net1225[22], net1225[23], net1225[24],
     net1225[25], net1225[26], net1225[27], net1225[28], net1225[29],
     net1225[30], net1225[31], net1225[32], net1225[33], net1225[34],
     net1225[35], net1225[36], net1225[37], net1225[38], net1225[39],
     net1225[40], net1225[41], net1225[42], net1225[43], net1225[44],
     net1225[45], net1225[46], net1225[47]}, {net1224[0], net1224[1],
     net1224[2], net1224[3], net1224[4], net1224[5], net1224[6],
     net1224[7], net1224[8], net1224[9], net1224[10], net1224[11],
     net1224[12], net1224[13], net1224[14], net1224[15], net1224[16],
     net1224[17], net1224[18], net1224[19], net1224[20], net1224[21],
     net1224[22], net1224[23], net1224[24], net1224[25], net1224[26],
     net1224[27], net1224[28], net1224[29], net1224[30], net1224[31],
     net1224[32], net1224[33], net1224[34], net1224[35], net1224[36],
     net1224[37], net1224[38], net1224[39], net1224[40], net1224[41],
     net1224[42], net1224[43], net1224[44], net1224[45], net1224[46],
     net1224[47]}, {net1223[0], net1223[1], net1223[2], net1223[3],
     net1223[4], net1223[5], net1223[6], net1223[7], net1223[8],
     net1223[9], net1223[10], net1223[11], net1223[12], net1223[13],
     net1223[14], net1223[15], net1223[16], net1223[17], net1223[18],
     net1223[19], net1223[20], net1223[21], net1223[22], net1223[23],
     net1223[24], net1223[25], net1223[26], net1223[27], net1223[28],
     net1223[29], net1223[30], net1223[31], net1223[32], net1223[33],
     net1223[34], net1223[35], net1223[36], net1223[37], net1223[38],
     net1223[39], net1223[40], net1223[41], net1223[42], net1223[43],
     net1223[44], net1223[45], net1223[46], net1223[47]}, {net1228[0],
     net1228[1], net1228[2], net1228[3], net1228[4], net1228[5],
     net1228[6], net1228[7], net1228[8], net1228[9], net1228[10],
     net1228[11], net1228[12], net1228[13], net1228[14], net1228[15],
     net1228[16], net1228[17], net1228[18], net1228[19], net1228[20],
     net1228[21], net1228[22], net1228[23], net1228[24], net1228[25],
     net1228[26], net1228[27], net1228[28], net1228[29], net1228[30],
     net1228[31], net1228[32], net1228[33], net1228[34], net1228[35],
     net1228[36], net1228[37], net1228[38], net1228[39], net1228[40],
     net1228[41], net1228[42], net1228[43], net1228[44], net1228[45],
     net1228[46], net1228[47]}, {net1242[0], net1242[1], net1242[2],
     net1242[3], net1242[4], net1242[5], net1242[6], net1242[7],
     net1242[8], net1242[9], net1242[10], net1242[11], net1242[12],
     net1242[13], net1242[14], net1242[15], net1242[16], net1242[17],
     net1242[18], net1242[19], net1242[20], net1242[21], net1242[22],
     net1242[23], net1242[24], net1242[25], net1242[26], net1242[27],
     net1242[28], net1242[29], net1242[30], net1242[31], net1242[32],
     net1242[33], net1242[34], net1242[35], net1242[36], net1242[37],
     net1242[38], net1242[39], net1242[40], net1242[41], net1242[42],
     net1242[43], net1242[44], net1242[45], net1242[46], net1242[47]},
     {net1241[0], net1241[1], net1241[2], net1241[3], net1241[4],
     net1241[5], net1241[6], net1241[7], net1241[8], net1241[9],
     net1241[10], net1241[11], net1241[12], net1241[13], net1241[14],
     net1241[15], net1241[16], net1241[17], net1241[18], net1241[19],
     net1241[20], net1241[21], net1241[22], net1241[23], net1241[24],
     net1241[25], net1241[26], net1241[27], net1241[28], net1241[29],
     net1241[30], net1241[31], net1241[32], net1241[33], net1241[34],
     net1241[35], net1241[36], net1241[37], net1241[38], net1241[39],
     net1241[40], net1241[41], net1241[42], net1241[43], net1241[44],
     net1241[45], net1241[46], net1241[47]}, {net1221[0], net1221[1],
     net1221[2], net1221[3], net1221[4], net1221[5], net1221[6],
     net1221[7], net1221[8], net1221[9], net1221[10], net1221[11],
     net1221[12], net1221[13], net1221[14], net1221[15], net1221[16],
     net1221[17], net1221[18], net1221[19], net1221[20], net1221[21],
     net1221[22], net1221[23], net1221[24], net1221[25], net1221[26],
     net1221[27], net1221[28], net1221[29], net1221[30], net1221[31],
     net1221[32], net1221[33], net1221[34], net1221[35], net1221[36],
     net1221[37], net1221[38], net1221[39], net1221[40], net1221[41],
     net1221[42], net1221[43], net1221[44], net1221[45], net1221[46],
     net1221[47]}, {net1220[0], net1220[1], net1220[2], net1220[3],
     net1220[4], net1220[5], net1220[6], net1220[7], net1220[8],
     net1220[9], net1220[10], net1220[11], net1220[12], net1220[13],
     net1220[14], net1220[15], net1220[16], net1220[17], net1220[18],
     net1220[19], net1220[20], net1220[21], net1220[22], net1220[23],
     net1220[24], net1220[25], net1220[26], net1220[27], net1220[28],
     net1220[29], net1220[30], net1220[31], net1220[32], net1220[33],
     net1220[34], net1220[35], net1220[36], net1220[37], net1220[38],
     net1220[39], net1220[40], net1220[41], net1220[42], net1220[43],
     net1220[44], net1220[45], net1220[46], net1220[47]}, {net1219[0],
     net1219[1], net1219[2], net1219[3], net1219[4], net1219[5],
     net1219[6], net1219[7], net1219[8], net1219[9], net1219[10],
     net1219[11], net1219[12], net1219[13], net1219[14], net1219[15],
     net1219[16], net1219[17], net1219[18], net1219[19], net1219[20],
     net1219[21], net1219[22], net1219[23], net1219[24], net1219[25],
     net1219[26], net1219[27], net1219[28], net1219[29], net1219[30],
     net1219[31], net1219[32], net1219[33], net1219[34], net1219[35],
     net1219[36], net1219[37], net1219[38], net1219[39], net1219[40],
     net1219[41], net1219[42], net1219[43], net1219[44], net1219[45],
     net1219[46], net1219[47]}, {net1218[0], net1218[1], net1218[2],
     net1218[3], net1218[4], net1218[5], net1218[6], net1218[7],
     net1218[8], net1218[9], net1218[10], net1218[11], net1218[12],
     net1218[13], net1218[14], net1218[15], net1218[16], net1218[17],
     net1218[18], net1218[19], net1218[20], net1218[21], net1218[22],
     net1218[23], net1218[24], net1218[25], net1218[26], net1218[27],
     net1218[28], net1218[29], net1218[30], net1218[31], net1218[32],
     net1218[33], net1218[34], net1218[35], net1218[36], net1218[37],
     net1218[38], net1218[39], net1218[40], net1218[41], net1218[42],
     net1218[43], net1218[44], net1218[45], net1218[46], net1218[47]},
     {net1217[0], net1217[1], net1217[2], net1217[3], net1217[4],
     net1217[5], net1217[6], net1217[7], net1217[8], net1217[9],
     net1217[10], net1217[11], net1217[12], net1217[13], net1217[14],
     net1217[15], net1217[16], net1217[17], net1217[18], net1217[19],
     net1217[20], net1217[21], net1217[22], net1217[23], net1217[24],
     net1217[25], net1217[26], net1217[27], net1217[28], net1217[29],
     net1217[30], net1217[31], net1217[32], net1217[33], net1217[34],
     net1217[35], net1217[36], net1217[37], net1217[38], net1217[39],
     net1217[40], net1217[41], net1217[42], net1217[43], net1217[44],
     net1217[45], net1217[46], net1217[47]}, {net1199[0], net1199[1],
     net1199[2], net1199[3], net1199[4], net1199[5], net1199[6],
     net1199[7], net1199[8], net1199[9], net1199[10], net1199[11],
     net1199[12], net1199[13], net1199[14], net1199[15], net1199[16],
     net1199[17], net1199[18], net1199[19], net1199[20], net1199[21],
     net1199[22], net1199[23], net1199[24], net1199[25], net1199[26],
     net1199[27], net1199[28], net1199[29], net1199[30], net1199[31],
     net1199[32], net1199[33], net1199[34], net1199[35], net1199[36],
     net1199[37], net1199[38], net1199[39], net1199[40], net1199[41],
     net1199[42], net1199[43], net1199[44], net1199[45], net1199[46],
     net1199[47]}, {net1200[0], net1200[1], net1200[2], net1200[3],
     net1200[4], net1200[5], net1200[6], net1200[7], net1200[8],
     net1200[9], net1200[10], net1200[11], net1200[12], net1200[13],
     net1200[14], net1200[15], net1200[16], net1200[17], net1200[18],
     net1200[19], net1200[20], net1200[21], net1200[22], net1200[23],
     net1200[24], net1200[25], net1200[26], net1200[27], net1200[28],
     net1200[29], net1200[30], net1200[31], net1200[32], net1200[33],
     net1200[34], net1200[35], net1200[36], net1200[37], net1200[38],
     net1200[39], net1200[40], net1200[41], net1200[42], net1200[43],
     net1200[44], net1200[45], net1200[46], net1200[47]}, {net1165[0],
     net1165[1], net1165[2], net1165[3], net1165[4], net1165[5],
     net1165[6], net1165[7], net1165[8], net1165[9], net1165[10],
     net1165[11], net1165[12], net1165[13], net1165[14], net1165[15],
     net1165[16], net1165[17], net1165[18], net1165[19], net1165[20],
     net1165[21], net1165[22], net1165[23], net1165[24], net1165[25],
     net1165[26], net1165[27], net1165[28], net1165[29], net1165[30],
     net1165[31], net1165[32], net1165[33], net1165[34], net1165[35],
     net1165[36], net1165[37], net1165[38], net1165[39], net1165[40],
     net1165[41], net1165[42], net1165[43], net1165[44], net1165[45],
     net1165[46], net1165[47]}, {net921[0], net921[1], net921[2],
     net921[3], net921[4], net921[5], net921[6], net921[7], net921[8],
     net921[9], net921[10], net921[11], net921[12], net921[13],
     net921[14], net921[15], net921[16], net921[17], net921[18],
     net921[19], net921[20], net921[21], net921[22], net921[23],
     net921[24], net921[25], net921[26], net921[27], net921[28],
     net921[29], net921[30], net921[31], net921[32], net921[33],
     net921[34], net921[35], net921[36], net921[37], net921[38],
     net921[39], net921[40], net921[41], net921[42], net921[43],
     net921[44], net921[45], net921[46], net921[47]}, {net967[0],
     net967[1], net967[2], net967[3], net967[4], net967[5], net967[6],
     net967[7], net967[8], net967[9], net967[10], net967[11],
     net967[12], net967[13], net967[14], net967[15], net967[16],
     net967[17], net967[18], net967[19], net967[20], net967[21],
     net967[22], net967[23], net967[24], net967[25], net967[26],
     net967[27], net967[28], net967[29], net967[30], net967[31],
     net967[32], net967[33], net967[34], net967[35], net967[36],
     net967[37], net967[38], net967[39], net967[40], net967[41],
     net967[42], net967[43], net967[44], net967[45], net967[46],
     net967[47]}, {net998[0], net998[1], net998[2], net998[3],
     net998[4], net998[5], net998[6], net998[7], net998[8], net998[9],
     net998[10], net998[11], net998[12], net998[13], net998[14],
     net998[15], net998[16], net998[17], net998[18], net998[19],
     net998[20], net998[21], net998[22], net998[23], net998[24],
     net998[25], net998[26], net998[27], net998[28], net998[29],
     net998[30], net998[31], net998[32], net998[33], net998[34],
     net998[35], net998[36], net998[37], net998[38], net998[39],
     net998[40], net998[41], net998[42], net998[43], net998[44],
     net998[45], net998[46], net998[47]}, {net1001[0], net1001[1],
     net1001[2], net1001[3], net1001[4], net1001[5], net1001[6],
     net1001[7], net1001[8], net1001[9], net1001[10], net1001[11],
     net1001[12], net1001[13], net1001[14], net1001[15], net1001[16],
     net1001[17], net1001[18], net1001[19], net1001[20], net1001[21],
     net1001[22], net1001[23], net1001[24], net1001[25], net1001[26],
     net1001[27], net1001[28], net1001[29], net1001[30], net1001[31],
     net1001[32], net1001[33], net1001[34], net1001[35], net1001[36],
     net1001[37], net1001[38], net1001[39], net1001[40], net1001[41],
     net1001[42], net1001[43], net1001[44], net1001[45], net1001[46],
     net1001[47]}, {net1000[0], net1000[1], net1000[2], net1000[3],
     net1000[4], net1000[5], net1000[6], net1000[7], net1000[8],
     net1000[9], net1000[10], net1000[11], net1000[12], net1000[13],
     net1000[14], net1000[15], net1000[16], net1000[17], net1000[18],
     net1000[19], net1000[20], net1000[21], net1000[22], net1000[23],
     net1000[24], net1000[25], net1000[26], net1000[27], net1000[28],
     net1000[29], net1000[30], net1000[31], net1000[32], net1000[33],
     net1000[34], net1000[35], net1000[36], net1000[37], net1000[38],
     net1000[39], net1000[40], net1000[41], net1000[42], net1000[43],
     net1000[44], net1000[45], net1000[46], net1000[47]}, {net999[0],
     net999[1], net999[2], net999[3], net999[4], net999[5], net999[6],
     net999[7], net999[8], net999[9], net999[10], net999[11],
     net999[12], net999[13], net999[14], net999[15], net999[16],
     net999[17], net999[18], net999[19], net999[20], net999[21],
     net999[22], net999[23], net999[24], net999[25], net999[26],
     net999[27], net999[28], net999[29], net999[30], net999[31],
     net999[32], net999[33], net999[34], net999[35], net999[36],
     net999[37], net999[38], net999[39], net999[40], net999[41],
     net999[42], net999[43], net999[44], net999[45], net999[46],
     net999[47]}, {net911[0], net911[1], net911[2], net911[3],
     net911[4], net911[5], net911[6], net911[7], net911[8], net911[9],
     net911[10], net911[11], net911[12], net911[13], net911[14],
     net911[15]}, {net1209[0], net1209[1], net1209[2], net1209[3],
     net1209[4], net1209[5], net1209[6], net1209[7], net1209[8],
     net1209[9], net1209[10], net1209[11], net1209[12], net1209[13],
     net1209[14], net1209[15], net1209[16], net1209[17], net1209[18],
     net1209[19], net1209[20], net1209[21], net1209[22], net1209[23]},
     {net1208[0], net1208[1], net1208[2], net1208[3], net1208[4],
     net1208[5], net1208[6], net1208[7], net1208[8], net1208[9],
     net1208[10], net1208[11], net1208[12], net1208[13], net1208[14],
     net1208[15], net1208[16], net1208[17], net1208[18], net1208[19],
     net1208[20], net1208[21], net1208[22], net1208[23]}, {net1207[0],
     net1207[1], net1207[2], net1207[3], net1207[4], net1207[5],
     net1207[6], net1207[7], net1207[8], net1207[9], net1207[10],
     net1207[11], net1207[12], net1207[13], net1207[14], net1207[15],
     net1207[16], net1207[17], net1207[18], net1207[19], net1207[20],
     net1207[21], net1207[22], net1207[23]}, {net1206[0], net1206[1],
     net1206[2], net1206[3], net1206[4], net1206[5], net1206[6],
     net1206[7], net1206[8], net1206[9], net1206[10], net1206[11],
     net1206[12], net1206[13], net1206[14], net1206[15], net1206[16],
     net1206[17], net1206[18], net1206[19], net1206[20], net1206[21],
     net1206[22], net1206[23]}, {net1205[0], net1205[1], net1205[2],
     net1205[3], net1205[4], net1205[5], net1205[6], net1205[7],
     net1205[8], net1205[9], net1205[10], net1205[11], net1205[12],
     net1205[13], net1205[14], net1205[15], net1205[16], net1205[17],
     net1205[18], net1205[19], net1205[20], net1205[21], net1205[22],
     net1205[23]}, {net1198[0], net1198[1], net1198[2], net1198[3],
     net1198[4], net1198[5], net1198[6], net1198[7], net1198[8],
     net1198[9], net1198[10], net1198[11], net1198[12], net1198[13],
     net1198[14], net1198[15], net1198[16], net1198[17], net1198[18],
     net1198[19], net1198[20], net1198[21], net1198[22], net1198[23]},
     {net1197[0], net1197[1], net1197[2], net1197[3], net1197[4],
     net1197[5], net1197[6], net1197[7], net1197[8], net1197[9],
     net1197[10], net1197[11], net1197[12], net1197[13], net1197[14],
     net1197[15], net1197[16], net1197[17], net1197[18], net1197[19],
     net1197[20], net1197[21], net1197[22], net1197[23]}, {net1222[0],
     net1222[1], net1222[2], net1222[3], net1222[4], net1222[5],
     net1222[6], net1222[7], net1222[8], net1222[9], net1222[10],
     net1222[11], net1222[12], net1222[13], net1222[14], net1222[15],
     net1222[16], net1222[17], net1222[18], net1222[19], net1222[20],
     net1222[21], net1222[22], net1222[23]}, {net986[0], net986[1],
     net986[2], net986[3], net986[4], net986[5], net986[6], net986[7],
     net986[8], net986[9], net986[10], net986[11], net986[12],
     net986[13], net986[14], net986[15], net986[16], net986[17],
     net986[18], net986[19], net986[20], net986[21], net986[22],
     net986[23]}, {net985[0], net985[1], net985[2], net985[3],
     net985[4], net985[5], net985[6], net985[7], net985[8], net985[9],
     net985[10], net985[11], net985[12], net985[13], net985[14],
     net985[15], net985[16], net985[17], net985[18], net985[19],
     net985[20], net985[21], net985[22], net985[23]}, {net984[0],
     net984[1], net984[2], net984[3], net984[4], net984[5], net984[6],
     net984[7], net984[8], net984[9], net984[10], net984[11],
     net984[12], net984[13], net984[14], net984[15], net984[16],
     net984[17], net984[18], net984[19], net984[20], net984[21],
     net984[22], net984[23]}, {net983[0], net983[1], net983[2],
     net983[3], net983[4], net983[5], net983[6], net983[7], net983[8],
     net983[9], net983[10], net983[11], net983[12], net983[13],
     net983[14], net983[15], net983[16], net983[17], net983[18],
     net983[19], net983[20], net983[21], net983[22], net983[23]},
     {net982[0], net982[1], net982[2], net982[3], net982[4], net982[5],
     net982[6], net982[7], net982[8], net982[9], net982[10],
     net982[11], net982[12], net982[13], net982[14], net982[15],
     net982[16], net982[17], net982[18], net982[19], net982[20],
     net982[21], net982[22], net982[23]}, {net981[0], net981[1],
     net981[2], net981[3], net981[4], net981[5], net981[6], net981[7],
     net981[8], net981[9], net981[10], net981[11], net981[12],
     net981[13], net981[14], net981[15], net981[16], net981[17],
     net981[18], net981[19], net981[20], net981[21], net981[22],
     net981[23]}, vdd_cntl_r[143:0], wl_r[143:0], {net1071[0],
     net1071[1], net1071[2], net1071[3], net1071[4], net1071[5],
     net1071[6], net1071[7], net1071[8], net1071[9], net1071[10]},
     {net1046[0], net1046[1], net1046[2], net1046[3], net1046[4],
     net1046[5], net1046[6], net1046[7], net1046[8], net1046[9],
     net1046[10]}, bm_bank30_init_o, bm_bank30_rcapmux_en_o,
     bm_bank30_sa_o[7:0], bm_bank30_sclk_o[1], {net952[0], net952[1]},
     bm_bank30_sdi_o[3:2], {bm_sdo_b3_o_0, bm_sdi_b2_o[0]},
     bm_bank30_sreb_o, {net948[0], net948[1]}, bm_wdummymux_en_o,
     slf_op_06_00[3:0], net1182, bs_en, net1176, ceb, end_of_startup,
     gclk[7:0], net1167, hiz_b, fabric_out_05_00_bicegate,
     fabric_out_13_10_ricegate, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr[2], last_rsr[3],
     slf_op_06_01[7:0], slf_op_06_02[7:0], slf_op_06_03[7:0],
     slf_op_06_04[7:0], slf_op_06_05[7:0], slf_op_06_06[7:0],
     slf_op_06_07[7:0], slf_op_06_08[7:0], md_spi_b, net1166, mode,
     mux_jtag_sel_b, padin_b[11], padin_b[23:13], padin_r[12:0],
     pll_sdo, prog, purst, net1164, r, sdio_mb, sdi_pad, sdo_enable,
     net1162, shift, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out,
     tclkio_mb, tclk, slf_op_06_09[7:0], slf_op_07_09[7:0],
     slf_op_08_09[7:0], slf_op_09_09[7:0], slf_op_10_09[7:0],
     slf_op_11_09[7:0], slf_op_12_09[7:0], slf_op_08_09[7:0],
     slf_op_09_09[7:0], slf_op_10_09[7:0], slf_op_11_09[7:0],
     slf_op_12_09[7:0], {slf_op_13_09[3], slf_op_13_09[2],
     slf_op_13_09[1], slf_op_13_09[0], slf_op_13_09[3],
     slf_op_13_09[2], slf_op_13_09[1], slf_op_13_09[0]},
     slf_op_07_09[7:0], slf_op_08_09[7:0], slf_op_09_09[7:0],
     slf_op_10_09[7:0], slf_op_11_09[7:0], slf_op_12_09[7:0], totdopad,
     trstb_pad, net1152, update);
quad_bl_ice1 i_bl_quad ( net1192, net1191, {net1190[0], net1190[1],
     net1190[2], net1190[3], net1190[4], net1190[5], net1190[6],
     net1190[7]}, bm_sck_b0_o, bm_sclkrw_b0_o[1:0], bm_sdi_b0_o[1:0],
     bm_sdo_b0_o[1:0], net1185, bm_sweb_b0_o[1:0], net1183, net1182,
     carry_io_01_0809, carry_io_02_0809, carry_io_04_0809,
     carry_io_05_0809, carry_io_06_0809, net1176, cf_b[143:0],
     cf_l[191:0], fabric_out_00_07_licegate, fabric_out_00_08,
     fabric_out_05_00_bicegate, fabric_out_06_00, fo_bypass,
     fo_dlyadj[2:0], fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, net1167,
     net1166, n_inter_01, n_inter_02, n_inter_04, n_inter_05,
     n_inter_06, padeb_b[10:0], padeb_b[12], padeb_l[11:0],
     padin_0008b_ck, padin_0600b_ck, pado_b[10:0], pado_b[12],
     pado_l[11:0], net1164, sdio_mb, net1162, slf_op_00_08[3:0],
     slf_op_01_08[7:0], slf_op_02_08[7:0], slf_op_03_08[7:0],
     slf_op_04_08[7:0], slf_op_05_08[7:0], slf_op_06_00[3:0],
     slf_op_06_01[7:0], slf_op_06_02[7:0], slf_op_06_03[7:0],
     slf_op_06_04[7:0], slf_op_06_05[7:0], slf_op_06_06[7:0],
     slf_op_06_07[7:0], slf_op_06_08[7:0], tclkio_mb, net1152,
     bl_bot[329:0], pgate_l[143:0], reset_b_l[143:0], {net1154[0],
     net1154[1], net1154[2], net1154[3], net1154[4], net1154[5],
     net1154[6], net1154[7], net1154[8], net1154[9], net1154[10],
     net1154[11], net1154[12], net1154[13], net1154[14], net1154[15]},
     {net1227[0], net1227[1], net1227[2], net1227[3], net1227[4],
     net1227[5], net1227[6], net1227[7], net1227[8], net1227[9],
     net1227[10], net1227[11], net1227[12], net1227[13], net1227[14],
     net1227[15], net1227[16], net1227[17], net1227[18], net1227[19],
     net1227[20], net1227[21], net1227[22], net1227[23], net1227[24],
     net1227[25], net1227[26], net1227[27], net1227[28], net1227[29],
     net1227[30], net1227[31], net1227[32], net1227[33], net1227[34],
     net1227[35], net1227[36], net1227[37], net1227[38], net1227[39],
     net1227[40], net1227[41], net1227[42], net1227[43], net1227[44],
     net1227[45], net1227[46], net1227[47]}, {net1226[0], net1226[1],
     net1226[2], net1226[3], net1226[4], net1226[5], net1226[6],
     net1226[7], net1226[8], net1226[9], net1226[10], net1226[11],
     net1226[12], net1226[13], net1226[14], net1226[15], net1226[16],
     net1226[17], net1226[18], net1226[19], net1226[20], net1226[21],
     net1226[22], net1226[23], net1226[24], net1226[25], net1226[26],
     net1226[27], net1226[28], net1226[29], net1226[30], net1226[31],
     net1226[32], net1226[33], net1226[34], net1226[35], net1226[36],
     net1226[37], net1226[38], net1226[39], net1226[40], net1226[41],
     net1226[42], net1226[43], net1226[44], net1226[45], net1226[46],
     net1226[47]}, {net1225[0], net1225[1], net1225[2], net1225[3],
     net1225[4], net1225[5], net1225[6], net1225[7], net1225[8],
     net1225[9], net1225[10], net1225[11], net1225[12], net1225[13],
     net1225[14], net1225[15], net1225[16], net1225[17], net1225[18],
     net1225[19], net1225[20], net1225[21], net1225[22], net1225[23],
     net1225[24], net1225[25], net1225[26], net1225[27], net1225[28],
     net1225[29], net1225[30], net1225[31], net1225[32], net1225[33],
     net1225[34], net1225[35], net1225[36], net1225[37], net1225[38],
     net1225[39], net1225[40], net1225[41], net1225[42], net1225[43],
     net1225[44], net1225[45], net1225[46], net1225[47]}, {net1224[0],
     net1224[1], net1224[2], net1224[3], net1224[4], net1224[5],
     net1224[6], net1224[7], net1224[8], net1224[9], net1224[10],
     net1224[11], net1224[12], net1224[13], net1224[14], net1224[15],
     net1224[16], net1224[17], net1224[18], net1224[19], net1224[20],
     net1224[21], net1224[22], net1224[23], net1224[24], net1224[25],
     net1224[26], net1224[27], net1224[28], net1224[29], net1224[30],
     net1224[31], net1224[32], net1224[33], net1224[34], net1224[35],
     net1224[36], net1224[37], net1224[38], net1224[39], net1224[40],
     net1224[41], net1224[42], net1224[43], net1224[44], net1224[45],
     net1224[46], net1224[47]}, {net1223[0], net1223[1], net1223[2],
     net1223[3], net1223[4], net1223[5], net1223[6], net1223[7],
     net1223[8], net1223[9], net1223[10], net1223[11], net1223[12],
     net1223[13], net1223[14], net1223[15], net1223[16], net1223[17],
     net1223[18], net1223[19], net1223[20], net1223[21], net1223[22],
     net1223[23], net1223[24], net1223[25], net1223[26], net1223[27],
     net1223[28], net1223[29], net1223[30], net1223[31], net1223[32],
     net1223[33], net1223[34], net1223[35], net1223[36], net1223[37],
     net1223[38], net1223[39], net1223[40], net1223[41], net1223[42],
     net1223[43], net1223[44], net1223[45], net1223[46], net1223[47]},
     {net1228[0], net1228[1], net1228[2], net1228[3], net1228[4],
     net1228[5], net1228[6], net1228[7], net1228[8], net1228[9],
     net1228[10], net1228[11], net1228[12], net1228[13], net1228[14],
     net1228[15], net1228[16], net1228[17], net1228[18], net1228[19],
     net1228[20], net1228[21], net1228[22], net1228[23], net1228[24],
     net1228[25], net1228[26], net1228[27], net1228[28], net1228[29],
     net1228[30], net1228[31], net1228[32], net1228[33], net1228[34],
     net1228[35], net1228[36], net1228[37], net1228[38], net1228[39],
     net1228[40], net1228[41], net1228[42], net1228[43], net1228[44],
     net1228[45], net1228[46], net1228[47]}, {net1242[0], net1242[1],
     net1242[2], net1242[3], net1242[4], net1242[5], net1242[6],
     net1242[7], net1242[8], net1242[9], net1242[10], net1242[11],
     net1242[12], net1242[13], net1242[14], net1242[15], net1242[16],
     net1242[17], net1242[18], net1242[19], net1242[20], net1242[21],
     net1242[22], net1242[23], net1242[24], net1242[25], net1242[26],
     net1242[27], net1242[28], net1242[29], net1242[30], net1242[31],
     net1242[32], net1242[33], net1242[34], net1242[35], net1242[36],
     net1242[37], net1242[38], net1242[39], net1242[40], net1242[41],
     net1242[42], net1242[43], net1242[44], net1242[45], net1242[46],
     net1242[47]}, {net1241[0], net1241[1], net1241[2], net1241[3],
     net1241[4], net1241[5], net1241[6], net1241[7], net1241[8],
     net1241[9], net1241[10], net1241[11], net1241[12], net1241[13],
     net1241[14], net1241[15], net1241[16], net1241[17], net1241[18],
     net1241[19], net1241[20], net1241[21], net1241[22], net1241[23],
     net1241[24], net1241[25], net1241[26], net1241[27], net1241[28],
     net1241[29], net1241[30], net1241[31], net1241[32], net1241[33],
     net1241[34], net1241[35], net1241[36], net1241[37], net1241[38],
     net1241[39], net1241[40], net1241[41], net1241[42], net1241[43],
     net1241[44], net1241[45], net1241[46], net1241[47]}, {net1221[0],
     net1221[1], net1221[2], net1221[3], net1221[4], net1221[5],
     net1221[6], net1221[7], net1221[8], net1221[9], net1221[10],
     net1221[11], net1221[12], net1221[13], net1221[14], net1221[15],
     net1221[16], net1221[17], net1221[18], net1221[19], net1221[20],
     net1221[21], net1221[22], net1221[23], net1221[24], net1221[25],
     net1221[26], net1221[27], net1221[28], net1221[29], net1221[30],
     net1221[31], net1221[32], net1221[33], net1221[34], net1221[35],
     net1221[36], net1221[37], net1221[38], net1221[39], net1221[40],
     net1221[41], net1221[42], net1221[43], net1221[44], net1221[45],
     net1221[46], net1221[47]}, {net1220[0], net1220[1], net1220[2],
     net1220[3], net1220[4], net1220[5], net1220[6], net1220[7],
     net1220[8], net1220[9], net1220[10], net1220[11], net1220[12],
     net1220[13], net1220[14], net1220[15], net1220[16], net1220[17],
     net1220[18], net1220[19], net1220[20], net1220[21], net1220[22],
     net1220[23], net1220[24], net1220[25], net1220[26], net1220[27],
     net1220[28], net1220[29], net1220[30], net1220[31], net1220[32],
     net1220[33], net1220[34], net1220[35], net1220[36], net1220[37],
     net1220[38], net1220[39], net1220[40], net1220[41], net1220[42],
     net1220[43], net1220[44], net1220[45], net1220[46], net1220[47]},
     {net1219[0], net1219[1], net1219[2], net1219[3], net1219[4],
     net1219[5], net1219[6], net1219[7], net1219[8], net1219[9],
     net1219[10], net1219[11], net1219[12], net1219[13], net1219[14],
     net1219[15], net1219[16], net1219[17], net1219[18], net1219[19],
     net1219[20], net1219[21], net1219[22], net1219[23], net1219[24],
     net1219[25], net1219[26], net1219[27], net1219[28], net1219[29],
     net1219[30], net1219[31], net1219[32], net1219[33], net1219[34],
     net1219[35], net1219[36], net1219[37], net1219[38], net1219[39],
     net1219[40], net1219[41], net1219[42], net1219[43], net1219[44],
     net1219[45], net1219[46], net1219[47]}, {net1218[0], net1218[1],
     net1218[2], net1218[3], net1218[4], net1218[5], net1218[6],
     net1218[7], net1218[8], net1218[9], net1218[10], net1218[11],
     net1218[12], net1218[13], net1218[14], net1218[15], net1218[16],
     net1218[17], net1218[18], net1218[19], net1218[20], net1218[21],
     net1218[22], net1218[23], net1218[24], net1218[25], net1218[26],
     net1218[27], net1218[28], net1218[29], net1218[30], net1218[31],
     net1218[32], net1218[33], net1218[34], net1218[35], net1218[36],
     net1218[37], net1218[38], net1218[39], net1218[40], net1218[41],
     net1218[42], net1218[43], net1218[44], net1218[45], net1218[46],
     net1218[47]}, {net1217[0], net1217[1], net1217[2], net1217[3],
     net1217[4], net1217[5], net1217[6], net1217[7], net1217[8],
     net1217[9], net1217[10], net1217[11], net1217[12], net1217[13],
     net1217[14], net1217[15], net1217[16], net1217[17], net1217[18],
     net1217[19], net1217[20], net1217[21], net1217[22], net1217[23],
     net1217[24], net1217[25], net1217[26], net1217[27], net1217[28],
     net1217[29], net1217[30], net1217[31], net1217[32], net1217[33],
     net1217[34], net1217[35], net1217[36], net1217[37], net1217[38],
     net1217[39], net1217[40], net1217[41], net1217[42], net1217[43],
     net1217[44], net1217[45], net1217[46], net1217[47]}, {net1199[0],
     net1199[1], net1199[2], net1199[3], net1199[4], net1199[5],
     net1199[6], net1199[7], net1199[8], net1199[9], net1199[10],
     net1199[11], net1199[12], net1199[13], net1199[14], net1199[15],
     net1199[16], net1199[17], net1199[18], net1199[19], net1199[20],
     net1199[21], net1199[22], net1199[23], net1199[24], net1199[25],
     net1199[26], net1199[27], net1199[28], net1199[29], net1199[30],
     net1199[31], net1199[32], net1199[33], net1199[34], net1199[35],
     net1199[36], net1199[37], net1199[38], net1199[39], net1199[40],
     net1199[41], net1199[42], net1199[43], net1199[44], net1199[45],
     net1199[46], net1199[47]}, {net1200[0], net1200[1], net1200[2],
     net1200[3], net1200[4], net1200[5], net1200[6], net1200[7],
     net1200[8], net1200[9], net1200[10], net1200[11], net1200[12],
     net1200[13], net1200[14], net1200[15], net1200[16], net1200[17],
     net1200[18], net1200[19], net1200[20], net1200[21], net1200[22],
     net1200[23], net1200[24], net1200[25], net1200[26], net1200[27],
     net1200[28], net1200[29], net1200[30], net1200[31], net1200[32],
     net1200[33], net1200[34], net1200[35], net1200[36], net1200[37],
     net1200[38], net1200[39], net1200[40], net1200[41], net1200[42],
     net1200[43], net1200[44], net1200[45], net1200[46], net1200[47]},
     {net1165[0], net1165[1], net1165[2], net1165[3], net1165[4],
     net1165[5], net1165[6], net1165[7], net1165[8], net1165[9],
     net1165[10], net1165[11], net1165[12], net1165[13], net1165[14],
     net1165[15], net1165[16], net1165[17], net1165[18], net1165[19],
     net1165[20], net1165[21], net1165[22], net1165[23], net1165[24],
     net1165[25], net1165[26], net1165[27], net1165[28], net1165[29],
     net1165[30], net1165[31], net1165[32], net1165[33], net1165[34],
     net1165[35], net1165[36], net1165[37], net1165[38], net1165[39],
     net1165[40], net1165[41], net1165[42], net1165[43], net1165[44],
     net1165[45], net1165[46], net1165[47]}, {net1250[0], net1250[1],
     net1250[2], net1250[3], net1250[4], net1250[5], net1250[6],
     net1250[7], net1250[8], net1250[9], net1250[10], net1250[11],
     net1250[12], net1250[13], net1250[14], net1250[15]}, {net1115[0],
     net1115[1], net1115[2], net1115[3], net1115[4], net1115[5],
     net1115[6], net1115[7], net1115[8], net1115[9], net1115[10],
     net1115[11], net1115[12], net1115[13], net1115[14], net1115[15],
     net1115[16], net1115[17], net1115[18], net1115[19], net1115[20],
     net1115[21], net1115[22], net1115[23], net1115[24], net1115[25],
     net1115[26], net1115[27], net1115[28], net1115[29], net1115[30],
     net1115[31], net1115[32], net1115[33], net1115[34], net1115[35],
     net1115[36], net1115[37], net1115[38], net1115[39], net1115[40],
     net1115[41], net1115[42], net1115[43], net1115[44], net1115[45],
     net1115[46], net1115[47]}, {net1216[0], net1216[1], net1216[2],
     net1216[3], net1216[4], net1216[5], net1216[6], net1216[7],
     net1216[8], net1216[9], net1216[10], net1216[11], net1216[12],
     net1216[13], net1216[14], net1216[15], net1216[16], net1216[17],
     net1216[18], net1216[19], net1216[20], net1216[21], net1216[22],
     net1216[23], net1216[24], net1216[25], net1216[26], net1216[27],
     net1216[28], net1216[29], net1216[30], net1216[31], net1216[32],
     net1216[33], net1216[34], net1216[35], net1216[36], net1216[37],
     net1216[38], net1216[39], net1216[40], net1216[41], net1216[42],
     net1216[43], net1216[44], net1216[45], net1216[46], net1216[47]},
     {net1215[0], net1215[1], net1215[2], net1215[3], net1215[4],
     net1215[5], net1215[6], net1215[7], net1215[8], net1215[9],
     net1215[10], net1215[11], net1215[12], net1215[13], net1215[14],
     net1215[15], net1215[16], net1215[17], net1215[18], net1215[19],
     net1215[20], net1215[21], net1215[22], net1215[23], net1215[24],
     net1215[25], net1215[26], net1215[27], net1215[28], net1215[29],
     net1215[30], net1215[31], net1215[32], net1215[33], net1215[34],
     net1215[35], net1215[36], net1215[37], net1215[38], net1215[39],
     net1215[40], net1215[41], net1215[42], net1215[43], net1215[44],
     net1215[45], net1215[46], net1215[47]}, {net1214[0], net1214[1],
     net1214[2], net1214[3], net1214[4], net1214[5], net1214[6],
     net1214[7], net1214[8], net1214[9], net1214[10], net1214[11],
     net1214[12], net1214[13], net1214[14], net1214[15], net1214[16],
     net1214[17], net1214[18], net1214[19], net1214[20], net1214[21],
     net1214[22], net1214[23], net1214[24], net1214[25], net1214[26],
     net1214[27], net1214[28], net1214[29], net1214[30], net1214[31],
     net1214[32], net1214[33], net1214[34], net1214[35], net1214[36],
     net1214[37], net1214[38], net1214[39], net1214[40], net1214[41],
     net1214[42], net1214[43], net1214[44], net1214[45], net1214[46],
     net1214[47]}, {net1213[0], net1213[1], net1213[2], net1213[3],
     net1213[4], net1213[5], net1213[6], net1213[7], net1213[8],
     net1213[9], net1213[10], net1213[11], net1213[12], net1213[13],
     net1213[14], net1213[15], net1213[16], net1213[17], net1213[18],
     net1213[19], net1213[20], net1213[21], net1213[22], net1213[23],
     net1213[24], net1213[25], net1213[26], net1213[27], net1213[28],
     net1213[29], net1213[30], net1213[31], net1213[32], net1213[33],
     net1213[34], net1213[35], net1213[36], net1213[37], net1213[38],
     net1213[39], net1213[40], net1213[41], net1213[42], net1213[43],
     net1213[44], net1213[45], net1213[46], net1213[47]}, {net1212[0],
     net1212[1], net1212[2], net1212[3], net1212[4], net1212[5],
     net1212[6], net1212[7], net1212[8], net1212[9], net1212[10],
     net1212[11], net1212[12], net1212[13], net1212[14], net1212[15],
     net1212[16], net1212[17], net1212[18], net1212[19], net1212[20],
     net1212[21], net1212[22], net1212[23], net1212[24], net1212[25],
     net1212[26], net1212[27], net1212[28], net1212[29], net1212[30],
     net1212[31], net1212[32], net1212[33], net1212[34], net1212[35],
     net1212[36], net1212[37], net1212[38], net1212[39], net1212[40],
     net1212[41], net1212[42], net1212[43], net1212[44], net1212[45],
     net1212[46], net1212[47]}, {net1209[0], net1209[1], net1209[2],
     net1209[3], net1209[4], net1209[5], net1209[6], net1209[7],
     net1209[8], net1209[9], net1209[10], net1209[11], net1209[12],
     net1209[13], net1209[14], net1209[15], net1209[16], net1209[17],
     net1209[18], net1209[19], net1209[20], net1209[21], net1209[22],
     net1209[23]}, {net1208[0], net1208[1], net1208[2], net1208[3],
     net1208[4], net1208[5], net1208[6], net1208[7], net1208[8],
     net1208[9], net1208[10], net1208[11], net1208[12], net1208[13],
     net1208[14], net1208[15], net1208[16], net1208[17], net1208[18],
     net1208[19], net1208[20], net1208[21], net1208[22], net1208[23]},
     {net1207[0], net1207[1], net1207[2], net1207[3], net1207[4],
     net1207[5], net1207[6], net1207[7], net1207[8], net1207[9],
     net1207[10], net1207[11], net1207[12], net1207[13], net1207[14],
     net1207[15], net1207[16], net1207[17], net1207[18], net1207[19],
     net1207[20], net1207[21], net1207[22], net1207[23]}, {net1206[0],
     net1206[1], net1206[2], net1206[3], net1206[4], net1206[5],
     net1206[6], net1206[7], net1206[8], net1206[9], net1206[10],
     net1206[11], net1206[12], net1206[13], net1206[14], net1206[15],
     net1206[16], net1206[17], net1206[18], net1206[19], net1206[20],
     net1206[21], net1206[22], net1206[23]}, {net1205[0], net1205[1],
     net1205[2], net1205[3], net1205[4], net1205[5], net1205[6],
     net1205[7], net1205[8], net1205[9], net1205[10], net1205[11],
     net1205[12], net1205[13], net1205[14], net1205[15], net1205[16],
     net1205[17], net1205[18], net1205[19], net1205[20], net1205[21],
     net1205[22], net1205[23]}, {net1198[0], net1198[1], net1198[2],
     net1198[3], net1198[4], net1198[5], net1198[6], net1198[7],
     net1198[8], net1198[9], net1198[10], net1198[11], net1198[12],
     net1198[13], net1198[14], net1198[15], net1198[16], net1198[17],
     net1198[18], net1198[19], net1198[20], net1198[21], net1198[22],
     net1198[23]}, {net1197[0], net1197[1], net1197[2], net1197[3],
     net1197[4], net1197[5], net1197[6], net1197[7], net1197[8],
     net1197[9], net1197[10], net1197[11], net1197[12], net1197[13],
     net1197[14], net1197[15], net1197[16], net1197[17], net1197[18],
     net1197[19], net1197[20], net1197[21], net1197[22], net1197[23]},
     {net1222[0], net1222[1], net1222[2], net1222[3], net1222[4],
     net1222[5], net1222[6], net1222[7], net1222[8], net1222[9],
     net1222[10], net1222[11], net1222[12], net1222[13], net1222[14],
     net1222[15], net1222[16], net1222[17], net1222[18], net1222[19],
     net1222[20], net1222[21], net1222[22], net1222[23]}, {net1103[0],
     net1103[1], net1103[2], net1103[3], net1103[4], net1103[5],
     net1103[6], net1103[7], net1103[8], net1103[9], net1103[10],
     net1103[11], net1103[12], net1103[13], net1103[14], net1103[15],
     net1103[16], net1103[17], net1103[18], net1103[19], net1103[20],
     net1103[21], net1103[22], net1103[23]}, {net1171[0], net1171[1],
     net1171[2], net1171[3], net1171[4], net1171[5], net1171[6],
     net1171[7], net1171[8], net1171[9], net1171[10], net1171[11],
     net1171[12], net1171[13], net1171[14], net1171[15], net1171[16],
     net1171[17], net1171[18], net1171[19], net1171[20], net1171[21],
     net1171[22], net1171[23]}, {net1231[0], net1231[1], net1231[2],
     net1231[3], net1231[4], net1231[5], net1231[6], net1231[7],
     net1231[8], net1231[9], net1231[10], net1231[11], net1231[12],
     net1231[13], net1231[14], net1231[15], net1231[16], net1231[17],
     net1231[18], net1231[19], net1231[20], net1231[21], net1231[22],
     net1231[23]}, {net1196[0], net1196[1], net1196[2], net1196[3],
     net1196[4], net1196[5], net1196[6], net1196[7], net1196[8],
     net1196[9], net1196[10], net1196[11], net1196[12], net1196[13],
     net1196[14], net1196[15], net1196[16], net1196[17], net1196[18],
     net1196[19], net1196[20], net1196[21], net1196[22], net1196[23]},
     {net1170[0], net1170[1], net1170[2], net1170[3], net1170[4],
     net1170[5], net1170[6], net1170[7], net1170[8], net1170[9],
     net1170[10], net1170[11], net1170[12], net1170[13], net1170[14],
     net1170[15], net1170[16], net1170[17], net1170[18], net1170[19],
     net1170[20], net1170[21], net1170[22], net1170[23]}, {net1195[0],
     net1195[1], net1195[2], net1195[3], net1195[4], net1195[5],
     net1195[6], net1195[7], net1195[8], net1195[9], net1195[10],
     net1195[11], net1195[12], net1195[13], net1195[14], net1195[15],
     net1195[16], net1195[17], net1195[18], net1195[19], net1195[20],
     net1195[21], net1195[22], net1195[23]}, vdd_cntl_l[143:0],
     wl_l[143:0], {net1138[0], net1138[1], net1138[2], net1138[3],
     net1138[4], net1138[5], net1138[6], net1138[7], net1138[8],
     net1138[9], net1138[10]}, {net1232[0], net1232[1], net1232[2],
     net1232[3], net1232[4], net1232[5], net1232[6], net1232[7],
     net1232[8], net1232[9], net1232[10]}, net1151, net1150,
     {net1149[0], net1149[1], net1149[2], net1149[3], net1149[4],
     net1149[5], net1149[6], net1149[7]}, bm_sck_b0_i, {net1147[0],
     net1147[1]}, {net1146[0], net1146[1]}, {bm_sdo_b1_o_0,
     bm_sdi_b0_o[0]}, net1144, {net1143[0], net1143[1]}, net1142,
     slf_op_07_00[3:0], net1140, net1139, gclk[7:0], net1136,
     fabric_out_05_00_bicegate, fabric_out_00_07_licegate,
     jtag_rowtest_mode_rowu0_b, last_rsr[0], net1135, padin_b[10:0],
     padin_b[12], padin_l[11:0], pll_lock_out, prog, purst, net1132,
     slf_op_07_01[7:0], slf_op_07_02[7:0], slf_op_07_03[7:0],
     slf_op_07_04[7:0], slf_op_07_05[7:0], slf_op_07_06[7:0],
     slf_op_07_07[7:0], slf_op_07_08[7:0], sdio_ml, net1124, tclkio_ml,
     {slf_op_00_09[3], slf_op_00_09[2], slf_op_00_09[1],
     slf_op_00_09[0], slf_op_00_09[3], slf_op_00_09[2],
     slf_op_00_09[1], slf_op_00_09[0]}, slf_op_01_09[7:0],
     slf_op_02_09[7:0], slf_op_03_09[7:0], slf_op_04_09[7:0],
     slf_op_05_09[7:0], slf_op_01_09[7:0], slf_op_02_09[7:0],
     slf_op_03_09[7:0], slf_op_04_09[7:0], slf_op_05_09[7:0],
     slf_op_06_09[7:0], slf_op_07_09[7:0], slf_op_01_09[7:0],
     slf_op_02_09[7:0], slf_op_03_09[7:0], slf_op_04_09[7:0],
     slf_op_05_09[7:0], slf_op_06_09[7:0], net1102);
bram_bank_logic_bot I21 ( .bm_sdo_i({bm_sdo_b2_o[1], bm_sdo_b2_o_0}),
     .bm_sclk_i(bm_bank30_sclk_o[1]), .bm_sclkrw_i(bm_bank30_sclkrw_o),
     .bm_sweb_i(bm_bank30_sweb_o), .bm_sdo_o(bm_bank30_sdo_i[3:2]),
     .bm_sweb_o({net948[0], net948[1]}), .bm_sclkrw_o({net952[0],
     net952[1]}), .bm_banksel_i(bm_bank30_banksel_o[3:2]));
bram_bank_logic_bot I63 ( .bm_sdo_i({bm_sdo_b0_o[1], bm_sdo_b0_o_0}),
     .bm_sclk_i(bm_sck_b0_i), .bm_sclkrw_i(net1273),
     .bm_sweb_i(net1274), .bm_sdo_o({net1275[0], net1275[1]}),
     .bm_sweb_o({net1143[0], net1143[1]}), .bm_sclkrw_o({net1147[0],
     net1147[1]}), .bm_banksel_i(bm_bank10_banksel_o[1:0]));
bram_hbuffer_dff_2xbank I_bram_buf1 ( .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_banksel_o(bm_bank30_banksel_o[3:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sweb_o(bm_bank30_sweb_o), .bm_sreb_o(bm_bank30_sreb_o),
     .bm_sclk_o(bm_bank30_sclk_o[1:0]), .bm_sa_o(bm_bank30_sa_o[7:0]),
     .bm_init_o(bm_bank30_init_o), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclkrw_o(bm_bank30_sclkrw_o), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sdo_o(bm_sdo_o[3:0]), .bm_sdi_o(bm_bank30_sdi_o[3:0]),
     .bm_rcapmux_en_o(bm_bank30_rcapmux_en_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_banksel_i(bm_banksel_i[3:0]),
     .bm_sdo_i(bm_bank30_sdo_i[3:0]));
bram_hbuffer_1xbank I2 ( .bm_sa_o({net1149[0], net1149[1], net1149[2],
     net1149[3], net1149[4], net1149[5], net1149[6], net1149[7]}),
     .bm_wdummymux_en_o(net1142), .bm_sweb_i(bm_bank30_sweb_o),
     .bm_sreb_i(bm_bank30_sreb_o), .bm_sdi_i(bm_bank30_sdi_o[1:0]),
     .bm_sclk_i(bm_bank30_sclk_o[0]), .bm_init_i(bm_bank30_init_o),
     .bm_banksel_o(bm_bank10_banksel_o[1:0]),
     .bm_rcapmux_en_i(bm_bank30_rcapmux_en_o),
     .bm_wdummymux_en_i(bm_wdummymux_en_o), .bm_sweb_o(net1274),
     .bm_sreb_o(net1144), .bm_sdi_o({net1146[0], net1146[1]}),
     .bm_sclk_o(bm_sck_b0_i), .bm_init_o(net1151),
     .bm_sa_i(bm_bank30_sa_o[7:0]), .bm_rcapmux_en_o(net1150),
     .bm_sclkrw_i(bm_bank30_sclkrw_o), .bm_sclkrw_o(net1273),
     .bm_sdo_i({net1275[0], net1275[1]}),
     .bm_banksel_i(bm_bank30_banksel_o[1:0]),
     .bm_sdo_o(bm_bank30_sdo_i[1:0]));

endmodule
// Library - leafcell, Cell - clkmux4to1, View - schematic
// LAST TIME SAVED: Jun 30 10:55:11 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module clkmux4to1 ( mout, cbit, .cdsNet0(min[0]), .cdsNet0(min[1]),
     .cdsNet0(min[2]), .cdsNet0(min[3]) );
output  mout;


input [3:0]  min;
input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cbit_b;



txgate_hvt I4 ( .in(net_2_0), .out(net52), .pp(cbit[1]),
     .nn(cbit_b[1]));
txgate_hvt I3 ( .in(net_2_1), .out(net52), .pp(cbit_b[1]),
     .nn(cbit[1]));
txgate_hvt I6 ( .in(min[2]), .out(net_2_1), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I5 ( .in(min[3]), .out(net_2_1), .pp(cbit_b[0]),
     .nn(cbit[0]));
txgate_hvt Itg20 ( .in(min[0]), .out(net_2_0), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I7 ( .in(min[1]), .out(net_2_0), .pp(cbit_b[0]),
     .nn(cbit[0]));
inv_hvt I2 ( .A(net046), .Y(mout));
inv_hvt I1_1_ ( .A(cbit[1]), .Y(cbit_b[1]));
inv_hvt I1_0_ ( .A(cbit[0]), .Y(cbit_b[0]));
inv_hvt I0 ( .A(net52), .Y(net046));

endmodule
// Library - sbtlibn65lp, Cell - vddp_tiehigh, View - schematic
// LAST TIME SAVED: Jun 21 10:52:52 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module vddp_tiehigh ( vddp_tieh );
inout  vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M8 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net9), .S(vddp_));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_rows, View - schematic
// LAST TIME SAVED: Jul 27 16:24:09 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module ml_testdec_rows ( dec_bias, dec_det, vddp_tieh, wp, wr );
inout  dec_bias, dec_det;

input  vddp_tieh, wp, wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M8 ( .D(dec_det), .B(GND_), .G(wr), .S(gnd_));
nch  M6 ( .D(dec_det), .B(GND_), .G(net20), .S(gnd_));
nch  M5 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(net20));
nch  M7 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(wr));
nch_25  M12 ( .D(net20), .B(gnd_), .G(vddp_tieh), .S(wp));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_rowsx108_1f, View - schematic
// LAST TIME SAVED: Dec 23 16:24:55 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module ml_testdec_rowsx108_1f ( dec_det_buf, dec_bias, dec_det, wp, wr
     );
output  dec_det_buf;

inout  dec_bias, dec_det;


input [107:0]  wr;
input [107:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(dec_det), .Y(net25));
inv_hvt I27 ( .A(net25), .Y(dec_det_buf));
vddp_tiehigh I25 ( .vddp_tieh(vddp_tiel));
ml_testdec_rows Itestdec_rows_107_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[107]), .wp(wp[107]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_106_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[106]), .wp(wp[106]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_105_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[105]), .wp(wp[105]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_104_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[104]), .wp(wp[104]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_103_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[103]), .wp(wp[103]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_102_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[102]), .wp(wp[102]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_101_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[101]), .wp(wp[101]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_100_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[100]), .wp(wp[100]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_99_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[99]), .wp(wp[99]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_98_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[98]), .wp(wp[98]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_97_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[97]), .wp(wp[97]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_96_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[96]), .wp(wp[96]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_95_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[95]), .wp(wp[95]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_94_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[94]), .wp(wp[94]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_93_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[93]), .wp(wp[93]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_92_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[92]), .wp(wp[92]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_91_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[91]), .wp(wp[91]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_90_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[90]), .wp(wp[90]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_89_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[89]), .wp(wp[89]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_88_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[88]), .wp(wp[88]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_87_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[87]), .wp(wp[87]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_86_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[86]), .wp(wp[86]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_85_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[85]), .wp(wp[85]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_84_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[84]), .wp(wp[84]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_83_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[83]), .wp(wp[83]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_82_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[82]), .wp(wp[82]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_81_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[81]), .wp(wp[81]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_80_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[80]), .wp(wp[80]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_79_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[79]), .wp(wp[79]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_78_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[78]), .wp(wp[78]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_77_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[77]), .wp(wp[77]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_76_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[76]), .wp(wp[76]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_75_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[75]), .wp(wp[75]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_74_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[74]), .wp(wp[74]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_73_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[73]), .wp(wp[73]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_72_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[72]), .wp(wp[72]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_71_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[71]), .wp(wp[71]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_70_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[70]), .wp(wp[70]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_69_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[69]), .wp(wp[69]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_68_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[68]), .wp(wp[68]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_67_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[67]), .wp(wp[67]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_66_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[66]), .wp(wp[66]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_65_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[65]), .wp(wp[65]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_64_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[64]), .wp(wp[64]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_63_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[63]), .wp(wp[63]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_62_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[62]), .wp(wp[62]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_61_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[61]), .wp(wp[61]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_60_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[60]), .wp(wp[60]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_59_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[59]), .wp(wp[59]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_58_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[58]), .wp(wp[58]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_57_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[57]), .wp(wp[57]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_56_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[56]), .wp(wp[56]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_55_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[55]), .wp(wp[55]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_54_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[54]), .wp(wp[54]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_53_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[53]), .wp(wp[53]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_52_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[52]), .wp(wp[52]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_51_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[51]), .wp(wp[51]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_50_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[50]), .wp(wp[50]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_49_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[49]), .wp(wp[49]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_48_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[48]), .wp(wp[48]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_47_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[47]), .wp(wp[47]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_46_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[46]), .wp(wp[46]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_45_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[45]), .wp(wp[45]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_44_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[44]), .wp(wp[44]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_43_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[43]), .wp(wp[43]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_42_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[42]), .wp(wp[42]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_41_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[41]), .wp(wp[41]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_40_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[40]), .wp(wp[40]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_39_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[39]), .wp(wp[39]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_38_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[38]), .wp(wp[38]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_37_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[37]), .wp(wp[37]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_36_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[36]), .wp(wp[36]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_35_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[35]), .wp(wp[35]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_34_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[34]), .wp(wp[34]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_33_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[33]), .wp(wp[33]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_32_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[32]), .wp(wp[32]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_31_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[31]), .wp(wp[31]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_30_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[30]), .wp(wp[30]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_29_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[29]), .wp(wp[29]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_28_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[28]), .wp(wp[28]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_27_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[27]), .wp(wp[27]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_26_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[26]), .wp(wp[26]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_25_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[25]), .wp(wp[25]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_24_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[24]), .wp(wp[24]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_23_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[23]), .wp(wp[23]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_22_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[22]), .wp(wp[22]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_21_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[21]), .wp(wp[21]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_20_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[20]), .wp(wp[20]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_19_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[19]), .wp(wp[19]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_18_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[18]), .wp(wp[18]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_17_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[17]), .wp(wp[17]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_16_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[16]), .wp(wp[16]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_15_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[15]), .wp(wp[15]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_14_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[14]), .wp(wp[14]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_13_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[13]), .wp(wp[13]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_12_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[12]), .wp(wp[12]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_11_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[11]), .wp(wp[11]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_10_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[10]), .wp(wp[10]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_9_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[9]), .wp(wp[9]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_8_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[8]), .wp(wp[8]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_7_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[7]), .wp(wp[7]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_6_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[6]), .wp(wp[6]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_5_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[5]), .wp(wp[5]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_4_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[4]), .wp(wp[4]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_3_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[3]), .wp(wp[3]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_2_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[2]), .wp(wp[2]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_1_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[1]), .wp(wp[1]),
     .dec_bias(dec_bias));
ml_testdec_rows Itestdec_rows_0_ ( .dec_det(dec_det),
     .vddp_tieh(vddp_tiel), .wr(wr[0]), .wp(wp[0]),
     .dec_bias(dec_bias));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd2vdd25, View - schematic
// LAST TIME SAVED: Jun 11 16:25:15 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
nch_25  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));
pch_25  M0 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
pch_25  M1 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
pch_25  M2 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
pch_25  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));

endmodule
// Library - tsmcN40, Cell - nor2_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:25 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nor2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  M2 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  M1 ( .D(net15), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(net15));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_columns, View - schematic
// LAST TIME SAVED: Jun 24 12:15:49 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module ml_testdec_columns ( bl, vdd_drv, dec_det_even_25,
     dec_det_odd_25 );
inout  vdd_drv;

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(vdd_drv), .B(gnd_), .G(dec_det_even_25), .S(bl[0]));
nch_25  M4 ( .D(vdd_drv), .B(gnd_), .G(dec_det_odd_25), .S(bl[1]));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_columnsx330_1f, View -
//schematic
// LAST TIME SAVED: Dec 28 17:38:01 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module ml_testdec_columnsx330_1f ( bl, bl_dummyl, bl_dummyr, bl_test,
     dec_det_buf, testdec_even_b_25, testdec_odd_b_25 );

input  dec_det_buf, testdec_even_b_25, testdec_odd_b_25;

inout [327:0]  bl;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I134 ( .A(dec_det_buf), .Y(net40));
inv_hvt I55 ( .A(net40), .Y(net36));
ml_ls_vdd2vdd25 I144 ( .in(net36), .sup(vddp_), .out_vddio_b(net38),
     .out_vddio(dec_det_25), .in_b(net40));
nor2_25 I26 ( .A(testdec_odd_b_25), .Y(dec_det_odd_25), .Gb(GND_),
     .G(GND_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
nor2_25 I59 ( .A(testdec_even_b_25), .Y(dec_det_even_25), .Gb(GND_),
     .G(GND_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
rppolywo  R1 ( .MINUS(vdd_drv), .PLUS(vdd_));
rppolywo  R2 ( .MINUS(vdd_drv), .PLUS(vdd_));
rppolywo  R3 ( .MINUS(vdd_drv), .PLUS(vdd_));
rppolywo  R0 ( .MINUS(vdd_drv), .PLUS(vdd_));
ml_testdec_columns Itestdec_columns_dml ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyl[1:0]));
ml_testdec_columns Itestdec_columns_163_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[327:326]));
ml_testdec_columns Itestdec_columns_162_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[325:324]));
ml_testdec_columns Itestdec_columns_161_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[323:322]));
ml_testdec_columns Itestdec_columns_160_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[321:320]));
ml_testdec_columns Itestdec_columns_159_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[319:318]));
ml_testdec_columns Itestdec_columns_158_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[317:316]));
ml_testdec_columns Itestdec_columns_157_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[315:314]));
ml_testdec_columns Itestdec_columns_156_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[313:312]));
ml_testdec_columns Itestdec_columns_155_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[311:310]));
ml_testdec_columns Itestdec_columns_154_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[309:308]));
ml_testdec_columns Itestdec_columns_153_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[307:306]));
ml_testdec_columns Itestdec_columns_152_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[305:304]));
ml_testdec_columns Itestdec_columns_151_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[303:302]));
ml_testdec_columns Itestdec_columns_150_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[301:300]));
ml_testdec_columns Itestdec_columns_149_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[299:298]));
ml_testdec_columns Itestdec_columns_148_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[297:296]));
ml_testdec_columns Itestdec_columns_147_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[295:294]));
ml_testdec_columns Itestdec_columns_146_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[293:292]));
ml_testdec_columns Itestdec_columns_145_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[291:290]));
ml_testdec_columns Itestdec_columns_144_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[289:288]));
ml_testdec_columns Itestdec_columns_143_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[287:286]));
ml_testdec_columns Itestdec_columns_142_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[285:284]));
ml_testdec_columns Itestdec_columns_141_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[283:282]));
ml_testdec_columns Itestdec_columns_140_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[281:280]));
ml_testdec_columns Itestdec_columns_139_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[279:278]));
ml_testdec_columns Itestdec_columns_138_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[277:276]));
ml_testdec_columns Itestdec_columns_137_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[275:274]));
ml_testdec_columns Itestdec_columns_136_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[273:272]));
ml_testdec_columns Itestdec_columns_135_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[271:270]));
ml_testdec_columns Itestdec_columns_134_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[269:268]));
ml_testdec_columns Itestdec_columns_133_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[267:266]));
ml_testdec_columns Itestdec_columns_132_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[265:264]));
ml_testdec_columns Itestdec_columns_131_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[263:262]));
ml_testdec_columns Itestdec_columns_130_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[261:260]));
ml_testdec_columns Itestdec_columns_129_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[259:258]));
ml_testdec_columns Itestdec_columns_128_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[257:256]));
ml_testdec_columns Itestdec_columns_127_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[255:254]));
ml_testdec_columns Itestdec_columns_126_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[253:252]));
ml_testdec_columns Itestdec_columns_125_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[251:250]));
ml_testdec_columns Itestdec_columns_124_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[249:248]));
ml_testdec_columns Itestdec_columns_123_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[247:246]));
ml_testdec_columns Itestdec_columns_122_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[245:244]));
ml_testdec_columns Itestdec_columns_121_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[243:242]));
ml_testdec_columns Itestdec_columns_120_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[241:240]));
ml_testdec_columns Itestdec_columns_119_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[239:238]));
ml_testdec_columns Itestdec_columns_118_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[237:236]));
ml_testdec_columns Itestdec_columns_117_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[235:234]));
ml_testdec_columns Itestdec_columns_116_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[233:232]));
ml_testdec_columns Itestdec_columns_115_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[231:230]));
ml_testdec_columns Itestdec_columns_114_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[229:228]));
ml_testdec_columns Itestdec_columns_113_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[227:226]));
ml_testdec_columns Itestdec_columns_112_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[225:224]));
ml_testdec_columns Itestdec_columns_111_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[223:222]));
ml_testdec_columns Itestdec_columns_110_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[221:220]));
ml_testdec_columns Itestdec_columns_109_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[219:218]));
ml_testdec_columns Itestdec_columns_108_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[217:216]));
ml_testdec_columns Itestdec_columns_107_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[215:214]));
ml_testdec_columns Itestdec_columns_106_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[213:212]));
ml_testdec_columns Itestdec_columns_105_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[211:210]));
ml_testdec_columns Itestdec_columns_104_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[209:208]));
ml_testdec_columns Itestdec_columns_103_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[207:206]));
ml_testdec_columns Itestdec_columns_102_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[205:204]));
ml_testdec_columns Itestdec_columns_101_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[203:202]));
ml_testdec_columns Itestdec_columns_100_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[201:200]));
ml_testdec_columns Itestdec_columns_99_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[199:198]));
ml_testdec_columns Itestdec_columns_98_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[197:196]));
ml_testdec_columns Itestdec_columns_97_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[195:194]));
ml_testdec_columns Itestdec_columns_96_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[193:192]));
ml_testdec_columns Itestdec_columns_95_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[191:190]));
ml_testdec_columns Itestdec_columns_94_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[189:188]));
ml_testdec_columns Itestdec_columns_93_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[187:186]));
ml_testdec_columns Itestdec_columns_92_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[185:184]));
ml_testdec_columns Itestdec_columns_91_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[183:182]));
ml_testdec_columns Itestdec_columns_90_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[181:180]));
ml_testdec_columns Itestdec_columns_89_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[179:178]));
ml_testdec_columns Itestdec_columns_88_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[177:176]));
ml_testdec_columns Itestdec_columns_87_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[175:174]));
ml_testdec_columns Itestdec_columns_86_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[173:172]));
ml_testdec_columns Itestdec_columns_85_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[171:170]));
ml_testdec_columns Itestdec_columns_84_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[169:168]));
ml_testdec_columns Itestdec_columns_83_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[167:166]));
ml_testdec_columns Itestdec_columns_82_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[165:164]));
ml_testdec_columns Itestdec_columns_81_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[163:162]));
ml_testdec_columns Itestdec_columns_80_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[161:160]));
ml_testdec_columns Itestdec_columns_79_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[159:158]));
ml_testdec_columns Itestdec_columns_78_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[157:156]));
ml_testdec_columns Itestdec_columns_77_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[155:154]));
ml_testdec_columns Itestdec_columns_76_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[153:152]));
ml_testdec_columns Itestdec_columns_75_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[151:150]));
ml_testdec_columns Itestdec_columns_74_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[149:148]));
ml_testdec_columns Itestdec_columns_73_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[147:146]));
ml_testdec_columns Itestdec_columns_72_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[145:144]));
ml_testdec_columns Itestdec_columns_71_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[143:142]));
ml_testdec_columns Itestdec_columns_70_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[141:140]));
ml_testdec_columns Itestdec_columns_69_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[139:138]));
ml_testdec_columns Itestdec_columns_68_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[137:136]));
ml_testdec_columns Itestdec_columns_67_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[135:134]));
ml_testdec_columns Itestdec_columns_66_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[133:132]));
ml_testdec_columns Itestdec_columns_65_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[131:130]));
ml_testdec_columns Itestdec_columns_64_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[129:128]));
ml_testdec_columns Itestdec_columns_63_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[127:126]));
ml_testdec_columns Itestdec_columns_62_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[125:124]));
ml_testdec_columns Itestdec_columns_61_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[123:122]));
ml_testdec_columns Itestdec_columns_60_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[121:120]));
ml_testdec_columns Itestdec_columns_59_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[119:118]));
ml_testdec_columns Itestdec_columns_58_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[117:116]));
ml_testdec_columns Itestdec_columns_57_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[115:114]));
ml_testdec_columns Itestdec_columns_56_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[113:112]));
ml_testdec_columns Itestdec_columns_55_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[111:110]));
ml_testdec_columns Itestdec_columns_54_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[109:108]));
ml_testdec_columns Itestdec_columns_53_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[107:106]));
ml_testdec_columns Itestdec_columns_52_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[105:104]));
ml_testdec_columns Itestdec_columns_51_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[103:102]));
ml_testdec_columns Itestdec_columns_50_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[101:100]));
ml_testdec_columns Itestdec_columns_49_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[99:98]));
ml_testdec_columns Itestdec_columns_48_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[97:96]));
ml_testdec_columns Itestdec_columns_47_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[95:94]));
ml_testdec_columns Itestdec_columns_46_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[93:92]));
ml_testdec_columns Itestdec_columns_45_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[91:90]));
ml_testdec_columns Itestdec_columns_44_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[89:88]));
ml_testdec_columns Itestdec_columns_43_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[87:86]));
ml_testdec_columns Itestdec_columns_42_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[85:84]));
ml_testdec_columns Itestdec_columns_41_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[83:82]));
ml_testdec_columns Itestdec_columns_40_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[81:80]));
ml_testdec_columns Itestdec_columns_39_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[79:78]));
ml_testdec_columns Itestdec_columns_38_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[77:76]));
ml_testdec_columns Itestdec_columns_37_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[75:74]));
ml_testdec_columns Itestdec_columns_36_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[73:72]));
ml_testdec_columns Itestdec_columns_35_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[71:70]));
ml_testdec_columns Itestdec_columns_34_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[69:68]));
ml_testdec_columns Itestdec_columns_33_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[67:66]));
ml_testdec_columns Itestdec_columns_32_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[65:64]));
ml_testdec_columns Itestdec_columns_31_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[63:62]));
ml_testdec_columns Itestdec_columns_30_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[61:60]));
ml_testdec_columns Itestdec_columns_29_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[59:58]));
ml_testdec_columns Itestdec_columns_28_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[57:56]));
ml_testdec_columns Itestdec_columns_27_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[55:54]));
ml_testdec_columns Itestdec_columns_26_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[53:52]));
ml_testdec_columns Itestdec_columns_25_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[51:50]));
ml_testdec_columns Itestdec_columns_24_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[49:48]));
ml_testdec_columns Itestdec_columns_23_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[47:46]));
ml_testdec_columns Itestdec_columns_22_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[45:44]));
ml_testdec_columns Itestdec_columns_21_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[43:42]));
ml_testdec_columns Itestdec_columns_20_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[41:40]));
ml_testdec_columns Itestdec_columns_19_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[39:38]));
ml_testdec_columns Itestdec_columns_18_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[37:36]));
ml_testdec_columns Itestdec_columns_17_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[35:34]));
ml_testdec_columns Itestdec_columns_16_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[33:32]));
ml_testdec_columns Itestdec_columns_15_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[31:30]));
ml_testdec_columns Itestdec_columns_14_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[29:28]));
ml_testdec_columns Itestdec_columns_13_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[27:26]));
ml_testdec_columns Itestdec_columns_12_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[25:24]));
ml_testdec_columns Itestdec_columns_11_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[23:22]));
ml_testdec_columns Itestdec_columns_10_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[21:20]));
ml_testdec_columns Itestdec_columns_9_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[19:18]));
ml_testdec_columns Itestdec_columns_8_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[17:16]));
ml_testdec_columns Itestdec_columns_7_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[15:14]));
ml_testdec_columns Itestdec_columns_6_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[13:12]));
ml_testdec_columns Itestdec_columns_5_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[11:10]));
ml_testdec_columns Itestdec_columns_4_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[9:8]));
ml_testdec_columns Itestdec_columns_3_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[7:6]));
ml_testdec_columns Itestdec_columns_2_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[5:4]));
ml_testdec_columns Itestdec_columns_1_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[3:2]));
ml_testdec_columns Itestdec_columns_0_ ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[1:0]));
ml_testdec_columns Itestdec_columns_dmr ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyr[1:0]));
ml_testdec_columns Itestdec_columns_tst ( .vdd_drv(vdd_drv),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_test[1:0]));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tielow, View - schematic
// LAST TIME SAVED: Jul 20 11:25:32 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module vdd_tielow ( gnd_tiel );
inout  gnd_tiel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(gnd_tiel), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(net9), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - NVCM_40nm, Cell - cell_1x1, View - schematic
// LAST TIME SAVED: Oct 15 17:03:11 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module cell_1x1 ( bl, wp, wr );
inout  bl;

input  wp, wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nchx  WR_CELL ( .D(net08), .G(wr), .S(bl));
nchx  WP_CELL ( .D(net011), .G(wp), .S(net08));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x1, View - schematic
// LAST TIME SAVED: Jul 12 16:56:42 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nvcm_cell_2x1 ( bl, wp, wr );

input  wp, wr;

inout [1:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cell_1x1 I11 ( .wp(wp), .wr(wr), .bl(bl[0]));
cell_1x1 I12 ( .wp(wp), .wr(wr), .bl(bl[1]));

endmodule
// Library - leafcell, Cell - buffer500um, View - schematic
// LAST TIME SAVED: May 13 11:02:42 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module buffer500um ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_2x8, View - schematic
// LAST TIME SAVED: Feb 26 14:36:29 2008
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nvcm_cell_2x8 ( bl, wp, wr );


inout [1:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m7 ( .bl(bl[1:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_2x1 m6 ( .bl(bl[1:0]), .wr(wr[6]), .wp(wp[6]));
nvcm_cell_2x1 m5 ( .bl(bl[1:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_2x1 m4 ( .bl(bl[1:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_2x1 m3 ( .bl(bl[1:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_2x1 m2 ( .bl(bl[1:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_1x8, View - schematic
// LAST TIME SAVED: Jul  8 17:57:53 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nvcm_cell_1x8 ( bl, wp, wr );

input  wp, wr;

inout [7:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cell_1x1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
cell_1x1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));
cell_1x1 m2 ( .wp(wp), .wr(wr), .bl(bl[2]));
cell_1x1 m3 ( .wp(wp), .wr(wr), .bl(bl[3]));
cell_1x1 m4 ( .wp(wp), .wr(wr), .bl(bl[4]));
cell_1x1 m5 ( .wp(wp), .wr(wr), .bl(bl[5]));
cell_1x1 m6 ( .wp(wp), .wr(wr), .bl(bl[6]));
cell_1x1 m7 ( .wp(wp), .wr(wr), .bl(bl[7]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_8x8, View - schematic
// LAST TIME SAVED: Jun 24 17:57:01 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nvcm_cell_8x8 ( bl, wp, wr );


inout [7:0]  bl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 m0 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 m1 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 m2 ( .bl(bl[7:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_1x8 m3 ( .bl(bl[7:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_1x8 m7 ( .bl(bl[7:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_1x8 m4 ( .bl(bl[7:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_1x8 m5 ( .bl(bl[7:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_1x8 m6 ( .bl(bl[7:0]), .wr(wr[6]), .wp(wp[6]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_16x8, View - schematic
// LAST TIME SAVED: Jun 24 17:57:26 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nvcm_cell_16x8 ( bl, wp, wr );


inout [15:0]  bl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_8x8 m0 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[7:0]));
nvcm_cell_8x8 m1 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[15:8]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_336x8, View - schematic
// LAST TIME SAVED: Dec 30 14:06:16 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nvcm_cell_336x8 ( bl, bl_dummyl, bl_dummyr, bl_test, wp, wr );


inout [5:0]  bl_dummyr;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [327:0]  bl;

input [7:0]  wp;
input [7:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x8 Invcm_cell_2x8 ( .wp(wp[7:0]), .wr(wr[7:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_16x8 Invcm_cell_16x8_19_ ( .wp(wp[7:0]), .bl(bl[319:304]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_18_ ( .wp(wp[7:0]), .bl(bl[303:288]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_17_ ( .wp(wp[7:0]), .bl(bl[287:272]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_16_ ( .wp(wp[7:0]), .bl(bl[271:256]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_15_ ( .wp(wp[7:0]), .bl(bl[255:240]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_14_ ( .wp(wp[7:0]), .bl(bl[239:224]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_13_ ( .wp(wp[7:0]), .bl(bl[223:208]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_12_ ( .wp(wp[7:0]), .bl(bl[207:192]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_11_ ( .wp(wp[7:0]), .bl(bl[191:176]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_10_ ( .wp(wp[7:0]), .bl(bl[175:160]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_9_ ( .wp(wp[7:0]), .bl(bl[159:144]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_8_ ( .wp(wp[7:0]), .bl(bl[143:128]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_7_ ( .wp(wp[7:0]), .bl(bl[127:112]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_6_ ( .wp(wp[7:0]), .bl(bl[111:96]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_5_ ( .wp(wp[7:0]), .bl(bl[95:80]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_4_ ( .wp(wp[7:0]), .bl(bl[79:64]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_3_ ( .wp(wp[7:0]), .bl(bl[63:48]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_2_ ( .wp(wp[7:0]), .bl(bl[47:32]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_1_ ( .wp(wp[7:0]), .bl(bl[31:16]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_0_ ( .wp(wp[7:0]), .bl(bl[15:0]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_20_ ( .wp(wp[7:0]), .bl({bl_dummyr[5:0],
     bl_test[1:0], bl[327:320]}), .wr(wr[7:0]));

endmodule
// Library - NVCM_40nm, Cell - nvcm_cell_338x112_1f, View - schematic
// LAST TIME SAVED: Dec 28 17:18:26 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module nvcm_cell_338x112_1f ( bl, bl_dummyl, bl_dummyr, bl_test, wp,
     wp_dummyb, wp_dummyt, wr, wr_dummyb, wr_dummyt );


inout [1:0]  bl_dummyr;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [327:0]  bl;

input [1:0]  wp_dummyb;
input [1:0]  wr_dummyb;
input [1:0]  wr_dummyt;
input [107:0]  wp;
input [1:0]  wp_dummyt;
input [107:0]  wr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_336x8 Invcm_cell_336x8_11_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[101:94]), .wp(wp[101:94]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_10_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[93:86]), .wp(wp[93:86]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_9_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[85:78]), .wp(wp[85:78]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_8_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[77:70]), .wp(wp[77:70]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_7_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[69:62]), .wp(wp[69:62]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_6_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[61:54]), .wp(wp[61:54]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_5_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[53:46]), .wp(wp[53:46]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_4_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[45:38]), .wp(wp[45:38]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_3_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[37:30]), .wp(wp[37:30]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_2_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[29:22]), .wp(wp[29:22]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_1_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[21:14]), .wp(wp[21:14]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_0_ ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr(wr[13:6]), .wp(wp[13:6]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_t ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr({wr[5:0], wr_dummyt[1:0]}), .wp({wp[5:0], wp_dummyt[1:0]}),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8 Invcm_cell_336x8_b ( .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl(bl[327:0]), .bl_test(bl_test[1:0]),
     .wr({wr_dummyb[1:0], wr[107:102]}), .wp({wp_dummyb[1:0],
     wp[107:102]}), .bl_dummyl(bl_dummyl[1:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_testdec_bgen, View - schematic
// LAST TIME SAVED: Jul 15 18:50:47 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module ml_testdec_bgen ( dec_ok, dec_bias, dec_det, testdec_en_b,
     testdec_prec_b );
output  dec_ok;

inout  dec_bias, dec_det;

input  testdec_en_b, testdec_prec_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M4 ( .D(dec_det), .B(GND_), .G(testdec_en_b), .S(gnd_));
pch_hvt  M0 ( .D(dec_det), .B(vdd_), .G(testdec_prec_b), .S(vdd_));
inv_hvt I134 ( .A(dec_det), .Y(dec_ok));
nch  M13 ( .D(dec_bias), .B(GND_), .G(testdec_en_b), .S(gnd_));
nch  M6 ( .D(dec_bias), .B(GND_), .G(dec_bias), .S(gnd_));
nch  M7 ( .D(dec_bias_p), .B(GND_), .G(dec_bias), .S(gnd_));
nch  M14 ( .D(ngate), .B(GND_), .G(dec_bias), .S(gnd_));
nch  M15 ( .D(ngate), .B(GND_), .G(testdec_en_b), .S(gnd_));
nch  M10 ( .D(dec_bias_sup), .B(GND_), .G(ngate), .S(dec_bias));
pch  M19 ( .D(ngate), .B(vdd_), .G(testdec_en_b), .S(net76));
pch  M16 ( .D(net76), .B(vdd_), .G(testdec_en_b), .S(vdd_));
pch  M18_1_ ( .D(dec_bias_sup), .B(vdd_), .G(testdec_en_b), .S(vdd_));
pch  M18_0_ ( .D(dec_bias_sup), .B(vdd_), .G(testdec_en_b), .S(vdd_));
pch  M9_2_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));
pch  M9_1_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));
pch  M9_0_ ( .D(dec_det), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));
pch  M8 ( .D(dec_bias_p), .B(vdd_), .G(dec_bias_p), .S(dec_bias_sup));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_yp3_x8, View - schematic
// LAST TIME SAVED: Jul 13 16:32:00 2010
// NETLIST TIME: May  5 11:56:44 2011
`timescale 1ns / 1ns 

module ml_ymux_yp3_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M17 ( .D(bl[5]), .B(GND_), .G(yp3_25[5]), .S(bl_out));
nch_25  M16 ( .D(bl[6]), .B(GND_), .G(yp3_25[6]), .S(bl_out));
nch_25  M18 ( .D(bl[4]), .B(GND_), .G(yp3_25[4]), .S(bl_out));
nch_25  M19 ( .D(bl[3]), .B(GND_), .G(yp3_25[3]), .S(bl_out));
nch_25  M26 ( .D(bl[0]), .B(GND_), .G(yp3_b_25[0]), .S(vblinhi_rde));
nch_25  M0 ( .D(bl[1]), .B(GND_), .G(yp3_b_25[1]), .S(vblinhi_rdo));
nch_25  M3 ( .D(bl[3]), .B(GND_), .G(yp3_b_25[3]), .S(vblinhi_rdo));
nch_25  M2 ( .D(bl[2]), .B(GND_), .G(yp3_b_25[2]), .S(vblinhi_rde));
nch_25  M4 ( .D(bl[4]), .B(GND_), .G(yp3_b_25[4]), .S(vblinhi_rde));
nch_25  M6 ( .D(bl[5]), .B(GND_), .G(yp3_b_25[5]), .S(vblinhi_rdo));
nch_25  M22 ( .D(bl[0]), .B(GND_), .G(yp3_25[0]), .S(bl_out));
nch_25  M20 ( .D(bl[2]), .B(GND_), .G(yp3_25[2]), .S(bl_out));
nch_25  M21 ( .D(bl[1]), .B(GND_), .G(yp3_25[1]), .S(bl_out));
nch_25  M8 ( .D(bl[7]), .B(GND_), .G(yp3_b_25[7]), .S(vblinhi_rdo));
nch_25  M15 ( .D(bl[7]), .B(GND_), .G(yp3_25[7]), .S(bl_out));
nch_25  M7 ( .D(bl[6]), .B(GND_), .G(yp3_b_25[6]), .S(vblinhi_rde));
pch_25  M5_7_ ( .D(bl[7]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_6_ ( .D(bl[6]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_5_ ( .D(bl[5]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_4_ ( .D(bl[4]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_3_ ( .D(bl[3]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_2_ ( .D(bl[2]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_1_ ( .D(bl[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_0_ ( .D(bl[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x8, View - schematic
// LAST TIME SAVED: May  4 13:03:21 2008
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_dummy, View - schematic
// LAST TIME SAVED: Jun 23 14:12:41 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_dummy ( bl_dummyr, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, pgminhi_dmmy_b_25, vdd_tieh );
inout  vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo;

input  pgminhi_dmmy_b_25, vdd_tieh;

inout [1:0]  bl_dummyr;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(bl_dummyr[1]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rdo));
nch_25  M2 ( .D(bl_dummyr[0]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rde));
pch_25  M8 ( .D(bl_dummyr[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M0 ( .D(bl_dummyr[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));

endmodule
// Library - leafcell, Cell - cfg4pllreset, View - schematic
// LAST TIME SAVED: Jul  7 08:09:12 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module cfg4pllreset ( out, in, prog );
output  out;

input  in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2 I1 ( .A(net012), .B(prog), .Y(net8));
inv I2 ( .A(in), .Y(net012));
inv I3 ( .A(net8), .Y(out));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_yp2_8, View - schematic
// LAST TIME SAVED: Jun 23 14:36:38 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_yp2_8 ( bl, bl_out, vblinhi_rde, vblinhi_rdo, yp2,
     yp2_b_25 );
inout  bl_out, vblinhi_rde, vblinhi_rdo;


inout [7:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M6 ( .D(bl[6]), .B(GND_), .G(yp2[6]), .S(bl_out));
nch_hvt  M7 ( .D(bl[7]), .B(GND_), .G(yp2[7]), .S(bl_out));
nch_hvt  M0 ( .D(bl[1]), .B(GND_), .G(yp2[1]), .S(bl_out));
nch_hvt  M5 ( .D(bl[5]), .B(GND_), .G(yp2[5]), .S(bl_out));
nch_hvt  M4 ( .D(bl[4]), .B(GND_), .G(yp2[4]), .S(bl_out));
nch_hvt  M3 ( .D(bl[3]), .B(GND_), .G(yp2[3]), .S(bl_out));
nch_hvt  M2 ( .D(bl[0]), .B(GND_), .G(yp2[0]), .S(bl_out));
nch_hvt  M1 ( .D(bl[2]), .B(GND_), .G(yp2[2]), .S(bl_out));
nch_25  M14 ( .D(bl[7]), .B(GND_), .G(yp2_b_25[7]), .S(vblinhi_rdo));
nch_25  M13 ( .D(bl[6]), .B(GND_), .G(yp2_b_25[6]), .S(vblinhi_rde));
nch_25  M8 ( .D(bl[1]), .B(GND_), .G(yp2_b_25[1]), .S(vblinhi_rdo));
nch_25  M20 ( .D(bl[0]), .B(GND_), .G(yp2_b_25[0]), .S(vblinhi_rde));
nch_25  M12 ( .D(bl[5]), .B(GND_), .G(yp2_b_25[5]), .S(vblinhi_rdo));
nch_25  M11 ( .D(bl[4]), .B(GND_), .G(yp2_b_25[4]), .S(vblinhi_rde));
nch_25  M10 ( .D(bl[3]), .B(GND_), .G(yp2_b_25[3]), .S(vblinhi_rdo));
nch_25  M9 ( .D(bl[2]), .B(GND_), .G(yp2_b_25[2]), .S(vblinhi_rde));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x64, View - schematic
// LAST TIME SAVED: Feb 26 14:34:16 2008
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_x64 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp2, yp2_b_25, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [63:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
input [7:0]  yp3_25;
input [7:0]  yp3_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  bl_med;



ml_ymux_yp2_8 Iml_ymux_yp2_x8 ( .bl(bl_med[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[0]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_2 ( .vdd_tieh(vdd_tieh), .bl(bl[23:16]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[2]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_3 ( .vdd_tieh(vdd_tieh), .bl(bl[31:24]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[3]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_6 ( .vdd_tieh(vdd_tieh), .bl(bl[55:48]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[6]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_7 ( .vdd_tieh(vdd_tieh), .bl(bl[63:56]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[7]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_5 ( .vdd_tieh(vdd_tieh), .bl(bl[47:40]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[5]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_4 ( .vdd_tieh(vdd_tieh), .bl(bl[39:32]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[4]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_1 ( .vdd_tieh(vdd_tieh), .bl(bl[15:8]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[1]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_bls_x328_1f, View - schematic
// LAST TIME SAVED: Jan 17 11:59:56 2011
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_bls_x328_1f ( bl, bl_dummyl, bl_dummyr, bl_out, bl_test,
     vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh,
     pgminhi_dmmy_b_25, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test, yp_test_25, yp_test_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25;

inout [327:0]  bl;
inout [1:0]  bl_test;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;

input [7:0]  yp2;
input [7:0]  yp3_b_25;
input [5:0]  yp1_b_25;
input [1:0]  yp_test_b_25;
input [1:0]  yp_test;
input [7:0]  yp2_b_25;
input [1:0]  yp_test_25;
input [5:0]  yp1;
input [7:0]  yp3_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:5]  blx8_out;

wire  [4:0]  blx64_out;



nch_hvt  M21 ( .D(net224), .B(GND_), .G(yp_test[1]), .S(bl_out));
nch_hvt  M19 ( .D(net228), .B(GND_), .G(yp_test[1]), .S(net224));
nch_hvt  M23 ( .D(net232), .B(GND_), .G(yp_test[0]), .S(bl_out));
nch_hvt  M28 ( .D(net236), .B(GND_), .G(yp1[5]), .S(bl_out));
nch_hvt  M0 ( .D(blx64_out[2]), .B(GND_), .G(yp1[2]), .S(bl_out));
nch_hvt  M22 ( .D(net244), .B(GND_), .G(yp_test[0]), .S(net232));
nch_hvt  M24 ( .D(blx64_out[0]), .B(GND_), .G(yp1[0]), .S(bl_out));
nch_hvt  M30 ( .D(blx8_out[5]), .B(GND_), .G(yp1[5]), .S(net236));
nch_hvt  M3 ( .D(blx64_out[4]), .B(GND_), .G(yp1[4]), .S(bl_out));
nch_hvt  M4 ( .D(blx64_out[3]), .B(GND_), .G(yp1[3]), .S(bl_out));
nch_hvt  M2 ( .D(blx64_out[1]), .B(GND_), .G(yp1[1]), .S(bl_out));
pch_25  M7 ( .D(bl_test[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M8 ( .D(bl_test[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
nch_25  M1 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[0]),
     .S(blx64_out[0]));
nch_25  M26 ( .D(vblinhi_rdo), .B(GND_), .G(yp_test_b_25[1]),
     .S(bl_test[1]));
nch_25  M25 ( .D(bl_test[1]), .B(GND_), .G(yp_test_25[1]), .S(net228));
nch_25  M18 ( .D(vblinhi_rde), .B(GND_), .G(yp_test_b_25[0]),
     .S(bl_test[0]));
nch_25  M11 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[5]),
     .S(blx8_out[5]));
nch_25  M17 ( .D(bl_test[0]), .B(GND_), .G(yp_test_25[0]), .S(net244));
nch_25  M6 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[2]),
     .S(blx64_out[2]));
nch_25  M5 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[1]),
     .S(blx64_out[1]));
nch_25  M10 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[4]),
     .S(blx64_out[4]));
nch_25  M9 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[3]),
     .S(blx64_out[3]));
ml_ymux_bls_x8 Iml_ymux_bls_x8 ( .bl_out(blx8_out[5]),
     .bl(bl[327:320]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_r ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyr[1:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_l ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyl[1:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_0 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[0]), .bl(bl[63:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_2 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[2]), .bl(bl[191:128]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_4 ( .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]), .bl(bl[319:256]),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .bl_out(blx64_out[4]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo));
ml_ymux_bls_x64 Iml_ymux_bls_x64_1 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[1]), .bl(bl[127:64]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_3 ( .yp2(yp2[7:0]), .bl_out(blx64_out[3]),
     .bl(bl[255:192]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .yp2_b_25(yp2_b_25[7:0]), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));

endmodule
// Library - tsmcN40, Cell - inv_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:17 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module inv_25 ( OUT, G, Gb, IN, P, Pb );
output  OUT;

input  G, Gb, IN, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(OUT), .B(Gb), .G(IN), .S(G));
pch_25  M1 ( .D(OUT), .B(Pb), .G(IN), .S(P));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_sup_25, View - schematic
// LAST TIME SAVED: Jul 23 11:45:41 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module oai21x2_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
nch_25  M4 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
nch_25  M7 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));
pch_25  M2 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
pch_25  M0 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));
pch_25  M3 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd25_nor2, View - schematic
// LAST TIME SAVED: Sep 14 15:26:13 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ls_vdd25_nor2 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_25 I79 ( .A(in), .Y(out_vddio_b), .Gb(gnd_), .G(gnd_), .Pb(sup),
     .P(sup), .B(out_vddio));
nor2_25 I151 ( .A(out_vddio_b), .Y(out_vddio), .Gb(gnd_), .G(gnd_),
     .Pb(sup), .P(sup), .B(in_b));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yptest, View - schematic
// LAST TIME SAVED: Jul 21 11:48:14 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yptest ( yp_test_25, yp_test_b_25, yp_test,
     yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25, ysup_25 );
output  yp_test_25, yp_test_b_25;

input  yp_test, yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25,
     ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I181 ( .A(yp_test), .Y(net40));
inv_25 I182 ( .IN(net028), .OUT(yp_test_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));
oai21x2_sup_25 I180 ( .A1(yp_test_b_low_ysup_25), .Y(yp_test_b_25),
     .A0(net37), .B0(yp_test_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(yp_test), .sup(ysup_25),
     .out_vddio_b(net028), .out_vddio(net37), .in_b(net40));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_yp3_sup_25, View - schematic
// LAST TIME SAVED: Jul 23 14:26:50 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module oai21x2_yp3_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M12 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
nch_25  M1 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
nch_25  M0 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));
pch_25  M4 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
pch_25  M6 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));
pch_25  M5 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yp3, View - schematic
// LAST TIME SAVED: Jul 23 14:27:58 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp3 ( yp3_25, yp3_b_25, yp3_b_high_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, ysup_25 );
output  yp3_25, yp3_b_25;

input  yp3_b_high_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



oai21x2_yp3_sup_25 I209 ( .A1(yp3_b_low_ysup_25), .Y(yp3_b_25),
     .A0(net069), .B0(yp3_b_high_b_ysup_25), .ysup_25(ysup_25));
inv_hvt I201 ( .A(yp3_sel), .Y(net075));
inv_hvt I101 ( .A(net075), .Y(net070));
inv_25 I204 ( .IN(yp3_25_b), .OUT(yp3_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd25_nor2 I192 ( .in(net070), .sup(ysup_25),
     .out_vddio_b(yp3_25_b), .out_vddio(net069), .in_b(net075));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_yp21, View - schematic
// LAST TIME SAVED: Jul 21 11:47:41 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp21 ( yp21, yp21_b_25, yp21_b_low_b, yp21_sel,
     ysup_25 );
output  yp21, yp21_b_25;

input  yp21_b_low_b, yp21_sel, ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I213 ( .IN(yp21_b_25_b), .OUT(yp21_b_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
nand2_hvt I206 ( .A(yp21_sel_b), .Y(net50), .B(yp21_b_low_b));
inv_hvt I207 ( .A(net50), .Y(net68));
inv_hvt I208 ( .A(yp21_sel), .Y(yp21_sel_b));
inv_hvt I209 ( .A(yp21_sel_b), .Y(yp21));
ml_ls_vdd25_nor2 I194 ( .in(net68), .sup(ysup_25),
     .out_vddio_b(yp21_b_25_b), .out_vddio(net72), .in_b(net50));

endmodule
// Library - leafcell, Cell - delay150to600ps, View - schematic
// LAST TIME SAVED: Apr 24 15:51:58 2009
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module delay150to600ps ( dly600psout, dlyout, cbit, dlyin );
output  dly600psout, dlyout;

input  dlyin;

input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  min;



delay150ps I0 ( .in(dlyin), .out(min[0]));
delay150ps I4 ( .in(min[2]), .out(dly600psout));
delay150ps I3 ( .in(min[1]), .out(min[2]));
delay150ps I2 ( .in(min[0]), .out(min[1]));
mux4plldly I1 ( .min({dly600psout, min[2:0]}), .cbit(cbit[1:0]),
     .mout(dlyout));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_vblinhi_pgm_drv, View -
//schematic
// LAST TIME SAVED: Jul 29 15:49:55 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_vblinhi_pgm_drv ( vblinhi_pgm_25, ysup_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25 );
inout  vblinhi_pgm_25, ysup_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd_), .B(GND_), .G(en_blinhi_pgm_b_ysup_25),
     .S(vblinhi_pgm_25));
pch_25  M5 ( .D(net10), .B(ysup_25), .G(en_blinhi_pgm_b_ysup_25),
     .S(ysup_25));
pch_25  M0 ( .D(net10), .B(vblinhi_pgm_25), .G(en_blinhi_pgm_b),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_1f, View - schematic
// LAST TIME SAVED: Dec 28 15:35:42 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_1f ( yp1, yp1_b_25, yp2, yp2_b_25, yp3_25,
     yp3_b_25, yp_test_25, yp_test_b_25, vblinhi_pgm_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b, yp1_sel,
     yp2_b_low_b, yp2_sel, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, yp_test,
     ysup_25 );

inout  vblinhi_pgm_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b,
     yp2_b_low_b, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, ysup_25;

output [7:0]  yp3_b_25;
output [7:0]  yp3_25;
output [7:0]  yp2;
output [5:0]  yp1;
output [1:0]  yp_test_25;
output [1:0]  yp_test_b_25;
output [7:0]  yp2_b_25;
output [5:0]  yp1_b_25;

input [7:0]  yp3_sel;
input [5:0]  yp1_sel;
input [7:0]  yp2_sel;
input [1:0]  yp_test;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_1_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1]), .yp_test(yp_test[1]),
     .yp_test_25(yp_test_25[1]));
ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_0_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[0]), .yp_test(yp_test[0]),
     .yp_test_25(yp_test_25[0]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_7_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[7]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[7]), .yp3_25(yp3_25[7]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_6_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[6]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[6]), .yp3_25(yp3_25[6]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_5_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[5]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[5]), .yp3_25(yp3_25[5]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_4_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[4]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[4]), .yp3_25(yp3_25[4]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_3_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[3]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[3]), .yp3_25(yp3_25[3]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_2_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[2]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[2]), .yp3_25(yp3_25[2]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_1_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[1]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[1]), .yp3_25(yp3_25[1]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_0_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[0]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[0]), .yp3_25(yp3_25[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_7_ ( .yp21_sel(yp2_sel[7]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[7]), .yp21(yp2[7]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_6_ ( .yp21_sel(yp2_sel[6]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[6]), .yp21(yp2[6]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_5_ ( .yp21_sel(yp2_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[5]), .yp21(yp2[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_4_ ( .yp21_sel(yp2_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[4]), .yp21(yp2[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_3_ ( .yp21_sel(yp2_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[3]), .yp21(yp2[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_2_ ( .yp21_sel(yp2_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[2]), .yp21(yp2[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_1_ ( .yp21_sel(yp2_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[1]), .yp21(yp2[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_0_ ( .yp21_sel(yp2_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[0]), .yp21(yp2[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_5_ ( .yp21_sel(yp1_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[5]), .yp21(yp1[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_4_ ( .yp21_sel(yp1_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[4]), .yp21(yp1[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_3_ ( .yp21_sel(yp1_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[3]), .yp21(yp1[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_2_ ( .yp21_sel(yp1_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[2]), .yp21(yp1[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_1_ ( .yp21_sel(yp1_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[1]), .yp21(yp1[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_0_ ( .yp21_sel(yp1_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[0]), .yp21(yp1[0]));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_1_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_0_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_a_clkdly, View - schematic
// LAST TIME SAVED: Jul 15 18:44:33 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_pump_a_clkdly ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I206 ( .A(in), .Y(net66));
inv_hvt I205 ( .A(net66), .Y(net70));
inv_hvt I207 ( .A(net70), .Y(out));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(net66), .S(vdd_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_logic_8f_sbb, View -
//schematic
// LAST TIME SAVED: Jul 15 18:44:43 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_8f_sbb ( out_hv_winv, out_hv_woinv, in );
output  out_hv_winv, out_hv_woinv;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_pump_a_clkdly I141 ( .in(net262), .out(net270));
ml_pump_a_clkdly I219 ( .in(net266), .out(net268));
ml_ls_vdd2vdd25 I144 ( .in(net266), .sup(vddp_),
     .out_vddio_b(out_hv_winv), .out_vddio(net279), .in_b(net258));
ml_ls_vdd2vdd25 I148 ( .in(net262), .sup(vddp_),
     .out_vddio_b(out_hv_woinv), .out_vddio(net274), .in_b(net255));
nor2_hvt I140 ( .A(net268), .B(in), .Y(net255));
nor2_hvt I227 ( .A(net264), .B(net270), .Y(net258));
inv_hvt I225 ( .A(net258), .Y(net266));
inv_hvt I134 ( .A(in), .Y(net264));
inv_hvt I226 ( .A(net255), .Y(net262));

endmodule
// Library - sbtlibn65lp, Cell - oai2211x2_hvt, View - schematic
// LAST TIME SAVED: Jul 23 15:48:12 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module oai2211x2_hvt ( Y, A0, A1, B0, B1, C0, D0 );
output  Y;

input  A0, A1, B0, B1, C0, D0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M10 ( .D(net040), .B(GND_), .G(A1), .S(net024));
nch_hvt  M13 ( .D(net040), .B(GND_), .G(A0), .S(net024));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
nch_hvt  M11 ( .D(Y), .B(GND_), .G(C0), .S(net044));
nch_hvt  M0 ( .D(net044), .B(GND_), .G(D0), .S(net040));
nch_hvt  M1 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
pch_hvt  M12 ( .D(Y), .B(VDD_), .G(D0), .S(vdd_));
pch_hvt  M2 ( .D(Y), .B(VDD_), .G(C0), .S(vdd_));
pch_hvt  M18 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M8 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M19 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M7 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - sbtlibn65lp, Cell - anor31_hvt, View - schematic
// LAST TIME SAVED: Jul 23 15:32:42 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module anor31_hvt ( Y, A, B, C, D );
output  Y;

input  A, B, C, D;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(Y), .B(gnd_), .G(A), .S(net23));
nch_hvt  M6 ( .D(net030), .B(gnd_), .G(C), .S(gnd_));
nch_hvt  M5 ( .D(net23), .B(gnd_), .G(B), .S(net030));
nch_hvt  M7 ( .D(Y), .B(gnd_), .G(D), .S(gnd_));
pch_hvt  M3 ( .D(Y), .B(vdd_), .G(D), .S(net35));
pch_hvt  M4 ( .D(net35), .B(vdd_), .G(A), .S(vdd_));
pch_hvt  M0 ( .D(net35), .B(vdd_), .G(B), .S(vdd_));
pch_hvt  M2 ( .D(net35), .B(vdd_), .G(C), .S(vdd_));

endmodule
// Library - sbtlibn65lp, Cell - oai22x2_hvt, View - schematic
// LAST TIME SAVED: Jul 23 15:55:46 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module oai22x2_hvt ( Y, A0, A1, B0, B1 );
output  Y;

input  A0, A1, B0, B1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(Y), .B(GND_), .G(A0), .S(net024));
nch_hvt  M4 ( .D(Y), .B(GND_), .G(A1), .S(net024));
nch_hvt  M1 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M0 ( .D(Y), .B(VDD_), .G(A0), .S(net017));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_logic_1f, View - schematic
// LAST TIME SAVED: Dec 30 13:06:02 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_1f ( dec_trim, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, s_rd, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25, yp1_sel,
     yp2_sel, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, yp21_b_low_b, yp_test, vdd_tieh,
     fsm_blkadd, fsm_coladd, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     tm_allbank_sel, tm_tcol, ysup_25 );
output  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp21_b_low_b;

inout  vdd_tieh;

input  fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h,
     fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec,
     fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis, tm_allbank_sel,
     tm_tcol, ysup_25;

output [3:0]  sb25_high_25;
output [3:0]  sb25_gnd_25;
output [7:0]  yp3_sel;
output [3:0]  sbhv_high_25;
output [7:5]  dec_trim;
output [7:0]  yp2_sel;
output [5:0]  yp1_sel;
output [3:0]  s_rd;
output [3:0]  sbhv_gnd_25;
output [1:0]  yp_test;

input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefpgm;
input [9:0]  fsm_coladd;
input [1:0]  fsm_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp2_sel_b;

wire  [7:0]  yp3_sel_b;

wire  [7:5]  dec_trim_b;

wire  [3:0]  sb25low_b;

wire  [5:0]  yp1_sel_b;

wire  [1:0]  yp_test_b;

wire  [3:0]  s_rd_b;

wire  [2:0]  tdec;

wire  [3:0]  sbhvlow_b;

wire  [1:0]  xadd_b;

wire  [1:0]  xadd;

wire  [9:0]  yadd;

wire  [9:0]  yadd_b;

wire  [3:0]  net561;

wire  [2:0]  tdec_b;



inv_25 I104 ( .IN(net302), .OUT(en_blinhi_pgm_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I285 ( .IN(net311), .OUT(yp3_b_low_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I284 ( .IN(net306), .OUT(yp3_b_high_odd_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I283 ( .IN(net316), .OUT(yp3_b_high_even_b_ysup_25),
     .P(ysup_25), .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
ml_core_ctrl_logic_8f_sbb Isb25_3_ ( .in(sb25low_b[3]),
     .out_hv_woinv(sb25_gnd_25[3]), .out_hv_winv(sb25_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isb25_2_ ( .in(sb25low_b[2]),
     .out_hv_woinv(sb25_gnd_25[2]), .out_hv_winv(sb25_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isb25_1_ ( .in(sb25low_b[1]),
     .out_hv_woinv(sb25_gnd_25[1]), .out_hv_winv(sb25_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isb25_0_ ( .in(sb25low_b[0]),
     .out_hv_woinv(sb25_gnd_25[0]), .out_hv_winv(sb25_high_25[0]));
ml_core_ctrl_logic_8f_sbb Isbhv_3_ ( .in(sbhvlow_b[3]),
     .out_hv_woinv(sbhv_gnd_25[3]), .out_hv_winv(sbhv_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isbhv_2_ ( .in(sbhvlow_b[2]),
     .out_hv_woinv(sbhv_gnd_25[2]), .out_hv_winv(sbhv_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isbhv_1_ ( .in(sbhvlow_b[1]),
     .out_hv_woinv(sbhv_gnd_25[1]), .out_hv_winv(sbhv_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isbhv_0_ ( .in(sbhvlow_b[0]),
     .out_hv_woinv(sbhv_gnd_25[0]), .out_hv_winv(sbhv_high_25[0]));
ml_ls_vdd25_nor2 I106 ( .in(net343), .sup(ysup_25),
     .out_vddio_b(net301), .out_vddio(net302), .in_b(en_blinhi_pgm_b));
ml_ls_vdd25_nor2 I68 ( .in(net576), .sup(ysup_25),
     .out_vddio_b(net306), .out_vddio(net307), .in_b(net308));
ml_ls_vdd25_nor2 I192 ( .in(net396), .sup(ysup_25),
     .out_vddio_b(net311), .out_vddio(net312), .in_b(net544));
ml_ls_vdd25_nor2 I65 ( .in(net571), .sup(ysup_25),
     .out_vddio_b(net316), .out_vddio(net317), .in_b(net318));
exor2_hvt I151_3_ ( .A(net561[0]), .Y(sb25low_b[3]), .B(pgm_hvact_b));
exor2_hvt I151_2_ ( .A(net561[1]), .Y(sb25low_b[2]), .B(pgm_hvact_b));
exor2_hvt I151_1_ ( .A(net561[2]), .Y(sb25low_b[1]), .B(pgm_hvact_b));
exor2_hvt I151_0_ ( .A(net561[3]), .Y(sb25low_b[0]), .B(pgm_hvact_b));
mux2_hvt I152 ( .in1(net504), .in0(net514), .out(ensb25_dec),
     .sel(pgm_hvact));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(tdec[2]), .sel(ref_pgm));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(tdec[1]), .sel(ref_pgm));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(tdec[0]), .sel(ref_pgm));
oai21x2_hvt I55 ( .A1(sa_bl_to_blsa), .Y(net331), .A0(blk_dec),
     .B0(ymux_dis_b));
nor3_hvt I324 ( .B(fsm_tm_testdec), .Y(net335), .A(fsm_tm_allbl_l),
     .C(fsm_tm_allbl_h));
nor3_hvt I321 ( .B(fsm_tm_allbl_h), .Y(net339), .A(nvcmen_buf_b),
     .C(yp3_b_high_b));
nor4_hvt I326 ( .B(fsm_tm_allbl_l), .Y(net343), .D(nvcmen_buf_b),
     .A(net384), .C(fsm_tm_allbl_l));
nor4_hvt I327 ( .B(fsm_tm_allbl_h), .Y(ymux_dis_b), .D(net405),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_h));
nand3_hvt I227 ( .Y(net352), .B(pgm_hvact), .C(fsm_tm_allwl_h),
     .A(fsm_lshven));
nand3_hvt I236_3_ ( .Y(s_rd_b[3]), .B(xadd[0]), .C(en_rdp),
     .A(xadd[1]));
nand3_hvt I236_2_ ( .Y(s_rd_b[2]), .B(xadd_b[0]), .C(en_rdp),
     .A(xadd[1]));
nand3_hvt I236_1_ ( .Y(s_rd_b[1]), .B(xadd[0]), .C(en_rdp),
     .A(xadd_b[1]));
nand3_hvt I236_0_ ( .Y(s_rd_b[0]), .B(xadd_b[0]), .C(en_rdp),
     .A(xadd_b[1]));
nand3_hvt I230 ( .Y(pgm_hvact_b), .B(fsm_pgm), .C(net502),
     .A(fsm_lshven));
nand3_hvt I232 ( .Y(net364), .B(sa_bl_to_blsa), .C(tm_allwl_l_b),
     .A(fsm_vpxaset));
nand3_hvt I233 ( .Y(net368), .B(net492), .C(nvcmen_buf), .A(net387));
nand3_hvt I234_7_ ( .Y(dec_trim_b[7]), .B(tdec[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I234_6_ ( .Y(dec_trim_b[6]), .B(tdec[1]), .C(tdec_b[0]),
     .A(tdec[2]));
nand3_hvt I234_5_ ( .Y(dec_trim_b[5]), .B(tdec_b[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I231_7_ ( .Y(yp2_sel_b[7]), .B(yadd[4]), .C(yadd[3]),
     .A(yadd[5]));
nand3_hvt I231_6_ ( .Y(yp2_sel_b[6]), .B(yadd[4]), .C(yadd_b[3]),
     .A(yadd[5]));
nand3_hvt I231_5_ ( .Y(yp2_sel_b[5]), .B(yadd_b[4]), .C(yadd[3]),
     .A(yadd[5]));
nand3_hvt I231_4_ ( .Y(yp2_sel_b[4]), .B(yadd_b[4]), .C(yadd_b[3]),
     .A(yadd[5]));
nand3_hvt I231_3_ ( .Y(yp2_sel_b[3]), .B(yadd[4]), .C(yadd[3]),
     .A(yadd_b[5]));
nand3_hvt I231_2_ ( .Y(yp2_sel_b[2]), .B(yadd[4]), .C(yadd_b[3]),
     .A(yadd_b[5]));
nand3_hvt I231_1_ ( .Y(yp2_sel_b[1]), .B(yadd_b[4]), .C(yadd[3]),
     .A(yadd_b[5]));
nand3_hvt I231_0_ ( .Y(yp2_sel_b[0]), .B(yadd_b[4]), .C(yadd_b[3]),
     .A(yadd_b[5]));
nand2_hvt I299 ( .A(fsm_tm_rd_mode), .Y(one_blk_sel_b), .B(blk_dec));
nand2_hvt I301 ( .A(pgm_hvact), .Y(net384), .B(pgm_hvact));
nand2_hvt I293 ( .A(fsm_lshven), .Y(net387), .B(pgm_hvact));
nand2_hvt I297 ( .A(blk_dec_b), .Y(blk_dec), .B(tm_pgm_rd_allblk_n));
nand2_hvt I296 ( .A(blk_dec), .Y(net393), .B(fsm_pgmien));
nand2_hvt I294 ( .A(net387), .Y(net396), .B(net335));
nand2_hvt I298 ( .A(all_blk_sel_b), .Y(sa_bl_to_blsa),
     .B(one_blk_sel_b));
nand2_hvt I300 ( .A(tm_allwl_l_b), .Y(net503), .B(blk_dec));
nand2_hvt I295 ( .A(fsm_nvcmen), .Y(net405), .B(fsm_lshven));
nand2_hvt I291_1_ ( .A(yadd[0]), .Y(yp_test_b[1]), .B(ymux_test_en));
nand2_hvt I291_0_ ( .A(yadd_b[0]), .Y(yp_test_b[0]), .B(ymux_test_en));
nand2_hvt I245 ( .A(rd_and_vfy), .Y(all_blk_sel_b), .B(net536));
nand4_hvt I306 ( .D(fsm_blkadd[0]), .A(fsm_blkadd[3]),
     .C(fsm_blkadd[1]), .Y(blk_dec_b), .B(fsm_blkadd[2]));
nand4_hvt I307_5_ ( .D(yadd[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[5]), .B(yadd[8]));
nand4_hvt I307_4_ ( .D(yadd_b[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[4]), .B(yadd[8]));
nand4_hvt I304_7_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[7]), .B(yadd[2]));
nand4_hvt I304_6_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[6]), .B(yadd[2]));
nand4_hvt I304_5_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[5]), .B(yadd[2]));
nand4_hvt I304_4_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[4]), .B(yadd[2]));
nand4_hvt I304_3_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[3]), .B(yadd_b[2]));
nand4_hvt I304_2_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[2]), .B(yadd_b[2]));
nand4_hvt I304_1_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[1]), .B(yadd_b[2]));
nand4_hvt I304_0_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[0]), .B(yadd_b[2]));
nand4_hvt I239 ( .D(fsm_tm_rprd), .Y(net429), .B(fsm_lshven),
     .C(nvcmen_buf), .A(rd_and_vfy));
nand4_hvt I308 ( .D(fsm_lshven), .A(tm_allwl_l_b), .C(pgm_hvact),
     .Y(net436), .B(blk_dec));
nor2_hvt I316_5_ ( .A(yp1_sel_b[5]), .B(tm_tcol), .Y(yp1_sel[5]));
nor2_hvt I316_4_ ( .A(yp1_sel_b[4]), .B(tm_tcol), .Y(yp1_sel[4]));
nor2_hvt I310 ( .A(fsm_pgmvfy), .B(fsm_pgm), .Y(net443));
nor2_hvt I315 ( .A(net331), .B(net530), .Y(ymux_test_en));
nor2_hvt I312 ( .A(net579), .B(net532), .Y(net449));
nor2_hvt I319 ( .A(fsm_rd), .B(fsm_pgmvfy), .Y(net452));
nor2_hvt I328 ( .A(net331), .B(tm_tcol), .Y(ymux_en_core));
nor2_hvt I317_3_ ( .A(yp1_sel_b[3]), .B(tm_tcol), .Y(yp1_sel[3]));
nor2_hvt I317_2_ ( .A(yp1_sel_b[2]), .B(tm_tcol), .Y(yp1_sel[2]));
nor2_hvt I317_1_ ( .A(yp1_sel_b[1]), .B(tm_tcol), .Y(yp1_sel[1]));
nor2_hvt I317_0_ ( .A(yp1_sel_b[0]), .B(tm_tcol), .Y(yp1_sel[0]));
nor2_hvt I313 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I318 ( .A(fsm_tm_rd_mode), .B(fsm_pgmvfy), .Y(net464));
anor21_hvt I119_1_ ( .A(fsm_rowadd[1]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I119_0_ ( .A(fsm_rowadd[0]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
anor21_hvt I109 ( .A(pgm_hvact), .B(fsm_tm_allwl_h), .Y(net505),
     .C(nvcmen_buf_b));
inv_hvt I271_9_ ( .A(yadd[9]), .Y(yadd_b[9]));
inv_hvt I272_9_ ( .A(vdd_tieh), .Y(yadd[9]));
inv_hvt I247 ( .A(net452), .Y(rd_and_vfy));
inv_hvt I265 ( .A(net464), .Y(net484));
inv_hvt I323 ( .A(fsm_tm_allbl_l), .Y(yp3_b_high_b));
inv_hvt I237_3_ ( .A(s_rd_b[3]), .Y(s_rd[3]));
inv_hvt I237_2_ ( .A(s_rd_b[2]), .Y(s_rd[2]));
inv_hvt I237_1_ ( .A(s_rd_b[1]), .Y(s_rd[1]));
inv_hvt I237_0_ ( .A(s_rd_b[0]), .Y(s_rd[0]));
inv_hvt I252_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I252_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I200 ( .A(fsm_tm_testdec), .Y(net492));
inv_hvt I261 ( .A(net393), .Y(sa_bl_to_pgm_glb));
inv_hvt I271_8_ ( .A(yadd_b[8]), .Y(yadd[8]));
inv_hvt I271_7_ ( .A(yadd_b[7]), .Y(yadd[7]));
inv_hvt I271_6_ ( .A(yadd_b[6]), .Y(yadd[6]));
inv_hvt I271_5_ ( .A(yadd_b[5]), .Y(yadd[5]));
inv_hvt I271_4_ ( .A(yadd_b[4]), .Y(yadd[4]));
inv_hvt I271_3_ ( .A(yadd_b[3]), .Y(yadd[3]));
inv_hvt I271_2_ ( .A(yadd_b[2]), .Y(yadd[2]));
inv_hvt I271_1_ ( .A(yadd_b[1]), .Y(yadd[1]));
inv_hvt I271_0_ ( .A(yadd_b[0]), .Y(yadd[0]));
inv_hvt I268 ( .A(net579), .Y(vddp_rd_overw));
inv_hvt I260 ( .A(nvcmen_buf_b), .Y(nvcmen_buf));
inv_hvt I254 ( .A(net576), .Y(net308));
inv_hvt I278 ( .A(fsm_pgmvfy), .Y(net502));
inv_hvt I281 ( .A(net503), .Y(net504));
inv_hvt I279 ( .A(net505), .Y(net506));
inv_hvt I251 ( .A(net352), .Y(net508));
inv_hvt I258 ( .A(net368), .Y(yp21_b_low_b));
inv_hvt I263 ( .A(fsm_nvcmen), .Y(nvcmen_buf_b));
inv_hvt I280 ( .A(net364), .Y(net514));
inv_hvt I264 ( .A(tm_allbank_sel), .Y(tm_pgm_rd_allblk_n));
inv_hvt I250 ( .A(net436), .Y(net518));
inv_hvt I241 ( .A(net429), .Y(en_rdp));
inv_hvt I255 ( .A(net343), .Y(en_blinhi_pgm_b));
inv_hvt I249 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I277 ( .A(pgm_hvact_b), .Y(pgm_hvact));
inv_hvt I266 ( .A(net443), .Y(ref_pgm));
inv_hvt I259 ( .A(tm_tcol), .Y(net530));
inv_hvt I267 ( .A(fsm_multibl_read), .Y(net532));
inv_hvt I262 ( .A(all_blk_sel_b), .Y(net534));
inv_hvt I272_8_ ( .A(fsm_coladd[8]), .Y(yadd_b[8]));
inv_hvt I272_7_ ( .A(fsm_coladd[7]), .Y(yadd_b[7]));
inv_hvt I272_6_ ( .A(fsm_coladd[6]), .Y(yadd_b[6]));
inv_hvt I272_5_ ( .A(fsm_coladd[5]), .Y(yadd_b[5]));
inv_hvt I272_4_ ( .A(fsm_coladd[4]), .Y(yadd_b[4]));
inv_hvt I272_3_ ( .A(fsm_coladd[3]), .Y(yadd_b[3]));
inv_hvt I272_2_ ( .A(fsm_coladd[2]), .Y(yadd_b[2]));
inv_hvt I272_1_ ( .A(fsm_coladd[1]), .Y(yadd_b[1]));
inv_hvt I272_0_ ( .A(fsm_coladd[0]), .Y(yadd_b[0]));
inv_hvt I201 ( .A(fsm_tm_rd_mode), .Y(net536));
inv_hvt I270_2_ ( .A(tdec[2]), .Y(tdec_b[2]));
inv_hvt I270_1_ ( .A(tdec[1]), .Y(tdec_b[1]));
inv_hvt I270_0_ ( .A(tdec[0]), .Y(tdec_b[0]));
inv_hvt I273_7_ ( .A(yp2_sel_b[7]), .Y(yp2_sel[7]));
inv_hvt I273_6_ ( .A(yp2_sel_b[6]), .Y(yp2_sel[6]));
inv_hvt I273_5_ ( .A(yp2_sel_b[5]), .Y(yp2_sel[5]));
inv_hvt I273_4_ ( .A(yp2_sel_b[4]), .Y(yp2_sel[4]));
inv_hvt I273_3_ ( .A(yp2_sel_b[3]), .Y(yp2_sel[3]));
inv_hvt I273_2_ ( .A(yp2_sel_b[2]), .Y(yp2_sel[2]));
inv_hvt I273_1_ ( .A(yp2_sel_b[1]), .Y(yp2_sel[1]));
inv_hvt I273_0_ ( .A(yp2_sel_b[0]), .Y(yp2_sel[0]));
inv_hvt I256_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I256_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I256_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I257 ( .A(net396), .Y(net544));
inv_hvt I274_7_ ( .A(yp3_sel_b[7]), .Y(yp3_sel[7]));
inv_hvt I274_6_ ( .A(yp3_sel_b[6]), .Y(yp3_sel[6]));
inv_hvt I274_5_ ( .A(yp3_sel_b[5]), .Y(yp3_sel[5]));
inv_hvt I274_4_ ( .A(yp3_sel_b[4]), .Y(yp3_sel[4]));
inv_hvt I274_3_ ( .A(yp3_sel_b[3]), .Y(yp3_sel[3]));
inv_hvt I274_2_ ( .A(yp3_sel_b[2]), .Y(yp3_sel[2]));
inv_hvt I274_1_ ( .A(yp3_sel_b[1]), .Y(yp3_sel[1]));
inv_hvt I274_0_ ( .A(yp3_sel_b[0]), .Y(yp3_sel[0]));
inv_hvt I253 ( .A(net571), .Y(net318));
inv_hvt I275_1_ ( .A(yp_test_b[1]), .Y(yp_test[1]));
inv_hvt I275_0_ ( .A(yp_test_b[0]), .Y(yp_test[0]));
oai2211x2_hvt I86_3_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[3]), .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai2211x2_hvt I86_2_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[2]), .A0(yadd[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
oai2211x2_hvt I86_1_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[1]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd[6]));
oai2211x2_hvt I86_0_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net449),
     .Y(yp1_sel_b[0]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
anor31_hvt I155_3_ ( .A(ensb25_dec), .D(net506), .B(xadd[1]),
     .Y(net561[0]), .C(xadd[0]));
anor31_hvt I155_2_ ( .A(ensb25_dec), .D(net506), .B(xadd[1]),
     .Y(net561[1]), .C(xadd_b[0]));
anor31_hvt I155_1_ ( .A(ensb25_dec), .D(net506), .B(xadd_b[1]),
     .Y(net561[2]), .C(xadd[0]));
anor31_hvt I155_0_ ( .A(ensb25_dec), .D(net506), .B(xadd_b[1]),
     .Y(net561[3]), .C(xadd_b[0]));
anor31_hvt I121_3_ ( .A(net518), .D(net508), .B(xadd[1]),
     .Y(sbhvlow_b[3]), .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net518), .D(net508), .B(xadd[1]),
     .Y(sbhvlow_b[2]), .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net518), .D(net508), .B(xadd_b[1]),
     .Y(sbhvlow_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net518), .D(net508), .B(xadd_b[1]),
     .Y(sbhvlow_b[0]), .C(xadd_b[0]));
anor31_hvt I107 ( .A(fsm_tm_testdec), .D(net339), .B(nvcmen_buf),
     .Y(net571), .C(yadd[0]));
anor31_hvt I108 ( .A(fsm_tm_testdec), .D(net339), .B(nvcmen_buf),
     .Y(net576), .C(yadd_b[0]));
oai22x2_hvt I93 ( .A1(net534), .Y(net579), .A0(net484),
     .B0(fsm_nv_rri_trim), .B1(fsm_nv_sisi_ui));

endmodule
// Library - NVCM_40nm, Cell - ml_dff_nvcm, View - schematic
// LAST TIME SAVED: Jun 21 11:02:43 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_dff_nvcm ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I132 ( .A(clk_b), .Y(clk_buf));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I146 ( .A(net57), .Y(Q));
inv_hvt I147 ( .A(net60), .Y(QN));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net64), .Y(net57));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net64), .Y(net53));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net60), .Y(net57));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net53));
nor2_hvt I129 ( .A(net57), .B(R), .Y(net60));
nor2_hvt I125 ( .A(net53), .B(R), .Y(net64));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_resref_40nm, View - schematic
// LAST TIME SAVED: Sep 11 14:49:31 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_sa_resref_40nm ( bl_in, bl_out, ref );
inout  bl_in, bl_out;

inout [3:0]  ref;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R9 ( .MINUS(ref[3]), .PLUS(ref[2]), .BULK(gnd_));
rppolywo_m  R11 ( .MINUS(ref[1]), .PLUS(ref[0]), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(net41), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(ref[2]), .PLUS(ref[1]), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(ref[0]), .PLUS(net41), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(ref[3]), .BULK(gnd_));

endmodule
// Library - leafcell, Cell - pll_finedly, View - schematic
// LAST TIME SAVED: May 11 17:26:27 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pll_finedly ( pll_fbout, cbit, pll_fbin );
output  pll_fbout;

input  pll_fbin;

input [3:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  min;



delay150to600ps I6 ( .dly600psout(net40), .cbit(cbit[1:0]),
     .dlyin(net44), .dlyout(min[2]));
delay150to600ps I5 ( .dly600psout(net44), .cbit(cbit[1:0]),
     .dlyin(net52), .dlyout(min[1]));
delay150to600ps I4 ( .dly600psout(net48), .cbit(cbit[1:0]),
     .dlyin(net40), .dlyout(min[3]));
delay150to600ps I0 ( .dly600psout(net52), .cbit(cbit[1:0]),
     .dlyin(pll_fbin), .dlyout(min[0]));
mux4plldly I1 ( .min(min[3:0]), .cbit(cbit[3:2]), .mout(pll_fbout));

endmodule
// Library - ice1chip, Cell - pll_bufwrap_ice1f, View - schematic
// LAST TIME SAVED: Apr  8 12:23:22 2011
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pll_bufwrap_ice1f ( f_out, f_in );
output  f_out;

input  f_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



fabric_buf_ice8p I6 ( .f_in(f_in), .f_out(f_out));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_restop_40nm, View - schematic
// LAST TIME SAVED: Sep 16 19:06:55 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_sa_restop_40nm ( bl_bot, bl_top );
inout  bl_bot, bl_top;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R24 ( .MINUS(bl_top), .PLUS(net66), .BULK(gnd_));
rppolywo_m  R23 ( .MINUS(net66), .PLUS(bl_bot), .BULK(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_resbot_40nm, View - schematic
// LAST TIME SAVED: Sep 16 11:24:37 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_sa_resbot_40nm ( bl_in, bl_out, in_dec, sa_ngate );
inout  bl_in, bl_out, in_dec;


input [4:1]  sa_ngate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M9 ( .D(net026), .B(GND_), .G(sa_ngate[2]), .S(gnd_));
nch_hvt  M20 ( .D(in_dec), .B(GND_), .G(sa_ngate[1]), .S(gnd_));
nch_hvt  M10 ( .D(net072), .B(GND_), .G(sa_ngate[3]), .S(gnd_));
nch_hvt  M11 ( .D(net132), .B(GND_), .G(sa_ngate[4]), .S(gnd_));
rppolywo_m  R15 ( .MINUS(bl_in), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(bl_in), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(net026), .PLUS(in_dec), .BULK(gnd_));
rppolywo_m  R12 ( .MINUS(bl_in), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(in_dec), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R9 ( .MINUS(bl_out), .PLUS(net132), .BULK(gnd_));
rppolywo_m  R8 ( .MINUS(net072), .PLUS(net026), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(net132), .PLUS(net072), .BULK(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_gwlgnd_nor2, View - schematic
// LAST TIME SAVED: Jul 10 13:02:38 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_gwlgnd_nor2 ( gwl_gnd_25, gwl_b_sup_25, gwl_b_25,
     gwl_b_gnden_25 );
output  gwl_gnd_25;

inout  gwl_b_sup_25;

input  gwl_b_25, gwl_b_gnden_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(net14), .B(GND_), .G(gwl_b_gnden_25), .S(GND_));
nch_25  M0 ( .D(gwl_gnd_25), .B(GND_), .G(gwl_b_25), .S(net14));
pch_25  M2 ( .D(gwl_gnd_25), .B(gwl_b_sup_25), .G(gwl_b_25),
     .S(gwl_b_sup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp, View - schematic
// LAST TIME SAVED: Nov 30 17:03:56 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp ( wp, gwl_gnd_rp_25, ngate_25, gwl_b_25,
     gwl_gnd_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv );
output  wp;

inout  gwl_gnd_rp_25, ngate_25;

input  gwl_b_25, gwl_gnd_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M11 ( .D(net18), .B(GND_), .G(s_b_25), .S(gwl_gnd_25));
nch_25  M12 ( .D(wp), .B(GND_), .G(ngate_25), .S(net18));
nch_25  M10 ( .D(net18), .B(GND_), .G(gwl_b_25), .S(gwl_gnd_25));
pch_25  M0 ( .D(gwl_gnd_rp_25), .B(gwp_hv), .G(s_rd_b_hv), .S(wp));
pch_25  M6 ( .D(wp), .B(gwp_hv), .G(s_b_hv), .S(gwp_hv));

endmodule
// Library - tsmcN40, Cell - nand2_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:22 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module nand2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(Y), .B(Gb), .G(A), .S(net16));
nch_25  M3 ( .D(net16), .B(Gb), .G(B), .S(G));
pch_25  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M2 ( .D(Y), .B(Pb), .G(B), .S(P));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp, View - schematic
// LAST TIME SAVED: Aug 27 14:09:22 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_b_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(out_ref), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M2 ( .D(out_div), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M8 ( .D(out_ref), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M5 ( .D(out_div), .B(GND_), .G(saen_b_25), .S(gnd_));
pch_25  M4_1_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M3 ( .D(out_ref), .B(vddp_), .G(in_ref), .S(net65));
pch_25  M6 ( .D(out_div), .B(vddp_), .G(in_div), .S(net65));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_top, View - schematic
// LAST TIME SAVED: Sep 15 18:21:46 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp_top ( sa_out, vdd_tieh, in_div, in_ref, saen_25
     );
output  sa_out;

inout  vdd_tieh;

input  in_div, in_ref, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M6 ( .D(sa_out_b_25), .B(gnd_), .G(saen_b_25), .S(gnd_));
nch_25  M0 ( .D(net053), .B(gnd_), .G(saen_25), .S(gnd_));
nch_25  M5 ( .D(sa_out_b_25), .B(gnd_), .G(out_div2), .S(gnd_));
nch_25  M1 ( .D(sa_bias), .B(gnd_), .G(vdd_tieh), .S(net45));
rppolywo_m  R0 ( .MINUS(net039), .PLUS(net45), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net053), .PLUS(net039), .BULK(gnd_));
pch_25  M43 ( .D(sa_bias), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M4_1_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M7 ( .D(sa_out_b_25), .B(vddp_), .G(out_div2), .S(net089));
pch_25  M3 ( .D(net089), .B(vddp_), .G(sa_bias), .S(vddp_));
nand2_25 I80 ( .G(gnd_), .Pb(vdd_), .A(net051), .Y(net038), .P(vdd_),
     .B(saen_25), .Gb(gnd_));
inv_25 I89 ( .IN(sa_out_b_25), .OUT(net051), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I91 ( .IN(saen_25), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net038), .OUT(sa_out), .P(vdd_), .Pb(vdd_), .G(gnd_),
     .Gb(gnd_));
ml_core_sa_comp Icore_sa_comp0 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp Icore_sa_comp1 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref2), .in_div(in_div2),
     .out_ref(out_ref), .out_div(out_div2));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa, View - schematic
// LAST TIME SAVED: Dec  7 15:20:54 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_sa ( nv_dataout, blsa, vdd_tieh, vddp_tieh, vpxa,
     dec_ok, dec_trim, fsm_rst_b, fsm_sample, fsm_tm_ref,
     fsm_tm_testdec, sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, tm_testdec_wr );
output  nv_dataout;

inout  blsa, vdd_tieh, vddp_tieh, vpxa;

input  dec_ok, fsm_rst_b, fsm_sample, fsm_tm_testdec, saen_25,
     saen_b_vpxa, saprd_b_vpxa, testdec_en_b, tm_testdec_wr;

input [1:0]  fsm_tm_ref;
input [4:1]  sa_ngate;
input [7:5]  dec_trim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  ref;



ml_dff_nvcm I132 ( .R(net273), .D(net274), .CLK(fsm_sample),
     .QN(net276), .Q(nv_dataout));
nch  WR_CELL ( .D(net0159), .B(GND_), .G(testdec_b), .S(net167));
rppolywo_m  R9 ( .MINUS(net171), .PLUS(net175), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net0137), .PLUS(net171), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net220), .PLUS(net0137), .BULK(gnd_));
ml_core_sa_resref_40nm Irref_bot ( .bl_in(net142), .bl_out(net236),
     .ref(ref[3:0]));
ml_core_sa_restop_40nm Irref_top ( .bl_top(net0221), .bl_bot(net0159));
ml_core_sa_resbot_40nm Irsen_bot ( .bl_in(blsa), .bl_out(net175),
     .sa_ngate(sa_ngate[4:1]), .in_dec(net197));
pch  M0 ( .D(net167), .B(vdd_), .G(testdec_en_b), .S(vdd_));
nor2_hvt I214 ( .B(high_res_b), .Y(net214), .A(fsm_tm_testdec));
nor3_hvt I102 ( .B(dec_trim[6]), .Y(high_res_b), .A(dec_trim[5]),
     .C(dec_trim[7]));
mux2_hvt I206 ( .in1(blsa), .in0(net197), .out(in_div),
     .sel(testdec_b));
mux2_hvt I270 ( .in1(ref[1]), .in0(ref[0]), .out(net185),
     .sel(fsm_tm_ref[0]));
mux2_hvt I271 ( .in1(ref[3]), .in0(ref[2]), .out(net184),
     .sel(fsm_tm_ref[0]));
mux2_hvt I279 ( .in1(net0195), .in0(ref[2]), .out(in_ref),
     .sel(testdec_b));
mux2_hvt I234 ( .in1(dec_ok), .in0(sa_out), .out(net274),
     .sel(tm_testdec_wr));
mux2_hvt I272 ( .in1(net184), .in0(net185), .out(net0195),
     .sel(fsm_tm_ref[1]));
inv_hvt I247 ( .A(fsm_rst_b), .Y(net273));
inv_hvt I208 ( .A(fsm_tm_testdec), .Y(testdec_b));
inv_hvt I248 ( .A(net214), .Y(net226));
nch_hvt  M23 ( .D(net220), .B(GND_), .G(dec_trim[7]), .S(gnd_));
nch_hvt  M16 ( .D(net175), .B(GND_), .G(net226), .S(gnd_));
nch_hvt  M13 ( .D(net228), .B(GND_), .G(vdd_tieh), .S(net240));
nch_hvt  M18 ( .D(net151), .B(GND_), .G(vdd_tieh), .S(net142));
nch_hvt  M21 ( .D(net0137), .B(GND_), .G(dec_trim[6]), .S(gnd_));
nch_hvt  M19 ( .D(net236), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M20 ( .D(net171), .B(GND_), .G(dec_trim[5]), .S(gnd_));
nch_hvt  M12 ( .D(net240), .B(GND_), .G(vdd_tieh), .S(net151));
nch_25  M22 ( .D(net167), .B(GND_), .G(vddp_tieh), .S(net228));
vdd_tielow I204 ( .gnd_tiel(gnd_tlow));
ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 ( .gwl_b_gnden_25(vddp_tieh),
     .gwl_b_sup_25(vpxa), .gwl_b_25(saen_b_vpxa),
     .gwl_gnd_25(gwl_gnd_25_ref));
ml_rock_lwldrv_wp Irock_lwldrv_wp ( .gwl_gnd_rp_25(gwl_gnd_25_ref),
     .s_rd_b_hv(saprd_b_vpxa), .gwl_gnd_25(gwl_gnd_25_ref),
     .s_b_hv(gwl_gnd_25_ref), .gwp_hv(gwl_gnd_25_ref),
     .gwl_b_25(gnd_tlow), .ngate_25(vpxa), .s_b_25(saprd_b_vpxa),
     .wp(net0221));
ml_core_sa_comp_top Icore_sa_comp_top ( .vdd_tieh(vdd_tieh),
     .saen_25(saen_25), .in_ref(in_ref), .in_div(in_div),
     .sa_out(sa_out));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_top, View - schematic
// LAST TIME SAVED: Sep 11 13:36:38 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_sa_top ( nv_dataout, bl_out, bl_pgm_glb, vdd_tieh,
     vddp_tieh, vpxa, dec_ok, dec_trim, fsm_rst_b, fsm_sample,
     fsm_tm_ref, fsm_tm_testdec, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     tm_dma, tm_testdec_wr );
output  nv_dataout;

inout  bl_out, bl_pgm_glb, vdd_tieh, vddp_tieh, vpxa;

input  dec_ok, fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, tm_dma, tm_testdec_wr;

input [1:0]  fsm_tm_ref;
input [4:1]  sa_ngate;
input [7:5]  dec_trim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(net073), .Y(net048));
inv_hvt I45 ( .A(net048), .Y(nv_dataout));
nch_hvt  M2 ( .D(bl_out), .B(GND_), .G(sa_bl_to_blsa), .S(net71));
nch_hvt  M1 ( .D(bl_out), .B(GND_), .G(sa_bl_to_pgm_glb),
     .S(bl_pgm_glb));
nch_hvt  M4 ( .D(net71), .B(GND_), .G(tm_dma), .S(gnd_));
ml_core_sa Iml_core_sa ( .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .vddp_tieh(vddp_tieh),
     .vdd_tieh(vdd_tieh), .sa_ngate(sa_ngate[4:1]), .dec_ok(dec_ok),
     .testdec_en_b(testdec_en_b), .tm_testdec_wr(tm_testdec_wr),
     .fsm_tm_testdec(fsm_tm_testdec), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .dec_trim(dec_trim[7:5]), .nv_dataout(net073), .vpxa(vpxa),
     .blsa(net71));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_core_40nm, View - schematic
// LAST TIME SAVED: Jul 15 18:30:49 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_hv_ls_inv_core_40nm ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net26), .G(sel_25), .S(net26));
pch_25  M5 ( .D(net19), .B(net22), .G(sel_b_25), .S(net22));
pch_25  M7 ( .D(net26), .B(in_hv), .G(net19), .S(in_hv));
pch_25  M6 ( .D(net22), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(net19), .B(GND_), .G(vddp_tieh), .S(net37));
nch_25  M15 ( .D(net37), .B(GND_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(GND_), .G(vddp_tieh), .S(net29));
nch_25  M14 ( .D(net29), .B(GND_), .G(sel_25), .S(gnd_));

endmodule
// Library - leafcell, Cell - pllmate_40lp, View - schematic
// LAST TIME SAVED: Nov  3 07:32:44 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pllmate_40lp ( pll_bypass, pll_cbit, pll_fb, pll_fse, pll_out1,
     pll_out2, pll_ref, pll_reset, pll_sdo, cbit, fo_dlyadj,
     fo_pll_bypass, fo_pll_sck, fo_pll_sdi, fo_pllfb, fo_pllref,
     fo_pllreset, pad_pllref, pllout_in, prog );
output  pll_bypass, pll_fb, pll_fse, pll_out1, pll_out2, pll_ref,
     pll_reset, pll_sdo;

input  fo_pll_bypass, fo_pll_sck, fo_pll_sdi, fo_pllfb, fo_pllref,
     fo_pllreset, pad_pllref, pllout_in, prog;

output [16:0]  pll_cbit;

input [7:0]  fo_dlyadj;
input [36:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [25:0]  q;

wire  [25:0]  net137;

wire  [24:17]  obit;

wire  [1:0]  net165;

wire  [3:0]  net114;

wire  [3:0]  net119;

wire  [1:0]  net157;



pllcfg_sr26_40lp I_pllcfg_sr ( .q(q[25:0]), .reset(prog),
     .pll_sdi(fo_pll_sdi), .pll_sck(fo_pll_sck));
fabric_buf_ice8p I_BUF4PLL_SDO ( .f_in(net176), .f_out(pll_sdo));
tiehi I_tiehi ( .tiehi(net100));
tielo I_tielo ( .tielo(pll_tielo));
mux4plldly I14 ( .min({pll_tielo, pll_tielo, pll_tielo, pllout2_d1}),
     .cbit({pll_tielo, pll_tielo}), .mout(pllout2_d2));
mux4plldly I15 ( .min({pll_tielo, pll_tielo, pll_tielo, pllout2_d2}),
     .cbit({pll_tielo, pll_tielo}), .mout(net107));
delay150ps I12 ( .in(net108), .out(pllout2_d1));
oa4plldly_40lp I_oa4plldly_fb_3_ ( .cbit(cbit[29]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[3]), .out(net114[0]));
oa4plldly_40lp I_oa4plldly_fb_2_ ( .cbit(cbit[28]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[2]), .out(net114[1]));
oa4plldly_40lp I_oa4plldly_fb_1_ ( .cbit(cbit[27]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[1]), .out(net114[2]));
oa4plldly_40lp I_oa4plldly_fb_0_ ( .cbit(cbit[26]), .fda_en(cbit[30]),
     .prog(prog), .in(fo_dlyadj[0]), .out(net114[3]));
oa4plldly_40lp I_oa4plldly_out_3_ ( .cbit(cbit[34]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[7]), .out(net119[0]));
oa4plldly_40lp I_oa4plldly_out_2_ ( .cbit(cbit[33]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[6]), .out(net119[1]));
oa4plldly_40lp I_oa4plldly_out_1_ ( .cbit(cbit[32]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[5]), .out(net119[2]));
oa4plldly_40lp I_oa4plldly_out_0_ ( .cbit(cbit[31]), .fda_en(cbit[35]),
     .prog(prog), .in(fo_dlyadj[4]), .out(net119[3]));
nand2_hvt I9_1_ ( .A(obit[24]), .Y(net157[0]), .B(net140));
nand2_hvt I9_0_ ( .A(obit[23]), .Y(net157[1]), .B(net140));
nand2_hvt I2_1_ ( .A(obit[20]), .B(net140), .Y(net165[0]));
nand2_hvt I2_0_ ( .A(obit[19]), .B(net140), .Y(net165[1]));
pllphase_sr_40lp I_pllphase_sr ( .tielo(pll_tielo), .tiehi(net100),
     .f_out(f_out), .cbit(obit[21]), .f_dvd2(f_dvd2),
     .f_dvd4_p0(f_dvd4_p0), .f_dvd4_p90(f_dvd4_p90), .sr(pll_reset),
     .CLK(pllout_in));
mux2_hvt I_MUX4ShftCbit_25_ ( .in1(q[25]), .in0(cbit[36]),
     .out(net137[0]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_24_ ( .in1(q[24]), .in0(cbit[24]),
     .out(net137[1]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_23_ ( .in1(q[23]), .in0(cbit[23]),
     .out(net137[2]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_22_ ( .in1(q[22]), .in0(cbit[22]),
     .out(net137[3]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_21_ ( .in1(q[21]), .in0(cbit[21]),
     .out(net137[4]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_20_ ( .in1(q[20]), .in0(cbit[20]),
     .out(net137[5]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_19_ ( .in1(q[19]), .in0(cbit[19]),
     .out(net137[6]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_18_ ( .in1(q[18]), .in0(cbit[18]),
     .out(net137[7]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_17_ ( .in1(q[17]), .in0(cbit[17]),
     .out(net137[8]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_16_ ( .in1(q[16]), .in0(cbit[16]),
     .out(net137[9]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_15_ ( .in1(q[15]), .in0(cbit[15]),
     .out(net137[10]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_14_ ( .in1(q[14]), .in0(cbit[14]),
     .out(net137[11]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_13_ ( .in1(q[13]), .in0(cbit[13]),
     .out(net137[12]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_12_ ( .in1(q[12]), .in0(cbit[12]),
     .out(net137[13]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_11_ ( .in1(q[11]), .in0(cbit[11]),
     .out(net137[14]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_10_ ( .in1(q[10]), .in0(cbit[10]),
     .out(net137[15]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_9_ ( .in1(q[9]), .in0(cbit[9]),
     .out(net137[16]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_8_ ( .in1(q[8]), .in0(cbit[8]),
     .out(net137[17]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_7_ ( .in1(q[7]), .in0(cbit[7]),
     .out(net137[18]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_6_ ( .in1(q[6]), .in0(cbit[6]),
     .out(net137[19]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_5_ ( .in1(q[5]), .in0(cbit[5]),
     .out(net137[20]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_4_ ( .in1(q[4]), .in0(cbit[4]),
     .out(net137[21]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_3_ ( .in1(q[3]), .in0(cbit[3]),
     .out(net137[22]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_2_ ( .in1(q[2]), .in0(cbit[2]),
     .out(net137[23]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_1_ ( .in1(q[1]), .in0(cbit[1]),
     .out(net137[24]), .sel(net178));
mux2_hvt I_MUX4ShftCbit_0_ ( .in1(q[0]), .in0(cbit[0]),
     .out(net137[25]), .sel(net178));
inv_hvt I0 ( .A(pll_bypass), .Y(net140));
clkmux2buffer I_MUX4PLLRef ( .in1(fo_pllref_buf), .in0(pad_pllref),
     .out(pll_ref), .sel(obit[22]));
clkbuffer500um BUF_PLL_OUT1 ( .in(net189), .out(pll_out1));
clkbuffer500um BUF_PLL_OUT2 ( .in(net107), .out(pll_out2));
clkbuffer500um I_BUF4PLL_FB ( .in(net186), .out(pll_fb));
clkbuffer200u Ifo_pllfb_buf ( .in(fo_pllfb), .out(fo_pllfb_buf));
clkbuffer200u Ifo_pllref_buf ( .in(fo_pllref), .out(fo_pllref_buf));
clkmux4to1 I7 ( net158, {net157[0], net157[1]}, f_dvd4_p0, f_dvd4_p90,
     f_dvd2, f_out);
clkmux4to1 I_mux4PhaseOut ( net108, {net165[0], net165[1]}, f_dvd4_p0,
     f_dvd4_p90, f_dvd2, f_out);
clkmux4to1 I_clkmux4finedly ( net172, obit[18:17], pllout_in,
     f_dvd4_p0, f_dvd4_p0, fo_pllfb_buf);
buffer500um I_BUF4PLL_BYPASS ( .in(fo_pll_bypass), .out(pll_bypass));
bram_bufferx4 I3 ( .in(q[25]), .out(net176));
bram_bufferx4 I_cbit23_buffer ( .in(cbit[25]), .out(net178));
bram_bufferx4 I_cbit_buffer_25_ ( .in(net137[0]), .out(pll_fse));
bram_bufferx4 I_cbit_buffer_24_ ( .in(net137[1]), .out(obit[24]));
bram_bufferx4 I_cbit_buffer_23_ ( .in(net137[2]), .out(obit[23]));
bram_bufferx4 I_cbit_buffer_22_ ( .in(net137[3]), .out(obit[22]));
bram_bufferx4 I_cbit_buffer_21_ ( .in(net137[4]), .out(obit[21]));
bram_bufferx4 I_cbit_buffer_20_ ( .in(net137[5]), .out(obit[20]));
bram_bufferx4 I_cbit_buffer_19_ ( .in(net137[6]), .out(obit[19]));
bram_bufferx4 I_cbit_buffer_18_ ( .in(net137[7]), .out(obit[18]));
bram_bufferx4 I_cbit_buffer_17_ ( .in(net137[8]), .out(obit[17]));
bram_bufferx4 I_cbit_buffer_16_ ( .in(net137[9]), .out(pll_cbit[16]));
bram_bufferx4 I_cbit_buffer_15_ ( .in(net137[10]), .out(pll_cbit[15]));
bram_bufferx4 I_cbit_buffer_14_ ( .in(net137[11]), .out(pll_cbit[14]));
bram_bufferx4 I_cbit_buffer_13_ ( .in(net137[12]), .out(pll_cbit[13]));
bram_bufferx4 I_cbit_buffer_12_ ( .in(net137[13]), .out(pll_cbit[12]));
bram_bufferx4 I_cbit_buffer_11_ ( .in(net137[14]), .out(pll_cbit[11]));
bram_bufferx4 I_cbit_buffer_10_ ( .in(net137[15]), .out(pll_cbit[10]));
bram_bufferx4 I_cbit_buffer_9_ ( .in(net137[16]), .out(pll_cbit[9]));
bram_bufferx4 I_cbit_buffer_8_ ( .in(net137[17]), .out(pll_cbit[8]));
bram_bufferx4 I_cbit_buffer_7_ ( .in(net137[18]), .out(pll_cbit[7]));
bram_bufferx4 I_cbit_buffer_6_ ( .in(net137[19]), .out(pll_cbit[6]));
bram_bufferx4 I_cbit_buffer_5_ ( .in(net137[20]), .out(pll_cbit[5]));
bram_bufferx4 I_cbit_buffer_4_ ( .in(net137[21]), .out(pll_cbit[4]));
bram_bufferx4 I_cbit_buffer_3_ ( .in(net137[22]), .out(pll_cbit[3]));
bram_bufferx4 I_cbit_buffer_2_ ( .in(net137[23]), .out(pll_cbit[2]));
bram_bufferx4 I_cbit_buffer_1_ ( .in(net137[24]), .out(pll_cbit[1]));
bram_bufferx4 I_cbit_buffer_0_ ( .in(net137[25]), .out(pll_cbit[0]));
cfg4pllreset I_cfg4pllreset ( .prog(prog), .in(fo_pllreset),
     .out(pll_reset));
pll_finedly I11 ( .cbit({net114[0], net114[1], net114[2], net114[3]}),
     .pll_fbin(net172), .pll_fbout(net186));
pll_finedly I_pll_finedly ( .cbit({net119[0], net119[1], net119[2],
     net119[3]}), .pll_fbin(net158), .pll_fbout(net189));

endmodule
// Library - NVCM_40nm, Cell - ml_s_b_hv_sw, View - schematic
// LAST TIME SAVED: Sep  7 10:32:39 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_s_b_hv_sw ( sbout_hv, ssup_hv, sbout_gnd_25, sbout_high_25,
     vddp_tieh );
inout  sbout_hv, ssup_hv;

input  sbout_gnd_25, sbout_high_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_core_40nm Iml_hv_ls_inv_core_40nm ( .sel_b_25(net62),
     .sel_25(sbout_high_25), .out_b_hv(sbout_hv_b), .in_hv(ssup_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M23 ( .D(sbout_hv), .B(GND_), .G(vddp_tieh), .S(net34));
nch_25  M7 ( .D(net34), .B(GND_), .G(sbout_gnd_25), .S(gnd_));
inv_25 I114 ( .IN(sbout_high_25), .OUT(net62), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M0 ( .D(net46), .B(ssup_hv), .G(sbout_hv_b), .S(ssup_hv));
pch_25  M2 ( .D(sbout_hv), .B(net46), .G(sbout_gnd_25), .S(net46));

endmodule
// Library - NVCM_40nm, Cell - ml_wp_ctrl, View - schematic
// LAST TIME SAVED: Jul 27 15:30:44 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_wp_ctrl ( s_b_25, s_b_hv, sb25sup_25, sbhvsup_hv, vddp_tieh,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25 );
inout  sb25sup_25, sbhvsup_hv, vddp_tieh;


inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [3:0]  sbhv_gnd_25;
input [3:0]  sb25_high_25;
input [3:0]  sb25_gnd_25;
input [3:0]  sbhv_high_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_s_b_hv_sw Iml_s_b_25_sw_3_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[3]),
     .sbout_hv(s_b_25[3]), .sbout_high_25(sb25_high_25[3]));
ml_s_b_hv_sw Iml_s_b_25_sw_2_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[2]),
     .sbout_hv(s_b_25[2]), .sbout_high_25(sb25_high_25[2]));
ml_s_b_hv_sw Iml_s_b_25_sw_1_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[1]),
     .sbout_hv(s_b_25[1]), .sbout_high_25(sb25_high_25[1]));
ml_s_b_hv_sw Iml_s_b_25_sw_0_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[0]),
     .sbout_hv(s_b_25[0]), .sbout_high_25(sb25_high_25[0]));
ml_s_b_hv_sw Iml_s_b_hv_sw_3_ ( .sbout_high_25(sbhv_high_25[3]),
     .sbout_hv(s_b_hv[3]), .sbout_gnd_25(sbhv_gnd_25[3]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_2_ ( .sbout_high_25(sbhv_high_25[2]),
     .sbout_hv(s_b_hv[2]), .sbout_gnd_25(sbhv_gnd_25[2]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_1_ ( .sbout_high_25(sbhv_high_25[1]),
     .sbout_hv(s_b_hv[1]), .sbout_gnd_25(sbhv_gnd_25[1]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_0_ ( .sbout_high_25(sbhv_high_25[0]),
     .sbout_hv(s_b_hv[0]), .sbout_gnd_25(sbhv_gnd_25[0]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_core_ctrl_top_1f, View - schematic
// LAST TIME SAVED: Dec 29 14:16:08 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_ctrl_top_1f ( gwl_b_gnden_25, nv_dataout, s_rd, yp1,
     yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25, yp_test, yp_test_25,
     yp_test_b_25, bl_out, bl_pgm_glb, s_b_25, s_b_hv, sb25sup_25,
     sbhvsup_hv, vblinhi_pgm_25, vdd_tieh, vpxa, ysup_25, dec_ok,
     fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, testdec_en_b, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );
output  gwl_b_gnden_25, nv_dataout;

inout  bl_out, bl_pgm_glb, sb25sup_25, sbhvsup_hv, vblinhi_pgm_25,
     vdd_tieh, vpxa, ysup_25;

input  dec_ok, fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [7:0]  yp2;
output [5:0]  yp1_b_25;
output [1:0]  yp_test_25;
output [7:0]  yp3_b_25;
output [1:0]  yp_test_b_25;
output [7:0]  yp2_b_25;
output [1:0]  yp_test;
output [5:0]  yp1;
output [7:0]  yp3_25;
output [3:0]  s_rd;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [2:0]  fsm_trim_rrefrd;
input [9:0]  fsm_coladd;
input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefpgm;
input [1:0]  fsm_tm_ref;
input [3:0]  fsm_blkadd;
input [4:1]  sa_ngate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp2_sel;

wire  [3:0]  sb25_gnd_25;

wire  [3:0]  sbhv_gnd_25;

wire  [3:0]  sbhv_high_25;

wire  [5:0]  yp1_sel;

wire  [3:0]  sb25_high_25;

wire  [7:5]  dec_trim;

wire  [7:0]  yp3_sel;



ml_ymux_ctrl_1f Iml_ymux_ctrl_1f ( .yp1_b_25(yp1_b_25[5:0]),
     .yp1(yp1[5:0]), .yp1_sel(yp1_sel[5:0]), .yp2(yp2[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2_sel(yp2_sel[7:0]),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_sel(yp3_sel[7:0]), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test(yp_test[1:0]),
     .yp2_b_low_b(yp21_b_low_b), .yp1_b_low_b(yp21_b_low_b),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .yp_test_25(yp_test_25[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_core_ctrl_logic_1f Icore_ctrl_logic_1f (
     .fsm_coladd(fsm_coladd[9:0]), .yp1_sel(yp1_sel[5:0]),
     .vdd_tieh(vdd_tieh), .fsm_tm_rprd(fsm_tm_rprd), .s_rd(s_rd[3:0]),
     .tm_allbank_sel(tm_allbank_sel), .yp2_sel(yp2_sel[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_tm_allwl_l(tm_allwl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25), .tm_tcol(tm_tcol),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_allbl_l(tm_allbl_l), .fsm_pgm(fsm_pgm),
     .fsm_tm_allbl_h(tm_allbl_h), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_nvcmen(fsm_nvcmen), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_blkadd(fsm_blkadd[3:0]),
     .yp_test(yp_test[1:0]), .yp21_b_low_b(yp21_b_low_b),
     .yp3_sel(yp3_sel[7:0]), .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .sbhv_high_25(sbhv_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sb25_gnd_25(sb25_gnd_25[3:0]),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .dec_trim(dec_trim[7:5]));
pch_hvt  M0 ( .D(vdd_tieh), .B(vdd_), .G(net223), .S(vdd_));
pch_25  M4 ( .D(vddp_tieh), .B(vddp_), .G(net223), .S(vddp_));
nch_hvt  M3 ( .D(net223), .B(GND_), .G(net223), .S(gnd_));
inv_25 I38 ( .IN(net240), .OUT(gwl_b_gnden_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I30 ( .IN(fsm_gwlbdis_b_25), .OUT(net240), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_core_sa_top Icore_sa_top ( .fsm_tm_ref(fsm_tm_ref[1:0]),
     .saprd_b_vpxa(saprd_b_vpxa), .vddp_tieh(vddp_tieh),
     .vdd_tieh(vdd_tieh), .sa_ngate(sa_ngate[4:1]), .dec_ok(dec_ok),
     .testdec_en_b(testdec_en_b), .tm_dma(tm_dma),
     .fsm_tm_testdec(fsm_tm_testdec), .tm_testdec_wr(tm_testdec_wr),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .dec_trim(dec_trim[7:5]), .nv_dataout(nv_dataout), .vpxa(vpxa),
     .bl_pgm_glb(bl_pgm_glb), .bl_out(bl_out));
ml_wp_ctrl Iml_wp_ctrl ( .vddp_tieh(vddp_tieh),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .sbhv_high_25(sbhv_high_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_gnd_25(sb25_gnd_25[3:0]), .s_b_25(s_b_25[3:0]),
     .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp_x4, View - schematic
// LAST TIME SAVED: Nov 30 17:14:06 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x4 ( wp, gwl_b_sup_25, ngate_25, gwl_b_25,
     gwl_b_gnden_25, gwp_hv, s_b_25, s_b_hv, s_rd_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_25, gwl_b_gnden_25, gwp_hv;

output [3:0]  wp;

input [3:0]  s_b_25;
input [3:0]  s_rd_b_hv;
input [3:0]  s_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwl_b_25(gwl_b_25), .gwl_gnd_25(gwl_gnd_25));
ml_rock_lwldrv_wp Iml_lwldrv_1 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[1]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[1]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[1]), .wp(wp[1]));
ml_rock_lwldrv_wp Iml_lwldrv_2 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[2]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[2]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[2]), .wp(wp[2]));
ml_rock_lwldrv_wp Iml_lwldrv_3 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[3]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[3]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3]), .wp(wp[3]));
ml_rock_lwldrv_wp Iml_lwldrv_0 ( .gwl_gnd_rp_25(rp_float),
     .s_rd_b_hv(s_rd_b_hv[0]), .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[0]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[0]), .wp(wp[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wp_x108_1f, View -
//schematic
// LAST TIME SAVED: Dec 29 14:15:11 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x108_1f ( wp, gwl_b_sup_25, ngate_25, s_b_25,
     s_b_hv, gwl_b_25, gwl_b_gnden_25, gwp_hv, s_rd_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_gnden_25;

output [107:0]  wp;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [26:0]  gwp_hv;
input [26:0]  gwl_b_25;
input [3:0]  s_rd_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_26_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[26]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[107:104]),
     .gwl_b_25(gwl_b_25[26]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_25_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[25]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[103:100]),
     .gwl_b_25(gwl_b_25[25]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_24_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[24]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[99:96]),
     .gwl_b_25(gwl_b_25[24]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_23_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[23]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[95:92]),
     .gwl_b_25(gwl_b_25[23]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_22_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[22]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[91:88]),
     .gwl_b_25(gwl_b_25[22]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_21_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[21]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[87:84]),
     .gwl_b_25(gwl_b_25[21]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_20_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[20]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[83:80]),
     .gwl_b_25(gwl_b_25[20]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_19_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[19]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[79:76]),
     .gwl_b_25(gwl_b_25[19]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_18_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[18]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[75:72]),
     .gwl_b_25(gwl_b_25[18]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_17_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[17]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[71:68]),
     .gwl_b_25(gwl_b_25[17]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_16_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[16]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[67:64]),
     .gwl_b_25(gwl_b_25[16]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_15_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[15]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[63:60]),
     .gwl_b_25(gwl_b_25[15]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_14_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[14]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[59:56]),
     .gwl_b_25(gwl_b_25[14]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_13_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[13]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[55:52]),
     .gwl_b_25(gwl_b_25[13]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_12_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[12]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[51:48]),
     .gwl_b_25(gwl_b_25[12]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_11_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[11]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[47:44]),
     .gwl_b_25(gwl_b_25[11]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_10_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[10]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[43:40]),
     .gwl_b_25(gwl_b_25[10]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_9_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[9]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[39:36]),
     .gwl_b_25(gwl_b_25[9]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_8_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[8]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[35:32]),
     .gwl_b_25(gwl_b_25[8]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_7_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[7]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[31:28]),
     .gwl_b_25(gwl_b_25[7]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_6_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[6]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[27:24]),
     .gwl_b_25(gwl_b_25[6]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_5_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[5]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[23:20]),
     .gwl_b_25(gwl_b_25[5]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_4_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[4]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[19:16]),
     .gwl_b_25(gwl_b_25[4]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_3_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[3]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[15:12]),
     .gwl_b_25(gwl_b_25[3]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_2_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[2]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[11:8]),
     .gwl_b_25(gwl_b_25[2]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_1_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[1]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[7:4]),
     .gwl_b_25(gwl_b_25[1]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_0_ (
     .s_rd_b_hv(s_rd_b_hv[3:0]), .gwl_b_gnden_25(gwl_b_gnden_25),
     .gwl_b_sup_25(gwl_b_sup_25), .gwp_hv(gwp_hv[0]),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]), .wp(wp[3:0]),
     .gwl_b_25(gwl_b_25[0]), .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_338x112_top_1f, View - schematic
// LAST TIME SAVED: Dec 29 14:19:40 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_338x112_top_1f ( nv_dataout, s_rd, bl_pgm_glb,
     gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde,
     vblinhi_rdo, vpxa, ysup_25, fsm_blkadd, fsm_coladd,
     fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25,
     s_rd_b_hv, sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa,
     testdec_en_b, testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );
output  nv_dataout;

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  s_rd;

input [1:0]  fsm_rowadd;
input [107:0]  wr;
input [9:0]  fsm_coladd;
input [26:0]  gwl_b_25;
input [2:0]  fsm_trim_rrefrd;
input [26:0]  gwp_hv;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [4:1]  sa_ngate;
input [1:0]  fsm_tm_ref;
input [3:0]  s_rd_b_hv;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp3_b_25;

wire  [1:0]  bl_dummyl;

wire  [5:0]  yp1;

wire  [107:0]  wp;

wire  [7:0]  yp2_b_25;

wire  [1:0]  bl_dummyr;

wire  [327:0]  bl;

wire  [7:0]  yp3;

wire  [5:0]  yp1_b_25;

wire  [1:0]  yp_test_25;

wire  [1:0]  bl_test;

wire  [3:0]  s_b_hv;

wire  [1:0]  yp_test_b_25;

wire  [1:0]  yp_test;

wire  [7:0]  yp2;

wire  [3:0]  s_b_25;



ml_testdec_rowsx108_1f Iml_testdec_rowsx108_1f (
     .dec_det_buf(dec_det_buf), .dec_bias(dec_bias), .dec_det(dec_det),
     .wr(wr[107:0]), .wp(wp[107:0]));
ml_testdec_columnsx330_1f Iml_testdec_columnsx330_1f ( .bl(bl[327:0]),
     .dec_det_buf(dec_det_buf), .bl_test(bl_test[1:0]),
     .bl_dummyl(bl_dummyl[1:0]), .bl_dummyr(bl_dummyr[1:0]),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25));
vdd_tielow I47 ( .gnd_tiel(net148));
nvcm_cell_338x112_1f Invcm_cell_338x112_1f ( .wr_dummyt({net148,
     net148}), .wr_dummyb({net148, net148}), .wp_dummyt({net148,
     net148}), .wp_dummyb({net148, net148}), .bl_test(bl_test[1:0]),
     .bl_dummyr(bl_dummyr[1:0]), .bl_dummyl(bl_dummyl[1:0]),
     .bl(bl[327:0]), .wp(wp[107:0]), .wr(wr[107:0]));
ml_testdec_bgen Itestdec_bgen ( .dec_ok(dec_ok_l),
     .testdec_en_b(testdec_en_b), .testdec_prec_b(testdec_prec_b),
     .dec_bias(dec_bias), .dec_det(dec_det));
ml_ymux_bls_x328_1f Iml_ymux_bls_x328_1f (
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_25(yp_test_25[1:0]),
     .yp_test(yp_test[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .yp2_b_25(yp2_b_25[7:0]),
     .vblinhi_rdo(vblinhi_rdo), .bl_dummyr(bl_dummyr[1:0]),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyl(bl_dummyl[1:0]), .bl_test(bl_test[1:0]),
     .bl_out(bl_out), .bl(bl[327:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vdd_tieh(vdd_tieh),
     .yp1(yp1[5:0]), .yp2(yp2[7:0]), .yp1_b_25(yp1_b_25[5:0]));
ml_core_ctrl_top_1f Icore_ctrl_top_1f ( .yp1(yp1[5:0]),
     .yp1_b_25(yp1_b_25[5:0]), .dec_ok(dec_ok_l),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .s_rd(s_rd[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .sa_ngate(sa_ngate[4:1]), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .fsm_coladd(fsm_coladd[9:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .gwl_b_gnden_25(gwl_b_gnden_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .vdd_tieh(vdd_tieh), .tm_testdec_wr(tm_testdec_wr),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_blkadd(fsm_blkadd[3:0]), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .nv_dataout(nv_dataout), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_pgm_25(vblinhi_pgm_25),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .bl_out(bl_out),
     .yp_test(yp_test[1:0]));
ml_rock_lwldrv_wp_x108_1f Iml_rock_lwldrv_wp_x108_1f (
     .gwp_hv(gwp_hv[26:0]), .gwl_b_25(gwl_b_25[26:0]),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .ngate_25(ngate_25),
     .gwl_b_sup_25(gwl_b_sup_25), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .gwl_b_gnden_25(gwl_b_gnden_25), .wp(wp[107:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_bank_1_1f, View - schematic
// LAST TIME SAVED: Dec 30 15:03:13 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_bank_1_1f ( nv_dataout, s_rd, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  s_rd;
output [8:4]  nv_dataout;

input [2:0]  fsm_trim_rrefrd;
input [26:0]  gwl_b_25;
input [1:0]  fsm_tm_ref;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [7:0]  fsm_rowadd;
input [26:0]  gwp_hv;
input [4:1]  sa_ngate;
input [3:0]  s_rd_b_hv;
input [107:0]  wr;
input [9:0]  fsm_coladd;
input [3:0]  fsm_blkadd_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net530;

wire  [3:0]  net524;

wire  [3:0]  net297;

wire  [3:0]  net355;

wire  [3:0]  net523;

wire  [3:0]  net529;



ml_core_338x112_top_1f Iblk_4 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net523[0], net523[1], net523[2],
     net523[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .sa_ngate(sa_ngate[4:1]), .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[4]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f Iblk_7 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net530[0], net530[1], net530[2],
     net530[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .sa_ngate(sa_ngate[4:1]), .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd[1], fsm_blkadd[0]}), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .ysup_25(ysup_25), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .testdec_odd_b_25(testdec_odd_b_25),
     .vpxa(vpxa), .testdec_even_b_25(testdec_even_b_25),
     .saen_b_vpxa(saen_b_vpxa), .vblinhi_rdo(vblinhi_rdo),
     .saen_25(saen_25), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[7]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f blk_6 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net355[0], net355[1], net355[2],
     net355[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .sa_ngate(sa_ngate[4:1]), .tm_allbank_sel(tm_allbank_sel),
     .nv_dataout(nv_dataout[6]), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nvcmen(fsm_nvcmen), .fsm_pgm(fsm_pgm),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_rd(fsm_rd), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rowadd(fsm_rowadd[1:0]), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rst_b(fsm_rst_b), .fsm_sample(fsm_sample),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .ngate_25(ngate_25),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .saen_25(saen_25), .vblinhi_rdo(vblinhi_rdo),
     .saen_b_vpxa(saen_b_vpxa), .testdec_even_b_25(testdec_even_b_25),
     .vpxa(vpxa), .testdec_odd_b_25(testdec_odd_b_25),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ysup_25(ysup_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd[2], fsm_blkadd[1],
     fsm_blkadd_b[0]}), .tm_testdec_wr(tm_testdec_wr),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_338x112_top_1f Iblk_5 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net297[0], net297[1], net297[2],
     net297[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .sa_ngate(sa_ngate[4:1]), .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[5]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f Iblk_8 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net529[0], net529[1], net529[2],
     net529[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .sa_ngate(sa_ngate[4:1]), .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[8]),
     .fsm_coladd(fsm_coladd[9:0]));
inv_hvt I66_3_ ( .A(net523[0]), .Y(net524[0]));
inv_hvt I66_2_ ( .A(net523[1]), .Y(net524[1]));
inv_hvt I66_1_ ( .A(net523[2]), .Y(net524[2]));
inv_hvt I66_0_ ( .A(net523[3]), .Y(net524[3]));
inv_hvt I6_3_ ( .A(net524[0]), .Y(s_rd[3]));
inv_hvt I6_2_ ( .A(net524[1]), .Y(s_rd[2]));
inv_hvt I6_1_ ( .A(net524[2]), .Y(s_rd[1]));
inv_hvt I6_0_ ( .A(net524[3]), .Y(s_rd[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_core_bank_0_1f, View - schematic
// LAST TIME SAVED: Dec 30 14:58:14 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_core_bank_0_1f ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_ref, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv,
     sa_ngate, saen_25, saen_b_vpxa, saprd_b_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen,
     fsm_ymuxdis, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, testdec_en_b, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  nv_dataout;

input [9:0]  fsm_coladd;
input [1:0]  fsm_tm_ref;
input [3:0]  s_rd_b_hv;
input [2:0]  fsm_trim_rrefrd;
input [107:0]  wr;
input [26:0]  gwp_hv;
input [7:0]  fsm_rowadd;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefpgm;
input [26:0]  gwl_b_25;
input [4:1]  sa_ngate;
input [3:0]  fsm_blkadd_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net378;

wire  [3:0]  net320;

wire  [3:0]  net431;

wire  [3:0]  net432;



ml_core_338x112_top_1f Iblk_2 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net320[0], net320[1], net320[2],
     net320[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[2]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f blk_1 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net431[0], net431[1], net431[2],
     net431[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[1]),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_tm_trow(fsm_tm_trow),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_rd(fsm_rd),
     .bl_pgm_glb(bl_pgm_glb), .fsm_rowadd(fsm_rowadd[1:0]),
     .gwl_b_sup_25(gwl_b_sup_25), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .ngate_25(ngate_25), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .saen_25(saen_25), .vblinhi_rdo(vblinhi_rdo),
     .saen_b_vpxa(saen_b_vpxa), .testdec_even_b_25(testdec_even_b_25),
     .vpxa(vpxa), .testdec_odd_b_25(testdec_odd_b_25),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ysup_25(ysup_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd[0]}), .tm_testdec_wr(tm_testdec_wr),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_338x112_top_1f Iblk_0 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net432[0], net432[1], net432[2],
     net432[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[0]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_338x112_top_1f Iblk_3 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_b_25(gwl_b_25[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .saprd_b_vpxa(saprd_b_vpxa),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rd({net378[0], net378[1], net378[2],
     net378[3]}), .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .tm_allbank_sel(tm_allbank_sel), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .tm_testdec_wr(tm_testdec_wr), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd_b[2], fsm_blkadd[1], fsm_blkadd[0]}),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .vblinhi_rde(vblinhi_rde), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .sbhvsup_hv(sbhvsup_hv), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .sb25sup_25(sb25sup_25), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[3]),
     .fsm_coladd(fsm_coladd[9:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr, View - schematic
// LAST TIME SAVED: Jul 28 11:15:51 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr ( wr, gwl_wr_25, s_25, wr_sup_25 );
output  wr;

input  gwl_wr_25, s_25, wr_sup_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I59 ( .A(gwl_wr_25), .Y(net27), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(s_25));
inv_25 I38 ( .IN(net27), .OUT(wr), .P(wr_sup_25), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr_x4, View - schematic
// LAST TIME SAVED: Jan 21 18:09:38 2008
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x4 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  gwl_wr_25, wr_sup_25;

output [3:0]  wr;

input [3:0]  s_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr Iml_lwldrv_2 ( .gwl_wr_25(gwl_wr_25), .wr(wr[2]),
     .s_25(s_25[2]), .wr_sup_25(wr_sup_25));
ml_rock_lwldrv_wr Iml_lwldrv_1 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[1]), .wr(wr[1]));
ml_rock_lwldrv_wr Iml_lwldrv_3 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3]), .wr(wr[3]));
ml_rock_lwldrv_wr Iml_lwldrv_0 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[0]), .wr(wr[0]));

endmodule
// Library - leafcell, Cell - pinlatbuf12p, View - schematic
// LAST TIME SAVED: Dec 24 09:07:59 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pinlatbuf12p ( cout, cbit, icegate, pad_in, prog );
output  cout;

input  cbit, icegate, pad_in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I_txgate_lvt_2 ( .in(cout), .out(net13), .pp(net046),
     .nn(net17));
txgate_lvt I_txgate_lvt_1 ( .in(pad_in), .out(net13), .pp(net17),
     .nn(net046));
nand2_lvt I_nand2_lvt ( .A(net19), .Y(net044), .B(net13));
nand2_lvt I5 ( .A(icegate), .Y(net046), .B(cbit));
inv_lvt I6 ( .A(net046), .Y(net17));
inv_lvt I24 ( .A(prog), .Y(net19));
inv_lvt I_inv_lvt ( .A(net044), .Y(cout));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_wr_x108_1f, View -
//schematic
// LAST TIME SAVED: Dec 29 14:33:23 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x108_1f ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  wr_sup_25;

output [107:0]  wr;

input [26:0]  gwl_wr_25;
input [3:0]  s_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_26_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[107:104]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[26]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_25_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[103:100]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[25]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_24_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[99:96]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[24]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_23_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[95:92]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[23]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_22_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[91:88]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[22]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_21_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[87:84]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[21]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_20_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[83:80]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[20]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_19_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[79:76]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[19]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_18_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[75:72]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[18]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_17_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[71:68]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[17]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_16_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[67:64]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[16]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_15_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[63:60]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[15]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_14_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[59:56]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[14]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_13_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[55:52]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[13]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_12_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[51:48]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[12]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_11_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[47:44]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[11]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_10_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[43:40]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[10]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_9_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[39:36]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[9]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_8_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[35:32]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[8]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_7_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[31:28]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[7]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_6_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[27:24]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[6]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_5_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[23:20]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[5]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_4_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[19:16]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[4]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_3_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[15:12]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[3]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_2_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[11:8]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[2]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_1_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[7:4]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[1]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_0_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[3:0]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[0]));

endmodule
// Library - tsmcN40, Cell - nor3_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:26 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module nor3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(Y), .B(Gb), .G(B), .S(G));
nch_25  M5 ( .D(Y), .B(Gb), .G(C), .S(G));
nch_25  M4 ( .D(Y), .B(Gb), .G(A), .S(G));
pch_25  M0 ( .D(net16), .B(Pb), .G(B), .S(net12));
pch_25  M1 ( .D(net12), .B(Pb), .G(A), .S(P));
pch_25  M2 ( .D(Y), .B(Pb), .G(C), .S(net16));

endmodule
// Library - tsmcN40, Cell - nand3_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:23 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module nand3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(net21), .B(Gb), .G(C), .S(G));
nch_25  M3 ( .D(Y), .B(Gb), .G(A), .S(net25));
nch_25  M4 ( .D(net25), .B(Gb), .G(B), .S(net21));
pch_25  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(P));
pch_25  M2 ( .D(Y), .B(Pb), .G(C), .S(P));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vddp2vpxa, View - schematic
// LAST TIME SAVED: Jul 28 11:31:26 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_ls_vddp2vpxa ( out_33, out_b_33, sup, in_25, in_b_25 );
output  out_33, out_b_33;

inout  sup;

input  in_25, in_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(out_33), .B(gnd_), .G(in_b_25), .S(gnd_));
nch_25  M7 ( .D(out_b_33), .B(gnd_), .G(in_25), .S(gnd_));
pch_25  M1 ( .D(out_b_33), .B(sup), .G(in_25), .S(net60));
pch_25  M2 ( .D(out_33), .B(sup), .G(in_b_25), .S(net56));
pch_25  M3 ( .D(net56), .B(sup), .G(out_b_33), .S(sup));
pch_25  M5 ( .D(net60), .B(sup), .G(out_33), .S(sup));

endmodule
// Library - NVCM_40nm, Cell - ml_rock_lwldrv_gwhv, View - schematic
// LAST TIME SAVED: Jul 13 15:44:38 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rock_lwldrv_gwhv ( gwp_hv, gwp_sup_hv, gwl_25, gwl_25_b,
     vddp_tieh );
output  gwp_hv;

inout  gwp_sup_hv;

input  gwl_25, gwl_25_b, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M10 ( .D(net0129), .B(gnd_), .G(vddp_tieh), .S(net050));
nch_25  M12 ( .D(gwp_hv), .B(gnd_), .G(vddp_tieh), .S(net034));
nch_25  M11 ( .D(net034), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M13 ( .D(net050), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M14 ( .D(net054), .B(gnd_), .G(vddp_tieh), .S(net058));
nch_25  M15 ( .D(net058), .B(gnd_), .G(gwl_25), .S(gnd_));
pch_25  M6 ( .D(net067), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M16 ( .D(gwp_hv), .B(net067), .G(gwl_25_b), .S(net067));
pch_25  M5 ( .D(net054), .B(net087), .G(gwl_25), .S(net087));
pch_25  M8 ( .D(net087), .B(gwp_sup_hv), .G(net0129), .S(gwp_sup_hv));
pch_25  M9 ( .D(net091), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M7 ( .D(net0129), .B(net091), .G(gwl_25_b), .S(net091));

endmodule
// Library - NVCM_40nm, Cell - ml_gwl_drv, View - schematic
// LAST TIME SAVED: Aug  2 17:23:15 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_gwl_drv ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25,
     radd_1_25, radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );
output  gwl_b_25, gwl_wr_25, gwp_hv;

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25, radd_1_25,
     radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I133 ( .IN(gwl_wp_25), .OUT(gwl_wp_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I100 ( .IN(out_33), .OUT(gwl_b_25), .P(gwl_b_sup_25),
     .Pb(gwl_b_sup_25), .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(gwlb_25), .OUT(gwlb_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nor3_25 I123 ( .B(net76), .A(net68), .C(net84), .Y(dec_sel_25),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nand3_25 I44 ( .B(radd_4_25), .A(radd_5_25), .Y(net76), .C(radd_3_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I122 ( .B(radd_1_25), .A(radd_2_25), .Y(net84), .C(radd_0_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I121 ( .B(gwlgrpsel_25), .A(gwlgrpsel_25), .Y(net68),
     .C(radd_6_25), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nor2_25 I128 ( .A(wr_frcen_25), .Y(net056), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(dec_sel_25));
nor2_25 I127 ( .A(wr_dis_25), .Y(gwl_wr_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(net056));
nor2_25 I129 ( .A(dec_sel_25), .Y(net096), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_en_25));
nor2_25 I130 ( .A(net096), .Y(gwlb_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_dis_25));
nor2_25 I131 ( .A(dec_sel_25), .Y(net058), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_frcen_25));
nor2_25 I132 ( .A(net058), .Y(gwl_wp_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_dis_25));
ml_ls_vddp2vpxa I99 ( .in_25(gwlb_25), .sup(gwl_b_sup_25),
     .in_b_25(gwlb_b_25), .out_33(out_33), .out_b_33(net053));
ml_rock_lwldrv_gwhv Iml_rock_lwldrv_gwhv ( .gwp_sup_hv(gwp_sup_hv),
     .vddp_tieh(vddp_tieh), .gwp_hv(gwp_hv), .gwl_25(gwl_wp_25),
     .gwl_25_b(gwl_wp_b_25));

endmodule
// Library - NVCM_40nm, Cell - ml_gwl_drv_x27_1f, View - schematic
// LAST TIME SAVED: Dec 29 15:02:09 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_gwl_drv_x27_1f ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25,
     gnv2_b_25, gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25,
     gnv5_b_25, gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1,
     gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25, gnv2_b_25,
     gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25, gnv5_b_25,
     gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1, gwl_misc_25,
     gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

output [26:0]  gwp_hv;
output [26:0]  gwl_b_25;
output [26:0]  gwl_wr_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_gwl_drv Igwl_drv_25_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[25]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[25]), .gwl_wr_25(gwl_wr_25[25]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_24_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[24]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[24]), .gwl_wr_25(gwl_wr_25[24]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_23_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[23]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[23]), .gwl_wr_25(gwl_wr_25[23]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_22_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[22]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[22]), .gwl_wr_25(gwl_wr_25[22]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_21_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[21]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[21]), .gwl_wr_25(gwl_wr_25[21]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_20_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[20]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[20]), .gwl_wr_25(gwl_wr_25[20]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_19_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[19]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[19]), .gwl_wr_25(gwl_wr_25[19]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_18_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[18]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[18]), .gwl_wr_25(gwl_wr_25[18]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_17_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[17]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[17]), .gwl_wr_25(gwl_wr_25[17]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_16_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[16]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[16]), .gwl_wr_25(gwl_wr_25[16]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_b_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_misc_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[26]),
     .radd_0_25(vddp_tieh), .radd_1_25(vddp_tieh),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_misc_25),
     .gwp_hv(gwp_hv[26]), .gwl_wr_25(gwl_wr_25[26]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_15_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[15]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[15]), .gwl_wr_25(gwl_wr_25[15]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_14_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[14]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[14]), .gwl_wr_25(gwl_wr_25[14]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_13_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[13]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[13]), .gwl_wr_25(gwl_wr_25[13]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_12_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[12]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[12]), .gwl_wr_25(gwl_wr_25[12]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_11_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[11]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[11]), .gwl_wr_25(gwl_wr_25[11]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_10_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[10]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[10]), .gwl_wr_25(gwl_wr_25[10]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_9_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[9]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[9]), .gwl_wr_25(gwl_wr_25[9]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_8_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[8]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[8]),
     .gwl_wr_25(gwl_wr_25[8]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_7_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[7]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[7]),
     .gwl_wr_25(gwl_wr_25[7]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_6_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[6]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[6]),
     .gwl_wr_25(gwl_wr_25[6]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_5_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[5]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[5]),
     .gwl_wr_25(gwl_wr_25[5]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_4_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[4]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[4]),
     .gwl_wr_25(gwl_wr_25[4]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[3]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[3]),
     .gwl_wr_25(gwl_wr_25[3]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[2]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[2]),
     .gwl_wr_25(gwl_wr_25[2]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[1]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[1]),
     .gwl_wr_25(gwl_wr_25[1]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[0]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25),
     .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[0]), .gwl_wr_25(gwl_wr_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_1f, View - schematic
// LAST TIME SAVED: Dec 30 14:56:08 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_gwlwr_1f ( gwl_b_25, gwp_hv, wr, gwl_b_sup_25, gwp_sup_hv,
     gnv_25, gnv_b_25, gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25,
     gwl_red_25, gwlb_dis_25, gwlb_en_25, s_25, vddp_tieh, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, wr_sup_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wr_sup_25;

output [26:0]  gwl_b_25;
output [107:0]  wr;
output [26:0]  gwp_hv;

input [3:0]  s_25;
input [1:0]  gred_25;
input [1:0]  gred_b_25;
input [5:0]  gnv_b_25;
input [5:0]  gnv_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [26:0]  gwl_wr_25;



ml_rock_lwldrv_wr_x108_1f Iml_rock_lwldrv_wr_x108_1f (
     .gwl_wr_25(gwl_wr_25[26:0]), .wr(wr[107:0]),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3:0]));
ml_gwl_drv_x27_1f Igwl_drv_x27 ( .gwp_hv(gwp_hv[26:0]),
     .gwl_wr_25(gwl_wr_25[26:0]), .gwl_b_25(gwl_b_25[26:0]),
     .gwlb_en_25(gwlb_en_25), .gwlb_dis_25(gwlb_dis_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25_1(gred_b_25[1]), .gred_b_25_0(gred_b_25[0]),
     .gred_25_1(gred_25[1]), .gred_25_0(gred_25[0]),
     .gnv5_b_25(gnv_b_25[5]), .gnv5_25(gnv_25[5]),
     .gnv4_b_25(gnv_b_25[4]), .gnv4_25(gnv_25[4]),
     .gnv3_b_25(gnv_b_25[3]), .gnv3_25(gnv_25[3]),
     .gnv2_b_25(gnv_b_25[2]), .gnv2_25(gnv_25[2]),
     .gnv1_b_25(gnv_b_25[1]), .gnv1_25(gnv_25[1]),
     .gnv0_b_25(gnv_b_25[0]), .gnv0_25(gnv_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_rdhv_inv, View - schematic
// LAST TIME SAVED: Jul 27 12:11:18 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_rdhv_inv ( s_rd_b_hv, srdsup_hv, s_rdin_hv, vddp_tieh );
output  s_rd_b_hv;

inout  srdsup_hv;

input  s_rdin_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M1 ( .D(rd_in_25), .B(GND_), .G(vddp_tieh), .S(s_rdin_hv));
pch_25  M0 ( .D(net12), .B(srdsup_hv), .G(s_rdin_hv), .S(srdsup_hv));
pch_25  M3 ( .D(s_rd_b_hv), .B(net12), .G(rd_in_25), .S(net12));
nch_25  M21 ( .D(s_rd_b_hv), .B(GND_), .G(vddp_tieh), .S(net19));
nch_25  M29 ( .D(net19), .B(GND_), .G(rd_in_25), .S(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_invx3_enhance, View - schematic
// LAST TIME SAVED: Oct  1 12:05:13 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_hv_invx3_enhance ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh
     );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));
pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));

endmodule
// Library - ice8chip, Cell - pllclkbuf_n40, View - schematic
// LAST TIME SAVED: Nov  2 13:03:26 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pllclkbuf_n40 ( gclk_l2clktv, gclk_r2clktv, padin_clkl_out,
     padin_clkr_out, pll_bypass, pll_cbit, pll_fb, pll_fse,
     pll_lock_out, pll_ref, pll_reset, pll_sdo, cbit, fabric_clkl_in,
     fabric_clkr_in, fo_bypass, fo_dlyadj, fo_fb, fo_ref, fo_reset,
     fo_sck, fo_sdi, icegate, padin_clkl_in, padin_clkr_in,
     pll_lock_in, pll_out, prog );
output  padin_clkl_out, padin_clkr_out, pll_bypass, pll_fb, pll_fse,
     pll_lock_out, pll_ref, pll_reset, pll_sdo;

input  fabric_clkl_in, fabric_clkr_in, fo_bypass, fo_fb, fo_ref,
     fo_reset, fo_sck, fo_sdi, icegate, padin_clkl_in, padin_clkr_in,
     pll_lock_in, pll_out, prog;

output [1:0]  gclk_l2clktv;
output [16:0]  pll_cbit;
output [1:0]  gclk_r2clktv;

input [7:0]  fo_dlyadj;
input [40:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



fabric_buf_ice8p I_GBUF_R_1_ ( .f_in(fabric_clkr_in),
     .f_out(gclk_r2clktv[1]));
fabric_buf_ice8p I_GBUF_R_0_ ( .f_in(padin_clkr_gate),
     .f_out(gclk_r2clktv[0]));
fabric_buf_ice8p I_GBUF_L_1_ ( .f_in(fabric_clkl_in),
     .f_out(gclk_l2clktv[1]));
fabric_buf_ice8p I_GBUF_L_0_ ( .f_in(padin_clkl_gate),
     .f_out(gclk_l2clktv[0]));
fabric_buf_ice8p I_buf4pll_lock ( .f_in(pll_lock_in),
     .f_out(pll_lock_out));
pllmate_40lp I_pllmate ( .pll_cbit(pll_cbit[16:0]), .cbit({cbit[40],
     cbit[35], cbit[34], cbit[33], cbit[32], cbit[31], cbit[30],
     cbit[29], cbit[28], cbit[27], cbit[26], cbit[25], cbit[24],
     cbit[23], cbit[22], cbit[21], cbit[20], cbit[19], cbit[18],
     cbit[17], cbit[16], cbit[15], cbit[14], cbit[13], cbit[12],
     cbit[11], cbit[10], cbit[9], cbit[8], cbit[7], cbit[6], cbit[5],
     cbit[4], cbit[3], cbit[2], cbit[1], cbit[0]}),
     .fo_dlyadj(fo_dlyadj[7:0]), .pll_out2(superpll_out2),
     .pll_out1(superpll_out1), .prog(prog), .pllout_in(pll_out),
     .pad_pllref(padin_clkl_in), .pll_bypass(pll_bypass),
     .fo_pllreset(fo_reset), .fo_pllref(fo_ref), .fo_pllfb(fo_fb),
     .pll_sdo(pll_sdo), .pll_reset(pll_reset), .pll_ref(pll_ref),
     .pll_fse(pll_fse), .pll_fb(pll_fb), .fo_pll_sck(fo_sck),
     .fo_pll_sdi(fo_sdi), .fo_pll_bypass(fo_bypass));
clkmux2buffer I_PadPLLMux_R ( .in1(superpll_out2), .in0(padin_clkr_in),
     .out(padin_clkr_out), .sel(cbit[38]));
clkmux2buffer I_PadPLLMux_L ( .in1(superpll_out1), .in0(padin_clkl_in),
     .out(padin_clkl_out), .sel(cbit[36]));
pinlatbuf12p I_GBUF_CLKGAT_L ( .pad_in(padin_clkl_out),
     .icegate(icegate), .cbit(cbit[37]), .cout(padin_clkl_gate),
     .prog(prog));
pinlatbuf12p I_GBUF_CLKGAT_R ( .pad_in(padin_clkr_out),
     .icegate(icegate), .cbit(cbit[39]), .cout(padin_clkr_gate),
     .prog(prog));

endmodule
// Library - NVCM_40nm, Cell - ml_lshv_6v_switch_enhance, View -
//schematic
// LAST TIME SAVED: Oct  1 12:06:46 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_lshv_6v_switch_enhance ( out_b_hv, out_hv, in_hv, sel_25,
     sel_b_25, vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M0 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
pch_25  M1 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_hotsw_enhance, View -
//schematic
// LAST TIME SAVED: Jun 30 18:50:37 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw_enhance ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3_enhance Ihv_invx3 ( .vddp_tieh(vddp_tieh),
     .out_b_hv(out_b_hv), .sel_25(sel_25), .in_hv(in_hv),
     .sel_hv(sel_hv));
ml_lshv_6v_switch_enhance Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_hotswitch_enhance, View -
//schematic
// LAST TIME SAVED: Sep  8 10:25:27 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_hv_hotswitch_enhance ( hv_in_hv, hv_out_hv, selhv_25,
     vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net042));
nch_25  M2 ( .D(net031), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
nch_25  M4 ( .D(net031), .B(GND_), .G(selhv_25), .S(net042));
inv_25 I112 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M6 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_hotswitch_enhance, View -
//schematic
// LAST TIME SAVED: Apr 30 11:28:27 2008
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch_enhance ( hvin_a_hv, hvin_b_hv, out_hv,
     sel_hv_a_25, sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch_enhance Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tiehigh, View - schematic
// LAST TIME SAVED: May 13 15:28:20 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module vdd_tiehigh ( vdd_tieh );
inout  vdd_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(vdd_tieh), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_logic, View - schematic
// LAST TIME SAVED: Sep 14 11:51:05 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_logic ( gnv, gred, gwl_misc, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, s, sa_trim, saen, testdec_en_b, testdec_even_b,
     testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd, fsm_coladd, fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rprd, fsm_tm_trow,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr );
output  gwl_misc, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, saen, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [3:0]  s;
output [2:0]  sa_trim;
output [5:0]  gnv;
output [1:0]  gred;

input [2:0]  fsm_trim_rrefpgm;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [0:0]  fsm_coladd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  net390;

wire  [3:0]  s_b;

wire  [5:0]  gnv_b;

wire  [2:0]  sa_trim_b;

wire  [1:0]  xadd_b;

wire  [1:0]  gred_b;

wire  [1:0]  xadd;

wire  [1:0]  net386;



anor21_hvt I109_1_ ( .A(net386[0]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I109_0_ ( .A(net386[1]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
nor4_hvt I287 ( .B(fsm_nvcmen_b), .Y(net216), .D(testdec_wp),
     .A(fsm_wren_b), .C(net331));
nor4_hvt I286 ( .B(fsm_pgmvfy), .Y(net211), .D(fsm_tm_allwl_h),
     .A(fsm_pgmvfy), .C(fsm_rd));
nor4_hvt I282 ( .B(fsm_tm_allbl_l), .Y(net0258), .D(net282),
     .A(fsm_tm_allbl_l), .C(fsm_nvcmen_b));
nor4_hvt I284 ( .B(pgm_hvpulse), .Y(wrsup_2vdd), .D(fsm_nvcmen_b),
     .A(pgm_hvpulse), .C(testdec_wr));
nor4_hvt I285 ( .B(fsm_nvcmen_b), .Y(net226), .D(fsm_wpen_b),
     .A(testdec_wr), .C(fsm_tm_allwl_l));
nand2_hvt I302 ( .A(net0341), .Y(net307), .B(tm_testdec));
nand2_hvt I297 ( .A(tm_testdec_wr), .Y(testwr_wpgnd_b),
     .B(tm_testdec));
nand2_hvt I269 ( .A(net355), .Y(testdec_even_b), .B(testdec_en));
nand2_hvt I268 ( .A(testdec_en), .Y(testdec_odd_b), .B(fsm_coladd[0]));
nand2_hvt I267 ( .A(fsm_rd), .Y(net0266), .B(tm_testdec));
nand3_hvt I298 ( .Y(net282), .B(net341), .C(fsm_lshven), .A(fsm_pgm));
nand3_hvt I299 ( .Y(net0278), .B(fsm_rd), .C(fsm_ymuxdis),
     .A(tm_testdec));
nand3_hvt I293 ( .Y(net286), .B(fsm_pgm), .C(fsm_tm_allwl_h),
     .A(fsm_wren));
nand3_hvt I288 ( .Y(net274), .B(fsm_tm_allwl_h), .C(fsm_tm_allwl_h),
     .A(stress2));
nand3_hvt I292 ( .Y(net292), .B(tm_allwl_l_b), .C(net307),
     .A(fsm_nvcmen));
nand3_hvt I303 ( .Y(gwlb_dis), .B(fsm_nvcmen), .C(testwr_wpgnd_b),
     .A(net0332));
inv_hvt I307_5_ ( .A(fsm_rowadd[7]), .Y(gnv_b[5]));
inv_hvt I307_4_ ( .A(fsm_rowadd[6]), .Y(gnv_b[4]));
inv_hvt I307_3_ ( .A(fsm_rowadd[5]), .Y(gnv_b[3]));
inv_hvt I307_2_ ( .A(fsm_rowadd[4]), .Y(gnv_b[2]));
inv_hvt I307_1_ ( .A(fsm_rowadd[3]), .Y(gnv_b[1]));
inv_hvt I307_0_ ( .A(fsm_rowadd[2]), .Y(gnv_b[0]));
inv_hvt I238 ( .A(net0274), .Y(gwl_misc));
inv_hvt I234 ( .A(testdec_en), .Y(testdec_en_b));
inv_hvt I240 ( .A(gwlbsup_vddp), .Y(net202));
inv_hvt I236 ( .A(net0300), .Y(testdec_prec_b));
inv_hvt I305_1_ ( .A(gred_b[1]), .Y(gred[1]));
inv_hvt I305_0_ ( .A(gred_b[0]), .Y(gred[0]));
inv_hvt I314_2_ ( .A(sa_trim_b[2]), .Y(sa_trim[2]));
inv_hvt I314_1_ ( .A(sa_trim_b[1]), .Y(sa_trim[1]));
inv_hvt I314_0_ ( .A(sa_trim_b[0]), .Y(sa_trim[0]));
inv_hvt I315_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I315_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I306_5_ ( .A(gnv_b[5]), .Y(gnv[5]));
inv_hvt I306_4_ ( .A(gnv_b[4]), .Y(gnv[4]));
inv_hvt I306_3_ ( .A(gnv_b[3]), .Y(gnv[3]));
inv_hvt I306_2_ ( .A(gnv_b[2]), .Y(gnv[2]));
inv_hvt I306_1_ ( .A(gnv_b[1]), .Y(gnv[1]));
inv_hvt I306_0_ ( .A(gnv_b[0]), .Y(gnv[0]));
inv_hvt I261 ( .A(pgm_hvpulse), .Y(net0390));
inv_hvt I291 ( .A(net0428), .Y(net331));
inv_hvt I263 ( .A(net282), .Y(pgm_hvpulse));
inv_hvt I250 ( .A(fsm_coladd[0]), .Y(net355));
inv_hvt I255 ( .A(net307), .Y(testdec_wp));
inv_hvt I248 ( .A(net246), .Y(net359));
inv_hvt I252 ( .A(fsm_wren), .Y(fsm_wren_b));
inv_hvt I241 ( .A(gwlbsup_vpxa), .Y(net204));
inv_hvt I244 ( .A(net0278), .Y(net0300));
inv_hvt I264 ( .A(fsm_pgmvfy), .Y(net341));
inv_hvt I246_2_ ( .A(net390[0]), .Y(sa_trim_b[2]));
inv_hvt I246_1_ ( .A(net390[1]), .Y(sa_trim_b[1]));
inv_hvt I246_0_ ( .A(net390[2]), .Y(sa_trim_b[0]));
inv_hvt I254 ( .A(net292), .Y(net365));
inv_hvt I242 ( .A(gwphv_vddp), .Y(net206));
inv_hvt I249 ( .A(net0266), .Y(testdec_en));
inv_hvt I266 ( .A(net0388), .Y(net0327));
inv_hvt I243 ( .A(gwphv_vppint), .Y(net200));
inv_hvt I256 ( .A(net286), .Y(net0343));
inv_hvt I258 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I257 ( .A(tm_testdec_wr), .Y(net0341));
inv_hvt I259 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I304_1_ ( .A(fsm_rowadd[3]), .Y(gred_b[1]));
inv_hvt I304_0_ ( .A(fsm_rowadd[2]), .Y(gred_b[0]));
inv_hvt I253 ( .A(net196), .Y(net351));
inv_hvt I251 ( .A(fsm_wpen), .Y(fsm_wpen_b));
inv_hvt I262 ( .A(fsm_pgm), .Y(fsm_pgm_b));
inv_hvt I309 ( .A(net211), .Y(wp_frcen));
inv_hvt I310 ( .A(net216), .Y(wr_dis));
inv_hvt I308 ( .A(net226), .Y(wp_dis));
inv_hvt I311 ( .A(net274), .Y(wr_frcen));
inv_hvt I312 ( .A(testwr_wpgnd_b), .Y(testdec_wr));
inv_hvt I147_3_ ( .A(s_b[3]), .Y(s[3]));
inv_hvt I147_2_ ( .A(s_b[2]), .Y(s[2]));
inv_hvt I147_1_ ( .A(s_b[1]), .Y(s[1]));
inv_hvt I147_0_ ( .A(s_b[0]), .Y(s[0]));
nor2_hvt I272 ( .A(net0258), .B(tm_testdec), .Y(pgminhi_dmmy_b));
nor2_hvt I279 ( .A(fsm_pgm), .B(fsm_pgmvfy), .Y(net0388));
nor2_hvt I313 ( .A(net0288), .B(net0390), .Y(gwlb_en));
nor2_hvt I274 ( .A(net359), .B(net201), .Y(gwphv_vddp));
nor2_hvt I273 ( .A(fsm_nvcmen_b), .B(tm_dma), .Y(saen));
nor2_hvt I278 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I300 ( .A(fsm_pgmdisc), .B(fsm_pgmhv), .Y(net0231));
nor2_hvt I316 ( .A(net207), .B(net246), .Y(gwphv_vppint));
nor2_hvt I275 ( .A(net0232), .B(fsm_nvcmen_b), .Y(net246));
nor2_hvt I276 ( .A(net203), .B(net351), .Y(gwlbsup_vpxa));
nor2_hvt I296 ( .A(fsm_pgmvfy), .B(fsm_pgm_b), .Y(stress2));
nor2_hvt I277 ( .A(net196), .B(net205), .Y(gwlbsup_vddp));
nor3_hvt I290 ( .B(fsm_tm_allwl_l), .Y(net0428), .A(fsm_tm_allwl_l),
     .C(fsm_tm_allwl_l));
nor3_hvt I324 ( .B(fsm_tm_allwl_h), .Y(net0288), .A(fsm_tm_allwl_h),
     .C(fsm_tm_allwl_h));
nor3_hvt I295 ( .B(fsm_tm_trow), .Y(net0274), .A(fsm_nv_rri_trim),
     .C(fsm_nv_sisi_ui));
nor3_hvt I294 ( .B(fsm_tm_rprd), .Y(net196), .A(fsm_tm_rprd),
     .C(fsm_tm_rprd));
mux2_hvt I180_1_ ( .in1(fsm_rowadd[1]), .in0(fsm_rowadd[1]),
     .out(net386[0]), .sel(fsm_nv_rrow));
mux2_hvt I180_0_ ( .in1(fsm_rowadd[0]), .in0(fsm_rowadd[0]),
     .out(net386[1]), .sel(fsm_nv_rrow));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net390[0]), .sel(net0327));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net390[1]), .sel(net0327));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net390[2]), .sel(net0327));
mux2_hvt I221 ( .in1(fsm_wpen), .in0(fsm_wgnden), .out(net0332),
     .sel(pgm_hvpulse));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_pump_a_clkdly I230 ( .in(net0231), .out(net0232));
ml_pump_a_clkdly I208 ( .in(net200), .out(net201));
ml_pump_a_clkdly I202 ( .in(net202), .out(net203));
ml_pump_a_clkdly I198 ( .in(net204), .out(net205));
ml_pump_a_clkdly I207 ( .in(net206), .out(net207));
anor31_hvt I121_3_ ( .A(net365), .D(net0343), .B(xadd[1]), .Y(s_b[3]),
     .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net365), .D(net0343), .B(xadd[1]), .Y(s_b[2]),
     .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net365), .D(net0343), .B(xadd_b[1]),
     .Y(s_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net365), .D(net0343), .B(xadd_b[1]),
     .Y(s_b[0]), .C(xadd_b[0]));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_invx3, View - schematic
// LAST TIME SAVED: Jul 29 12:21:23 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_hv_invx3 ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));
pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_lshv_6v_switch, View - schematic
// LAST TIME SAVED: Jul 29 12:23:54 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_lshv_6v_switch ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M3 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M0 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_ls_inv_hotsw, View - schematic
// LAST TIME SAVED: Jul  1 14:28:58 2010
// NETLIST TIME: May  5 11:56:45 2011
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3 Ihv_invx3 ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));
ml_lshv_6v_switch Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_hv_hotswitch, View - schematic
// LAST TIME SAVED: Sep 10 14:28:35 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hv_hotswitch ( hv_in_hv, hv_out_hv, selhv_25, vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M3 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
nch_25  M4 ( .D(net15), .B(GND_), .G(selhv_25), .S(net12));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - ice1chip, Cell - pll_wrapbuf_ice1f, View - schematic
// LAST TIME SAVED: May  3 11:46:09 2011
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pll_wrapbuf_ice1f ( gclk_l2clktv[1:0], gclk_r2clktv[1:0],
     padin_clkl_out, padin_clkr_out, pll_bypass, pll_cbit[16:0],
     pll_fb, pll_fse, pll_lock_out, pll_ref, pll_reset, pll_sdo,
     cf_bbank[159], cf_bbank[135], cf_lbank[9:1], cf_lbank[33:25],
     cf_lbank[57:49], cf_lbank[81:73], cf_lbank[97], cf_lbank[99],
     cf_lbank[101], fabric_clkl_in, fabric_clkr_in, fo_bypass,
     fo_dlyadj[7:0], fo_fb, fo_ref, fo_reset, fo_sck, fo_sdi, icegate,
     padin_clkl_in, padin_clkr_in, pll_lock_in, pll_out, prog );
output  padin_clkl_out, padin_clkr_out, pll_bypass, pll_fb, pll_fse,
     pll_lock_out, pll_ref, pll_reset, pll_sdo;

input  fabric_clkl_in, fabric_clkr_in, fo_bypass, fo_fb, fo_ref,
     fo_reset, fo_sck, fo_sdi, icegate, padin_clkl_in, padin_clkr_in,
     pll_lock_in, pll_out, prog;

output [1:0]  gclk_r2clktv;
output [16:0]  pll_cbit;
output [1:0]  gclk_l2clktv;

input [7:0]  fo_dlyadj;
input [101:1]  cf_lbank;
input [159:135]  cf_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [40:0]  cbit;

wire  [1:0]  net129;

wire  [1:0]  net88;

wire  [1:0]  net82;

wire  [1:0]  net130;



pll_bufwrap_ice1f I8_1_ ( .f_in(net130[0]), .f_out(net82[0]));
pll_bufwrap_ice1f I8_0_ ( .f_in(net130[1]), .f_out(net82[1]));
pll_bufwrap_ice1f I15 ( .f_in(net145), .f_out(padin_clkr_out));
pll_bufwrap_ice1f I12_1_ ( .f_in(net88[0]), .f_out(gclk_l2clktv[1]));
pll_bufwrap_ice1f I12_0_ ( .f_in(net88[1]), .f_out(gclk_l2clktv[0]));
pll_bufwrap_ice1f I9_1_ ( .f_in(net129[0]), .f_out(net88[0]));
pll_bufwrap_ice1f I9_0_ ( .f_in(net129[1]), .f_out(net88[1]));
pll_bufwrap_ice1f I10 ( .f_in(fabric_clkl_in), .f_out(net142));
pll_bufwrap_ice1f I14 ( .f_in(net144), .f_out(padin_clkl_out));
pll_bufwrap_ice1f I11 ( .f_in(fabric_clkr_in), .f_out(net143));
pll_bufwrap_ice1f I13_1_ ( .f_in(net82[0]), .f_out(gclk_r2clktv[1]));
pll_bufwrap_ice1f I13_0_ ( .f_in(net82[1]), .f_out(gclk_r2clktv[0]));
pll_bufwrap_ice1f I16 ( .f_in(padin_clkl_in), .f_out(net124));
pll_bufwrap_ice1f I17 ( .f_in(padin_clkr_in), .f_out(net125));
bram_bufferx4 I25_39_ ( .in(cf_bbank[159]), .out(cbit[39]));
bram_bufferx4 I4_40_ ( .in(cf_lbank[101]), .out(cbit[40]));
bram_bufferx4 I4_26_ ( .in(cf_lbank[57]), .out(cbit[26]));
bram_bufferx4 I4_25_ ( .in(cf_lbank[56]), .out(cbit[25]));
bram_bufferx4 I4_24_ ( .in(cf_lbank[55]), .out(cbit[24]));
bram_bufferx4 I4_23_ ( .in(cf_lbank[54]), .out(cbit[23]));
bram_bufferx4 I4_22_ ( .in(cf_lbank[53]), .out(cbit[22]));
bram_bufferx4 I4_21_ ( .in(cf_lbank[52]), .out(cbit[21]));
bram_bufferx4 I4_20_ ( .in(cf_lbank[51]), .out(cbit[20]));
bram_bufferx4 I4_19_ ( .in(cf_lbank[50]), .out(cbit[19]));
bram_bufferx4 I4_18_ ( .in(cf_lbank[49]), .out(cbit[18]));
bram_bufferx4 I4_8_ ( .in(cf_lbank[9]), .out(cbit[8]));
bram_bufferx4 I4_7_ ( .in(cf_lbank[8]), .out(cbit[7]));
bram_bufferx4 I4_6_ ( .in(cf_lbank[7]), .out(cbit[6]));
bram_bufferx4 I4_5_ ( .in(cf_lbank[6]), .out(cbit[5]));
bram_bufferx4 I4_4_ ( .in(cf_lbank[5]), .out(cbit[4]));
bram_bufferx4 I4_3_ ( .in(cf_lbank[4]), .out(cbit[3]));
bram_bufferx4 I4_2_ ( .in(cf_lbank[3]), .out(cbit[2]));
bram_bufferx4 I4_1_ ( .in(cf_lbank[2]), .out(cbit[1]));
bram_bufferx4 I4_0_ ( .in(cf_lbank[1]), .out(cbit[0]));
bram_bufferx4 I4_36_ ( .in(cf_lbank[97]), .out(cbit[36]));
bram_bufferx4 I4_35_ ( .in(cf_lbank[81]), .out(cbit[35]));
bram_bufferx4 I4_34_ ( .in(cf_lbank[80]), .out(cbit[34]));
bram_bufferx4 I4_33_ ( .in(cf_lbank[79]), .out(cbit[33]));
bram_bufferx4 I4_32_ ( .in(cf_lbank[78]), .out(cbit[32]));
bram_bufferx4 I4_31_ ( .in(cf_lbank[77]), .out(cbit[31]));
bram_bufferx4 I4_30_ ( .in(cf_lbank[76]), .out(cbit[30]));
bram_bufferx4 I4_29_ ( .in(cf_lbank[75]), .out(cbit[29]));
bram_bufferx4 I4_28_ ( .in(cf_lbank[74]), .out(cbit[28]));
bram_bufferx4 I4_27_ ( .in(cf_lbank[73]), .out(cbit[27]));
bram_bufferx4 I4_38_ ( .in(cf_lbank[99]), .out(cbit[38]));
bram_bufferx4 I4_37_ ( .in(cf_bbank[135]), .out(cbit[37]));
bram_bufferx4 I4_17_ ( .in(cf_lbank[33]), .out(cbit[17]));
bram_bufferx4 I4_16_ ( .in(cf_lbank[32]), .out(cbit[16]));
bram_bufferx4 I4_15_ ( .in(cf_lbank[31]), .out(cbit[15]));
bram_bufferx4 I4_14_ ( .in(cf_lbank[30]), .out(cbit[14]));
bram_bufferx4 I4_13_ ( .in(cf_lbank[29]), .out(cbit[13]));
bram_bufferx4 I4_12_ ( .in(cf_lbank[28]), .out(cbit[12]));
bram_bufferx4 I4_11_ ( .in(cf_lbank[27]), .out(cbit[11]));
bram_bufferx4 I4_10_ ( .in(cf_lbank[26]), .out(cbit[10]));
bram_bufferx4 I4_9_ ( .in(cf_lbank[25]), .out(cbit[9]));
pllclkbuf_n40 I_pllclkbuf_cbuf_bot8p ( .fo_ref(fo_ref),
     .fo_sck(fo_sck), .fo_sdi(fo_sdi), .padin_clkl_in(net124),
     .padin_clkr_in(net125), .pll_lock_in(pll_lock_in),
     .pll_out(pll_out), .prog(prog), .gclk_l2clktv({net129[0],
     net129[1]}), .gclk_r2clktv({net130[0], net130[1]}),
     .pll_bypass(pll_bypass), .pll_cbit(pll_cbit[16:0]),
     .pll_fb(pll_fb), .pll_fse(pll_fse), .pll_lock_out(pll_lock_out),
     .pll_ref(pll_ref), .pll_reset(pll_reset), .pll_sdo(pll_sdo),
     .fo_bypass(fo_bypass), .fo_dlyadj(fo_dlyadj[7:0]), .fo_fb(fo_fb),
     .fabric_clkl_in(net142), .fabric_clkr_in(net143),
     .padin_clkl_out(net144), .padin_clkr_out(net145),
     .icegate(icegate), .fo_reset(fo_reset), .cbit(cbit[40:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_hotswitch, View - schematic
// LAST TIME SAVED: Jan 26 19:35:53 2008
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch ( hvin_a_hv, hvin_b_hv, out_hv, sel_hv_a_25,
     sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_bldrv, View - schematic
// LAST TIME SAVED: Nov 17 19:02:34 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_gwlwr_bldrv ( bgr, bl_pgm_glb, bl_frc_gnd, fsm_din, fsm_pgm,
     fsm_pgmien, fsm_trim_ipp, tm_dma );
inout  bgr, bl_pgm_glb;

input  bl_frc_gnd, fsm_din, fsm_pgm, fsm_pgmien, tm_dma;

input [3:0]  fsm_trim_ipp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net0115;

wire  [7:0]  net0152;

wire  [1:0]  net0160;

wire  [1:0]  net0180;

wire  [3:0]  net0172;

wire  [3:0]  net0156;



rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(gnd_), .PLUS(net0141), .BULK(GND_));
nch_25  M20 ( .D(net0173), .B(GND_), .G(pgm_inhi_bias),
     .S(bl_pgm_glb));
nch_25  M21 ( .D(pgm_inhi_bias), .B(GND_), .G(pgm_inhi_bias),
     .S(gnd_));
nch_25  M12_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[0]));
nch_25  M12_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[1]));
nch_25  M13_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[0]));
nch_25  M13_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[1]));
nch_25  M13_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[2]));
nch_25  M13_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[3]));
nch_25  M6 ( .D(net0164), .B(GND_), .G(net0164), .S(gnd_));
nch_25  M3 ( .D(dec_bias_p), .B(GND_), .G(bgr), .S(net0141));
nch_25  M10 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net089));
nch_25  M18_7_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[0]));
nch_25  M18_6_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[1]));
nch_25  M18_5_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[2]));
nch_25  M18_4_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[3]));
nch_25  M18_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[4]));
nch_25  M18_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[5]));
nch_25  M18_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[6]));
nch_25  M18_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[7]));
nch_25  M9 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net0135));
nch_25  M8 ( .D(net0164), .B(GND_), .G(pgmen_b_25), .S(gnd_));
nch_hvt  M36 ( .D(net0173), .B(GND_), .G(pgm_trim0_en), .S(net0107));
nch_hvt  M37 ( .D(net0107), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M31_7_ ( .D(net0115[0]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[0]));
nch_hvt  M31_6_ ( .D(net0115[1]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[1]));
nch_hvt  M31_5_ ( .D(net0115[2]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[2]));
nch_hvt  M31_4_ ( .D(net0115[3]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[3]));
nch_hvt  M31_3_ ( .D(net0115[4]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[4]));
nch_hvt  M31_2_ ( .D(net0115[5]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[5]));
nch_hvt  M31_1_ ( .D(net0115[6]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[6]));
nch_hvt  M31_0_ ( .D(net0115[7]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[7]));
nch_hvt  M19 ( .D(net0135), .B(GND_), .G(fsm_trim_ipp[0]),
     .S(net0131));
nch_hvt  M38_7_ ( .D(net0152[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_6_ ( .D(net0152[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_5_ ( .D(net0152[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_4_ ( .D(net0152[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_3_ ( .D(net0152[4]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_2_ ( .D(net0152[5]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_1_ ( .D(net0152[6]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_0_ ( .D(net0152[7]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_3_ ( .D(net0156[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_2_ ( .D(net0156[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_1_ ( .D(net0156[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_0_ ( .D(net0156[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_1_ ( .D(net0160[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_0_ ( .D(net0160[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M26 ( .D(net0131), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M33 ( .D(bl_pgm_glb), .B(GND_), .G(net0187), .S(gnd_));
nch_hvt  M30_3_ ( .D(net0172[0]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[0]));
nch_hvt  M30_2_ ( .D(net0172[1]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[1]));
nch_hvt  M30_1_ ( .D(net0172[2]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[2]));
nch_hvt  M30_0_ ( .D(net0172[3]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[3]));
nch_hvt  M34 ( .D(net089), .B(GND_), .G(pgm_trim0_en), .S(gnd_));
nch_hvt  M27_1_ ( .D(net0180[0]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[0]));
nch_hvt  M27_0_ ( .D(net0180[1]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[1]));
pch_25  M11 ( .D(pgm_inhi_bias), .B(vddp_), .G(vdd_tieh), .S(net0259));
pch_25  M14_1_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M14_0_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M5 ( .D(net0164), .B(vddp_), .G(dec_bias_p), .S(net0241));
pch_25  M7_1_ ( .D(net0241), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M7_0_ ( .D(net0241), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M4 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p), .S(net0241));
nor2_hvt I121 ( .A(net086), .B(fsm_pgmien_b_buf), .Y(pgm_trim0_en));
nor2_hvt I114 ( .B(tm_dma), .Y(net0116), .A(tm_dma));
nor4_hvt I105 ( .D(fsm_trim_ipp[0]), .B(fsm_trim_ipp[2]), .Y(net086),
     .A(fsm_trim_ipp[3]), .C(fsm_trim_ipp[1]));
nand2_hvt I71 ( .B(fsm_din), .A(fsm_pgmien), .Y(fsm_pgmien_b_buf));
inv_hvt I115 ( .A(net0116), .Y(net0187));
inv_hvt I58 ( .A(pgmen_b), .Y(pgmen));
inv_hvt I131 ( .A(fsm_pgm), .Y(pgmen_b));
inv_hvt I72 ( .A(fsm_pgmien_b_buf), .Y(fsm_pgmien_buf));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_ls_vdd2vdd25 I56 ( .in(pgmen), .sup(vddp_),
     .out_vddio_b(pgmen_b_25), .out_vddio(pgmen_25), .in_b(pgmen_b));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_wr_sup, View - schematic
// LAST TIME SAVED: Aug 10 11:01:54 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_wr_sup ( wr_sup_25, wrsup_2vdd, wrsup_2vdd_25 );
inout  wr_sup_25;

input  wrsup_2vdd, wrsup_2vdd_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_25  M5 ( .D(net17), .B(vddp_), .G(wrsup_2vdd_25), .S(vddp_));
pch_25  M0 ( .D(net17), .B(wr_sup_25), .G(wrsup_2vdd), .S(wr_sup_25));
nch_na25  M13 ( .D(vdd_), .B(GND_), .G(wrsup_2vdd_25), .S(wr_sup_25));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_ls25_1b, View - schematic
// LAST TIME SAVED: Oct  1 12:09:28 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25_1b ( out_25, in );
output  out_25;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I145 ( .A(in), .Y(net45));
inv_25 I153 ( .IN(out_b_25), .OUT(out_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I112 ( .in(in), .sup(vddp_), .out_vddio_b(out_b_25),
     .out_vddio(net025), .in_b(net45));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl_ls25, View - schematic
// LAST TIME SAVED: Sep  7 15:15:51 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25 ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25,
     gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25, s_25,
     testdec_even_b_25, testdec_odd_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, wrsup_2vdd_25, fsm_gwlbdis, gnv, gred,
     gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en, gwlbsup_vddp,
     gwlbsup_vpxa, gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, s,
     testdec_even_b, testdec_odd_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25,
     testdec_even_b_25, testdec_odd_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, wrsup_2vdd_25;

input  fsm_gwlbdis, gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, testdec_even_b, testdec_odd_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

output [5:0]  gnv_b_25;
output [3:0]  s_25;
output [5:0]  gnv_25;
output [1:0]  gred_25;
output [1:0]  gred_b_25;

input [5:0]  gnv;
input [3:0]  s;
input [1:0]  gred;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I_1_ ( .IN(gred_25[1]), .OUT(gred_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I_0_ ( .IN(gred_25[0]), .OUT(gred_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_5_ ( .IN(gnv_25[5]), .OUT(gnv_b_25[5]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_4_ ( .IN(gnv_25[4]), .OUT(gnv_b_25[4]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_3_ ( .IN(gnv_25[3]), .OUT(gnv_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_2_ ( .IN(gnv_25[2]), .OUT(gnv_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_1_ ( .IN(gnv_25[1]), .OUT(gnv_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I145_0_ ( .IN(gnv_25[0]), .OUT(gnv_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I143 ( .IN(net101), .OUT(fsm_gwlbdis_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_gwlwr_ctrl_ls25_1b I139 ( .in(gwlb_dis), .out_25(gwlb_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_frcen ( .in(wr_frcen),
     .out_25(wr_frcen_25));
ml_gwlwr_ctrl_ls25_1b I144 ( .in(gwlb_en), .out_25(gwlb_en_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vpp ( .in(gwphv_vppint),
     .out_25(gwphv_vppint_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwlb_vddp ( .in(gwlbsup_vddp),
     .out_25(gwlbsup_vddp_25));
ml_gwlwr_ctrl_ls25_1b ls25_gwlb_vpp ( .in(gwlbsup_vpxa),
     .out_25(gwlbsup_vpxa_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_vdd ( .in(wrsup_2vdd),
     .out_25(wrsup_2vdd_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_dis ( .in(wr_dis), .out_25(wr_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vddp ( .in(gwphv_vddp),
     .out_25(gwphv_vddp_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_frcen ( .in(wp_frcen),
     .out_25(wp_frcen_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_dis ( .in(wp_dis), .out_25(wp_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwl_red ( .in(gwl_red),
     .out_25(gwl_red_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_nvcm ( .in(gwl_nvcm),
     .out_25(gwl_nvcm_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_misc ( .in(gwl_misc),
     .out_25(gwl_misc_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_1_ ( .in(gred[1]),
     .out_25(gred_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_0_ ( .in(gred[0]),
     .out_25(gred_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_5_ ( .in(gnv[5]), .out_25(gnv_25[5]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_4_ ( .in(gnv[4]), .out_25(gnv_25[4]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_3_ ( .in(gnv[3]), .out_25(gnv_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_2_ ( .in(gnv[2]), .out_25(gnv_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_1_ ( .in(gnv[1]), .out_25(gnv_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_0_ ( .in(gnv[0]), .out_25(gnv_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_3_ ( .in(s[3]), .out_25(s_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_2_ ( .in(s[2]), .out_25(s_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_1_ ( .in(s[1]), .out_25(s_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_0_ ( .in(s[0]), .out_25(s_25[0]));
ml_gwlwr_ctrl_ls25_1b I136 ( .in(pgminhi_dmmy_b),
     .out_25(pgminhi_dmmy_b_25));
ml_gwlwr_ctrl_ls25_1b I140 ( .in(fsm_gwlbdis), .out_25(net101));
ml_gwlwr_ctrl_ls25_1b I137 ( .in(testdec_even_b),
     .out_25(testdec_even_b_25));
ml_gwlwr_ctrl_ls25_1b I138 ( .in(testdec_odd_b),
     .out_25(testdec_odd_b_25));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_npgate_gen, View - schematic
// LAST TIME SAVED: Sep  2 17:11:20 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_core_sa_npgate_gen ( sa_ngate, saen_25, saen_b_vpxa,
     saprd_b_vpxa, sdiode_en_vpxa, vpxa, fsm_tm_rprd, fsm_tm_sdiode,
     fsm_tm_testdec, saen, satrim, vddp_tieh );
output  saen_25, saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa;

inout  vpxa;

input  fsm_tm_rprd, fsm_tm_sdiode, fsm_tm_testdec, saen, vddp_tieh;

output [4:1]  sa_ngate;

input [2:0]  satrim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  ydec_b;

wire  [2:0]  ydec;

wire  [4:1]  trim;

wire  [7:0]  dec_trim;

wire  [7:0]  dec_trim_b;

wire  [3:0]  net48;



nand2_hvt I183 ( .Y(net037), .B(fsm_tm_rprd), .A(net078));
inv_25 I149 ( .IN(net052), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nor4_hvt I102 ( .D(fsm_tm_testdec), .C(dec_trim[7]), .A(dec_trim[5]),
     .B(dec_trim[6]), .Y(net47));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_4_ ( .Y(dec_trim_b[4]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_3_ ( .Y(dec_trim_b[3]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_2_ ( .Y(dec_trim_b[2]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nand3_hvt I37_1_ ( .Y(dec_trim_b[1]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_0_ ( .Y(dec_trim_b[0]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nor2_hvt I75_4_ ( .Y(net48[0]), .B(dec_trim[4]), .A(sa_high_res));
nor2_hvt I75_3_ ( .Y(net48[1]), .B(dec_trim[3]), .A(trim[4]));
nor2_hvt I75_2_ ( .Y(net48[2]), .B(dec_trim[2]), .A(trim[3]));
nor2_hvt I75_1_ ( .Y(net48[3]), .B(dec_trim[1]), .A(trim[2]));
inv_hvt I158_2_ ( .A(satrim[2]), .Y(ydec_b[2]));
inv_hvt I158_1_ ( .A(satrim[1]), .Y(ydec_b[1]));
inv_hvt I158_0_ ( .A(satrim[0]), .Y(ydec_b[0]));
inv_hvt I160_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I160_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I160_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I160_4_ ( .A(dec_trim_b[4]), .Y(dec_trim[4]));
inv_hvt I160_3_ ( .A(dec_trim_b[3]), .Y(dec_trim[3]));
inv_hvt I160_2_ ( .A(dec_trim_b[2]), .Y(dec_trim[2]));
inv_hvt I160_1_ ( .A(dec_trim_b[1]), .Y(dec_trim[1]));
inv_hvt I160_0_ ( .A(dec_trim_b[0]), .Y(dec_trim[0]));
inv_hvt I163 ( .A(net078), .Y(net080));
inv_hvt I162 ( .A(net076), .Y(net078));
inv_hvt I165 ( .A(net073), .Y(net071));
inv_hvt I166 ( .A(net075), .Y(net073));
inv_hvt I167 ( .A(fsm_tm_sdiode), .Y(net075));
inv_hvt I175 ( .A(net059), .Y(net061));
inv_hvt I176 ( .A(net037), .Y(net059));
inv_hvt I114 ( .A(net47), .Y(sa_high_res));
inv_hvt I161 ( .A(saen), .Y(net076));
inv_hvt I159_2_ ( .A(ydec_b[2]), .Y(ydec[2]));
inv_hvt I159_1_ ( .A(ydec_b[1]), .Y(ydec[1]));
inv_hvt I159_0_ ( .A(ydec_b[0]), .Y(ydec[0]));
inv_hvt I76_4_ ( .A(net48[0]), .Y(trim[4]));
inv_hvt I76_3_ ( .A(net48[1]), .Y(trim[3]));
inv_hvt I76_2_ ( .A(net48[2]), .Y(trim[2]));
inv_hvt I76_1_ ( .A(net48[3]), .Y(trim[1]));
inv_hvt I78_4_ ( .A(trim[4]), .Y(sa_ngate[4]));
inv_hvt I78_3_ ( .A(trim[3]), .Y(sa_ngate[3]));
inv_hvt I78_2_ ( .A(trim[2]), .Y(sa_ngate[2]));
inv_hvt I78_1_ ( .A(trim[1]), .Y(sa_ngate[1]));
ml_hv_invx3 I135 ( .sel_hv(net048), .sel_25(net048),
     .vddp_tieh(vddp_tieh), .out_b_hv(saen_b_vpxa), .in_hv(vpxa));
ml_hv_invx3 I168 ( .sel_hv(net0123), .sel_25(net0123),
     .vddp_tieh(vddp_tieh), .out_b_hv(sdiode_en_vpxa), .in_hv(vpxa));
ml_hv_invx3 I178 ( .sel_hv(net0109), .sel_25(net0109),
     .vddp_tieh(vddp_tieh), .out_b_hv(saprd_b_vpxa), .in_hv(vpxa));
ml_ls_vdd2vdd25 I136 ( .in(net053), .sup(vpxa), .out_vddio_b(net047),
     .out_vddio(net048), .in_b(net052));
ml_ls_vdd2vdd25 I137 ( .in(net078), .sup(vddp_), .out_vddio_b(net052),
     .out_vddio(net053), .in_b(net080));
ml_ls_vdd2vdd25 I172 ( .in(net0129), .sup(vpxa), .out_vddio_b(net0123),
     .out_vddio(net0124), .in_b(net0128));
ml_ls_vdd2vdd25 I173 ( .in(net073), .sup(vddp_), .out_vddio_b(net0128),
     .out_vddio(net0129), .in_b(net071));
ml_ls_vdd2vdd25 I180 ( .in(net0104), .sup(vpxa), .out_vddio_b(net0108),
     .out_vddio(net0109), .in_b(net0103));
ml_ls_vdd2vdd25 I181 ( .in(net059), .sup(vddp_), .out_vddio_b(net0103),
     .out_vddio(net0104), .in_b(net061));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_ctrl, View - schematic
// LAST TIME SAVED: Nov 22 16:36:48 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25, gred_25,
     gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25,
     gwlb_en_25, pgminhi_dmmy_b_25, s_25, s_rd_b_hv, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, bgr, bl_pgm_glb,
     gwl_b_sup_25, gwp_sup_hv, srdsup_hv, vddp_tieh, vpp_int, vpxa,
     wr_sup_25, fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rprd, fsm_tm_trow,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, s_rdin_hv, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25;

inout  bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv, srdsup_hv, vddp_tieh,
     vpp_int, vpxa, wr_sup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [3:0]  s_rd_b_hv;
output [3:0]  s_25;
output [1:0]  gred_b_25;
output [1:0]  gred_25;
output [5:0]  gnv_b_25;
output [4:1]  sa_ngate;
output [5:0]  gnv_25;

input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_trim_rrefpgm;
input [7:0]  fsm_rowadd;
input [0:0]  fsm_coladd;
input [3:0]  s_rdin_hv;
input [2:0]  fsm_trim_rrefrd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  gred;

wire  [2:0]  sa_trim;

wire  [5:0]  gnv;

wire  [3:0]  s;



vdd_tielow I204 ( .gnd_tiel(net0165));
nch_hvt  M2 ( .D(net0159), .B(GND_), .G(net0159), .S(gnd_));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net0159), .S(vddp_));
ml_rdhv_inv Iml_rdhv_inv_3_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[3]), .s_rd_b_hv(s_rd_b_hv[3]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_2_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[2]), .s_rd_b_hv(s_rd_b_hv[2]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_1_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[1]), .s_rd_b_hv(s_rd_b_hv[1]),
     .vddp_tieh(vddp_tieh));
ml_rdhv_inv Iml_rdhv_inv_0_ ( .srdsup_hv(srdsup_hv),
     .s_rdin_hv(s_rdin_hv[0]), .s_rd_b_hv(s_rd_b_hv[0]),
     .vddp_tieh(vddp_tieh));
ml_hvmux_hotswitch_enhance Ihvmux_gwpsup_hv ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwphv_vppint_25), .sel_hv_a_25(gwphv_vddp_25),
     .out_hv(gwp_sup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_gwlwr_ctrl_logic Igwlwr_ctrl_logic ( .fsm_tm_rprd(fsm_tm_rprd),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_pgmdisc(fsm_pgmdisc), .gwlb_en(gwlb_en),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_rd(fsm_rd), .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[0]), .wrsup_2vdd(wrsup_2vdd),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .testdec_prec_b(testdec_prec_b),
     .testdec_odd_b(testdec_odd_b), .testdec_even_b(testdec_even_b),
     .testdec_en_b(testdec_en_b), .saen(saen), .sa_trim(sa_trim[2:0]),
     .s(s[3:0]), .pgminhi_dmmy_b(net179), .gwphv_vppint(gwphv_vppint),
     .gwphv_vddp(gwphv_vddp), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vddp(gwlbsup_vddp), .gwlb_dis(gwlb_dis),
     .gwl_misc(gwl_misc), .gred(gred[1:0]), .gnv(gnv[5:0]));
ml_hvmux_hotswitch Ihvmux_gwlbsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwlbsup_vpxa_25), .sel_hv_a_25(gwlbsup_vddp_25),
     .out_hv(gwl_b_sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_gwlwr_bldrv Igwlwr_bldrv ( .fsm_din(fsm_din), .tm_dma(tm_dma),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .bl_frc_gnd(gnd_), .bgr(bgr),
     .bl_pgm_glb(bl_pgm_glb));
ml_gwlwr_ctrl_wr_sup Igwlwr_ctrl_wr_sup ( .wrsup_2vdd(wrsup_2vdd),
     .wrsup_2vdd_25(wrsup_2vdd_25), .wr_sup_25(wr_sup_25));
ml_gwlwr_ctrl_ls25 Igwlwr_ctrl_ls25 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_en(gwlb_en), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwlb_dis(gwlb_dis), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vpxa_25(gwlbsup_vpxa_25), .wrsup_2vdd_25(wrsup_2vdd_25),
     .wrsup_2vdd(wrsup_2vdd), .testdec_odd_b(testdec_odd_b),
     .testdec_even_b(testdec_even_b),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .pgminhi_dmmy_b(net179),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwphv_vddp(gwphv_vddp),
     .gwlbsup_vddp(gwlbsup_vddp), .gwphv_vppint(gwphv_vppint),
     .gwlbsup_vddp_25(gwlbsup_vddp_25),
     .gwphv_vppint_25(gwphv_vppint_25), .gwphv_vddp_25(gwphv_vddp_25),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .s(s[3:0]), .gwl_red(fsm_nv_rrow),
     .gwl_nvcm(fsm_nv_bstream), .gwl_misc(gwl_misc), .gred(gred[1:0]),
     .gnv(gnv[5:0]), .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]));
ml_core_sa_npgate_gen Icore_sa_npgate_gen ( .fsm_tm_sdiode(net0165),
     .saprd_b_vpxa(saprd_b_vpxa), .fsm_tm_rprd(fsm_tm_rprd),
     .sdiode_en_vpxa(sdiode_en_vpxa), .sa_ngate(sa_ngate[4:1]),
     .fsm_tm_testdec(tm_testdec), .satrim(sa_trim[2:0]),
     .vddp_tieh(vddp_tieh), .saen(saen), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .vpxa(vpxa));

endmodule
// Library - NVCM_40nm, Cell - ml_gwlwr_top_1f, View - schematic
// LAST TIME SAVED: Mar  7 17:51:21 2011
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_gwlwr_top_1f ( fsm_gwlbdis_b_25, gwl_b_25, gwl_b_sup_25,
     gwp_hv, pgminhi_dmmy_b_25, s_rd_b_hv, sa_ngate, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b, wr, bgr,
     bl_pgm_glb, srdsup_hv, vpp_int, vpxa, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     s_rdin_hv, tm_dma, tm_testdec, tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_b_sup_25, pgminhi_dmmy_b_25, saen_25,
     saen_b_vpxa, saprd_b_vpxa, sdiode_en_vpxa, testdec_en_b,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b;

inout  bgr, bl_pgm_glb, srdsup_hv, vpp_int, vpxa;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rprd, fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren,
     fsm_ymuxdis, tm_dma, tm_testdec, tm_testdec_wr;

output [107:0]  wr;
output [26:0]  gwl_b_25;
output [3:0]  s_rd_b_hv;
output [26:0]  gwp_hv;
output [4:1]  sa_ngate;

input [7:0]  fsm_rowadd;
input [3:0]  s_rdin_hv;
input [2:0]  fsm_trim_rrefpgm;
input [0:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_trim_ipp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_25;

wire  [1:0]  gred_b_25;

wire  [1:0]  gred_25;

wire  [5:0]  gnv_b_25;

wire  [5:0]  gnv_25;



ml_gwlwr_1f Igwlwr ( .gwp_hv(gwp_hv[26:0]), .gwl_b_25(gwl_b_25[26:0]),
     .wr(wr[107:0]), .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .wr_sup_25(wr_sup_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));
ml_gwlwr_ctrl Igwlwr_ctrl ( .saprd_b_vpxa(saprd_b_vpxa),
     .sdiode_en_vpxa(sdiode_en_vpxa), .srdsup_hv(srdsup_hv),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rdin_hv(s_rdin_hv[3:0]),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .sa_ngate(sa_ngate[4:1]),
     .testdec_en_b(testdec_en_b), .testdec_prec_b(testdec_prec_b),
     .fsm_pgmdisc(fsm_pgmdisc), .gwlb_en_25(gwlb_en_25),
     .fsm_din(fsm_din), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_allwl_l(fsm_tm_allwl_l), .fsm_tm_allwl_h(fsm_tm_allwl_h),
     .fsm_tm_allbl_l(fsm_tm_allbl_l), .fsm_tm_allbl_h(fsm_tm_allbl_h),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .s_25(s_25[3:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_red_25(gwl_red_25), .gwl_nvcm_25(gwl_nvcm_25),
     .gwl_misc_25(gwl_misc_25), .gred_b_25(gred_b_25[1:0]),
     .gred_25(gred_25[1:0]), .gnv_b_25(gnv_b_25[5:0]),
     .gnv_25(gnv_25[5:0]), .wr_sup_25(wr_sup_25), .vpxa(vpxa),
     .vpp_int(vpp_int), .vddp_tieh(vddp_tieh), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_core_1f, View - schematic
// LAST TIME SAVED: Dec 31 15:08:48 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_chip_nvcm_core_1f ( nv_dataout, s_rd, bgr, ngate_25,
     sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi, vpp_int, vpxa,
     ysup_25, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_multibl_read, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_ref,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_trim_ipp,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, s_rdin_hv, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi,
     vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [8:0]  nv_dataout;
output [3:0]  s_rd;

input [2:0]  fsm_trim_rrefpgm;
input [1:0]  fsm_tm_ref;
input [3:0]  fsm_trim_ipp;
input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_blkadd;
input [9:0]  fsm_coladd;
input [3:0]  s_rdin_hv;
input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [26:0]  gwl_b_25;

wire  [107:0]  wr;

wire  [3:0]  s_rd_b_hv;

wire  [26:0]  gwp_hv;

wire  [4:1]  sa_ngate;



ml_core_bank_1_1f Ibank_1 ( .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .gwl_b_25(gwl_b_25[26:0]), .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]),
     .fsm_tm_ref(fsm_tm_ref[1:0]), .tm_allbank_sel(tm_allbank_sel),
     .saprd_b_vpxa(saprd_b_vxpa), .gwl_b_sup_25(gwl_b_sup_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .ngate_25(ngate_25),
     .s_rd(s_rd[3:0]), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .bl_pgm_glb(bl_pgm_glb),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd(fsm_blkadd[3:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_rprd(fsm_tm_rprd), .nv_dataout(nv_dataout[8:4]));
ml_core_bank_0_1f Ibank_0 ( .sa_ngate(sa_ngate[4:1]),
     .testdec_prec_b(testdec_prec_b), .testdec_en_b(testdec_en_b),
     .gwl_b_25(gwl_b_25[26:0]), .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .saen_25(saen_25), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .saen_b_vpxa(saen_b_vpxa),
     .saprd_b_vpxa(saprd_b_vxpa), .gwl_b_sup_25(gwl_b_sup_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .fsm_tm_ref(fsm_tm_ref[1:0]),
     .fsm_nvcmen(fsm_nvcmen), .fsm_pgm(fsm_pgm),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd(fsm_blkadd[3:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_tm_trow(fsm_tm_trow), .ngate_25(ngate_25),
     .nv_dataout(nv_dataout[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .tm_allbank_sel(tm_allbank_sel));
ml_gwlwr_top_1f Igwlwr_top_1f ( .gwl_b_25(gwl_b_25[26:0]),
     .gwp_hv(gwp_hv[26:0]), .wr(wr[107:0]),
     .tm_testdec_wr(tm_testdec_wr), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wgnden(fsm_wgnden), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_tm_allbl_h(tm_allbl_h),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .saprd_b_vpxa(saprd_b_vxpa),
     .fsm_lshven(fsm_lshven), .fsm_wren(fsm_wren),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .testdec_en_b(testdec_en_b), .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .sdiode_en_vpxa(net335), .srdsup_hv(srdsup_hv), .vpxa(vpxa),
     .vpp_int(vpp_int), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr),
     .gwl_b_sup_25(gwl_b_sup_25), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rdin_hv(s_rdin_hv[3:0]), .tm_testdec(fsm_tm_testdec),
     .s_rd_b_hv(s_rd_b_hv[3:0]), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .sa_ngate(sa_ngate[4:1]), .testdec_prec_b(testdec_prec_b),
     .fsm_wpen(fsm_wpen), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_tm_allwl_l(tm_allwl_l), .fsm_tm_allbl_l(tm_allbl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .fsm_din(fsm_din), .tm_dma(tm_dma));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_buf, View - schematic
// LAST TIME SAVED: Sep 30 11:47:35 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_chip_buf ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(in), .Y(net120));
inv_hvt I45 ( .A(net120), .Y(out));

endmodule
// Library - xpmem, Cell - cram2x2, View - schematic
// LAST TIME SAVED: Jun 24 18:02:08 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module cram2x2 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [3:0]  q_b;
output [3:0]  q;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
input [1:0]  r_vdd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



eh_cram_cell_4 I_1_10 ( .q_b(q_b[1]), .q(q[1]), .wl(wl[0]), .bl(bl[1]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I_2_01 ( .q_b(q_b[2]), .q(q[2]), .wl(wl[1]), .bl(bl[0]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));
eh_cram_cell_4 I_0_00 ( .q_b(q_b[0]), .q(q[0]), .wl(wl[0]), .bl(bl[0]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I_3_11 ( .q_b(q_b[3]), .q(q[3]), .wl(wl[1]), .bl(bl[1]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_buf_hvsw_8f, View - schematic
// LAST TIME SAVED: Sep 10 14:09:50 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_chip_buf_hvsw_8f ( fsm_bgr_dis_buf, fsm_nvcmen_buf,
     fsm_pumpen_buf, fsm_tm_xforce_buf, fsm_tm_xvpxaint_buf,
     fsm_trim_vbg_buf, fsm_vrdwl_buf, fsm_bgr_dis, fsm_nvcmen,
     fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint, fsm_trim_vbg,
     fsm_vrdwl );
output  fsm_bgr_dis_buf, fsm_nvcmen_buf, fsm_pumpen_buf,
     fsm_tm_xforce_buf, fsm_tm_xvpxaint_buf;

input  fsm_bgr_dis, fsm_nvcmen, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint;

output [2:0]  fsm_vrdwl_buf;
output [3:0]  fsm_trim_vbg_buf;

input [2:0]  fsm_vrdwl;
input [3:0]  fsm_trim_vbg;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net256;



mux2_hvt I158 ( .in1(net153), .in0(net153), .out(net263),
     .sel(gnd_in));
mux2_hvt I206 ( .in1(gnd_in), .in0(gnd_in), .out(net161),
     .sel(gnd_in));
mux2_hvt I156 ( .in1(net161), .in0(net161), .out(net157),
     .sel(gnd_in));
mux2_hvt I157 ( .in1(net157), .in0(net157), .out(net153),
     .sel(gnd_in));
nor3_hvt I137 ( .B(net203), .Y(net199), .A(net203), .C(net203));
nor3_hvt I138 ( .B(net199), .Y(net195), .A(net199), .C(net199));
nor3_hvt I141 ( .B(net195), .Y(net191), .A(net195), .C(net195));
nor3_hvt I142 ( .B(net191), .Y(net187), .A(net191), .C(net191));
nor3_hvt I152 ( .B(net175), .Y(net171), .A(net175), .C(net175));
nor3_hvt I151 ( .B(net179), .Y(net175), .A(net179), .C(net179));
nor3_hvt I148 ( .B(net183), .Y(net179), .A(net183), .C(net183));
nor3_hvt I147 ( .B(net187), .Y(net183), .A(net187), .C(net187));
nor3_hvt I129 ( .B(net207), .Y(net203), .A(net207), .C(net207));
nor3_hvt I155 ( .B(net171), .Y(net262), .A(net171), .C(net171));
nand3_hvt I154 ( .Y(net261), .B(net212), .C(net212), .A(net212));
nand3_hvt I246 ( .Y(net244), .B(net248), .C(net248), .A(net248));
nand3_hvt I143 ( .Y(net228), .B(net232), .C(net232), .A(net232));
nand3_hvt I140 ( .Y(net232), .B(net236), .C(net236), .A(net236));
nand3_hvt I139 ( .Y(net236), .B(net240), .C(net240), .A(net240));
nand3_hvt I136 ( .Y(net240), .B(net244), .C(net244), .A(net244));
nand3_hvt I146 ( .Y(net224), .B(net228), .C(net228), .A(net228));
nand3_hvt I149 ( .Y(net220), .B(net224), .C(net224), .A(net224));
nand3_hvt I150 ( .Y(net216), .B(net220), .C(net220), .A(net220));
nand3_hvt I153 ( .Y(net212), .B(net216), .C(net216), .A(net216));
ml_chip_buf I120_3_ ( .in(vdd_spare), .out(net256[0]));
ml_chip_buf I120_2_ ( .in(vdd_spare), .out(net256[1]));
ml_chip_buf I120_1_ ( .in(vdd_spare), .out(net256[2]));
ml_chip_buf I120_0_ ( .in(vdd_spare), .out(net256[3]));
ml_chip_buf I159 ( .in(fsm_pumpen), .out(fsm_pumpen_buf));
ml_chip_buf I50_3_ ( .in(fsm_trim_vbg[3]), .out(fsm_trim_vbg_buf[3]));
ml_chip_buf I50_2_ ( .in(fsm_trim_vbg[2]), .out(fsm_trim_vbg_buf[2]));
ml_chip_buf I50_1_ ( .in(fsm_trim_vbg[1]), .out(fsm_trim_vbg_buf[1]));
ml_chip_buf I50_0_ ( .in(fsm_trim_vbg[0]), .out(fsm_trim_vbg_buf[0]));
ml_chip_buf I163 ( .in(fsm_bgr_dis), .out(fsm_bgr_dis_buf));
ml_chip_buf I49_2_ ( .in(fsm_vrdwl[2]), .out(fsm_vrdwl_buf[2]));
ml_chip_buf I49_1_ ( .in(fsm_vrdwl[1]), .out(fsm_vrdwl_buf[1]));
ml_chip_buf I49_0_ ( .in(fsm_vrdwl[0]), .out(fsm_vrdwl_buf[0]));
ml_chip_buf I53 ( .in(fsm_nvcmen), .out(fsm_nvcmen_buf));
ml_chip_buf I161 ( .in(fsm_tm_xvpxaint), .out(fsm_tm_xvpxaint_buf));
ml_chip_buf I160 ( .in(fsm_tm_xforce), .out(fsm_tm_xforce_buf));
vdd_tielow I135 ( .gnd_tiel(gnd_in));
vdd_tielow I145 ( .gnd_tiel(net248));
vdd_tielow I144 ( .gnd_tiel(net207));
vdd_tiehigh I117 ( .vdd_tieh(vdd_spare));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_buf, View - schematic
// LAST TIME SAVED: Oct  6 16:26:13 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_bgr_buf ( sa_out, en_25, inn, inp, sa_bias_25 );
inout  sa_out;

input  en_25, inn, inp, sa_bias_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M0 ( .D(sa_mirr_25), .B(GND_), .G(inp), .S(net436));
nch_na25  M1 ( .D(sa_out), .B(GND_), .G(inn), .S(net436));
nch_na25  M2 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_na25  M4 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_na25  M8 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_na25  M7 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M46 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M92 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M97 ( .D(tie_low), .B(GND_), .G(net0239), .S(GND_));
nch_25  M3 ( .D(net436), .B(GND_), .G(sa_bias_25), .S(GND_));
pch_25  M93 ( .D(net0123), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M95 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M94 ( .D(net0119), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M96 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M71 ( .D(sa_mirr_25), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M101 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M102 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M98 ( .D(net0239), .B(vddp_), .G(net0239), .S(vddp_));
pch_25  M10 ( .D(sa_mirr_25), .B(vddp_), .G(en_25), .S(vddp_));
pch_25  M91 ( .D(sa_out), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M25 ( .D(sa_out), .B(vddp_), .G(en_25), .S(vddp_));

endmodule
// Library - tsmcN40, Cell - nand4_25, View - schematic
// LAST TIME SAVED: Jan 25 22:28:24 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module nand4_25 ( Y, A, B, C, D, G, Gb, P, Pb );
output  Y;

input  A, B, C, D, G, Gb, P, Pb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M6 ( .D(net14), .B(Gb), .G(C), .S(net10));
nch_25  M7 ( .D(net10), .B(Gb), .G(D), .S(G));
nch_25  M4 ( .D(Y), .B(Gb), .G(A), .S(net18));
nch_25  M5 ( .D(net18), .B(Gb), .G(B), .S(net14));
pch_25  M2 ( .D(Y), .B(Pb), .G(C), .S(P));
pch_25  M1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(P));
pch_25  M3 ( .D(Y), .B(Pb), .G(D), .S(P));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ref_sw, View - schematic
// LAST TIME SAVED: Jul  9 15:54:44 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpp_ref_sw ( in, out, sel_b_25 );
inout  in, out;

input  sel_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I281 ( .IN(sel_b_25), .OUT(net122), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M12 ( .D(out), .B(GND_), .G(net122), .S(in));
pch_25  M14 ( .D(in), .B(vddp_), .G(sel_b_25), .S(out));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_res_100_ohm, View - schematic
// LAST TIME SAVED: May 28 16:29:33 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_bgr_res_100_ohm ( b, t );
inout  b, t;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo  R9 ( .MINUS(net7), .PLUS(net7));
rppolywo  R3 ( .MINUS(b), .PLUS(t));
rppolywo  R2 ( .MINUS(b), .PLUS(t));
rppolywo  R4 ( .MINUS(b), .PLUS(t));
rppolywo  R5 ( .MINUS(b), .PLUS(t));
rppolywo  R6 ( .MINUS(b), .PLUS(t));
rppolywo  R8 ( .MINUS(b), .PLUS(t));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr, View - schematic
// LAST TIME SAVED: Jan  3 16:50:37 2011
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_bgr ( bgr, bgr_bias, sa_bias_25, en_25 );
inout  bgr, bgr_bias, sa_bias_25;

input  en_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M75 ( .D(sa_mirr_25), .B(GND_), .G(in_pnpx8), .S(net436));
nch_na25  M60 ( .D(bgr_bias), .B(GND_), .G(in_pnpx1), .S(net436));
inv_25 I186 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nch_na25_macx  M76 ( .D(GND_), .G(tie_low), .S(GND_));
nch_na25_macx  M79 ( .D(GND_), .G(tie_low), .S(GND_));
nch_na25_macx  M78 ( .D(GND_), .G(tie_low), .S(GND_));
nch_na25_macx  M77 ( .D(GND_), .G(tie_low), .S(GND_));
pnp  QQ8 ( .C(GND_), .B(GND_), .E(net423));
pnp  QQ1 ( .C(GND_), .B(GND_), .E(in_pnpx1));
rppolywo  R4 ( .MINUS(sa_bias_25), .PLUS(net0209));
rppolywo  R0 ( .MINUS(net0209), .PLUS(net0303));
rppolywo  R3 ( .MINUS(in_pnpx1), .PLUS(bgr));
rppolywo  R1 ( .MINUS(in_pnpx8), .PLUS(bgr));
rppolywo  R2 ( .MINUS(net423), .PLUS(in_pnpx8));
rppolywo  R5 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R6 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R7 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R8 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R10 ( .MINUS(GND_), .PLUS(GND_));
rppolywo  R11 ( .MINUS(GND_), .PLUS(GND_));
nch_25  M97 ( .D(tie_low), .B(GND_), .G(net0309), .S(GND_));
nch_25  M82 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M58 ( .D(net0224), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M59 ( .D(net0224), .B(GND_), .G(en_b_25), .S(GND_));
nch_25  M85 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M100 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M96 ( .D(net0224), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M86 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M91 ( .D(GND_), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M94 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M23 ( .D(bgr), .B(GND_), .G(en_b_25), .S(GND_));
nch_25  M46 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M27 ( .D(sa_bias_25), .B(GND_), .G(en_b_25), .S(GND_));
nch_25  M92 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M81 ( .D(sa_bias_25), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M95 ( .D(net0224), .B(GND_), .G(sa_bias_25), .S(GND_));
nch_25  M93 ( .D(GND_), .B(GND_), .G(tie_low), .S(GND_));
nch_25  M3 ( .D(net436), .B(GND_), .G(sa_bias_25), .S(GND_));
pch_25  M88 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M22 ( .D(vddp_), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M62 ( .D(in_pnpx1), .B(vddp_), .G(net0224), .S(net0303));
pch_25  M83 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M98 ( .D(net0309), .B(vddp_), .G(net0309), .S(vddp_));
pch_25  M71 ( .D(sa_mirr_25), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M89 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M99 ( .D(net0323), .B(vddp_), .G(en_b_25), .S(vddp_));
pch_25  M74 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M40 ( .D(net0303), .B(vddp_), .G(en_b_25), .S(vddp_));
pch_25  M90 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M10 ( .D(sa_mirr_25), .B(vddp_), .G(en_25), .S(vddp_));
pch_25  M72 ( .D(net0224), .B(vddp_), .G(bgr_bias), .S(net0303));
pch_25  M80 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M73 ( .D(bgr), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M84 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M64 ( .D(bgr_bias), .B(vddp_), .G(sa_mirr_25), .S(vddp_));
pch_25  M87 ( .D(vddp_), .B(vddp_), .G(tie_low), .S(vddp_));
pch_25  M25 ( .D(bgr_bias), .B(vddp_), .G(en_25), .S(vddp_));

endmodule
// Library - NVCM_40nm, Cell - ml_bgr_top, View - schematic
// LAST TIME SAVED: Sep 10 14:19:39 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_bgr_top ( bgr_int, fsm_bgr_dis_buf, fsm_nvcmen_buf,
     fsm_trim_vbg_buf );
inout  bgr_int;

input  fsm_bgr_dis_buf, fsm_nvcmen_buf;

input [3:0]  fsm_trim_vbg_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net0169;

wire  [3:0]  net190;

wire  [3:0]  net192;

wire  [1:0]  net0170;

wire  [3:0]  net200;

wire  [3:0]  net201;

wire  [3:0]  bgrtrim_25;

wire  [15:0]  bgr_dec_b_25;

wire  [15:0]  vref;

wire  [3:0]  bgrtrim_b_25;



vdd_tiehigh I205 ( .vdd_tieh(net0167));
nand2_hvt I323 ( .B(fsm_nvcmen_buf), .A(net0281), .Y(net188));
ml_bgr_buf Iml_bgr_buf ( .sa_bias_25(sa_bias_25), .inp(bgr),
     .inn(vref[8]), .en_25(bgr_en_25), .sa_out(vref_reg));
nand4_25 I135_7_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[7]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_6_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[6]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_5_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[5]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_4_ ( .B(bgrtrim_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[4]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_3_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[3]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_2_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[2]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_1_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[1]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I135_0_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_25[3]),
     .Y(bgr_dec_b_25[0]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_15_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[15]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_14_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[14]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_13_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[13]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_12_ ( .B(bgrtrim_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[12]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_11_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[11]), .C(bgrtrim_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_10_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[10]), .C(bgrtrim_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_9_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[9]), .C(bgrtrim_b_25[1]), .D(bgrtrim_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
nand4_25 I184_8_ ( .B(bgrtrim_b_25[2]), .A(bgrtrim_b_25[3]),
     .Y(bgr_dec_b_25[8]), .C(bgrtrim_b_25[1]), .D(bgrtrim_b_25[0]),
     .P(vddp_), .G(gnd_), .Pb(vddp_), .Gb(gnd_));
pch_25  M6_1_ ( .D(net0169[0]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M6_0_ ( .D(net0169[1]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M7_1_ ( .D(net0170[0]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M7_0_ ( .D(net0170[1]), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M3 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M73 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M4 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M2 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M5 ( .D(net0155), .B(vddp_), .G(bgr_bias), .S(vddp_));
pch_25  M25 ( .D(net113), .B(vddp_), .G(bgr_en_b), .S(vddp_));
nch_na25_macx  M10 ( .D(gnd_), .G(vref_reg), .S(gnd_));
nch_na25_macx  M8 ( .D(gnd_), .G(vref_reg), .S(gnd_));
nch_na25_macx  M11 ( .D(gnd_), .G(bgr_int), .S(gnd_));
nch_na25_macx  M60 ( .D(net124), .G(vref_reg), .S(net0155));
nch_na25_macx  M0 ( .D(gnd_), .G(vref_reg), .S(gnd_));
ml_vpp_ref_sw I169 ( .in(bgr_int), .out(net0238), .sel_b_25(bgr_en_b));
ml_vpp_ref_sw I170 ( .in(bgr_int), .out(vref_vdd),
     .sel_b_25(bgr_en_25));
ml_vpp_ref_sw ref_sw_7_ ( .in(net0238), .out(vref[7]),
     .sel_b_25(bgr_dec_b_25[7]));
ml_vpp_ref_sw ref_sw_6_ ( .in(net0238), .out(vref[6]),
     .sel_b_25(bgr_dec_b_25[6]));
ml_vpp_ref_sw ref_sw_5_ ( .in(net0238), .out(vref[5]),
     .sel_b_25(bgr_dec_b_25[5]));
ml_vpp_ref_sw ref_sw_4_ ( .in(net0238), .out(vref[4]),
     .sel_b_25(bgr_dec_b_25[4]));
ml_vpp_ref_sw ref_sw_3_ ( .in(net0238), .out(vref[3]),
     .sel_b_25(bgr_dec_b_25[3]));
ml_vpp_ref_sw ref_sw_2_ ( .in(net0238), .out(vref[2]),
     .sel_b_25(bgr_dec_b_25[2]));
ml_vpp_ref_sw ref_sw_1_ ( .in(net0238), .out(vref[1]),
     .sel_b_25(bgr_dec_b_25[1]));
ml_vpp_ref_sw ref_sw_0_ ( .in(net0238), .out(vref[0]),
     .sel_b_25(bgr_dec_b_25[0]));
ml_vpp_ref_sw ref_sw_15_ ( .in(net0238), .out(vref[15]),
     .sel_b_25(bgr_dec_b_25[15]));
ml_vpp_ref_sw ref_sw_14_ ( .in(net0238), .out(vref[14]),
     .sel_b_25(bgr_dec_b_25[14]));
ml_vpp_ref_sw ref_sw_13_ ( .in(net0238), .out(vref[13]),
     .sel_b_25(bgr_dec_b_25[13]));
ml_vpp_ref_sw ref_sw_12_ ( .in(net0238), .out(vref[12]),
     .sel_b_25(bgr_dec_b_25[12]));
ml_vpp_ref_sw ref_sw_11_ ( .in(net0238), .out(vref[11]),
     .sel_b_25(bgr_dec_b_25[11]));
ml_vpp_ref_sw ref_sw_10_ ( .in(net0238), .out(vref[10]),
     .sel_b_25(bgr_dec_b_25[10]));
ml_vpp_ref_sw ref_sw_9_ ( .in(net0238), .out(vref[9]),
     .sel_b_25(bgr_dec_b_25[9]));
ml_vpp_ref_sw ref_sw_8_ ( .in(net0238), .out(vref[8]),
     .sel_b_25(bgr_dec_b_25[8]));
rppolywo  R0 ( .MINUS(vref[15]), .PLUS(net0147));
rppolywo  R8 ( .MINUS(gnd_), .PLUS(vref[0]));
rppolywo  R2 ( .MINUS(net0147), .PLUS(net124));
ml_bgr_res_100_ohm I90 ( .t(vref[8]), .b(vref[7]));
ml_bgr_res_100_ohm I91 ( .t(vref[7]), .b(vref[6]));
ml_bgr_res_100_ohm I92 ( .t(vref[6]), .b(vref[5]));
ml_bgr_res_100_ohm I93 ( .t(vref[4]), .b(vref[3]));
ml_bgr_res_100_ohm I94 ( .t(vref[5]), .b(vref[4]));
ml_bgr_res_100_ohm I95 ( .t(vref[1]), .b(vref[0]));
ml_bgr_res_100_ohm I97 ( .t(vref[2]), .b(vref[1]));
ml_bgr_res_100_ohm I100 ( .t(vref[3]), .b(vref[2]));
ml_bgr_res_100_ohm I101 ( .t(vref[13]), .b(vref[14]));
ml_bgr_res_100_ohm I102 ( .t(vref[14]), .b(vref[15]));
ml_bgr_res_100_ohm I104 ( .t(vref[11]), .b(vref[12]));
ml_bgr_res_100_ohm I105 ( .t(vref[12]), .b(vref[13]));
ml_bgr_res_100_ohm I106 ( .t(vref[10]), .b(vref[11]));
ml_bgr_res_100_ohm I107 ( .t(vref[9]), .b(vref[10]));
ml_bgr_res_100_ohm I108 ( .t(vref[8]), .b(vref[9]));
ml_bgr Iml_bgr ( .bgr_bias(bgr_bias), .sa_bias_25(sa_bias_25),
     .en_25(bgr_en_25), .bgr(bgr));
inv_25 I186 ( .IN(net195), .OUT(bgr_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I139 ( .IN(net196), .OUT(bgr_en_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I198_3_ ( .IN(net201[0]), .OUT(bgrtrim_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_2_ ( .IN(net201[1]), .OUT(bgrtrim_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_1_ ( .IN(net201[2]), .OUT(bgrtrim_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I198_0_ ( .IN(net201[3]), .OUT(bgrtrim_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_3_ ( .IN(net200[0]), .OUT(bgrtrim_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_2_ ( .IN(net200[1]), .OUT(bgrtrim_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_1_ ( .IN(net200[2]), .OUT(bgrtrim_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I195_0_ ( .IN(net200[3]), .OUT(bgrtrim_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I192 ( .IN(net0313), .OUT(bgr2vdd_25_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I189 ( .IN(net0312), .OUT(bgr2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I88_3_ ( .A(fsm_trim_vbg_buf[3]), .Y(net190[0]));
inv_hvt I88_2_ ( .A(fsm_trim_vbg_buf[2]), .Y(net190[1]));
inv_hvt I88_1_ ( .A(fsm_trim_vbg_buf[1]), .Y(net190[2]));
inv_hvt I88_0_ ( .A(fsm_trim_vbg_buf[0]), .Y(net190[3]));
inv_hvt I167 ( .A(net188), .Y(net186));
inv_hvt I183 ( .A(net0167), .Y(net0326));
inv_hvt I168 ( .A(fsm_bgr_dis_buf), .Y(net0281));
inv_hvt I174 ( .A(net0326), .Y(vref_vdd));
inv_hvt I87_3_ ( .A(net190[0]), .Y(net192[0]));
inv_hvt I87_2_ ( .A(net190[1]), .Y(net192[1]));
inv_hvt I87_1_ ( .A(net190[2]), .Y(net192[2]));
inv_hvt I87_0_ ( .A(net190[3]), .Y(net192[3]));
ml_ls_vdd2vdd25 I80_3_ ( .in(net192[0]), .sup(vddp_),
     .out_vddio_b(net200[0]), .out_vddio(net201[0]), .in_b(net190[0]));
ml_ls_vdd2vdd25 I80_2_ ( .in(net192[1]), .sup(vddp_),
     .out_vddio_b(net200[1]), .out_vddio(net201[1]), .in_b(net190[1]));
ml_ls_vdd2vdd25 I80_1_ ( .in(net192[2]), .sup(vddp_),
     .out_vddio_b(net200[2]), .out_vddio(net201[2]), .in_b(net190[2]));
ml_ls_vdd2vdd25 I80_0_ ( .in(net192[3]), .sup(vddp_),
     .out_vddio_b(net200[3]), .out_vddio(net201[3]), .in_b(net190[3]));
ml_ls_vdd2vdd25 I177 ( .in(vref_vdd), .sup(vddp_),
     .out_vddio_b(net0312), .out_vddio(net0313), .in_b(net0326));
ml_ls_vdd2vdd25 I335 ( .in(net186), .sup(vddp_), .out_vddio_b(net195),
     .out_vddio(net196), .in_b(net188));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_buf, View - schematic
// LAST TIME SAVED: Sep  3 15:27:07 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_pump_vpxa_buf ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I38 ( .IN(in), .OUT(net15), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
inv_25 I195 ( .IN(net15), .OUT(out), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_pump, View - schematic
// LAST TIME SAVED: Aug 30 18:07:52 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpp_pump ( pump_in, clkin_25, en_25 );
inout  pump_in;

input  clkin_25, en_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));
nmoscap_25  C1 ( .MINUS(clk_b_25), .PLUS(s_3));
nch_na25  M1 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
nch_na25  M2 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
nch_na25  M3 ( .D(s_2), .B(GND_), .G(s_2), .S(s_3));
nch_na25  M22 ( .D(net23), .B(GND_), .G(net23), .S(s_0));
nch_na25  M4 ( .D(s_3), .B(GND_), .G(s_3), .S(pump_in));
pch_25  M0 ( .D(net23), .B(vddp_), .G(net64), .S(vddp_));
inv_25 I230 ( .IN(clkin_25), .OUT(net0124), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I232 ( .IN(net088), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I233 ( .IN(net0100), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I234 ( .IN(net094), .OUT(net0106), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I235 ( .IN(net0106), .OUT(net0100), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I236 ( .IN(clkin_25), .OUT(net094), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I237 ( .IN(net0124), .OUT(net088), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I231 ( .IN(en_25), .OUT(net64), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));

endmodule
// Library - NVCM_40nm, Cell - ml_ls_vdd2vdd25_vpxa, View - schematic
// LAST TIME SAVED: Nov  6 18:00:25 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25_vpxa ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
nch_25  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));
pch_25  M0 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
pch_25  M1 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
pch_25  M2 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
pch_25  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));

endmodule
// Library - ice8chip, Cell - cram_2x2x2_ice8p, View - schematic
// LAST TIME SAVED: Jun 24 17:55:16 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module cram_2x2x2_ice8p ( q, q_b, bl, pgate_l, pgate_r, r_gnd_l,
     r_gnd_r, reset_l, reset_r, wl_l, wl_r );



output [7:0]  q_b;
output [7:0]  q;

inout [3:0]  bl;

input [1:0]  r_gnd_r;
input [1:0]  pgate_l;
input [1:0]  reset_r;
input [1:0]  wl_r;
input [1:0]  reset_l;
input [1:0]  pgate_r;
input [1:0]  r_gnd_l;
input [1:0]  wl_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 I_mem_r ( .bl(bl[3:2]), .q_b(q_b[7:4]), .reset(reset_r[1:0]),
     .q(q[7:4]), .wl(wl_r[1:0]), .r_vdd(r_gnd_r[1:0]),
     .pgate(pgate_r[1:0]));
cram2x2 I_mem_l ( .bl(bl[1:0]), .q_b(q_b[3:0]), .reset(reset_l[1:0]),
     .q(q[3:0]), .wl(wl_l[1:0]), .r_vdd(r_gnd_l[1:0]),
     .pgate(pgate_l[1:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_hv2vddp_sw, View - schematic
// LAST TIME SAVED: Nov 30 14:58:28 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hv2vddp_sw ( out_hv, hv2vddp, vddp_tieh, vpxa );
inout  out_hv;

input  hv2vddp, vddp_tieh, vpxa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_ls_vdd2vdd25_vpxa I64 ( .in(net44), .sup(vddp_),
     .out_vddio_b(net060), .out_vddio(net37), .in_b(net46));
pch_25  M1 ( .D(net27), .B(out_hv), .G(sw_vpp_b), .S(out_hv));
pch_25  M0 ( .D(net27), .B(vddp_), .G(sw_vddp_b), .S(vddp_));
inv_25 I62 ( .IN(net37), .OUT(sw_vddp_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I71 ( .IN(net060), .OUT(net035), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I65 ( .A(hv2vddp), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(sw_vddp_b),
     .sel_25(net035), .out_b_hv(sw_vpp_b), .in_hv(out_hv),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ref, View - schematic
// LAST TIME SAVED: Oct  8 16:18:32 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpp_ref ( vref_25, bgr, pumpen_25, vppwl_25 );
inout  vref_25;

input  bgr, pumpen_25;

input [2:0]  vppwl_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_b_25;

wire  [7:0]  red_dec_25;



nand3_25 I44_7_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[7]),
     .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_6_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[6]),
     .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_5_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[5]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_4_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[4]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_3_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[3]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_2_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[2]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_1_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[1]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_0_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[0]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nch_25  M10 ( .D(net163), .B(GND_), .G(bgr), .S(gnd_));
nch_25  M14 ( .D(net0113), .B(GND_), .G(vppref_en_b_25), .S(gnd_));
nch_25  M15 ( .D(ctrl_gate_25), .B(GND_), .G(vppref_en_b_25),
     .S(gnd_));
nch_25  M8 ( .D(ctrl_gate_25), .B(GND_), .G(bgr_mirror_25),
     .S(net163));
nch_25  M13 ( .D(net0113), .B(GND_), .G(bgr), .S(net163));
nch_na25  M0 ( .D(net179), .B(GND_), .G(ctrl_gate_25),
     .S(bgr_mirror_25));
nmoscap_25  C3 ( .MINUS(net0129), .PLUS(net0113));
nmoscap_25  C2 ( .MINUS(gnd_), .PLUS(ctrl_gate_25));
rppolywo_m  R14 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R15 ( .MINUS(net104), .PLUS(net0216), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net0216), .PLUS(net139), .BULK(GND_));
rppolywo_m  R19 ( .MINUS(net139), .PLUS(net0213), .BULK(GND_));
rppolywo_m  R22 ( .MINUS(net0213), .PLUS(net98), .BULK(GND_));
rppolywo_m  R25 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R24 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(net0100), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(net0100), .PLUS(net0100), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(net0100), .PLUS(net0193), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net0193), .PLUS(net110), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(bgr_mirror_25), .PLUS(net0129), .BULK(GND_));
pch_25  M1 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(net175));
pch_25  M18 ( .D(net179), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
pch_25  M5 ( .D(ctrl_gate_25), .B(vddp_), .G(net0113), .S(net175));
pch_25  M6 ( .D(net0113), .B(vddp_), .G(net0113), .S(net175));
pch_25  M7 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
inv_25 I38 ( .IN(pumpen_25), .OUT(vppref_en_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_2_ ( .IN(vppwl_25[2]), .OUT(vppwl_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_1_ ( .IN(vppwl_25[1]), .OUT(vppwl_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_0_ ( .IN(vppwl_25[0]), .OUT(vppwl_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_vpp_ref_sw I281 ( .in(net0213), .out(vref_25),
     .sel_b_25(red_dec_25[6]));
ml_vpp_ref_sw I287 ( .in(net0216), .out(vref_25),
     .sel_b_25(red_dec_25[4]));
ml_vpp_ref_sw I283 ( .in(net98), .out(vref_25),
     .sel_b_25(red_dec_25[7]));
ml_vpp_ref_sw I290 ( .in(net0193), .out(vref_25),
     .sel_b_25(red_dec_25[0]));
ml_vpp_ref_sw I288 ( .in(net104), .out(vref_25),
     .sel_b_25(red_dec_25[3]));
ml_vpp_ref_sw I284 ( .in(net139), .out(vref_25),
     .sel_b_25(red_dec_25[5]));
ml_vpp_ref_sw I291 ( .in(net110), .out(vref_25),
     .sel_b_25(red_dec_25[1]));
ml_vpp_ref_sw I292 ( .in(net113), .out(vref_25),
     .sel_b_25(red_dec_25[2]));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_ctrl, View - schematic
// LAST TIME SAVED: Nov  6 18:30:47 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpp_ctrl ( pumpen_25, vpint_en, vpp_2_vdd, vppdisc_vpxa,
     vppwl_25, vpxa, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_vpgmwl_buf, fsm_wgnden );
output  pumpen_25, vpint_en, vpp_2_vdd, vppdisc_vpxa;

inout  vpxa;

input  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint, fsm_wgnden;

output [2:0]  vppwl_25;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  net082;

wire  [2:0]  net092;

wire  [2:0]  net038;

wire  [2:0]  net068;



ml_ls_vdd2vdd25_vpxa I173 ( .in(fsm_pgmdisc_buf), .sup(vpxa),
     .out_vddio_b(net088), .out_vddio(net048), .in_b(net0106));
ml_dff_nvcm I77 ( .CLK(net084), .QN(vpp_pumpen_b), .R(pgm_dis),
     .D(vdd_tieh), .Q(vpp_pumpen));
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(net0122));
inv_25 I95_2_ ( .IN(net068[0]), .OUT(vppwl_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_1_ ( .IN(net068[1]), .OUT(vppwl_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_0_ ( .IN(net068[2]), .OUT(vppwl_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I81 ( .IN(net073), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(net088), .OUT(vppdisc_vpxa), .P(vpxa), .Pb(vpxa),
     .G(gnd_), .Gb(gnd_));
nand3_hvt I79 ( .C(net086), .A(fsm_pgm_buf), .Y(pgm_dis),
     .B(fsm_nvcmen_buf));
nor2_hvt I111 ( .A(vpp_pumpen_b), .B(net080), .Y(net0133));
nor2_hvt I87 ( .A(vpp_pumpen), .Y(net036), .B(fsm_pgmdisc_buf));
nand4_hvt I75 ( .D(fsm_pgm_buf), .C(fsm_lshven_buf), .A(net0127),
     .Y(net046), .B(net0127));
inv_hvt I107 ( .A(net0122), .Y(net0124));
inv_hvt I109 ( .A(fsm_pgmvfy_buf), .Y(net0127));
inv_hvt I131 ( .A(net049), .Y(net080));
inv_hvt I110_2_ ( .A(net092[0]), .Y(net082[0]));
inv_hvt I110_1_ ( .A(net092[1]), .Y(net082[1]));
inv_hvt I110_0_ ( .A(net092[2]), .Y(net082[2]));
inv_hvt I76 ( .A(net046), .Y(net084));
inv_hvt I108 ( .A(fsm_pgmdisc_buf), .Y(net0122));
inv_hvt I78 ( .A(net0124), .Y(net086));
inv_hvt I113 ( .A(vpp_pumpen_b), .Y(vpint_en));
inv_hvt I91 ( .A(net036), .Y(net089));
inv_hvt I90 ( .A(net089), .Y(vpp_2_vdd));
inv_hvt I98_2_ ( .A(fsm_vpgmwl_buf[2]), .Y(net092[0]));
inv_hvt I98_1_ ( .A(fsm_vpgmwl_buf[1]), .Y(net092[1]));
inv_hvt I98_0_ ( .A(fsm_vpgmwl_buf[0]), .Y(net092[2]));
inv_hvt I112 ( .A(net0133), .Y(net0134));
inv_hvt I101 ( .A(fsm_pgmdisc_buf), .Y(net0106));
nand2_hvt I104 ( .A(fsm_tm_xforce), .Y(net049), .B(fsm_tm_xvppint));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
ml_ls_vdd2vdd25 I96_2_ ( .in(net082[0]), .sup(vddp_),
     .out_vddio_b(net068[0]), .out_vddio(net038[0]), .in_b(net092[0]));
ml_ls_vdd2vdd25 I96_1_ ( .in(net082[1]), .sup(vddp_),
     .out_vddio_b(net068[1]), .out_vddio(net038[1]), .in_b(net092[1]));
ml_ls_vdd2vdd25 I96_0_ ( .in(net082[2]), .sup(vddp_),
     .out_vddio_b(net068[2]), .out_vddio(net038[2]), .in_b(net092[2]));
ml_ls_vdd2vdd25 I84 ( .in(net0133), .sup(vddp_), .out_vddio_b(net073),
     .out_vddio(net074), .in_b(net0134));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_reg, View - schematic
// LAST TIME SAVED: Nov  8 10:29:35 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpp_reg ( slow_25, bgr, pbias_25, pump_in, vpp_int, vpxa,
     pumpen_25, vppdisc_vpxa, vref_25 );
output  slow_25;

inout  bgr, pbias_25, pump_in, vpp_int, vpxa;

input  pumpen_25, vppdisc_vpxa, vref_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I211 ( .IN(en_buf_b_25), .OUT(en_buf_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I212 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R5 ( .MINUS(net0165), .PLUS(vpp_int), .BULK(GND_));
rppolywo_m  R6 ( .MINUS(gnd_), .PLUS(net0178), .BULK(GND_));
rppolywo_m  R14 ( .MINUS(net0271), .PLUS(vdd_), .BULK(GND_));
rppolywo_m  R15 ( .MINUS(net0271), .PLUS(vdd_), .BULK(GND_));
rppolywo_m  R16 ( .MINUS(net0271), .PLUS(vdd_), .BULK(GND_));
rppolywo_m  R11 ( .MINUS(vdd_), .PLUS(net0271), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(vdd_), .PLUS(net0271), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(pump_gate), .PLUS(pump_in), .BULK(GND_));
rppolywo_m  R7 ( .MINUS(net0178), .PLUS(net0175), .BULK(GND_));
rppolywo_m  R13 ( .MINUS(vdd_), .PLUS(net0271), .BULK(GND_));
pch_25  M31 ( .D(net0203), .B(net0165), .G(dis_pgate_25), .S(net0165));
pch_25  M2 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
pch_25  M9 ( .D(net0200), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
pch_25  M8_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
pch_25  M8_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0200));
pch_25  M14 ( .D(pump_opamp_out), .B(net125), .G(vref_25), .S(net125));
pch_25  M18 ( .D(net122), .B(vpp_int), .G(net122), .S(vpp_int));
pch_25  M13 ( .D(net124), .B(net125), .G(vdiv), .S(net125));
pch_25  M32 ( .D(dis_pgate_25), .B(vpxa), .G(dis_pgate_25), .S(vpxa));
pch_25  M33 ( .D(dis_pgate_25), .B(vpxa), .G(vppdisc_vpxa), .S(vpxa));
pch_25  M12 ( .D(net125), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M19 ( .D(net134), .B(net122), .G(net134), .S(net122));
pch_25  M21 ( .D(net138), .B(net134), .G(net138), .S(net134));
pch_25  M23 ( .D(net142), .B(net138), .G(net142), .S(net138));
pch_25  M24 ( .D(vdiv), .B(net142), .G(vdiv), .S(net142));
pch_25  M25 ( .D(net0224), .B(vdiv), .G(net0224), .S(vdiv));
nch_25  M40 ( .D(net0264), .B(GND_), .G(vppdisc_vpxa), .S(gnd_));
nch_25  M16 ( .D(net124), .B(GND_), .G(net124), .S(net155));
nch_25  M17 ( .D(net155), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M6 ( .D(vpp_int), .B(GND_), .G(en_buf_25), .S(net168));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
nch_25  M20 ( .D(slow_25), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M7 ( .D(net168), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M4 ( .D(dis_pgate_25), .B(GND_), .G(net0208), .S(net0264));
nch_25  M41 ( .D(net0224), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M15 ( .D(pump_opamp_out), .B(GND_), .G(net124), .S(net155));
nch_25  M0 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net0175));
nch_na25  M11 ( .D(net0199), .B(GND_), .G(vppdisc_vpxa), .S(net0271));
nch_na25  M22 ( .D(vpp_int), .B(GND_), .G(pump_gate), .S(pump_in));
nch_na25  M1 ( .D(GND_), .B(GND_), .G(pump_gate), .S(GND_));
nch_na25  M10 ( .D(net0203), .B(GND_), .G(net0208), .S(net0199));
nch_na25  M5 ( .D(pump_opamp_out), .B(GND_), .G(vpp_int),
     .S(pump_opamp_out));
vddp_tiehigh I261 ( .vddp_tieh(net0208));

endmodule
// Library - NVCM_40nm, Cell - ml_vpp_vco, View - schematic
// LAST TIME SAVED: Aug 25 11:10:03 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpp_vco ( clk_25_0, clk_25_1, pbias_25, slow_25, en_25,
     freq_25 );
output  clk_25_0, clk_25_1;

inout  pbias_25, slow_25;

input  en_25;

input [1:0]  freq_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:1]  freq_b_25;



nch_na25  M4 ( .D(GND_), .B(GND_), .G(net173), .S(GND_));
nch_na25  M15 ( .D(GND_), .B(GND_), .G(net185), .S(GND_));
nch_na25  M16 ( .D(GND_), .B(GND_), .G(net193), .S(GND_));
nch_na25  M2 ( .D(GND_), .B(GND_), .G(net189), .S(GND_));
nch_25  M5 ( .D(net173), .B(GND_), .G(net185), .S(net177));
nch_25  M6 ( .D(net177), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M13 ( .D(net181), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M14 ( .D(net185), .B(GND_), .G(net193), .S(net181));
nch_25  M8 ( .D(net189), .B(GND_), .G(net173), .S(net201));
nch_25  M17 ( .D(net193), .B(GND_), .G(net195), .S(net197));
nch_25  M18 ( .D(net197), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M1 ( .D(net201), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M23 ( .D(pbias_osc_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M24 ( .D(slow_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M25 ( .D(nbias_osc_25), .B(GND_), .G(en_25), .S(slow_25));
nand2_25 I96 ( .G(GND_), .Pb(vddp_), .A(net189), .Y(net195), .P(vddp_),
     .B(en_25), .Gb(GND_));
nand2_25 I205 ( .G(GND_), .Pb(vddp_), .A(net185), .Y(net0205),
     .P(vddp_), .B(en_25), .Gb(GND_));
pch_25  M7 ( .D(net173), .B(vddp_), .G(net185), .S(net236));
pch_25  M10 ( .D(net236), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M9 ( .D(net248), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M3 ( .D(net189), .B(vddp_), .G(net173), .S(net248));
pch_25  M11 ( .D(net256), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M12 ( .D(net185), .B(vddp_), .G(net193), .S(net256));
pch_25  M19 ( .D(net193), .B(vddp_), .G(net195), .S(net260));
pch_25  M20 ( .D(net260), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M22 ( .D(pbias_osc_25), .B(vddp_), .G(en_b_25), .S(net228));
pch_25  M26_1_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M26_0_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_1_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_0_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M28 ( .D(net212), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M29 ( .D(nbias_osc_25), .B(vddp_), .G(freq_25[0]), .S(net212));
pch_25  M30 ( .D(nbias_osc_25), .B(vddp_), .G(freq_b_25[1]),
     .S(net208));
pch_25  M21 ( .D(net228), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
inv_25 I201 ( .IN(net195), .OUT(clk_25_0), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(net0205), .OUT(clk_25_1), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I188 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I199 ( .IN(freq_25[1]), .OUT(freq_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));

endmodule
// Library - NVCM_40nm, Cell - ml_vppint_top, View - schematic
// LAST TIME SAVED: Nov  6 18:24:09 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vppint_top ( vpint_en, vpp_int, vpxa, bgr, fsm_lshven_buf,
     fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf, fsm_pgmvfy_buf,
     fsm_tm_xforce, fsm_tm_xvppint, fsm_vpgmwl_buf, fsm_wgnden_buf );
output  vpint_en;

inout  vpp_int, vpxa;

input  bgr, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_wgnden_buf;

input [2:0]  fsm_vpgmwl_buf;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_25;

wire  [1:0]  freq_25;



ml_pump_vpxa_buf I95 ( .in(clkin_0_25), .out(net52));
ml_pump_vpxa_buf I81 ( .in(clkin_1_25), .out(net061));
ml_vpp_pump Ivpp_pump_0 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(clkin_1_25));
ml_vpp_pump Ivpp_pump_1 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net061));
ml_vpp_pump Ivpp_pump_2 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net52));
inv_25 I38 ( .IN(vddp_tieh), .OUT(freq_25[1]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I91 ( .IN(vddp_tieh), .OUT(freq_25[0]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpp_int));
ml_hv2vddp_sw Ivpxa_2vddp_sw ( .vpxa(vpxa), .hv2vddp(vpp_2_vdd),
     .vddp_tieh(vddp_tieh), .out_hv(vpp_int));
ml_vpp_ref Ivpp_ref ( .vref_25(vref_25), .vppwl_25(vppwl_25[2:0]),
     .pumpen_25(pumpen_25), .bgr(bgr));
ml_vpp_ctrl Ivpp_ctrl ( .vppdisc_vpxa(vppdisc_vpxa), .vpxa(vpxa),
     .vpint_en(vpint_en), .fsm_pgmvfy_buf(fsm_pgmvfy_buf),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .fsm_wgnden(fsm_wgnden_buf),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf), .vppwl_25(vppwl_25[2:0]),
     .vpp_2_vdd(vpp_2_vdd), .pumpen_25(pumpen_25));
ml_vpp_reg Ivpp_reg ( .vpxa(vpxa), .vppdisc_vpxa(vppdisc_vpxa),
     .bgr(bgr), .slow_25(slow_25), .pbias_25(pbias_25),
     .vref_25(vref_25), .pumpen_25(pumpen_25), .pump_in(pump_in),
     .vpp_int(vpp_int));
ml_vpp_vco Ivpp_vco ( .clk_25_1(clkin_1_25), .pbias_25(pbias_25),
     .slow_25(slow_25), .freq_25(freq_25[1:0]), .en_25(pumpen_25),
     .clk_25_0(clkin_0_25));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_3.3v, View - schematic
// LAST TIME SAVED: Aug 30 18:07:58 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_pump_vpxa_3_3v ( out, clkin_25, en_25 );
inout  out;

input  clkin_25, en_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C1 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C2 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C3 ( .MINUS(clk_25), .PLUS(s_2));
nch_na25  M1 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
nch_na25  M2 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
nch_na25  M3 ( .D(s_2), .B(GND_), .G(s_2), .S(out));
nch_na25  M4 ( .D(net73), .B(GND_), .G(net73), .S(s_0));
pch_25  M6 ( .D(net73), .B(vddp_), .G(net114), .S(vddp_));
inv_25 I230 ( .IN(clkin_25), .OUT(net120), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I231 ( .IN(en_25), .OUT(net114), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I232 ( .IN(net78), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I233 ( .IN(net90), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I234 ( .IN(net84), .OUT(net96), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I235 ( .IN(net96), .OUT(net90), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I236 ( .IN(clkin_25), .OUT(net84), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I237 ( .IN(net120), .OUT(net78), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));

endmodule
// Library - sbtlibn65lp, Cell - ml_dlatch_25, View - schematic
// LAST TIME SAVED: Aug 30 17:06:09 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_dlatch_25 ( Q_25, D_25, EN_25, R_25 );
output  Q_25;

input  D_25, EN_25, R_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_25 I161 ( .A(net52), .Y(Q_25), .Gb(GND_), .G(GND_), .Pb(vddp_),
     .P(vddp_), .B(R_25));
inv_25 I156 ( .IN(EN_25), .OUT(EN_B_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nch_25  M0 ( .D(net52), .B(GND_), .G(D_25), .S(net48));
nch_25  M1 ( .D(net48), .B(GND_), .G(EN_25), .S(GND_));
nch_25  M5 ( .D(net40), .B(GND_), .G(EN_B_25), .S(GND_));
nch_25  M6 ( .D(net52), .B(GND_), .G(Q_25), .S(net40));
pch_25  M2 ( .D(net52), .B(vddp_), .G(Q_25), .S(net31));
pch_25  M8 ( .D(net31), .B(vddp_), .G(EN_25), .S(vddp_));
pch_25  M7 ( .D(net39), .B(vddp_), .G(EN_B_25), .S(vddp_));
pch_25  M3 ( .D(net52), .B(vddp_), .G(D_25), .S(net39));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_clk_reg, View - schematic
// LAST TIME SAVED: Aug 30 17:59:46 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_pump_clk_reg ( clk_out_25, clk_in_25, pump_chrg_25,
     pump_on_25 );
output  clk_out_25;

input  clk_in_25, pump_chrg_25, pump_on_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I78 ( .G(GND_), .Pb(vddp_), .A(pump_chrg_25), .Y(clk_freeze),
     .P(vddp_), .B(pump_on_25), .Gb(GND_));
inv_25 I72 ( .IN(net020), .OUT(clk_equal), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(vddp_tieh), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
exor2_25 I85 ( .A(clk_in_25), .Y(net020), .B(clk_out_25));
vddp_tiehigh I117 ( .vddp_tieh(vddp_tieh));
ml_dlatch_25 I63 ( .D_25(clk_in_25), .EN_25(clk_go), .R_25(net34),
     .Q_25(clk_out_25));
ml_dlatch_25 I64 ( .D_25(vddp_tieh), .EN_25(clk_equal),
     .R_25(clk_freeze), .Q_25(clk_go));

endmodule
// Library - NVCM_40nm, Cell - ml_pump_vpxa_x2, View - schematic
// LAST TIME SAVED: Sep  1 14:53:51 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_pump_vpxa_x2 ( vpxa_int, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, pumpen_25, vpxa_clk_25, vpxa_clk_b_25 );
inout  vpxa_int;

input  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25, pumpen_25,
     vpxa_clk_25, vpxa_clk_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_pump_vpxa_buf I80 ( .in(net43), .out(clkin_2_25));
ml_pump_vpxa_buf I79 ( .in(net47), .out(net22));
ml_pump_vpxa_buf I78 ( .in(net39), .out(clkin_0_25));
ml_pump_vpxa_buf I81 ( .in(net22), .out(clkin_1_25));
ml_pump_vpxa_3_3v Ivpxa_pump_0 ( .en_25(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_0_25));
ml_pump_vpxa_3_3v Ivpxa_pump_2 ( .en_25(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_2_25));
ml_pump_vpxa_3_3v Ivpxa_pump_1 ( .en_25(pumpen_25),
     .clkin_25(clkin_1_25), .out(vpxa_int));
ml_pump_clk_reg Iclk_reg_0 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_0_25), .pump_on_25(pumpen_25),
     .clk_out_25(net39));
ml_pump_clk_reg Iclk_reg_2 ( .clk_in_25(vpxa_clk_b_25),
     .pump_chrg_25(pump_chrg_2_25), .pump_on_25(pumpen_25),
     .clk_out_25(net43));
ml_pump_clk_reg Iclk_reg_1 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_1_25), .pump_on_25(pumpen_25),
     .clk_out_25(net47));

endmodule
// Library - ice1chip, Cell - ice1f_cram_row142col4, View - schematic
// LAST TIME SAVED: Mar 10 12:33:59 2011
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module ice1f_cram_row142col4 ( bl, pgate_l, pgate_r, reset_l, reset_r,
     vdd_cntl_l, vdd_cntl_r, wl_l, wl_r );


inout [3:0]  bl;

input [141:0]  wl_r;
input [141:0]  pgate_l;
input [141:0]  wl_l;
input [141:0]  reset_r;
input [141:0]  vdd_cntl_r;
input [141:0]  pgate_r;
input [141:0]  reset_l;
input [141:0]  vdd_cntl_l;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [567:0]  net35;

wire  [567:0]  net36;

wire  [141:0]  r_gnd_r;

wire  [141:0]  r_gnd_l;



pch_hvt  M0_141_ ( .D(r_gnd_r[141]), .B(vdd_), .G(vdd_cntl_r[141]),
     .S(vdd_));
pch_hvt  M0_140_ ( .D(r_gnd_r[140]), .B(vdd_), .G(vdd_cntl_r[140]),
     .S(vdd_));
pch_hvt  M0_139_ ( .D(r_gnd_r[139]), .B(vdd_), .G(vdd_cntl_r[139]),
     .S(vdd_));
pch_hvt  M0_138_ ( .D(r_gnd_r[138]), .B(vdd_), .G(vdd_cntl_r[138]),
     .S(vdd_));
pch_hvt  M0_137_ ( .D(r_gnd_r[137]), .B(vdd_), .G(vdd_cntl_r[137]),
     .S(vdd_));
pch_hvt  M0_136_ ( .D(r_gnd_r[136]), .B(vdd_), .G(vdd_cntl_r[136]),
     .S(vdd_));
pch_hvt  M0_135_ ( .D(r_gnd_r[135]), .B(vdd_), .G(vdd_cntl_r[135]),
     .S(vdd_));
pch_hvt  M0_134_ ( .D(r_gnd_r[134]), .B(vdd_), .G(vdd_cntl_r[134]),
     .S(vdd_));
pch_hvt  M0_133_ ( .D(r_gnd_r[133]), .B(vdd_), .G(vdd_cntl_r[133]),
     .S(vdd_));
pch_hvt  M0_132_ ( .D(r_gnd_r[132]), .B(vdd_), .G(vdd_cntl_r[132]),
     .S(vdd_));
pch_hvt  M0_131_ ( .D(r_gnd_r[131]), .B(vdd_), .G(vdd_cntl_r[131]),
     .S(vdd_));
pch_hvt  M0_130_ ( .D(r_gnd_r[130]), .B(vdd_), .G(vdd_cntl_r[130]),
     .S(vdd_));
pch_hvt  M0_129_ ( .D(r_gnd_r[129]), .B(vdd_), .G(vdd_cntl_r[129]),
     .S(vdd_));
pch_hvt  M0_128_ ( .D(r_gnd_r[128]), .B(vdd_), .G(vdd_cntl_r[128]),
     .S(vdd_));
pch_hvt  M0_127_ ( .D(r_gnd_r[127]), .B(vdd_), .G(vdd_cntl_r[127]),
     .S(vdd_));
pch_hvt  M0_126_ ( .D(r_gnd_r[126]), .B(vdd_), .G(vdd_cntl_r[126]),
     .S(vdd_));
pch_hvt  M0_125_ ( .D(r_gnd_r[125]), .B(vdd_), .G(vdd_cntl_r[125]),
     .S(vdd_));
pch_hvt  M0_124_ ( .D(r_gnd_r[124]), .B(vdd_), .G(vdd_cntl_r[124]),
     .S(vdd_));
pch_hvt  M0_123_ ( .D(r_gnd_r[123]), .B(vdd_), .G(vdd_cntl_r[123]),
     .S(vdd_));
pch_hvt  M0_122_ ( .D(r_gnd_r[122]), .B(vdd_), .G(vdd_cntl_r[122]),
     .S(vdd_));
pch_hvt  M0_121_ ( .D(r_gnd_r[121]), .B(vdd_), .G(vdd_cntl_r[121]),
     .S(vdd_));
pch_hvt  M0_120_ ( .D(r_gnd_r[120]), .B(vdd_), .G(vdd_cntl_r[120]),
     .S(vdd_));
pch_hvt  M0_119_ ( .D(r_gnd_r[119]), .B(vdd_), .G(vdd_cntl_r[119]),
     .S(vdd_));
pch_hvt  M0_118_ ( .D(r_gnd_r[118]), .B(vdd_), .G(vdd_cntl_r[118]),
     .S(vdd_));
pch_hvt  M0_117_ ( .D(r_gnd_r[117]), .B(vdd_), .G(vdd_cntl_r[117]),
     .S(vdd_));
pch_hvt  M0_116_ ( .D(r_gnd_r[116]), .B(vdd_), .G(vdd_cntl_r[116]),
     .S(vdd_));
pch_hvt  M0_115_ ( .D(r_gnd_r[115]), .B(vdd_), .G(vdd_cntl_r[115]),
     .S(vdd_));
pch_hvt  M0_114_ ( .D(r_gnd_r[114]), .B(vdd_), .G(vdd_cntl_r[114]),
     .S(vdd_));
pch_hvt  M0_113_ ( .D(r_gnd_r[113]), .B(vdd_), .G(vdd_cntl_r[113]),
     .S(vdd_));
pch_hvt  M0_112_ ( .D(r_gnd_r[112]), .B(vdd_), .G(vdd_cntl_r[112]),
     .S(vdd_));
pch_hvt  M0_111_ ( .D(r_gnd_r[111]), .B(vdd_), .G(vdd_cntl_r[111]),
     .S(vdd_));
pch_hvt  M0_110_ ( .D(r_gnd_r[110]), .B(vdd_), .G(vdd_cntl_r[110]),
     .S(vdd_));
pch_hvt  M0_109_ ( .D(r_gnd_r[109]), .B(vdd_), .G(vdd_cntl_r[109]),
     .S(vdd_));
pch_hvt  M0_108_ ( .D(r_gnd_r[108]), .B(vdd_), .G(vdd_cntl_r[108]),
     .S(vdd_));
pch_hvt  M0_107_ ( .D(r_gnd_r[107]), .B(vdd_), .G(vdd_cntl_r[107]),
     .S(vdd_));
pch_hvt  M0_106_ ( .D(r_gnd_r[106]), .B(vdd_), .G(vdd_cntl_r[106]),
     .S(vdd_));
pch_hvt  M0_105_ ( .D(r_gnd_r[105]), .B(vdd_), .G(vdd_cntl_r[105]),
     .S(vdd_));
pch_hvt  M0_104_ ( .D(r_gnd_r[104]), .B(vdd_), .G(vdd_cntl_r[104]),
     .S(vdd_));
pch_hvt  M0_103_ ( .D(r_gnd_r[103]), .B(vdd_), .G(vdd_cntl_r[103]),
     .S(vdd_));
pch_hvt  M0_102_ ( .D(r_gnd_r[102]), .B(vdd_), .G(vdd_cntl_r[102]),
     .S(vdd_));
pch_hvt  M0_101_ ( .D(r_gnd_r[101]), .B(vdd_), .G(vdd_cntl_r[101]),
     .S(vdd_));
pch_hvt  M0_100_ ( .D(r_gnd_r[100]), .B(vdd_), .G(vdd_cntl_r[100]),
     .S(vdd_));
pch_hvt  M0_99_ ( .D(r_gnd_r[99]), .B(vdd_), .G(vdd_cntl_r[99]),
     .S(vdd_));
pch_hvt  M0_98_ ( .D(r_gnd_r[98]), .B(vdd_), .G(vdd_cntl_r[98]),
     .S(vdd_));
pch_hvt  M0_97_ ( .D(r_gnd_r[97]), .B(vdd_), .G(vdd_cntl_r[97]),
     .S(vdd_));
pch_hvt  M0_96_ ( .D(r_gnd_r[96]), .B(vdd_), .G(vdd_cntl_r[96]),
     .S(vdd_));
pch_hvt  M0_95_ ( .D(r_gnd_r[95]), .B(vdd_), .G(vdd_cntl_r[95]),
     .S(vdd_));
pch_hvt  M0_94_ ( .D(r_gnd_r[94]), .B(vdd_), .G(vdd_cntl_r[94]),
     .S(vdd_));
pch_hvt  M0_93_ ( .D(r_gnd_r[93]), .B(vdd_), .G(vdd_cntl_r[93]),
     .S(vdd_));
pch_hvt  M0_92_ ( .D(r_gnd_r[92]), .B(vdd_), .G(vdd_cntl_r[92]),
     .S(vdd_));
pch_hvt  M0_91_ ( .D(r_gnd_r[91]), .B(vdd_), .G(vdd_cntl_r[91]),
     .S(vdd_));
pch_hvt  M0_90_ ( .D(r_gnd_r[90]), .B(vdd_), .G(vdd_cntl_r[90]),
     .S(vdd_));
pch_hvt  M0_89_ ( .D(r_gnd_r[89]), .B(vdd_), .G(vdd_cntl_r[89]),
     .S(vdd_));
pch_hvt  M0_88_ ( .D(r_gnd_r[88]), .B(vdd_), .G(vdd_cntl_r[88]),
     .S(vdd_));
pch_hvt  M0_87_ ( .D(r_gnd_r[87]), .B(vdd_), .G(vdd_cntl_r[87]),
     .S(vdd_));
pch_hvt  M0_86_ ( .D(r_gnd_r[86]), .B(vdd_), .G(vdd_cntl_r[86]),
     .S(vdd_));
pch_hvt  M0_85_ ( .D(r_gnd_r[85]), .B(vdd_), .G(vdd_cntl_r[85]),
     .S(vdd_));
pch_hvt  M0_84_ ( .D(r_gnd_r[84]), .B(vdd_), .G(vdd_cntl_r[84]),
     .S(vdd_));
pch_hvt  M0_83_ ( .D(r_gnd_r[83]), .B(vdd_), .G(vdd_cntl_r[83]),
     .S(vdd_));
pch_hvt  M0_82_ ( .D(r_gnd_r[82]), .B(vdd_), .G(vdd_cntl_r[82]),
     .S(vdd_));
pch_hvt  M0_81_ ( .D(r_gnd_r[81]), .B(vdd_), .G(vdd_cntl_r[81]),
     .S(vdd_));
pch_hvt  M0_80_ ( .D(r_gnd_r[80]), .B(vdd_), .G(vdd_cntl_r[80]),
     .S(vdd_));
pch_hvt  M0_79_ ( .D(r_gnd_r[79]), .B(vdd_), .G(vdd_cntl_r[79]),
     .S(vdd_));
pch_hvt  M0_78_ ( .D(r_gnd_r[78]), .B(vdd_), .G(vdd_cntl_r[78]),
     .S(vdd_));
pch_hvt  M0_77_ ( .D(r_gnd_r[77]), .B(vdd_), .G(vdd_cntl_r[77]),
     .S(vdd_));
pch_hvt  M0_76_ ( .D(r_gnd_r[76]), .B(vdd_), .G(vdd_cntl_r[76]),
     .S(vdd_));
pch_hvt  M0_75_ ( .D(r_gnd_r[75]), .B(vdd_), .G(vdd_cntl_r[75]),
     .S(vdd_));
pch_hvt  M0_74_ ( .D(r_gnd_r[74]), .B(vdd_), .G(vdd_cntl_r[74]),
     .S(vdd_));
pch_hvt  M0_73_ ( .D(r_gnd_r[73]), .B(vdd_), .G(vdd_cntl_r[73]),
     .S(vdd_));
pch_hvt  M0_72_ ( .D(r_gnd_r[72]), .B(vdd_), .G(vdd_cntl_r[72]),
     .S(vdd_));
pch_hvt  M0_71_ ( .D(r_gnd_r[71]), .B(vdd_), .G(vdd_cntl_r[71]),
     .S(vdd_));
pch_hvt  M0_70_ ( .D(r_gnd_r[70]), .B(vdd_), .G(vdd_cntl_r[70]),
     .S(vdd_));
pch_hvt  M0_69_ ( .D(r_gnd_r[69]), .B(vdd_), .G(vdd_cntl_r[69]),
     .S(vdd_));
pch_hvt  M0_68_ ( .D(r_gnd_r[68]), .B(vdd_), .G(vdd_cntl_r[68]),
     .S(vdd_));
pch_hvt  M0_67_ ( .D(r_gnd_r[67]), .B(vdd_), .G(vdd_cntl_r[67]),
     .S(vdd_));
pch_hvt  M0_66_ ( .D(r_gnd_r[66]), .B(vdd_), .G(vdd_cntl_r[66]),
     .S(vdd_));
pch_hvt  M0_65_ ( .D(r_gnd_r[65]), .B(vdd_), .G(vdd_cntl_r[65]),
     .S(vdd_));
pch_hvt  M0_64_ ( .D(r_gnd_r[64]), .B(vdd_), .G(vdd_cntl_r[64]),
     .S(vdd_));
pch_hvt  M0_63_ ( .D(r_gnd_r[63]), .B(vdd_), .G(vdd_cntl_r[63]),
     .S(vdd_));
pch_hvt  M0_62_ ( .D(r_gnd_r[62]), .B(vdd_), .G(vdd_cntl_r[62]),
     .S(vdd_));
pch_hvt  M0_61_ ( .D(r_gnd_r[61]), .B(vdd_), .G(vdd_cntl_r[61]),
     .S(vdd_));
pch_hvt  M0_60_ ( .D(r_gnd_r[60]), .B(vdd_), .G(vdd_cntl_r[60]),
     .S(vdd_));
pch_hvt  M0_59_ ( .D(r_gnd_r[59]), .B(vdd_), .G(vdd_cntl_r[59]),
     .S(vdd_));
pch_hvt  M0_58_ ( .D(r_gnd_r[58]), .B(vdd_), .G(vdd_cntl_r[58]),
     .S(vdd_));
pch_hvt  M0_57_ ( .D(r_gnd_r[57]), .B(vdd_), .G(vdd_cntl_r[57]),
     .S(vdd_));
pch_hvt  M0_56_ ( .D(r_gnd_r[56]), .B(vdd_), .G(vdd_cntl_r[56]),
     .S(vdd_));
pch_hvt  M0_55_ ( .D(r_gnd_r[55]), .B(vdd_), .G(vdd_cntl_r[55]),
     .S(vdd_));
pch_hvt  M0_54_ ( .D(r_gnd_r[54]), .B(vdd_), .G(vdd_cntl_r[54]),
     .S(vdd_));
pch_hvt  M0_53_ ( .D(r_gnd_r[53]), .B(vdd_), .G(vdd_cntl_r[53]),
     .S(vdd_));
pch_hvt  M0_52_ ( .D(r_gnd_r[52]), .B(vdd_), .G(vdd_cntl_r[52]),
     .S(vdd_));
pch_hvt  M0_51_ ( .D(r_gnd_r[51]), .B(vdd_), .G(vdd_cntl_r[51]),
     .S(vdd_));
pch_hvt  M0_50_ ( .D(r_gnd_r[50]), .B(vdd_), .G(vdd_cntl_r[50]),
     .S(vdd_));
pch_hvt  M0_49_ ( .D(r_gnd_r[49]), .B(vdd_), .G(vdd_cntl_r[49]),
     .S(vdd_));
pch_hvt  M0_48_ ( .D(r_gnd_r[48]), .B(vdd_), .G(vdd_cntl_r[48]),
     .S(vdd_));
pch_hvt  M0_47_ ( .D(r_gnd_r[47]), .B(vdd_), .G(vdd_cntl_r[47]),
     .S(vdd_));
pch_hvt  M0_46_ ( .D(r_gnd_r[46]), .B(vdd_), .G(vdd_cntl_r[46]),
     .S(vdd_));
pch_hvt  M0_45_ ( .D(r_gnd_r[45]), .B(vdd_), .G(vdd_cntl_r[45]),
     .S(vdd_));
pch_hvt  M0_44_ ( .D(r_gnd_r[44]), .B(vdd_), .G(vdd_cntl_r[44]),
     .S(vdd_));
pch_hvt  M0_43_ ( .D(r_gnd_r[43]), .B(vdd_), .G(vdd_cntl_r[43]),
     .S(vdd_));
pch_hvt  M0_42_ ( .D(r_gnd_r[42]), .B(vdd_), .G(vdd_cntl_r[42]),
     .S(vdd_));
pch_hvt  M0_41_ ( .D(r_gnd_r[41]), .B(vdd_), .G(vdd_cntl_r[41]),
     .S(vdd_));
pch_hvt  M0_40_ ( .D(r_gnd_r[40]), .B(vdd_), .G(vdd_cntl_r[40]),
     .S(vdd_));
pch_hvt  M0_39_ ( .D(r_gnd_r[39]), .B(vdd_), .G(vdd_cntl_r[39]),
     .S(vdd_));
pch_hvt  M0_38_ ( .D(r_gnd_r[38]), .B(vdd_), .G(vdd_cntl_r[38]),
     .S(vdd_));
pch_hvt  M0_37_ ( .D(r_gnd_r[37]), .B(vdd_), .G(vdd_cntl_r[37]),
     .S(vdd_));
pch_hvt  M0_36_ ( .D(r_gnd_r[36]), .B(vdd_), .G(vdd_cntl_r[36]),
     .S(vdd_));
pch_hvt  M0_35_ ( .D(r_gnd_r[35]), .B(vdd_), .G(vdd_cntl_r[35]),
     .S(vdd_));
pch_hvt  M0_34_ ( .D(r_gnd_r[34]), .B(vdd_), .G(vdd_cntl_r[34]),
     .S(vdd_));
pch_hvt  M0_33_ ( .D(r_gnd_r[33]), .B(vdd_), .G(vdd_cntl_r[33]),
     .S(vdd_));
pch_hvt  M0_32_ ( .D(r_gnd_r[32]), .B(vdd_), .G(vdd_cntl_r[32]),
     .S(vdd_));
pch_hvt  M0_31_ ( .D(r_gnd_r[31]), .B(vdd_), .G(vdd_cntl_r[31]),
     .S(vdd_));
pch_hvt  M0_30_ ( .D(r_gnd_r[30]), .B(vdd_), .G(vdd_cntl_r[30]),
     .S(vdd_));
pch_hvt  M0_29_ ( .D(r_gnd_r[29]), .B(vdd_), .G(vdd_cntl_r[29]),
     .S(vdd_));
pch_hvt  M0_28_ ( .D(r_gnd_r[28]), .B(vdd_), .G(vdd_cntl_r[28]),
     .S(vdd_));
pch_hvt  M0_27_ ( .D(r_gnd_r[27]), .B(vdd_), .G(vdd_cntl_r[27]),
     .S(vdd_));
pch_hvt  M0_26_ ( .D(r_gnd_r[26]), .B(vdd_), .G(vdd_cntl_r[26]),
     .S(vdd_));
pch_hvt  M0_25_ ( .D(r_gnd_r[25]), .B(vdd_), .G(vdd_cntl_r[25]),
     .S(vdd_));
pch_hvt  M0_24_ ( .D(r_gnd_r[24]), .B(vdd_), .G(vdd_cntl_r[24]),
     .S(vdd_));
pch_hvt  M0_23_ ( .D(r_gnd_r[23]), .B(vdd_), .G(vdd_cntl_r[23]),
     .S(vdd_));
pch_hvt  M0_22_ ( .D(r_gnd_r[22]), .B(vdd_), .G(vdd_cntl_r[22]),
     .S(vdd_));
pch_hvt  M0_21_ ( .D(r_gnd_r[21]), .B(vdd_), .G(vdd_cntl_r[21]),
     .S(vdd_));
pch_hvt  M0_20_ ( .D(r_gnd_r[20]), .B(vdd_), .G(vdd_cntl_r[20]),
     .S(vdd_));
pch_hvt  M0_19_ ( .D(r_gnd_r[19]), .B(vdd_), .G(vdd_cntl_r[19]),
     .S(vdd_));
pch_hvt  M0_18_ ( .D(r_gnd_r[18]), .B(vdd_), .G(vdd_cntl_r[18]),
     .S(vdd_));
pch_hvt  M0_17_ ( .D(r_gnd_r[17]), .B(vdd_), .G(vdd_cntl_r[17]),
     .S(vdd_));
pch_hvt  M0_16_ ( .D(r_gnd_r[16]), .B(vdd_), .G(vdd_cntl_r[16]),
     .S(vdd_));
pch_hvt  M0_15_ ( .D(r_gnd_r[15]), .B(vdd_), .G(vdd_cntl_r[15]),
     .S(vdd_));
pch_hvt  M0_14_ ( .D(r_gnd_r[14]), .B(vdd_), .G(vdd_cntl_r[14]),
     .S(vdd_));
pch_hvt  M0_13_ ( .D(r_gnd_r[13]), .B(vdd_), .G(vdd_cntl_r[13]),
     .S(vdd_));
pch_hvt  M0_12_ ( .D(r_gnd_r[12]), .B(vdd_), .G(vdd_cntl_r[12]),
     .S(vdd_));
pch_hvt  M0_11_ ( .D(r_gnd_r[11]), .B(vdd_), .G(vdd_cntl_r[11]),
     .S(vdd_));
pch_hvt  M0_10_ ( .D(r_gnd_r[10]), .B(vdd_), .G(vdd_cntl_r[10]),
     .S(vdd_));
pch_hvt  M0_9_ ( .D(r_gnd_r[9]), .B(vdd_), .G(vdd_cntl_r[9]),
     .S(vdd_));
pch_hvt  M0_8_ ( .D(r_gnd_r[8]), .B(vdd_), .G(vdd_cntl_r[8]),
     .S(vdd_));
pch_hvt  M0_7_ ( .D(r_gnd_r[7]), .B(vdd_), .G(vdd_cntl_r[7]),
     .S(vdd_));
pch_hvt  M0_6_ ( .D(r_gnd_r[6]), .B(vdd_), .G(vdd_cntl_r[6]),
     .S(vdd_));
pch_hvt  M0_5_ ( .D(r_gnd_r[5]), .B(vdd_), .G(vdd_cntl_r[5]),
     .S(vdd_));
pch_hvt  M0_4_ ( .D(r_gnd_r[4]), .B(vdd_), .G(vdd_cntl_r[4]),
     .S(vdd_));
pch_hvt  M0_3_ ( .D(r_gnd_r[3]), .B(vdd_), .G(vdd_cntl_r[3]),
     .S(vdd_));
pch_hvt  M0_2_ ( .D(r_gnd_r[2]), .B(vdd_), .G(vdd_cntl_r[2]),
     .S(vdd_));
pch_hvt  M0_1_ ( .D(r_gnd_r[1]), .B(vdd_), .G(vdd_cntl_r[1]),
     .S(vdd_));
pch_hvt  M0_0_ ( .D(r_gnd_r[0]), .B(vdd_), .G(vdd_cntl_r[0]),
     .S(vdd_));
pch_hvt  M3_141_ ( .D(r_gnd_l[141]), .B(vdd_), .G(vdd_cntl_l[141]),
     .S(vdd_));
pch_hvt  M3_140_ ( .D(r_gnd_l[140]), .B(vdd_), .G(vdd_cntl_l[140]),
     .S(vdd_));
pch_hvt  M3_139_ ( .D(r_gnd_l[139]), .B(vdd_), .G(vdd_cntl_l[139]),
     .S(vdd_));
pch_hvt  M3_138_ ( .D(r_gnd_l[138]), .B(vdd_), .G(vdd_cntl_l[138]),
     .S(vdd_));
pch_hvt  M3_137_ ( .D(r_gnd_l[137]), .B(vdd_), .G(vdd_cntl_l[137]),
     .S(vdd_));
pch_hvt  M3_136_ ( .D(r_gnd_l[136]), .B(vdd_), .G(vdd_cntl_l[136]),
     .S(vdd_));
pch_hvt  M3_135_ ( .D(r_gnd_l[135]), .B(vdd_), .G(vdd_cntl_l[135]),
     .S(vdd_));
pch_hvt  M3_134_ ( .D(r_gnd_l[134]), .B(vdd_), .G(vdd_cntl_l[134]),
     .S(vdd_));
pch_hvt  M3_133_ ( .D(r_gnd_l[133]), .B(vdd_), .G(vdd_cntl_l[133]),
     .S(vdd_));
pch_hvt  M3_132_ ( .D(r_gnd_l[132]), .B(vdd_), .G(vdd_cntl_l[132]),
     .S(vdd_));
pch_hvt  M3_131_ ( .D(r_gnd_l[131]), .B(vdd_), .G(vdd_cntl_l[131]),
     .S(vdd_));
pch_hvt  M3_130_ ( .D(r_gnd_l[130]), .B(vdd_), .G(vdd_cntl_l[130]),
     .S(vdd_));
pch_hvt  M3_129_ ( .D(r_gnd_l[129]), .B(vdd_), .G(vdd_cntl_l[129]),
     .S(vdd_));
pch_hvt  M3_128_ ( .D(r_gnd_l[128]), .B(vdd_), .G(vdd_cntl_l[128]),
     .S(vdd_));
pch_hvt  M3_127_ ( .D(r_gnd_l[127]), .B(vdd_), .G(vdd_cntl_l[127]),
     .S(vdd_));
pch_hvt  M3_126_ ( .D(r_gnd_l[126]), .B(vdd_), .G(vdd_cntl_l[126]),
     .S(vdd_));
pch_hvt  M3_125_ ( .D(r_gnd_l[125]), .B(vdd_), .G(vdd_cntl_l[125]),
     .S(vdd_));
pch_hvt  M3_124_ ( .D(r_gnd_l[124]), .B(vdd_), .G(vdd_cntl_l[124]),
     .S(vdd_));
pch_hvt  M3_123_ ( .D(r_gnd_l[123]), .B(vdd_), .G(vdd_cntl_l[123]),
     .S(vdd_));
pch_hvt  M3_122_ ( .D(r_gnd_l[122]), .B(vdd_), .G(vdd_cntl_l[122]),
     .S(vdd_));
pch_hvt  M3_121_ ( .D(r_gnd_l[121]), .B(vdd_), .G(vdd_cntl_l[121]),
     .S(vdd_));
pch_hvt  M3_120_ ( .D(r_gnd_l[120]), .B(vdd_), .G(vdd_cntl_l[120]),
     .S(vdd_));
pch_hvt  M3_119_ ( .D(r_gnd_l[119]), .B(vdd_), .G(vdd_cntl_l[119]),
     .S(vdd_));
pch_hvt  M3_118_ ( .D(r_gnd_l[118]), .B(vdd_), .G(vdd_cntl_l[118]),
     .S(vdd_));
pch_hvt  M3_117_ ( .D(r_gnd_l[117]), .B(vdd_), .G(vdd_cntl_l[117]),
     .S(vdd_));
pch_hvt  M3_116_ ( .D(r_gnd_l[116]), .B(vdd_), .G(vdd_cntl_l[116]),
     .S(vdd_));
pch_hvt  M3_115_ ( .D(r_gnd_l[115]), .B(vdd_), .G(vdd_cntl_l[115]),
     .S(vdd_));
pch_hvt  M3_114_ ( .D(r_gnd_l[114]), .B(vdd_), .G(vdd_cntl_l[114]),
     .S(vdd_));
pch_hvt  M3_113_ ( .D(r_gnd_l[113]), .B(vdd_), .G(vdd_cntl_l[113]),
     .S(vdd_));
pch_hvt  M3_112_ ( .D(r_gnd_l[112]), .B(vdd_), .G(vdd_cntl_l[112]),
     .S(vdd_));
pch_hvt  M3_111_ ( .D(r_gnd_l[111]), .B(vdd_), .G(vdd_cntl_l[111]),
     .S(vdd_));
pch_hvt  M3_110_ ( .D(r_gnd_l[110]), .B(vdd_), .G(vdd_cntl_l[110]),
     .S(vdd_));
pch_hvt  M3_109_ ( .D(r_gnd_l[109]), .B(vdd_), .G(vdd_cntl_l[109]),
     .S(vdd_));
pch_hvt  M3_108_ ( .D(r_gnd_l[108]), .B(vdd_), .G(vdd_cntl_l[108]),
     .S(vdd_));
pch_hvt  M3_107_ ( .D(r_gnd_l[107]), .B(vdd_), .G(vdd_cntl_l[107]),
     .S(vdd_));
pch_hvt  M3_106_ ( .D(r_gnd_l[106]), .B(vdd_), .G(vdd_cntl_l[106]),
     .S(vdd_));
pch_hvt  M3_105_ ( .D(r_gnd_l[105]), .B(vdd_), .G(vdd_cntl_l[105]),
     .S(vdd_));
pch_hvt  M3_104_ ( .D(r_gnd_l[104]), .B(vdd_), .G(vdd_cntl_l[104]),
     .S(vdd_));
pch_hvt  M3_103_ ( .D(r_gnd_l[103]), .B(vdd_), .G(vdd_cntl_l[103]),
     .S(vdd_));
pch_hvt  M3_102_ ( .D(r_gnd_l[102]), .B(vdd_), .G(vdd_cntl_l[102]),
     .S(vdd_));
pch_hvt  M3_101_ ( .D(r_gnd_l[101]), .B(vdd_), .G(vdd_cntl_l[101]),
     .S(vdd_));
pch_hvt  M3_100_ ( .D(r_gnd_l[100]), .B(vdd_), .G(vdd_cntl_l[100]),
     .S(vdd_));
pch_hvt  M3_99_ ( .D(r_gnd_l[99]), .B(vdd_), .G(vdd_cntl_l[99]),
     .S(vdd_));
pch_hvt  M3_98_ ( .D(r_gnd_l[98]), .B(vdd_), .G(vdd_cntl_l[98]),
     .S(vdd_));
pch_hvt  M3_97_ ( .D(r_gnd_l[97]), .B(vdd_), .G(vdd_cntl_l[97]),
     .S(vdd_));
pch_hvt  M3_96_ ( .D(r_gnd_l[96]), .B(vdd_), .G(vdd_cntl_l[96]),
     .S(vdd_));
pch_hvt  M3_95_ ( .D(r_gnd_l[95]), .B(vdd_), .G(vdd_cntl_l[95]),
     .S(vdd_));
pch_hvt  M3_94_ ( .D(r_gnd_l[94]), .B(vdd_), .G(vdd_cntl_l[94]),
     .S(vdd_));
pch_hvt  M3_93_ ( .D(r_gnd_l[93]), .B(vdd_), .G(vdd_cntl_l[93]),
     .S(vdd_));
pch_hvt  M3_92_ ( .D(r_gnd_l[92]), .B(vdd_), .G(vdd_cntl_l[92]),
     .S(vdd_));
pch_hvt  M3_91_ ( .D(r_gnd_l[91]), .B(vdd_), .G(vdd_cntl_l[91]),
     .S(vdd_));
pch_hvt  M3_90_ ( .D(r_gnd_l[90]), .B(vdd_), .G(vdd_cntl_l[90]),
     .S(vdd_));
pch_hvt  M3_89_ ( .D(r_gnd_l[89]), .B(vdd_), .G(vdd_cntl_l[89]),
     .S(vdd_));
pch_hvt  M3_88_ ( .D(r_gnd_l[88]), .B(vdd_), .G(vdd_cntl_l[88]),
     .S(vdd_));
pch_hvt  M3_87_ ( .D(r_gnd_l[87]), .B(vdd_), .G(vdd_cntl_l[87]),
     .S(vdd_));
pch_hvt  M3_86_ ( .D(r_gnd_l[86]), .B(vdd_), .G(vdd_cntl_l[86]),
     .S(vdd_));
pch_hvt  M3_85_ ( .D(r_gnd_l[85]), .B(vdd_), .G(vdd_cntl_l[85]),
     .S(vdd_));
pch_hvt  M3_84_ ( .D(r_gnd_l[84]), .B(vdd_), .G(vdd_cntl_l[84]),
     .S(vdd_));
pch_hvt  M3_83_ ( .D(r_gnd_l[83]), .B(vdd_), .G(vdd_cntl_l[83]),
     .S(vdd_));
pch_hvt  M3_82_ ( .D(r_gnd_l[82]), .B(vdd_), .G(vdd_cntl_l[82]),
     .S(vdd_));
pch_hvt  M3_81_ ( .D(r_gnd_l[81]), .B(vdd_), .G(vdd_cntl_l[81]),
     .S(vdd_));
pch_hvt  M3_80_ ( .D(r_gnd_l[80]), .B(vdd_), .G(vdd_cntl_l[80]),
     .S(vdd_));
pch_hvt  M3_79_ ( .D(r_gnd_l[79]), .B(vdd_), .G(vdd_cntl_l[79]),
     .S(vdd_));
pch_hvt  M3_78_ ( .D(r_gnd_l[78]), .B(vdd_), .G(vdd_cntl_l[78]),
     .S(vdd_));
pch_hvt  M3_77_ ( .D(r_gnd_l[77]), .B(vdd_), .G(vdd_cntl_l[77]),
     .S(vdd_));
pch_hvt  M3_76_ ( .D(r_gnd_l[76]), .B(vdd_), .G(vdd_cntl_l[76]),
     .S(vdd_));
pch_hvt  M3_75_ ( .D(r_gnd_l[75]), .B(vdd_), .G(vdd_cntl_l[75]),
     .S(vdd_));
pch_hvt  M3_74_ ( .D(r_gnd_l[74]), .B(vdd_), .G(vdd_cntl_l[74]),
     .S(vdd_));
pch_hvt  M3_73_ ( .D(r_gnd_l[73]), .B(vdd_), .G(vdd_cntl_l[73]),
     .S(vdd_));
pch_hvt  M3_72_ ( .D(r_gnd_l[72]), .B(vdd_), .G(vdd_cntl_l[72]),
     .S(vdd_));
pch_hvt  M3_71_ ( .D(r_gnd_l[71]), .B(vdd_), .G(vdd_cntl_l[71]),
     .S(vdd_));
pch_hvt  M3_70_ ( .D(r_gnd_l[70]), .B(vdd_), .G(vdd_cntl_l[70]),
     .S(vdd_));
pch_hvt  M3_69_ ( .D(r_gnd_l[69]), .B(vdd_), .G(vdd_cntl_l[69]),
     .S(vdd_));
pch_hvt  M3_68_ ( .D(r_gnd_l[68]), .B(vdd_), .G(vdd_cntl_l[68]),
     .S(vdd_));
pch_hvt  M3_67_ ( .D(r_gnd_l[67]), .B(vdd_), .G(vdd_cntl_l[67]),
     .S(vdd_));
pch_hvt  M3_66_ ( .D(r_gnd_l[66]), .B(vdd_), .G(vdd_cntl_l[66]),
     .S(vdd_));
pch_hvt  M3_65_ ( .D(r_gnd_l[65]), .B(vdd_), .G(vdd_cntl_l[65]),
     .S(vdd_));
pch_hvt  M3_64_ ( .D(r_gnd_l[64]), .B(vdd_), .G(vdd_cntl_l[64]),
     .S(vdd_));
pch_hvt  M3_63_ ( .D(r_gnd_l[63]), .B(vdd_), .G(vdd_cntl_l[63]),
     .S(vdd_));
pch_hvt  M3_62_ ( .D(r_gnd_l[62]), .B(vdd_), .G(vdd_cntl_l[62]),
     .S(vdd_));
pch_hvt  M3_61_ ( .D(r_gnd_l[61]), .B(vdd_), .G(vdd_cntl_l[61]),
     .S(vdd_));
pch_hvt  M3_60_ ( .D(r_gnd_l[60]), .B(vdd_), .G(vdd_cntl_l[60]),
     .S(vdd_));
pch_hvt  M3_59_ ( .D(r_gnd_l[59]), .B(vdd_), .G(vdd_cntl_l[59]),
     .S(vdd_));
pch_hvt  M3_58_ ( .D(r_gnd_l[58]), .B(vdd_), .G(vdd_cntl_l[58]),
     .S(vdd_));
pch_hvt  M3_57_ ( .D(r_gnd_l[57]), .B(vdd_), .G(vdd_cntl_l[57]),
     .S(vdd_));
pch_hvt  M3_56_ ( .D(r_gnd_l[56]), .B(vdd_), .G(vdd_cntl_l[56]),
     .S(vdd_));
pch_hvt  M3_55_ ( .D(r_gnd_l[55]), .B(vdd_), .G(vdd_cntl_l[55]),
     .S(vdd_));
pch_hvt  M3_54_ ( .D(r_gnd_l[54]), .B(vdd_), .G(vdd_cntl_l[54]),
     .S(vdd_));
pch_hvt  M3_53_ ( .D(r_gnd_l[53]), .B(vdd_), .G(vdd_cntl_l[53]),
     .S(vdd_));
pch_hvt  M3_52_ ( .D(r_gnd_l[52]), .B(vdd_), .G(vdd_cntl_l[52]),
     .S(vdd_));
pch_hvt  M3_51_ ( .D(r_gnd_l[51]), .B(vdd_), .G(vdd_cntl_l[51]),
     .S(vdd_));
pch_hvt  M3_50_ ( .D(r_gnd_l[50]), .B(vdd_), .G(vdd_cntl_l[50]),
     .S(vdd_));
pch_hvt  M3_49_ ( .D(r_gnd_l[49]), .B(vdd_), .G(vdd_cntl_l[49]),
     .S(vdd_));
pch_hvt  M3_48_ ( .D(r_gnd_l[48]), .B(vdd_), .G(vdd_cntl_l[48]),
     .S(vdd_));
pch_hvt  M3_47_ ( .D(r_gnd_l[47]), .B(vdd_), .G(vdd_cntl_l[47]),
     .S(vdd_));
pch_hvt  M3_46_ ( .D(r_gnd_l[46]), .B(vdd_), .G(vdd_cntl_l[46]),
     .S(vdd_));
pch_hvt  M3_45_ ( .D(r_gnd_l[45]), .B(vdd_), .G(vdd_cntl_l[45]),
     .S(vdd_));
pch_hvt  M3_44_ ( .D(r_gnd_l[44]), .B(vdd_), .G(vdd_cntl_l[44]),
     .S(vdd_));
pch_hvt  M3_43_ ( .D(r_gnd_l[43]), .B(vdd_), .G(vdd_cntl_l[43]),
     .S(vdd_));
pch_hvt  M3_42_ ( .D(r_gnd_l[42]), .B(vdd_), .G(vdd_cntl_l[42]),
     .S(vdd_));
pch_hvt  M3_41_ ( .D(r_gnd_l[41]), .B(vdd_), .G(vdd_cntl_l[41]),
     .S(vdd_));
pch_hvt  M3_40_ ( .D(r_gnd_l[40]), .B(vdd_), .G(vdd_cntl_l[40]),
     .S(vdd_));
pch_hvt  M3_39_ ( .D(r_gnd_l[39]), .B(vdd_), .G(vdd_cntl_l[39]),
     .S(vdd_));
pch_hvt  M3_38_ ( .D(r_gnd_l[38]), .B(vdd_), .G(vdd_cntl_l[38]),
     .S(vdd_));
pch_hvt  M3_37_ ( .D(r_gnd_l[37]), .B(vdd_), .G(vdd_cntl_l[37]),
     .S(vdd_));
pch_hvt  M3_36_ ( .D(r_gnd_l[36]), .B(vdd_), .G(vdd_cntl_l[36]),
     .S(vdd_));
pch_hvt  M3_35_ ( .D(r_gnd_l[35]), .B(vdd_), .G(vdd_cntl_l[35]),
     .S(vdd_));
pch_hvt  M3_34_ ( .D(r_gnd_l[34]), .B(vdd_), .G(vdd_cntl_l[34]),
     .S(vdd_));
pch_hvt  M3_33_ ( .D(r_gnd_l[33]), .B(vdd_), .G(vdd_cntl_l[33]),
     .S(vdd_));
pch_hvt  M3_32_ ( .D(r_gnd_l[32]), .B(vdd_), .G(vdd_cntl_l[32]),
     .S(vdd_));
pch_hvt  M3_31_ ( .D(r_gnd_l[31]), .B(vdd_), .G(vdd_cntl_l[31]),
     .S(vdd_));
pch_hvt  M3_30_ ( .D(r_gnd_l[30]), .B(vdd_), .G(vdd_cntl_l[30]),
     .S(vdd_));
pch_hvt  M3_29_ ( .D(r_gnd_l[29]), .B(vdd_), .G(vdd_cntl_l[29]),
     .S(vdd_));
pch_hvt  M3_28_ ( .D(r_gnd_l[28]), .B(vdd_), .G(vdd_cntl_l[28]),
     .S(vdd_));
pch_hvt  M3_27_ ( .D(r_gnd_l[27]), .B(vdd_), .G(vdd_cntl_l[27]),
     .S(vdd_));
pch_hvt  M3_26_ ( .D(r_gnd_l[26]), .B(vdd_), .G(vdd_cntl_l[26]),
     .S(vdd_));
pch_hvt  M3_25_ ( .D(r_gnd_l[25]), .B(vdd_), .G(vdd_cntl_l[25]),
     .S(vdd_));
pch_hvt  M3_24_ ( .D(r_gnd_l[24]), .B(vdd_), .G(vdd_cntl_l[24]),
     .S(vdd_));
pch_hvt  M3_23_ ( .D(r_gnd_l[23]), .B(vdd_), .G(vdd_cntl_l[23]),
     .S(vdd_));
pch_hvt  M3_22_ ( .D(r_gnd_l[22]), .B(vdd_), .G(vdd_cntl_l[22]),
     .S(vdd_));
pch_hvt  M3_21_ ( .D(r_gnd_l[21]), .B(vdd_), .G(vdd_cntl_l[21]),
     .S(vdd_));
pch_hvt  M3_20_ ( .D(r_gnd_l[20]), .B(vdd_), .G(vdd_cntl_l[20]),
     .S(vdd_));
pch_hvt  M3_19_ ( .D(r_gnd_l[19]), .B(vdd_), .G(vdd_cntl_l[19]),
     .S(vdd_));
pch_hvt  M3_18_ ( .D(r_gnd_l[18]), .B(vdd_), .G(vdd_cntl_l[18]),
     .S(vdd_));
pch_hvt  M3_17_ ( .D(r_gnd_l[17]), .B(vdd_), .G(vdd_cntl_l[17]),
     .S(vdd_));
pch_hvt  M3_16_ ( .D(r_gnd_l[16]), .B(vdd_), .G(vdd_cntl_l[16]),
     .S(vdd_));
pch_hvt  M3_15_ ( .D(r_gnd_l[15]), .B(vdd_), .G(vdd_cntl_l[15]),
     .S(vdd_));
pch_hvt  M3_14_ ( .D(r_gnd_l[14]), .B(vdd_), .G(vdd_cntl_l[14]),
     .S(vdd_));
pch_hvt  M3_13_ ( .D(r_gnd_l[13]), .B(vdd_), .G(vdd_cntl_l[13]),
     .S(vdd_));
pch_hvt  M3_12_ ( .D(r_gnd_l[12]), .B(vdd_), .G(vdd_cntl_l[12]),
     .S(vdd_));
pch_hvt  M3_11_ ( .D(r_gnd_l[11]), .B(vdd_), .G(vdd_cntl_l[11]),
     .S(vdd_));
pch_hvt  M3_10_ ( .D(r_gnd_l[10]), .B(vdd_), .G(vdd_cntl_l[10]),
     .S(vdd_));
pch_hvt  M3_9_ ( .D(r_gnd_l[9]), .B(vdd_), .G(vdd_cntl_l[9]),
     .S(vdd_));
pch_hvt  M3_8_ ( .D(r_gnd_l[8]), .B(vdd_), .G(vdd_cntl_l[8]),
     .S(vdd_));
pch_hvt  M3_7_ ( .D(r_gnd_l[7]), .B(vdd_), .G(vdd_cntl_l[7]),
     .S(vdd_));
pch_hvt  M3_6_ ( .D(r_gnd_l[6]), .B(vdd_), .G(vdd_cntl_l[6]),
     .S(vdd_));
pch_hvt  M3_5_ ( .D(r_gnd_l[5]), .B(vdd_), .G(vdd_cntl_l[5]),
     .S(vdd_));
pch_hvt  M3_4_ ( .D(r_gnd_l[4]), .B(vdd_), .G(vdd_cntl_l[4]),
     .S(vdd_));
pch_hvt  M3_3_ ( .D(r_gnd_l[3]), .B(vdd_), .G(vdd_cntl_l[3]),
     .S(vdd_));
pch_hvt  M3_2_ ( .D(r_gnd_l[2]), .B(vdd_), .G(vdd_cntl_l[2]),
     .S(vdd_));
pch_hvt  M3_1_ ( .D(r_gnd_l[1]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  M3_0_ ( .D(r_gnd_l[0]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));
cram_2x2x2_ice8p I_mem2x2x2t_70_ ( .wl_r(wl_r[141:140]),
     .wl_l(wl_l[141:140]), .reset_r(reset_r[141:140]),
     .reset_l(reset_l[141:140]), .pgate_r(pgate_r[141:140]),
     .pgate_l(pgate_l[141:140]), .q_b({net35[0], net35[1], net35[2],
     net35[3], net35[4], net35[5], net35[6], net35[7]}), .q({net36[0],
     net36[1], net36[2], net36[3], net36[4], net36[5], net36[6],
     net36[7]}), .bl(bl[3:0]), .r_gnd_l(r_gnd_l[141:140]),
     .r_gnd_r(r_gnd_r[141:140]));
cram_2x2x2_ice8p I_mem2x2x2t_69_ ( .wl_r(wl_r[139:138]),
     .wl_l(wl_l[139:138]), .reset_r(reset_r[139:138]),
     .reset_l(reset_l[139:138]), .pgate_r(pgate_r[139:138]),
     .pgate_l(pgate_l[139:138]), .q_b({net35[8], net35[9], net35[10],
     net35[11], net35[12], net35[13], net35[14], net35[15]}),
     .q({net36[8], net36[9], net36[10], net36[11], net36[12],
     net36[13], net36[14], net36[15]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[139:138]), .r_gnd_r(r_gnd_r[139:138]));
cram_2x2x2_ice8p I_mem2x2x2t_68_ ( .wl_r(wl_r[137:136]),
     .wl_l(wl_l[137:136]), .reset_r(reset_r[137:136]),
     .reset_l(reset_l[137:136]), .pgate_r(pgate_r[137:136]),
     .pgate_l(pgate_l[137:136]), .q_b({net35[16], net35[17], net35[18],
     net35[19], net35[20], net35[21], net35[22], net35[23]}),
     .q({net36[16], net36[17], net36[18], net36[19], net36[20],
     net36[21], net36[22], net36[23]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[137:136]), .r_gnd_r(r_gnd_r[137:136]));
cram_2x2x2_ice8p I_mem2x2x2t_67_ ( .wl_r(wl_r[135:134]),
     .wl_l(wl_l[135:134]), .reset_r(reset_r[135:134]),
     .reset_l(reset_l[135:134]), .pgate_r(pgate_r[135:134]),
     .pgate_l(pgate_l[135:134]), .q_b({net35[24], net35[25], net35[26],
     net35[27], net35[28], net35[29], net35[30], net35[31]}),
     .q({net36[24], net36[25], net36[26], net36[27], net36[28],
     net36[29], net36[30], net36[31]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[135:134]), .r_gnd_r(r_gnd_r[135:134]));
cram_2x2x2_ice8p I_mem2x2x2t_66_ ( .wl_r(wl_r[133:132]),
     .wl_l(wl_l[133:132]), .reset_r(reset_r[133:132]),
     .reset_l(reset_l[133:132]), .pgate_r(pgate_r[133:132]),
     .pgate_l(pgate_l[133:132]), .q_b({net35[32], net35[33], net35[34],
     net35[35], net35[36], net35[37], net35[38], net35[39]}),
     .q({net36[32], net36[33], net36[34], net36[35], net36[36],
     net36[37], net36[38], net36[39]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[133:132]), .r_gnd_r(r_gnd_r[133:132]));
cram_2x2x2_ice8p I_mem2x2x2t_65_ ( .wl_r(wl_r[131:130]),
     .wl_l(wl_l[131:130]), .reset_r(reset_r[131:130]),
     .reset_l(reset_l[131:130]), .pgate_r(pgate_r[131:130]),
     .pgate_l(pgate_l[131:130]), .q_b({net35[40], net35[41], net35[42],
     net35[43], net35[44], net35[45], net35[46], net35[47]}),
     .q({net36[40], net36[41], net36[42], net36[43], net36[44],
     net36[45], net36[46], net36[47]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[131:130]), .r_gnd_r(r_gnd_r[131:130]));
cram_2x2x2_ice8p I_mem2x2x2t_64_ ( .wl_r(wl_r[129:128]),
     .wl_l(wl_l[129:128]), .reset_r(reset_r[129:128]),
     .reset_l(reset_l[129:128]), .pgate_r(pgate_r[129:128]),
     .pgate_l(pgate_l[129:128]), .q_b({net35[48], net35[49], net35[50],
     net35[51], net35[52], net35[53], net35[54], net35[55]}),
     .q({net36[48], net36[49], net36[50], net36[51], net36[52],
     net36[53], net36[54], net36[55]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[129:128]), .r_gnd_r(r_gnd_r[129:128]));
cram_2x2x2_ice8p I_mem2x2x2t_63_ ( .wl_r(wl_r[127:126]),
     .wl_l(wl_l[127:126]), .reset_r(reset_r[127:126]),
     .reset_l(reset_l[127:126]), .pgate_r(pgate_r[127:126]),
     .pgate_l(pgate_l[127:126]), .q_b({net35[56], net35[57], net35[58],
     net35[59], net35[60], net35[61], net35[62], net35[63]}),
     .q({net36[56], net36[57], net36[58], net36[59], net36[60],
     net36[61], net36[62], net36[63]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[127:126]), .r_gnd_r(r_gnd_r[127:126]));
cram_2x2x2_ice8p I_mem2x2x2t_62_ ( .wl_r(wl_r[125:124]),
     .wl_l(wl_l[125:124]), .reset_r(reset_r[125:124]),
     .reset_l(reset_l[125:124]), .pgate_r(pgate_r[125:124]),
     .pgate_l(pgate_l[125:124]), .q_b({net35[64], net35[65], net35[66],
     net35[67], net35[68], net35[69], net35[70], net35[71]}),
     .q({net36[64], net36[65], net36[66], net36[67], net36[68],
     net36[69], net36[70], net36[71]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[125:124]), .r_gnd_r(r_gnd_r[125:124]));
cram_2x2x2_ice8p I_mem2x2x2t_61_ ( .wl_r(wl_r[123:122]),
     .wl_l(wl_l[123:122]), .reset_r(reset_r[123:122]),
     .reset_l(reset_l[123:122]), .pgate_r(pgate_r[123:122]),
     .pgate_l(pgate_l[123:122]), .q_b({net35[72], net35[73], net35[74],
     net35[75], net35[76], net35[77], net35[78], net35[79]}),
     .q({net36[72], net36[73], net36[74], net36[75], net36[76],
     net36[77], net36[78], net36[79]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[123:122]), .r_gnd_r(r_gnd_r[123:122]));
cram_2x2x2_ice8p I_mem2x2x2t_60_ ( .wl_r(wl_r[121:120]),
     .wl_l(wl_l[121:120]), .reset_r(reset_r[121:120]),
     .reset_l(reset_l[121:120]), .pgate_r(pgate_r[121:120]),
     .pgate_l(pgate_l[121:120]), .q_b({net35[80], net35[81], net35[82],
     net35[83], net35[84], net35[85], net35[86], net35[87]}),
     .q({net36[80], net36[81], net36[82], net36[83], net36[84],
     net36[85], net36[86], net36[87]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[121:120]), .r_gnd_r(r_gnd_r[121:120]));
cram_2x2x2_ice8p I_mem2x2x2t_59_ ( .wl_r(wl_r[119:118]),
     .wl_l(wl_l[119:118]), .reset_r(reset_r[119:118]),
     .reset_l(reset_l[119:118]), .pgate_r(pgate_r[119:118]),
     .pgate_l(pgate_l[119:118]), .q_b({net35[88], net35[89], net35[90],
     net35[91], net35[92], net35[93], net35[94], net35[95]}),
     .q({net36[88], net36[89], net36[90], net36[91], net36[92],
     net36[93], net36[94], net36[95]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[119:118]), .r_gnd_r(r_gnd_r[119:118]));
cram_2x2x2_ice8p I_mem2x2x2t_58_ ( .wl_r(wl_r[117:116]),
     .wl_l(wl_l[117:116]), .reset_r(reset_r[117:116]),
     .reset_l(reset_l[117:116]), .pgate_r(pgate_r[117:116]),
     .pgate_l(pgate_l[117:116]), .q_b({net35[96], net35[97], net35[98],
     net35[99], net35[100], net35[101], net35[102], net35[103]}),
     .q({net36[96], net36[97], net36[98], net36[99], net36[100],
     net36[101], net36[102], net36[103]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[117:116]), .r_gnd_r(r_gnd_r[117:116]));
cram_2x2x2_ice8p I_mem2x2x2t_57_ ( .wl_r(wl_r[115:114]),
     .wl_l(wl_l[115:114]), .reset_r(reset_r[115:114]),
     .reset_l(reset_l[115:114]), .pgate_r(pgate_r[115:114]),
     .pgate_l(pgate_l[115:114]), .q_b({net35[104], net35[105],
     net35[106], net35[107], net35[108], net35[109], net35[110],
     net35[111]}), .q({net36[104], net36[105], net36[106], net36[107],
     net36[108], net36[109], net36[110], net36[111]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[115:114]), .r_gnd_r(r_gnd_r[115:114]));
cram_2x2x2_ice8p I_mem2x2x2t_56_ ( .wl_r(wl_r[113:112]),
     .wl_l(wl_l[113:112]), .reset_r(reset_r[113:112]),
     .reset_l(reset_l[113:112]), .pgate_r(pgate_r[113:112]),
     .pgate_l(pgate_l[113:112]), .q_b({net35[112], net35[113],
     net35[114], net35[115], net35[116], net35[117], net35[118],
     net35[119]}), .q({net36[112], net36[113], net36[114], net36[115],
     net36[116], net36[117], net36[118], net36[119]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[113:112]), .r_gnd_r(r_gnd_r[113:112]));
cram_2x2x2_ice8p I_mem2x2x2t_55_ ( .wl_r(wl_r[111:110]),
     .wl_l(wl_l[111:110]), .reset_r(reset_r[111:110]),
     .reset_l(reset_l[111:110]), .pgate_r(pgate_r[111:110]),
     .pgate_l(pgate_l[111:110]), .q_b({net35[120], net35[121],
     net35[122], net35[123], net35[124], net35[125], net35[126],
     net35[127]}), .q({net36[120], net36[121], net36[122], net36[123],
     net36[124], net36[125], net36[126], net36[127]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[111:110]), .r_gnd_r(r_gnd_r[111:110]));
cram_2x2x2_ice8p I_mem2x2x2t_54_ ( .wl_r(wl_r[109:108]),
     .wl_l(wl_l[109:108]), .reset_r(reset_r[109:108]),
     .reset_l(reset_l[109:108]), .pgate_r(pgate_r[109:108]),
     .pgate_l(pgate_l[109:108]), .q_b({net35[128], net35[129],
     net35[130], net35[131], net35[132], net35[133], net35[134],
     net35[135]}), .q({net36[128], net36[129], net36[130], net36[131],
     net36[132], net36[133], net36[134], net36[135]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[109:108]), .r_gnd_r(r_gnd_r[109:108]));
cram_2x2x2_ice8p I_mem2x2x2t_53_ ( .wl_r(wl_r[107:106]),
     .wl_l(wl_l[107:106]), .reset_r(reset_r[107:106]),
     .reset_l(reset_l[107:106]), .pgate_r(pgate_r[107:106]),
     .pgate_l(pgate_l[107:106]), .q_b({net35[136], net35[137],
     net35[138], net35[139], net35[140], net35[141], net35[142],
     net35[143]}), .q({net36[136], net36[137], net36[138], net36[139],
     net36[140], net36[141], net36[142], net36[143]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[107:106]), .r_gnd_r(r_gnd_r[107:106]));
cram_2x2x2_ice8p I_mem2x2x2t_52_ ( .wl_r(wl_r[105:104]),
     .wl_l(wl_l[105:104]), .reset_r(reset_r[105:104]),
     .reset_l(reset_l[105:104]), .pgate_r(pgate_r[105:104]),
     .pgate_l(pgate_l[105:104]), .q_b({net35[144], net35[145],
     net35[146], net35[147], net35[148], net35[149], net35[150],
     net35[151]}), .q({net36[144], net36[145], net36[146], net36[147],
     net36[148], net36[149], net36[150], net36[151]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[105:104]), .r_gnd_r(r_gnd_r[105:104]));
cram_2x2x2_ice8p I_mem2x2x2t_51_ ( .wl_r(wl_r[103:102]),
     .wl_l(wl_l[103:102]), .reset_r(reset_r[103:102]),
     .reset_l(reset_l[103:102]), .pgate_r(pgate_r[103:102]),
     .pgate_l(pgate_l[103:102]), .q_b({net35[152], net35[153],
     net35[154], net35[155], net35[156], net35[157], net35[158],
     net35[159]}), .q({net36[152], net36[153], net36[154], net36[155],
     net36[156], net36[157], net36[158], net36[159]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[103:102]), .r_gnd_r(r_gnd_r[103:102]));
cram_2x2x2_ice8p I_mem2x2x2t_50_ ( .wl_r(wl_r[101:100]),
     .wl_l(wl_l[101:100]), .reset_r(reset_r[101:100]),
     .reset_l(reset_l[101:100]), .pgate_r(pgate_r[101:100]),
     .pgate_l(pgate_l[101:100]), .q_b({net35[160], net35[161],
     net35[162], net35[163], net35[164], net35[165], net35[166],
     net35[167]}), .q({net36[160], net36[161], net36[162], net36[163],
     net36[164], net36[165], net36[166], net36[167]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[101:100]), .r_gnd_r(r_gnd_r[101:100]));
cram_2x2x2_ice8p I_mem2x2x2t_49_ ( .wl_r(wl_r[99:98]),
     .wl_l(wl_l[99:98]), .reset_r(reset_r[99:98]),
     .reset_l(reset_l[99:98]), .pgate_r(pgate_r[99:98]),
     .pgate_l(pgate_l[99:98]), .q_b({net35[168], net35[169],
     net35[170], net35[171], net35[172], net35[173], net35[174],
     net35[175]}), .q({net36[168], net36[169], net36[170], net36[171],
     net36[172], net36[173], net36[174], net36[175]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[99:98]), .r_gnd_r(r_gnd_r[99:98]));
cram_2x2x2_ice8p I_mem2x2x2t_48_ ( .wl_r(wl_r[97:96]),
     .wl_l(wl_l[97:96]), .reset_r(reset_r[97:96]),
     .reset_l(reset_l[97:96]), .pgate_r(pgate_r[97:96]),
     .pgate_l(pgate_l[97:96]), .q_b({net35[176], net35[177],
     net35[178], net35[179], net35[180], net35[181], net35[182],
     net35[183]}), .q({net36[176], net36[177], net36[178], net36[179],
     net36[180], net36[181], net36[182], net36[183]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[97:96]), .r_gnd_r(r_gnd_r[97:96]));
cram_2x2x2_ice8p I_mem2x2x2t_47_ ( .wl_r(wl_r[95:94]),
     .wl_l(wl_l[95:94]), .reset_r(reset_r[95:94]),
     .reset_l(reset_l[95:94]), .pgate_r(pgate_r[95:94]),
     .pgate_l(pgate_l[95:94]), .q_b({net35[184], net35[185],
     net35[186], net35[187], net35[188], net35[189], net35[190],
     net35[191]}), .q({net36[184], net36[185], net36[186], net36[187],
     net36[188], net36[189], net36[190], net36[191]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[95:94]), .r_gnd_r(r_gnd_r[95:94]));
cram_2x2x2_ice8p I_mem2x2x2t_46_ ( .wl_r(wl_r[93:92]),
     .wl_l(wl_l[93:92]), .reset_r(reset_r[93:92]),
     .reset_l(reset_l[93:92]), .pgate_r(pgate_r[93:92]),
     .pgate_l(pgate_l[93:92]), .q_b({net35[192], net35[193],
     net35[194], net35[195], net35[196], net35[197], net35[198],
     net35[199]}), .q({net36[192], net36[193], net36[194], net36[195],
     net36[196], net36[197], net36[198], net36[199]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[93:92]), .r_gnd_r(r_gnd_r[93:92]));
cram_2x2x2_ice8p I_mem2x2x2t_45_ ( .wl_r(wl_r[91:90]),
     .wl_l(wl_l[91:90]), .reset_r(reset_r[91:90]),
     .reset_l(reset_l[91:90]), .pgate_r(pgate_r[91:90]),
     .pgate_l(pgate_l[91:90]), .q_b({net35[200], net35[201],
     net35[202], net35[203], net35[204], net35[205], net35[206],
     net35[207]}), .q({net36[200], net36[201], net36[202], net36[203],
     net36[204], net36[205], net36[206], net36[207]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[91:90]), .r_gnd_r(r_gnd_r[91:90]));
cram_2x2x2_ice8p I_mem2x2x2t_44_ ( .wl_r(wl_r[89:88]),
     .wl_l(wl_l[89:88]), .reset_r(reset_r[89:88]),
     .reset_l(reset_l[89:88]), .pgate_r(pgate_r[89:88]),
     .pgate_l(pgate_l[89:88]), .q_b({net35[208], net35[209],
     net35[210], net35[211], net35[212], net35[213], net35[214],
     net35[215]}), .q({net36[208], net36[209], net36[210], net36[211],
     net36[212], net36[213], net36[214], net36[215]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[89:88]), .r_gnd_r(r_gnd_r[89:88]));
cram_2x2x2_ice8p I_mem2x2x2t_43_ ( .wl_r(wl_r[87:86]),
     .wl_l(wl_l[87:86]), .reset_r(reset_r[87:86]),
     .reset_l(reset_l[87:86]), .pgate_r(pgate_r[87:86]),
     .pgate_l(pgate_l[87:86]), .q_b({net35[216], net35[217],
     net35[218], net35[219], net35[220], net35[221], net35[222],
     net35[223]}), .q({net36[216], net36[217], net36[218], net36[219],
     net36[220], net36[221], net36[222], net36[223]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[87:86]), .r_gnd_r(r_gnd_r[87:86]));
cram_2x2x2_ice8p I_mem2x2x2t_42_ ( .wl_r(wl_r[85:84]),
     .wl_l(wl_l[85:84]), .reset_r(reset_r[85:84]),
     .reset_l(reset_l[85:84]), .pgate_r(pgate_r[85:84]),
     .pgate_l(pgate_l[85:84]), .q_b({net35[224], net35[225],
     net35[226], net35[227], net35[228], net35[229], net35[230],
     net35[231]}), .q({net36[224], net36[225], net36[226], net36[227],
     net36[228], net36[229], net36[230], net36[231]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[85:84]), .r_gnd_r(r_gnd_r[85:84]));
cram_2x2x2_ice8p I_mem2x2x2t_41_ ( .wl_r(wl_r[83:82]),
     .wl_l(wl_l[83:82]), .reset_r(reset_r[83:82]),
     .reset_l(reset_l[83:82]), .pgate_r(pgate_r[83:82]),
     .pgate_l(pgate_l[83:82]), .q_b({net35[232], net35[233],
     net35[234], net35[235], net35[236], net35[237], net35[238],
     net35[239]}), .q({net36[232], net36[233], net36[234], net36[235],
     net36[236], net36[237], net36[238], net36[239]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[83:82]), .r_gnd_r(r_gnd_r[83:82]));
cram_2x2x2_ice8p I_mem2x2x2t_40_ ( .wl_r(wl_r[81:80]),
     .wl_l(wl_l[81:80]), .reset_r(reset_r[81:80]),
     .reset_l(reset_l[81:80]), .pgate_r(pgate_r[81:80]),
     .pgate_l(pgate_l[81:80]), .q_b({net35[240], net35[241],
     net35[242], net35[243], net35[244], net35[245], net35[246],
     net35[247]}), .q({net36[240], net36[241], net36[242], net36[243],
     net36[244], net36[245], net36[246], net36[247]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[81:80]), .r_gnd_r(r_gnd_r[81:80]));
cram_2x2x2_ice8p I_mem2x2x2t_39_ ( .wl_r(wl_r[79:78]),
     .wl_l(wl_l[79:78]), .reset_r(reset_r[79:78]),
     .reset_l(reset_l[79:78]), .pgate_r(pgate_r[79:78]),
     .pgate_l(pgate_l[79:78]), .q_b({net35[248], net35[249],
     net35[250], net35[251], net35[252], net35[253], net35[254],
     net35[255]}), .q({net36[248], net36[249], net36[250], net36[251],
     net36[252], net36[253], net36[254], net36[255]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[79:78]), .r_gnd_r(r_gnd_r[79:78]));
cram_2x2x2_ice8p I_mem2x2x2t_38_ ( .wl_r(wl_r[77:76]),
     .wl_l(wl_l[77:76]), .reset_r(reset_r[77:76]),
     .reset_l(reset_l[77:76]), .pgate_r(pgate_r[77:76]),
     .pgate_l(pgate_l[77:76]), .q_b({net35[256], net35[257],
     net35[258], net35[259], net35[260], net35[261], net35[262],
     net35[263]}), .q({net36[256], net36[257], net36[258], net36[259],
     net36[260], net36[261], net36[262], net36[263]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[77:76]), .r_gnd_r(r_gnd_r[77:76]));
cram_2x2x2_ice8p I_mem2x2x2t_37_ ( .wl_r(wl_r[75:74]),
     .wl_l(wl_l[75:74]), .reset_r(reset_r[75:74]),
     .reset_l(reset_l[75:74]), .pgate_r(pgate_r[75:74]),
     .pgate_l(pgate_l[75:74]), .q_b({net35[264], net35[265],
     net35[266], net35[267], net35[268], net35[269], net35[270],
     net35[271]}), .q({net36[264], net36[265], net36[266], net36[267],
     net36[268], net36[269], net36[270], net36[271]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[75:74]), .r_gnd_r(r_gnd_r[75:74]));
cram_2x2x2_ice8p I_mem2x2x2t_36_ ( .wl_r(wl_r[73:72]),
     .wl_l(wl_l[73:72]), .reset_r(reset_r[73:72]),
     .reset_l(reset_l[73:72]), .pgate_r(pgate_r[73:72]),
     .pgate_l(pgate_l[73:72]), .q_b({net35[272], net35[273],
     net35[274], net35[275], net35[276], net35[277], net35[278],
     net35[279]}), .q({net36[272], net36[273], net36[274], net36[275],
     net36[276], net36[277], net36[278], net36[279]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[73:72]), .r_gnd_r(r_gnd_r[73:72]));
cram_2x2x2_ice8p I_mem2x2x2t_35_ ( .wl_r(wl_r[71:70]),
     .wl_l(wl_l[71:70]), .reset_r(reset_r[71:70]),
     .reset_l(reset_l[71:70]), .pgate_r(pgate_r[71:70]),
     .pgate_l(pgate_l[71:70]), .q_b({net35[280], net35[281],
     net35[282], net35[283], net35[284], net35[285], net35[286],
     net35[287]}), .q({net36[280], net36[281], net36[282], net36[283],
     net36[284], net36[285], net36[286], net36[287]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[71:70]), .r_gnd_r(r_gnd_r[71:70]));
cram_2x2x2_ice8p I_mem2x2x2t_34_ ( .wl_r(wl_r[69:68]),
     .wl_l(wl_l[69:68]), .reset_r(reset_r[69:68]),
     .reset_l(reset_l[69:68]), .pgate_r(pgate_r[69:68]),
     .pgate_l(pgate_l[69:68]), .q_b({net35[288], net35[289],
     net35[290], net35[291], net35[292], net35[293], net35[294],
     net35[295]}), .q({net36[288], net36[289], net36[290], net36[291],
     net36[292], net36[293], net36[294], net36[295]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[69:68]), .r_gnd_r(r_gnd_r[69:68]));
cram_2x2x2_ice8p I_mem2x2x2t_33_ ( .wl_r(wl_r[67:66]),
     .wl_l(wl_l[67:66]), .reset_r(reset_r[67:66]),
     .reset_l(reset_l[67:66]), .pgate_r(pgate_r[67:66]),
     .pgate_l(pgate_l[67:66]), .q_b({net35[296], net35[297],
     net35[298], net35[299], net35[300], net35[301], net35[302],
     net35[303]}), .q({net36[296], net36[297], net36[298], net36[299],
     net36[300], net36[301], net36[302], net36[303]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[67:66]), .r_gnd_r(r_gnd_r[67:66]));
cram_2x2x2_ice8p I_mem2x2x2t_32_ ( .wl_r(wl_r[65:64]),
     .wl_l(wl_l[65:64]), .reset_r(reset_r[65:64]),
     .reset_l(reset_l[65:64]), .pgate_r(pgate_r[65:64]),
     .pgate_l(pgate_l[65:64]), .q_b({net35[304], net35[305],
     net35[306], net35[307], net35[308], net35[309], net35[310],
     net35[311]}), .q({net36[304], net36[305], net36[306], net36[307],
     net36[308], net36[309], net36[310], net36[311]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[65:64]), .r_gnd_r(r_gnd_r[65:64]));
cram_2x2x2_ice8p I_mem2x2x2t_31_ ( .wl_r(wl_r[63:62]),
     .wl_l(wl_l[63:62]), .reset_r(reset_r[63:62]),
     .reset_l(reset_l[63:62]), .pgate_r(pgate_r[63:62]),
     .pgate_l(pgate_l[63:62]), .q_b({net35[312], net35[313],
     net35[314], net35[315], net35[316], net35[317], net35[318],
     net35[319]}), .q({net36[312], net36[313], net36[314], net36[315],
     net36[316], net36[317], net36[318], net36[319]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[63:62]), .r_gnd_r(r_gnd_r[63:62]));
cram_2x2x2_ice8p I_mem2x2x2t_30_ ( .wl_r(wl_r[61:60]),
     .wl_l(wl_l[61:60]), .reset_r(reset_r[61:60]),
     .reset_l(reset_l[61:60]), .pgate_r(pgate_r[61:60]),
     .pgate_l(pgate_l[61:60]), .q_b({net35[320], net35[321],
     net35[322], net35[323], net35[324], net35[325], net35[326],
     net35[327]}), .q({net36[320], net36[321], net36[322], net36[323],
     net36[324], net36[325], net36[326], net36[327]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[61:60]), .r_gnd_r(r_gnd_r[61:60]));
cram_2x2x2_ice8p I_mem2x2x2t_29_ ( .wl_r(wl_r[59:58]),
     .wl_l(wl_l[59:58]), .reset_r(reset_r[59:58]),
     .reset_l(reset_l[59:58]), .pgate_r(pgate_r[59:58]),
     .pgate_l(pgate_l[59:58]), .q_b({net35[328], net35[329],
     net35[330], net35[331], net35[332], net35[333], net35[334],
     net35[335]}), .q({net36[328], net36[329], net36[330], net36[331],
     net36[332], net36[333], net36[334], net36[335]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[59:58]), .r_gnd_r(r_gnd_r[59:58]));
cram_2x2x2_ice8p I_mem2x2x2t_28_ ( .wl_r(wl_r[57:56]),
     .wl_l(wl_l[57:56]), .reset_r(reset_r[57:56]),
     .reset_l(reset_l[57:56]), .pgate_r(pgate_r[57:56]),
     .pgate_l(pgate_l[57:56]), .q_b({net35[336], net35[337],
     net35[338], net35[339], net35[340], net35[341], net35[342],
     net35[343]}), .q({net36[336], net36[337], net36[338], net36[339],
     net36[340], net36[341], net36[342], net36[343]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[57:56]), .r_gnd_r(r_gnd_r[57:56]));
cram_2x2x2_ice8p I_mem2x2x2t_27_ ( .wl_r(wl_r[55:54]),
     .wl_l(wl_l[55:54]), .reset_r(reset_r[55:54]),
     .reset_l(reset_l[55:54]), .pgate_r(pgate_r[55:54]),
     .pgate_l(pgate_l[55:54]), .q_b({net35[344], net35[345],
     net35[346], net35[347], net35[348], net35[349], net35[350],
     net35[351]}), .q({net36[344], net36[345], net36[346], net36[347],
     net36[348], net36[349], net36[350], net36[351]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[55:54]), .r_gnd_r(r_gnd_r[55:54]));
cram_2x2x2_ice8p I_mem2x2x2t_26_ ( .wl_r(wl_r[53:52]),
     .wl_l(wl_l[53:52]), .reset_r(reset_r[53:52]),
     .reset_l(reset_l[53:52]), .pgate_r(pgate_r[53:52]),
     .pgate_l(pgate_l[53:52]), .q_b({net35[352], net35[353],
     net35[354], net35[355], net35[356], net35[357], net35[358],
     net35[359]}), .q({net36[352], net36[353], net36[354], net36[355],
     net36[356], net36[357], net36[358], net36[359]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[53:52]), .r_gnd_r(r_gnd_r[53:52]));
cram_2x2x2_ice8p I_mem2x2x2t_25_ ( .wl_r(wl_r[51:50]),
     .wl_l(wl_l[51:50]), .reset_r(reset_r[51:50]),
     .reset_l(reset_l[51:50]), .pgate_r(pgate_r[51:50]),
     .pgate_l(pgate_l[51:50]), .q_b({net35[360], net35[361],
     net35[362], net35[363], net35[364], net35[365], net35[366],
     net35[367]}), .q({net36[360], net36[361], net36[362], net36[363],
     net36[364], net36[365], net36[366], net36[367]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[51:50]), .r_gnd_r(r_gnd_r[51:50]));
cram_2x2x2_ice8p I_mem2x2x2t_24_ ( .wl_r(wl_r[49:48]),
     .wl_l(wl_l[49:48]), .reset_r(reset_r[49:48]),
     .reset_l(reset_l[49:48]), .pgate_r(pgate_r[49:48]),
     .pgate_l(pgate_l[49:48]), .q_b({net35[368], net35[369],
     net35[370], net35[371], net35[372], net35[373], net35[374],
     net35[375]}), .q({net36[368], net36[369], net36[370], net36[371],
     net36[372], net36[373], net36[374], net36[375]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[49:48]), .r_gnd_r(r_gnd_r[49:48]));
cram_2x2x2_ice8p I_mem2x2x2t_23_ ( .wl_r(wl_r[47:46]),
     .wl_l(wl_l[47:46]), .reset_r(reset_r[47:46]),
     .reset_l(reset_l[47:46]), .pgate_r(pgate_r[47:46]),
     .pgate_l(pgate_l[47:46]), .q_b({net35[376], net35[377],
     net35[378], net35[379], net35[380], net35[381], net35[382],
     net35[383]}), .q({net36[376], net36[377], net36[378], net36[379],
     net36[380], net36[381], net36[382], net36[383]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[47:46]), .r_gnd_r(r_gnd_r[47:46]));
cram_2x2x2_ice8p I_mem2x2x2t_22_ ( .wl_r(wl_r[45:44]),
     .wl_l(wl_l[45:44]), .reset_r(reset_r[45:44]),
     .reset_l(reset_l[45:44]), .pgate_r(pgate_r[45:44]),
     .pgate_l(pgate_l[45:44]), .q_b({net35[384], net35[385],
     net35[386], net35[387], net35[388], net35[389], net35[390],
     net35[391]}), .q({net36[384], net36[385], net36[386], net36[387],
     net36[388], net36[389], net36[390], net36[391]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[45:44]), .r_gnd_r(r_gnd_r[45:44]));
cram_2x2x2_ice8p I_mem2x2x2t_21_ ( .wl_r(wl_r[43:42]),
     .wl_l(wl_l[43:42]), .reset_r(reset_r[43:42]),
     .reset_l(reset_l[43:42]), .pgate_r(pgate_r[43:42]),
     .pgate_l(pgate_l[43:42]), .q_b({net35[392], net35[393],
     net35[394], net35[395], net35[396], net35[397], net35[398],
     net35[399]}), .q({net36[392], net36[393], net36[394], net36[395],
     net36[396], net36[397], net36[398], net36[399]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[43:42]), .r_gnd_r(r_gnd_r[43:42]));
cram_2x2x2_ice8p I_mem2x2x2t_20_ ( .wl_r(wl_r[41:40]),
     .wl_l(wl_l[41:40]), .reset_r(reset_r[41:40]),
     .reset_l(reset_l[41:40]), .pgate_r(pgate_r[41:40]),
     .pgate_l(pgate_l[41:40]), .q_b({net35[400], net35[401],
     net35[402], net35[403], net35[404], net35[405], net35[406],
     net35[407]}), .q({net36[400], net36[401], net36[402], net36[403],
     net36[404], net36[405], net36[406], net36[407]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[41:40]), .r_gnd_r(r_gnd_r[41:40]));
cram_2x2x2_ice8p I_mem2x2x2t_19_ ( .wl_r(wl_r[39:38]),
     .wl_l(wl_l[39:38]), .reset_r(reset_r[39:38]),
     .reset_l(reset_l[39:38]), .pgate_r(pgate_r[39:38]),
     .pgate_l(pgate_l[39:38]), .q_b({net35[408], net35[409],
     net35[410], net35[411], net35[412], net35[413], net35[414],
     net35[415]}), .q({net36[408], net36[409], net36[410], net36[411],
     net36[412], net36[413], net36[414], net36[415]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[39:38]), .r_gnd_r(r_gnd_r[39:38]));
cram_2x2x2_ice8p I_mem2x2x2t_18_ ( .wl_r(wl_r[37:36]),
     .wl_l(wl_l[37:36]), .reset_r(reset_r[37:36]),
     .reset_l(reset_l[37:36]), .pgate_r(pgate_r[37:36]),
     .pgate_l(pgate_l[37:36]), .q_b({net35[416], net35[417],
     net35[418], net35[419], net35[420], net35[421], net35[422],
     net35[423]}), .q({net36[416], net36[417], net36[418], net36[419],
     net36[420], net36[421], net36[422], net36[423]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[37:36]), .r_gnd_r(r_gnd_r[37:36]));
cram_2x2x2_ice8p I_mem2x2x2t_17_ ( .wl_r(wl_r[35:34]),
     .wl_l(wl_l[35:34]), .reset_r(reset_r[35:34]),
     .reset_l(reset_l[35:34]), .pgate_r(pgate_r[35:34]),
     .pgate_l(pgate_l[35:34]), .q_b({net35[424], net35[425],
     net35[426], net35[427], net35[428], net35[429], net35[430],
     net35[431]}), .q({net36[424], net36[425], net36[426], net36[427],
     net36[428], net36[429], net36[430], net36[431]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[35:34]), .r_gnd_r(r_gnd_r[35:34]));
cram_2x2x2_ice8p I_mem2x2x2t_16_ ( .wl_r(wl_r[33:32]),
     .wl_l(wl_l[33:32]), .reset_r(reset_r[33:32]),
     .reset_l(reset_l[33:32]), .pgate_r(pgate_r[33:32]),
     .pgate_l(pgate_l[33:32]), .q_b({net35[432], net35[433],
     net35[434], net35[435], net35[436], net35[437], net35[438],
     net35[439]}), .q({net36[432], net36[433], net36[434], net36[435],
     net36[436], net36[437], net36[438], net36[439]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[33:32]), .r_gnd_r(r_gnd_r[33:32]));
cram_2x2x2_ice8p I_mem2x2x2t_15_ ( .wl_r(wl_r[31:30]),
     .wl_l(wl_l[31:30]), .reset_r(reset_r[31:30]),
     .reset_l(reset_l[31:30]), .pgate_r(pgate_r[31:30]),
     .pgate_l(pgate_l[31:30]), .q_b({net35[440], net35[441],
     net35[442], net35[443], net35[444], net35[445], net35[446],
     net35[447]}), .q({net36[440], net36[441], net36[442], net36[443],
     net36[444], net36[445], net36[446], net36[447]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[31:30]), .r_gnd_r(r_gnd_r[31:30]));
cram_2x2x2_ice8p I_mem2x2x2t_14_ ( .wl_r(wl_r[29:28]),
     .wl_l(wl_l[29:28]), .reset_r(reset_r[29:28]),
     .reset_l(reset_l[29:28]), .pgate_r(pgate_r[29:28]),
     .pgate_l(pgate_l[29:28]), .q_b({net35[448], net35[449],
     net35[450], net35[451], net35[452], net35[453], net35[454],
     net35[455]}), .q({net36[448], net36[449], net36[450], net36[451],
     net36[452], net36[453], net36[454], net36[455]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[29:28]), .r_gnd_r(r_gnd_r[29:28]));
cram_2x2x2_ice8p I_mem2x2x2t_13_ ( .wl_r(wl_r[27:26]),
     .wl_l(wl_l[27:26]), .reset_r(reset_r[27:26]),
     .reset_l(reset_l[27:26]), .pgate_r(pgate_r[27:26]),
     .pgate_l(pgate_l[27:26]), .q_b({net35[456], net35[457],
     net35[458], net35[459], net35[460], net35[461], net35[462],
     net35[463]}), .q({net36[456], net36[457], net36[458], net36[459],
     net36[460], net36[461], net36[462], net36[463]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[27:26]), .r_gnd_r(r_gnd_r[27:26]));
cram_2x2x2_ice8p I_mem2x2x2t_12_ ( .wl_r(wl_r[25:24]),
     .wl_l(wl_l[25:24]), .reset_r(reset_r[25:24]),
     .reset_l(reset_l[25:24]), .pgate_r(pgate_r[25:24]),
     .pgate_l(pgate_l[25:24]), .q_b({net35[464], net35[465],
     net35[466], net35[467], net35[468], net35[469], net35[470],
     net35[471]}), .q({net36[464], net36[465], net36[466], net36[467],
     net36[468], net36[469], net36[470], net36[471]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[25:24]), .r_gnd_r(r_gnd_r[25:24]));
cram_2x2x2_ice8p I_mem2x2x2t_11_ ( .wl_r(wl_r[23:22]),
     .wl_l(wl_l[23:22]), .reset_r(reset_r[23:22]),
     .reset_l(reset_l[23:22]), .pgate_r(pgate_r[23:22]),
     .pgate_l(pgate_l[23:22]), .q_b({net35[472], net35[473],
     net35[474], net35[475], net35[476], net35[477], net35[478],
     net35[479]}), .q({net36[472], net36[473], net36[474], net36[475],
     net36[476], net36[477], net36[478], net36[479]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[23:22]), .r_gnd_r(r_gnd_r[23:22]));
cram_2x2x2_ice8p I_mem2x2x2t_10_ ( .wl_r(wl_r[21:20]),
     .wl_l(wl_l[21:20]), .reset_r(reset_r[21:20]),
     .reset_l(reset_l[21:20]), .pgate_r(pgate_r[21:20]),
     .pgate_l(pgate_l[21:20]), .q_b({net35[480], net35[481],
     net35[482], net35[483], net35[484], net35[485], net35[486],
     net35[487]}), .q({net36[480], net36[481], net36[482], net36[483],
     net36[484], net36[485], net36[486], net36[487]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[21:20]), .r_gnd_r(r_gnd_r[21:20]));
cram_2x2x2_ice8p I_mem2x2x2t_9_ ( .wl_r(wl_r[19:18]),
     .wl_l(wl_l[19:18]), .reset_r(reset_r[19:18]),
     .reset_l(reset_l[19:18]), .pgate_r(pgate_r[19:18]),
     .pgate_l(pgate_l[19:18]), .q_b({net35[488], net35[489],
     net35[490], net35[491], net35[492], net35[493], net35[494],
     net35[495]}), .q({net36[488], net36[489], net36[490], net36[491],
     net36[492], net36[493], net36[494], net36[495]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[19:18]), .r_gnd_r(r_gnd_r[19:18]));
cram_2x2x2_ice8p I_mem2x2x2t_8_ ( .wl_r(wl_r[17:16]),
     .wl_l(wl_l[17:16]), .reset_r(reset_r[17:16]),
     .reset_l(reset_l[17:16]), .pgate_r(pgate_r[17:16]),
     .pgate_l(pgate_l[17:16]), .q_b({net35[496], net35[497],
     net35[498], net35[499], net35[500], net35[501], net35[502],
     net35[503]}), .q({net36[496], net36[497], net36[498], net36[499],
     net36[500], net36[501], net36[502], net36[503]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[17:16]), .r_gnd_r(r_gnd_r[17:16]));
cram_2x2x2_ice8p I_mem2x2x2t_7_ ( .wl_r(wl_r[15:14]),
     .wl_l(wl_l[15:14]), .reset_r(reset_r[15:14]),
     .reset_l(reset_l[15:14]), .pgate_r(pgate_r[15:14]),
     .pgate_l(pgate_l[15:14]), .q_b({net35[504], net35[505],
     net35[506], net35[507], net35[508], net35[509], net35[510],
     net35[511]}), .q({net36[504], net36[505], net36[506], net36[507],
     net36[508], net36[509], net36[510], net36[511]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[15:14]), .r_gnd_r(r_gnd_r[15:14]));
cram_2x2x2_ice8p I_mem2x2x2t_6_ ( .wl_r(wl_r[13:12]),
     .wl_l(wl_l[13:12]), .reset_r(reset_r[13:12]),
     .reset_l(reset_l[13:12]), .pgate_r(pgate_r[13:12]),
     .pgate_l(pgate_l[13:12]), .q_b({net35[512], net35[513],
     net35[514], net35[515], net35[516], net35[517], net35[518],
     net35[519]}), .q({net36[512], net36[513], net36[514], net36[515],
     net36[516], net36[517], net36[518], net36[519]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[13:12]), .r_gnd_r(r_gnd_r[13:12]));
cram_2x2x2_ice8p I_mem2x2x2t_5_ ( .wl_r(wl_r[11:10]),
     .wl_l(wl_l[11:10]), .reset_r(reset_r[11:10]),
     .reset_l(reset_l[11:10]), .pgate_r(pgate_r[11:10]),
     .pgate_l(pgate_l[11:10]), .q_b({net35[520], net35[521],
     net35[522], net35[523], net35[524], net35[525], net35[526],
     net35[527]}), .q({net36[520], net36[521], net36[522], net36[523],
     net36[524], net36[525], net36[526], net36[527]}), .bl(bl[3:0]),
     .r_gnd_l(r_gnd_l[11:10]), .r_gnd_r(r_gnd_r[11:10]));
cram_2x2x2_ice8p I_mem2x2x2t_4_ ( .wl_r(wl_r[9:8]), .wl_l(wl_l[9:8]),
     .reset_r(reset_r[9:8]), .reset_l(reset_l[9:8]),
     .pgate_r(pgate_r[9:8]), .pgate_l(pgate_l[9:8]), .q_b({net35[528],
     net35[529], net35[530], net35[531], net35[532], net35[533],
     net35[534], net35[535]}), .q({net36[528], net36[529], net36[530],
     net36[531], net36[532], net36[533], net36[534], net36[535]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[9:8]), .r_gnd_r(r_gnd_r[9:8]));
cram_2x2x2_ice8p I_mem2x2x2t_3_ ( .wl_r(wl_r[7:6]), .wl_l(wl_l[7:6]),
     .reset_r(reset_r[7:6]), .reset_l(reset_l[7:6]),
     .pgate_r(pgate_r[7:6]), .pgate_l(pgate_l[7:6]), .q_b({net35[536],
     net35[537], net35[538], net35[539], net35[540], net35[541],
     net35[542], net35[543]}), .q({net36[536], net36[537], net36[538],
     net36[539], net36[540], net36[541], net36[542], net36[543]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[7:6]), .r_gnd_r(r_gnd_r[7:6]));
cram_2x2x2_ice8p I_mem2x2x2t_2_ ( .wl_r(wl_r[5:4]), .wl_l(wl_l[5:4]),
     .reset_r(reset_r[5:4]), .reset_l(reset_l[5:4]),
     .pgate_r(pgate_r[5:4]), .pgate_l(pgate_l[5:4]), .q_b({net35[544],
     net35[545], net35[546], net35[547], net35[548], net35[549],
     net35[550], net35[551]}), .q({net36[544], net36[545], net36[546],
     net36[547], net36[548], net36[549], net36[550], net36[551]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[5:4]), .r_gnd_r(r_gnd_r[5:4]));
cram_2x2x2_ice8p I_mem2x2x2t_1_ ( .wl_r(wl_r[3:2]), .wl_l(wl_l[3:2]),
     .reset_r(reset_r[3:2]), .reset_l(reset_l[3:2]),
     .pgate_r(pgate_r[3:2]), .pgate_l(pgate_l[3:2]), .q_b({net35[552],
     net35[553], net35[554], net35[555], net35[556], net35[557],
     net35[558], net35[559]}), .q({net36[552], net36[553], net36[554],
     net36[555], net36[556], net36[557], net36[558], net36[559]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[3:2]), .r_gnd_r(r_gnd_r[3:2]));
cram_2x2x2_ice8p I_mem2x2x2t_0_ ( .wl_r(wl_r[1:0]), .wl_l(wl_l[1:0]),
     .reset_r(reset_r[1:0]), .reset_l(reset_l[1:0]),
     .pgate_r(pgate_r[1:0]), .pgate_l(pgate_l[1:0]), .q_b({net35[560],
     net35[561], net35[562], net35[563], net35[564], net35[565],
     net35[566], net35[567]}), .q({net36[560], net36[561], net36[562],
     net36[563], net36[564], net36[565], net36[566], net36[567]}),
     .bl(bl[3:0]), .r_gnd_l(r_gnd_l[1:0]), .r_gnd_r(r_gnd_r[1:0]));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_osc, View - schematic
// LAST TIME SAVED: Sep  2 15:47:56 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpxa_osc ( vpxa_clk_25, bgr, freq_25, pumpen_25 );
output  vpxa_clk_25;

inout  bgr;

input  pumpen_25;

input [1:0]  freq_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  freq_buf_b_25;



rppolywo_m  R6 ( .MINUS(gnd_), .PLUS(net043), .BULK(GND_));
rppolywo_m  R7 ( .MINUS(net043), .PLUS(net044), .BULK(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
pch_25  M9 ( .D(net061), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
pch_25  M10 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
pch_25  M8_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
pch_25  M8_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net061));
nch_25  M12 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
nch_25  M11 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net044));
inv_25 I227 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I226 ( .IN(freq_25[0]), .OUT(freq_buf_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_vpp_vco Ivpx_vpp_vco ( .clk_25_1(net040), .pbias_25(pbias_25),
     .slow_25(net86), .freq_25({freq_25[1], freq_buf_b_25[0]}),
     .en_25(pumpen_25), .clk_25_0(vpxa_clk_25));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_ctrl, View - schematic
// LAST TIME SAVED: Sep  1 14:08:10 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpxa_ctrl ( pumpen, pumpen_25, vpxa_2_vdd, fsm_pumpen,
     fsm_tm_xforce, fsm_tm_xvpxaint );
output  pumpen, pumpen_25, vpxa_2_vdd;

input  fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I103 ( .A(vpxa_2_vdd), .B(net065), .Y(pumpen));
nand2_hvt I73 ( .A(fsm_tm_xvpxaint), .B(fsm_tm_xforce), .Y(net042));
inv_hvt I78 ( .A(pumpen), .Y(net075));
inv_hvt I77 ( .A(net042), .Y(net065));
inv_hvt I131 ( .A(fsm_pumpen), .Y(vpxa_2_vdd));
inv_25 I38 ( .IN(net045), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I173 ( .in(pumpen), .sup(vddp_), .out_vddio_b(net045),
     .out_vddio(net046), .in_b(net075));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff_25, View - schematic
// LAST TIME SAVED: Aug 30 17:06:17 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_dff_25 ( Q_25, Q_B_25, CLK_25, D_25, R_25 );
output  Q_25, Q_B_25;

input  CLK_25, D_25, R_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I96 ( .IN(Q_25), .OUT(Q_B_25), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I72 ( .IN(CLK_25), .OUT(net044), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I95 ( .IN(net044), .OUT(net038), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
ml_dlatch_25 Ilatch2 ( .D_25(net053), .EN_25(net038), .R_25(R_25),
     .Q_25(Q_25));
ml_dlatch_25 Ilatch1 ( .Q_25(net053), .EN_25(net044), .D_25(D_25),
     .R_25(R_25));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_n, View - schematic
// LAST TIME SAVED: Aug 30 15:13:05 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp_n ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M8 ( .D(out_ref), .B(GND_), .G(in_ref), .S(net049));
nch_25  M3 ( .D(out_div), .B(GND_), .G(in_div), .S(net049));
nch_25  M6_1_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
pch_25  M1 ( .D(out_ref), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M0 ( .D(out_div), .B(vddp_), .G(out_ref), .S(vddp_));
pch_25  M5 ( .D(out_div), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M7 ( .D(out_ref), .B(vddp_), .G(out_ref), .S(vddp_));

endmodule
// Library - NVCM_40nm, Cell - ml_core_sa_comp_top_n, View - schematic
// LAST TIME SAVED: Aug 30 15:12:30 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_core_sa_comp_top_n ( pump_chrg_25, in_div, in_ref, sa_bias,
     saen_25 );
output  pump_chrg_25;

input  in_div, in_ref, sa_bias, saen_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_25 I103 ( .G(gnd_), .Pb(vddp_), .A(saen_25), .Y(chrg_b_25),
     .P(vddp_), .B(net27), .Gb(gnd_));
nch_25  M6_1_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
inv_25 I102 ( .IN(chrg_b_25), .OUT(pump_chrg_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I104 ( .IN(out_div2), .OUT(net27), .P(vddp_), .Pb(vddp_),
     .G(net087), .Gb(gnd_));
ml_core_sa_comp_n Icore_sa_comp_n0 ( .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp_n Iml_core_sa_comp_n1 ( .out_div(out_div2),
     .out_ref(out_ref2), .in_div(in_div2), .in_ref(in_ref2),
     .sa_bias(sa_bias), .saen_25(saen_25));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_reg, View - schematic
// LAST TIME SAVED: Nov  6 18:01:31 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpxa_reg ( freq_25, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, vpxa_int, bgr, fsm_vrdwl, pumpen, vpxa_clk_25 );
output  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25;

inout  vpxa_int;

input  bgr, pumpen, vpxa_clk_25;

output [1:0]  freq_25;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vrdwl_b_vpxa;

wire  [2:0]  vrdwl_vpxa;

wire  [1:0]  freq_in_25;



ml_ls_vdd2vdd25_vpxa I191 ( .in(saen_25), .sup(vpxa_int),
     .out_vddio_b(saen_b_vpxa), .out_vddio(net0210), .in_b(saen_b_25));
ml_ls_vdd2vdd25_vpxa I87 ( .in(net171), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[2]), .out_vddio(vrdwl_b_vpxa[2]),
     .in_b(net175));
ml_ls_vdd2vdd25_vpxa I98 ( .in(net176), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[1]), .out_vddio(vrdwl_b_vpxa[1]),
     .in_b(net180));
ml_ls_vdd2vdd25_vpxa I99 ( .in(net181), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[0]), .out_vddio(vrdwl_b_vpxa[0]),
     .in_b(net185));
rppolywo_m  R29 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R28 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R27 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(in_div_0), .PLUS(net202), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net232), .PLUS(net223), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(net270), .PLUS(net226), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net226), .PLUS(net229), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(sa_bias), .PLUS(net232), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net202), .PLUS(net237), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(net237), .PLUS(net270), .BULK(GND_));
rppolywo_m  R30 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(gnd_), .PLUS(in_div_2), .BULK(GND_));
rppolywo_m  R31 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
nch_25  M2 ( .D(sa_bias), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M32 ( .D(net229), .B(GND_), .G(vrdwl_b_vpxa[2]), .S(net226));
nch_25  M0_3_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_2_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_1_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_0_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M7 ( .D(net270), .B(GND_), .G(vrdwl_b_vpxa[0]), .S(net237));
nch_25  M4 ( .D(net226), .B(GND_), .G(vrdwl_b_vpxa[1]), .S(net270));
nand2_25 I194 ( .G(GND_), .Pb(vddp_), .A(net0179), .Y(freq_in_25[1]),
     .P(vddp_), .B(net0234), .Gb(GND_));
nand2_25 I145 ( .G(GND_), .Pb(vddp_), .A(net0171), .Y(freq_in_25[0]),
     .P(vddp_), .B(net0179), .Gb(GND_));
nand3_25 I193 ( .B(pump_chrg_1_b_25), .A(pump_chrg_2_25), .Y(net0171),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I192 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0179),
     .C(pump_chrg_0_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I159 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0234),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
pch_25  M3 ( .D(net229), .B(vpxa_int), .G(saen_b_vpxa), .S(vpxa_int));
pch_25  M11_1_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M11_0_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M37 ( .D(net226), .B(vpxa_int), .G(vrdwl_vpxa[2]), .S(net229));
pch_25  M1 ( .D(net223), .B(vddp_), .G(saen_b_25), .S(vddp_));
pch_25  M5 ( .D(net270), .B(vpxa_int), .G(vrdwl_vpxa[1]), .S(net226));
pch_25  M6 ( .D(net237), .B(vpxa_int), .G(vrdwl_vpxa[0]), .S(net270));
pch_25  M8_1_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
pch_25  M8_0_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
inv_25 I196 ( .IN(net169), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I197 ( .IN(net168), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I195 ( .IN(pump_chrg_0_25), .OUT(pump_chrg_0_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
inv_25 I154 ( .IN(pump_chrg_1_25), .OUT(pump_chrg_1_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_dff_25 I125 ( .Q_B_25(net0187), .R_25(saen_b_25),
     .D_25(freq_in_25[1]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[1]));
ml_dff_25 I126 ( .Q_B_25(net0192), .R_25(saen_b_25),
     .D_25(freq_in_25[0]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[0]));
inv_hvt I85 ( .A(net171), .Y(net175));
inv_hvt I183 ( .A(fsm_vrdwl[2]), .Y(net171));
inv_hvt I83 ( .A(pumpen), .Y(net143));
inv_hvt I82 ( .A(net143), .Y(net145));
inv_hvt I184 ( .A(fsm_vrdwl[1]), .Y(net176));
inv_hvt I187 ( .A(fsm_vrdwl[0]), .Y(net181));
inv_hvt I186 ( .A(net181), .Y(net185));
inv_hvt I185 ( .A(net176), .Y(net180));
ml_ls_vdd2vdd25 I335 ( .in(net145), .sup(vddp_), .out_vddio_b(net168),
     .out_vddio(net169), .in_b(net143));
ml_core_sa_comp_top_n Icore_sa_comp_top_n2 (
     .pump_chrg_25(pump_chrg_2_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_2));
ml_core_sa_comp_top_n core_sa_comp_top_n0 (
     .pump_chrg_25(pump_chrg_0_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_0));
ml_core_sa_comp_top_n Icore_sa_comp_top_n1 (
     .pump_chrg_25(pump_chrg_1_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_1));

endmodule
// Library - NVCM_40nm, Cell - ml_hv2vdd_sw, View - schematic
// LAST TIME SAVED: Aug 30 15:14:40 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hv2vdd_sw ( out_hv, hv2vdd, vddp_tieh );
inout  out_hv;

input  hv2vdd, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M2 ( .D(vdd_), .B(GND_), .G(hv2vdd_25), .S(net27));
nch_na25  M0 ( .D(net27), .B(GND_), .G(vddp_tieh), .S(out_hv));
inv_25 I62 ( .IN(net40), .OUT(hv2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_hvt I71 ( .A(net46), .Y(net44));
inv_hvt I72 ( .A(hv2vdd), .Y(net46));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net40),
     .out_vddio(net37), .in_b(net46));

endmodule
// Library - NVCM_40nm, Cell - ml_vpxa_top, View - schematic
// LAST TIME SAVED: Nov  8 10:18:53 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_vpxa_top ( vpxa_int, bgr, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint, fsm_vrdwl );
inout  vpxa_int;

input  bgr, fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;

input [2:0]  fsm_vrdwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  freq_25;



nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpxa_int));
inv_25 I73 ( .IN(vpxa_clk_25), .OUT(vpxa_clk_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_pump_vpxa_x2 Ipump_vpxa_x3 ( .vpxa_clk_b_25(vpxa_clk_b_25),
     .vpxa_clk_25(vpxa_clk_25), .pumpen_25(pumpen_25),
     .pump_chrg_2_25(pump_chrg_2_25), .pump_chrg_1_25(pump_chrg_1_25),
     .pump_chrg_0_25(pump_chrg_0_25), .vpxa_int(vpxa_int));
ml_vpxa_osc Ivpxa_osc ( .freq_25(freq_25[1:0]), .bgr(bgr),
     .pumpen_25(pumpen_25), .vpxa_clk_25(vpxa_clk_25));
ml_vpxa_ctrl Ivpxa_ctrl ( .fsm_pumpen(fsm_pumpen), .pumpen(pumpen),
     .pumpen_25(pumpen_25), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .vpxa_2_vdd(vpxa_2_vdd));
vddp_tiehigh I118 ( .vddp_tieh(vddp_tieh));
ml_vpxa_reg Ivpxa_reg ( .pump_chrg_0_25(pump_chrg_0_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_2_25(pump_chrg_2_25),
     .freq_25(freq_25[1:0]), .vpxa_clk_25(vpxa_clk_25),
     .pumpen(pumpen), .fsm_vrdwl(fsm_vrdwl[2:0]), .bgr(bgr),
     .vpxa_int(vpxa_int));
ml_hv2vdd_sw Ivpxa_2vdd_sw ( .vddp_tieh(vddp_tieh),
     .hv2vdd(vpxa_2_vdd), .out_hv(vpxa_int));

endmodule
// Library - NVCM_40nm, Cell - ml_rdhv_gen, View - schematic
// LAST TIME SAVED: Jul 27 12:15:43 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_rdhv_gen ( s_rdin_hv, srdsup_hv, s_rdin, vddp_tieh );
output  s_rdin_hv;

inout  srdsup_hv;

input  s_rdin, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_s_b_hv_sw Iml_s_b_25_sw ( .sbout_high_25(s_rdin_high_25),
     .sbout_gnd_25(net31), .sbout_hv(s_rdin_hv), .ssup_hv(srdsup_hv),
     .vddp_tieh(vddp_tieh));
ml_ls_vdd2vdd25 Iml_ls_vdd2vdd25 ( .in(s_rdin), .sup(vddp_),
     .out_vddio_b(net31), .out_vddio(s_rdin_high_25), .in_b(net35));
inv_hvt I439 ( .A(s_rdin), .Y(net35));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_top_ctrl, View - schematic
// LAST TIME SAVED: Nov  5 16:32:34 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hvmux_top_ctrl ( bgrext_en, bgrint_en, en_vblinhi,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp, fsm_lshven,
     fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en );
output  bgrext_en, bgrint_en, en_vblinhi, ngate_vddp, ngate_vpxa,
     sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint,
     vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint, vpxaint_ext,
     vtmode, ysup25_2vdd, ysup25_2vddp;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor4_hvt I186 ( .D(fsm_tm_rprd), .C(fsm_rd), .A(fsm_tm_rd_mode),
     .B(fsm_pgmvfy), .Y(net0349));
nand4_hvt I322 ( .D(fsm_lshven), .A(fsm_pgm), .C(fsm_lshven),
     .Y(pgmpulse_b), .B(net0236));
nand4_hvt I35 ( .D(fsm_lshven), .C(net0318), .A(fsm_pgm), .Y(net0196),
     .B(net0327));
anor21_hvt I245 ( .A(net0189), .B(net0193), .Y(vppint_ext),
     .C(net0190));
anor21_hvt I109 ( .A(net0201), .B(net0199), .Y(vpxa_ext), .C(net0190));
nand3_hvt I288 ( .Y(net0193), .B(pmprd), .C(pmprd),
     .A(fsm_tm_xvppint));
nand3_hvt I291 ( .Y(net0201), .B(vddp_rd_b), .C(gnd_tiel),
     .A(fsm_tm_xforce));
nand3_hvt I292 ( .Y(net0213), .B(net0321), .C(net0196), .A(net0321));
nand3_hvt I290 ( .Y(net0199), .B(pmprd), .C(pmprd), .A(gnd_tiel));
nand3_hvt I289 ( .Y(net0189), .B(vpint_en), .C(fsm_tm_xvppint),
     .A(fsm_tm_xforce));
nor3_hvt I286 ( .B(net0240), .Y(rd_vddp), .A(net0240),
     .C(fsm_nvcmen_b));
nor3_hvt I285 ( .B(tm_testdec), .Y(en_vblinhi), .A(fsm_nvcmen_b),
     .C(tm_allbl_l));
mux2_hvt I260 ( .in1(fsm_wgnden), .in0(fsm_wpen), .out(net0217),
     .sel(pgmpulse_b));
nor2_hvt I272 ( .A(net75), .B(net93), .Y(ysup25_2vdd));
nor2_hvt I279 ( .A(net0251), .B(net0266), .Y(sbhvsup_vppint));
nor2_hvt I283 ( .A(vddp_rd_b), .B(net0258), .Y(vpxa_vppd));
nor2_hvt I271 ( .A(net87), .B(net73), .Y(ysup25_2vddp));
nor2_hvt I273 ( .A(net0349), .B(net0240), .Y(vddp_rd));
nor2_hvt I281 ( .A(net0324), .B(fsm_nvcmen_b), .Y(net0251));
nor2_hvt I276 ( .A(net0272), .B(rd_vddp), .Y(ngate_vpxa));
nor2_hvt I280 ( .A(net0268), .B(net0213), .Y(sb25sup_vpxa));
nor2_hvt I275 ( .A(net0331), .B(net0270), .Y(ngate_vddp));
nor2_hvt I274 ( .A(fsm_tm_rprd), .B(gnd_tiel), .Y(net0240));
nor2_hvt I278 ( .A(net0264), .B(net0311), .Y(sbhvsup_vddp));
nor2_hvt I282 ( .A(net0256), .B(vddp_rd), .Y(vpxa_vpxaint));
nor2_hvt I277 ( .A(net0325), .B(net0260), .Y(sb25sup_vddp));
inv_hvt I294 ( .A(net77), .Y(vtmode));
inv_hvt I323 ( .A(fsm_pgmvfy), .Y(net0236));
inv_hvt I319 ( .A(ngate_vpxa), .Y(net0339));
inv_hvt I304 ( .A(net0251), .Y(net0311));
inv_hvt I315 ( .A(vddp_rd), .Y(vddp_rd_b));
inv_hvt I318 ( .A(ysup25_2vdd), .Y(ysup25_2vdd_b));
inv_hvt I314 ( .A(vpxa_vppd), .Y(net0297));
inv_hvt I309 ( .A(net0277), .Y(bgrext_en));
inv_hvt I317 ( .A(fsm_pgmvfy), .Y(net0327));
inv_hvt I316 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I297 ( .A(ysup25_2vddp), .Y(ysup25_2vddp_b));
inv_hvt I298 ( .A(rd_vddp), .Y(net0331));
inv_hvt I310 ( .A(fsm_pumpen), .Y(net0190));
inv_hvt I307 ( .A(sbhvsup_vddp), .Y(net0309));
inv_hvt I305 ( .A(sb25sup_vpxa), .Y(net0323));
inv_hvt I308 ( .A(sbhvsup_vppint), .Y(net0313));
inv_hvt I296 ( .A(net93), .Y(net87));
inv_hvt I295 ( .A(net80), .Y(net93));
inv_hvt I321 ( .A(fsm_tm_rprd), .Y(net0318));
inv_hvt I303 ( .A(pgmpulse_b), .Y(net0324));
inv_hvt I306 ( .A(pgmpulse_b), .Y(pgmpulse));
inv_hvt I300 ( .A(sb25sup_vddp), .Y(net0329));
inv_hvt I302 ( .A(rd_vddp), .Y(net0321));
inv_hvt I301 ( .A(net0213), .Y(net0325));
inv_hvt I311 ( .A(net0286), .Y(vpxaint_ext));
inv_hvt I312 ( .A(fsm_tm_xforce), .Y(pmprd));
inv_hvt I299 ( .A(ngate_vddp), .Y(net0335));
inv_hvt I313 ( .A(vpxa_vpxaint), .Y(net0319));
inv_hvt I233 ( .A(fsm_nvcmen_b), .Y(fsm_nvcmen_buf));
nand2_hvt I268 ( .A(fsm_nvcmen_buf), .Y(net0277), .B(fsm_tm_xvbg));
nand2_hvt I266 ( .A(fsm_nvcmen), .Y(net80), .B(net0217));
nand2_hvt I269 ( .A(bgrext_en), .Y(bgrint_en), .B(fsm_tm_xforce));
nand2_hvt I267 ( .A(fsm_pumpen), .Y(net0286), .B(fsm_tm_xvpxaint));
nand2_hvt I104 ( .A(fsm_nvcmen), .Y(net77), .B(tm_wleqbl));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
ml_pump_a_clkdly I219 ( .in(ysup25_2vddp_b), .out(net75));
ml_pump_a_clkdly I227 ( .in(net0297), .out(net0256));
ml_pump_a_clkdly I226 ( .in(net0319), .out(net0258));
ml_pump_a_clkdly I209 ( .in(net0323), .out(net0260));
ml_pump_a_clkdly I184 ( .in(ysup25_2vdd_b), .out(net73));
ml_pump_a_clkdly I217 ( .in(net0313), .out(net0264));
ml_pump_a_clkdly I216 ( .in(net0309), .out(net0266));
ml_pump_a_clkdly I208 ( .in(net0329), .out(net0268));
ml_pump_a_clkdly I198 ( .in(net0339), .out(net0270));
ml_pump_a_clkdly I197 ( .in(net0335), .out(net0272));

endmodule
// Library - xpmem, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Aug 20 09:48:05 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_ls25, View - schematic
// LAST TIME SAVED: Sep  7 10:34:50 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hvmux_ls25 ( bgrext_en_25, bgrint_en_25, ngate_vddp_25,
     ngate_vpxa_25, sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25, bgrext_en, bgrint_en,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp );
output  bgrext_en_25, bgrint_en_25, ngate_vddp_25, ngate_vpxa_25,
     sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25;

input  bgrext_en, bgrint_en, ngate_vddp, ngate_vpxa, sb25sup_vddp,
     sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint, vppint_ext, vpxa_ext,
     vpxa_vppd, vpxa_vpxaint, vpxaint_ext, vtmode, ysup25_2vdd,
     ysup25_2vddp;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_25 I471 ( .IN(net0138), .OUT(bgrint_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I472 ( .IN(net0148), .OUT(bgrext_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I473 ( .IN(net0128), .OUT(vppint_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I474 ( .IN(net0123), .OUT(vpxa_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I475 ( .IN(net0158), .OUT(vpxaint_ext_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I476 ( .IN(net0133), .OUT(vpxa_vppd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I477 ( .IN(net0163), .OUT(vpxa_vpxaint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I406 ( .IN(net077), .OUT(ysup25_2vddp_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I463 ( .IN(net0168), .OUT(ysup25_2vdd_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I464 ( .IN(net0193), .OUT(vtmode_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I465 ( .IN(net0173), .OUT(ngate_vddp_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I466 ( .IN(net0183), .OUT(ngate_vpxa_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I467 ( .IN(net0188), .OUT(sb25sup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I468 ( .IN(net0153), .OUT(sb25sup_vpxa_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I469 ( .IN(net0203), .OUT(sbhvsup_vppint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I470 ( .IN(net0198), .OUT(sbhvsup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_hvt I457 ( .A(vpxa_vppd), .Y(net054));
inv_hvt I435 ( .A(vpxa_vpxaint), .Y(net0112));
inv_hvt I462 ( .A(bgrint_en), .Y(net058));
inv_hvt I461 ( .A(bgrext_en), .Y(net068));
inv_hvt I460 ( .A(vppint_ext), .Y(net066));
inv_hvt I455 ( .A(ysup25_2vddp), .Y(net0328));
inv_hvt I454 ( .A(ysup25_2vdd), .Y(net0312));
inv_hvt I447 ( .A(ngate_vpxa), .Y(net0318));
inv_hvt I439 ( .A(sbhvsup_vppint), .Y(net0326));
inv_hvt I446 ( .A(sb25sup_vddp), .Y(net0320));
inv_hvt I216 ( .A(ysup25_2vdd), .Y(net092));
inv_hvt I458 ( .A(vpxaint_ext), .Y(net060));
inv_hvt I442 ( .A(sbhvsup_vddp), .Y(net0324));
inv_hvt I443 ( .A(sb25sup_vpxa), .Y(net0322));
inv_hvt I450 ( .A(ngate_vddp), .Y(net0316));
inv_hvt I217 ( .A(net092), .Y(ysup25_2vdd_buf));
inv_hvt I451 ( .A(vtmode), .Y(net0314));
inv_hvt I459 ( .A(vpxa_ext), .Y(net082));
ml_ls_vdd2vdd25 I336 ( .in(vpxa_ext), .sup(vddp_),
     .out_vddio_b(net0123), .out_vddio(net0207), .in_b(net082));
ml_ls_vdd2vdd25 I337 ( .in(vppint_ext), .sup(vddp_),
     .out_vddio_b(net0128), .out_vddio(net0208), .in_b(net066));
ml_ls_vdd2vdd25 I338 ( .in(vpxa_vppd), .sup(vddp_),
     .out_vddio_b(net0133), .out_vddio(net0211), .in_b(net054));
ml_ls_vdd2vdd25 I339 ( .in(bgrint_en), .sup(vddp_),
     .out_vddio_b(net0138), .out_vddio(net0209), .in_b(net058));
ml_ls_vdd2vdd25 I332 ( .in(bgrext_en), .sup(vddp_),
     .out_vddio_b(net0148), .out_vddio(net0149), .in_b(net068));
ml_ls_vdd2vdd25 I238 ( .in(sb25sup_vpxa), .sup(vddp_),
     .out_vddio_b(net0153), .out_vddio(net0154), .in_b(net0322));
ml_ls_vdd2vdd25 I334 ( .in(vpxaint_ext), .sup(vddp_),
     .out_vddio_b(net0158), .out_vddio(net0214), .in_b(net060));
ml_ls_vdd2vdd25 I335 ( .in(vpxa_vpxaint), .sup(vddp_),
     .out_vddio_b(net0163), .out_vddio(net0206), .in_b(net0112));
ml_ls_vdd2vdd25 I212 ( .in(ysup25_2vdd), .sup(vddp_),
     .out_vddio_b(net0168), .out_vddio(net0169), .in_b(net0312));
ml_ls_vdd2vdd25 I226 ( .in(ngate_vddp), .sup(vddp_),
     .out_vddio_b(net0173), .out_vddio(net0174), .in_b(net0316));
ml_ls_vdd2vdd25 I203 ( .in(net0328), .sup(vddp_), .out_vddio_b(net077),
     .out_vddio(net078), .in_b(ysup25_2vddp));
ml_ls_vdd2vdd25 I221 ( .in(ngate_vpxa), .sup(vddp_),
     .out_vddio_b(net0183), .out_vddio(net0184), .in_b(net0318));
ml_ls_vdd2vdd25 I233 ( .in(sb25sup_vddp), .sup(vddp_),
     .out_vddio_b(net0188), .out_vddio(net0219), .in_b(net0320));
ml_ls_vdd2vdd25 I207 ( .in(vtmode), .sup(vddp_), .out_vddio_b(net0193),
     .out_vddio(net0194), .in_b(net0314));
ml_ls_vdd2vdd25 I260 ( .in(sbhvsup_vddp), .sup(vddp_),
     .out_vddio_b(net0198), .out_vddio(net0220), .in_b(net0324));
ml_ls_vdd2vdd25 I261 ( .in(sbhvsup_vppint), .sup(vddp_),
     .out_vddio_b(net0203), .out_vddio(net0204), .in_b(net0326));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_bgrxcvr, View - schematic
// LAST TIME SAVED: Sep  3 09:50:30 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hvmux_bgrxcvr ( bgr, bgr_int, bgrint_en_25, vpp,
     bgrext_en_25, vddp_tieh );
inout  bgr, bgr_int, bgrint_en_25, vpp;

input  bgrext_en_25, vddp_tieh;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M2 ( .D(vpp), .B(GND_), .G(vddp_tieh), .S(net53));
nch_25  M1 ( .D(net53), .B(GND_), .G(bgrext_en_25), .S(bgr));
nch_na25  M0 ( .D(bgr), .B(GND_), .G(bgrint_en_25), .S(bgr_int));

endmodule
// Library - NVCM_40nm, Cell - ml_ysup_25_switch, View - schematic
// LAST TIME SAVED: Sep  3 09:40:13 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_ysup_25_switch ( vdd, vddp, ysup_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25 );
inout  vdd, vddp, ysup_25;

input  ysup25_2vdd_25, ysup25_2vdd_buf, ysup25_2vddp_b_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd), .B(GND_), .G(ysup25_2vdd_25), .S(ysup_25));
pch_25  M5 ( .D(net73), .B(vddp), .G(ysup25_2vddp_b_25), .S(vddp));
pch_25  M0 ( .D(ysup_25), .B(ysup_25), .G(ysup25_2vdd_buf), .S(net73));

endmodule
// Library - NVCM_40nm, Cell - ml_ymux_ctrl_vblinhi, View - schematic
// LAST TIME SAVED: Nov  8 18:40:26 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_ymux_ctrl_vblinhi ( vblinhi, vpxa, en_vblinhi, vtmode,
     vtmode_25 );
inout  vblinhi, vpxa;

input  en_vblinhi, vtmode, vtmode_25;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M0_9_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_8_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_7_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_6_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_5_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_4_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_3_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_2_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_1_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_0_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
pch_hvt  M7_9_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_8_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_7_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_6_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_5_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_4_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_3_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_2_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_1_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_0_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
nch_25  M9 ( .D(net035), .B(GND_), .G(net035), .S(vblinhi));
nch_25  M8 ( .D(vpxa), .B(GND_), .G(vtmode_25), .S(net035));
nor2_hvt I191 ( .A(en_vblinhi), .B(vtmode_buf), .Y(ngate_inhi_lv));
inv_hvt I192 ( .A(net063), .Y(vtmode_buf));
inv_hvt I190 ( .A(vtmode), .Y(net063));
nand2_hvt I104 ( .A(net063), .Y(pgate_inhi_lv), .B(en_vblinhi));

endmodule
// Library - NVCM_40nm, Cell - ml_hvmux_top, View - schematic
// LAST TIME SAVED: Nov 24 19:40:38 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_hvmux_top ( s_rdin_hv, bgr, bgr_int, ngate_25, sb25sup_25,
     sbhvsup_hv, srdsup_hv, vblinhi, vpp, vpp_int, vpxa, vpxa_int,
     ysup_25, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen,
     fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, s_rd,
     tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );

inout  bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv,
     vblinhi, vpp, vpp_int, vpxa, vpxa_int, ysup_25;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l,
     tm_testdec, tm_wleqbl, vpint_en;

output [3:0]  s_rdin_hv;

input [3:0]  s_rd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_rdin;

wire  [3:0]  net294;



nch_hvt  M1 ( .D(net299), .B(GND_), .G(net299), .S(gnd_));
inv_hvt I210_3_ ( .A(s_rd[3]), .Y(net294[0]));
inv_hvt I210_2_ ( .A(s_rd[2]), .Y(net294[1]));
inv_hvt I210_1_ ( .A(s_rd[1]), .Y(net294[2]));
inv_hvt I210_0_ ( .A(s_rd[0]), .Y(net294[3]));
inv_hvt I211_3_ ( .A(net294[0]), .Y(s_rdin[3]));
inv_hvt I211_2_ ( .A(net294[1]), .Y(s_rdin[2]));
inv_hvt I211_1_ ( .A(net294[2]), .Y(s_rdin[1]));
inv_hvt I211_0_ ( .A(net294[3]), .Y(s_rdin[0]));
ml_rdhv_gen Iml_rdhv_inv_3_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[3]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[3]));
ml_rdhv_gen Iml_rdhv_inv_2_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[2]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[2]));
ml_rdhv_gen Iml_rdhv_inv_1_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[1]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[1]));
ml_rdhv_gen Iml_rdhv_inv_0_ ( .srdsup_hv(sbhvsup_hv),
     .s_rdin(s_rdin[0]), .vddp_tieh(vddp_tieh),
     .s_rdin_hv(s_rdin_hv[0]));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net299), .S(vddp_));
ml_hv_hotswitch_enhance Ixcvr_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(vppint_ext_25), .hv_in_hv(vpp_int), .hv_out_hv(vpp));
ml_hvmux_top_ctrl Ihvmux_top_ctrl ( .fsm_tm_rprd(fsm_tm_rprd),
     .vpint_en(vpint_en), .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl),
     .tm_testdec(tm_testdec), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_lshven(fsm_lshven), .ysup25_2vddp(ysup25_2vddp),
     .ysup25_2vdd(ysup25_2vdd), .vtmode(vtmode),
     .vpxaint_ext(vpxaint_ext), .vpxa_vpxaint(vpxa_vpxaint),
     .vpxa_vppd(vpxa_vppd), .vpxa_ext(vpxa_ext),
     .vppint_ext(vppint_ext), .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .en_vblinhi(en_vblinhi),
     .bgrint_en(bgrint_en), .bgrext_en(bgrext_en));
ml_hvmux_ls25 Ihvmux_ls25 ( .ysup25_2vddp(ysup25_2vddp),
     .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vppint_25(sbhvsup_vppint_25), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en), .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vtmode_25(vtmode_25),
     .vpxaint_ext_25(vpxaint_ext_25),
     .vpxa_vpxaint_25(vpxa_vpxaint_25), .vpxa_vppd_25(vpxa_vppd_25),
     .vpxa_ext_25(net309), .vppint_ext_25(vppint_ext_25),
     .sbhvsup_vddp_25(sbhvsup_vddp_25),
     .sb25sup_vpxa_25(sb25sup_vpxa_25),
     .sb25sup_vddp_25(sb25sup_vddp_25), .ngate_vpxa_25(ngate_vpxa_25),
     .ngate_vddp_25(ngate_vddp_25), .bgrint_en_25(bgrint_en_25),
     .bgrext_en_25(bgrext_en_25));
ml_hvmux_bgrxcvr Ixcvr_bgr ( .vddp_tieh(vddp_tieh),
     .bgrext_en_25(bgrext_en_25), .vpp(vpp),
     .bgrint_en_25(bgrint_en_25), .bgr_int(bgr_int), .bgr(bgr));
ml_hv_hotswitch Ixcvr_vpxa_int ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa_int), .hv_out_hv(vpp));
ml_hvmux_hotswitch I212 ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(srdsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sbhvsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(sbhvsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sb25sup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sb25sup_vpxa_25), .sel_hv_a_25(sb25sup_vddp_25),
     .out_hv(sb25sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_ngate ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(ngate_vpxa_25), .sel_hv_a_25(ngate_vddp_25),
     .out_hv(ngate_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_1_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vddp_), .hvin_a_hv(vpxa_int));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_0_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vddp_), .hvin_a_hv(vpxa_int));
ml_ysup_25_switch Isw_ysup25_1_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ysup_25_switch Isw_ysup25_0_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_1_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_0_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_hvsw_8f, View - schematic
// LAST TIME SAVED: Nov  6 17:49:25 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_chip_nvcm_hvsw_8f ( s_rdin_hv, bgr, ngate_25, sb25sup_25,
     sbhvsup_hv, srdsup_hv, vblinhi, vpp, vpp_int, vpxa, ysup_25,
     fsm_bgr_dis, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint,
     fsm_tm_xvpxaint, fsm_trim_vbg, fsm_vpgmwl, fsm_vrdwl, fsm_wgnden,
     fsm_wpen, s_rd, tm_allbl_l, tm_wleqbl );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, srdsup_hv, vblinhi, vpp,
     vpp_int, vpxa, ysup_25;

input  fsm_bgr_dis, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_wleqbl;

output [3:0]  s_rdin_hv;

input [2:0]  fsm_vrdwl;
input [3:0]  fsm_trim_vbg;
input [3:0]  s_rd;
input [2:0]  fsm_vpgmwl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  fsm_vrdw_buf;

wire  [3:0]  fsm_trim_vbg_buf;



ml_chip_buf_hvsw_8f Ichip_buf_top ( .fsm_bgr_dis(fsm_bgr_dis),
     .fsm_pumpen_buf(fsm_pumpen_buf),
     .fsm_vrdwl_buf(fsm_vrdw_buf[2:0]), .fsm_vrdwl(fsm_vrdwl[2:0]),
     .fsm_tm_xvpxaint_buf(net193),
     .fsm_tm_xforce_buf(fsm_tm_xforce_buf),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_bgr_dis_buf(fsm_bgr_dis_buf), .fsm_pumpen(fsm_pumpen),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]), .fsm_nvcmen(fsm_nvcmen),
     .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen_buf));
ml_bgr_top Ibgr_top ( .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .fsm_bgr_dis_buf(fsm_bgr_dis_buf), .bgr_int(bgr_int));
ml_vppint_top Ivppint_top ( .vpxa(vpxa),
     .fsm_vpgmwl_buf(fsm_vpgmwl[2:0]), .fsm_pgmdisc_buf(fsm_pgmdisc),
     .fsm_pgm_buf(fsm_pgm), .fsm_lshven_buf(fsm_lshven),
     .vpint_en(vpint_en), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmvfy_buf(fsm_pgmvfy), .fsm_wgnden_buf(fsm_wgnden),
     .fsm_nvcmen_buf(fsm_nvcmen), .bgr(bgr), .vpp_int(vpp_int),
     .fsm_tm_xvppint(fsm_tm_xvppint));
ml_vpxa_top Ivpxa_top ( .fsm_vrdwl(fsm_vrdw_buf[2:0]),
     .fsm_tm_xvpxaint(net193), .fsm_tm_xforce(fsm_tm_xforce_buf),
     .bgr(bgr), .vpxa_int(vpxa_int), .fsm_pumpen(fsm_pumpen_buf));
ml_hvmux_top Ihvmux_top ( .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_lshven(fsm_lshven), .bgr(bgr), .bgr_int(bgr_int),
     .ngate_25(ngate_25), .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .vpp(vpp), .vpp_int(vpp_int),
     .vpxa(vpxa), .ysup_25(ysup_25), .vblinhi(vblinhi),
     .tm_testdec(fsm_tm_testdec), .srdsup_hv(srdsup_hv),
     .s_rd(s_rd[3:0]), .fsm_tm_rprd(fsm_tm_rprd),
     .s_rdin_hv(s_rdin_hv[3:0]), .vpint_en(vpint_en),
     .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl), .vpxa_int(vpxa_int));

endmodule
// Library - NVCM_40nm, Cell - ml_chip_nvcm_1f, View - schematic
// LAST TIME SAVED: Dec 30 15:10:46 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_chip_nvcm_1f ( nv_dataout, vpp, fsm_bgr_dis, fsm_blkadd,
     fsm_blkadd_b, fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven,
     fsm_multibl_read, fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rowadd, fsm_rst_b,
     fsm_sample, fsm_tm_rd_mode, fsm_tm_ref, fsm_tm_rprd,
     fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxaint, fsm_trim_ipp, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_trim_vbg, fsm_vpgmwl, fsm_vpxaset, fsm_vrdwl,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr, tm_wleqbl );

inout  vpp;

input  fsm_bgr_dis, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_rprd, fsm_tm_testdec, fsm_tm_trow,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxaint,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl;

output [8:0]  nv_dataout;

input [3:0]  fsm_blkadd_b;
input [2:0]  fsm_trim_rrefpgm;
input [9:0]  fsm_coladd;
input [3:0]  fsm_trim_vbg;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_vrdwl;
input [1:0]  fsm_tm_ref;
input [2:0]  fsm_vpgmwl;
input [7:0]  fsm_rowadd;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_rdin_hv;

wire  [3:0]  s_rd;



ml_chip_nvcm_core_1f Iml_chip_nvcm_core_1f (
     .fsm_tm_ref(fsm_tm_ref[1:0]), .fsm_wren(fsm_wren),
     .fsm_tm_rprd(fsm_tm_rprd), .s_rdin_hv(s_rdin_hv[3:0]),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout(nv_dataout[8:0]),
     .fsm_pgmhv(fsm_pgmhv), .fsm_gwlbdis(fsm_gwlbdis),
     .vpp_int(vpp_int), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_pgm(fsm_pgm),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_din(fsm_din), .fsm_rd(fsm_rd), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_rst_b(fsm_rst_b),
     .fsm_sample(fsm_sample), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_pgmdisc(fsm_pgmdisc),
     .tm_allbl_h(tm_allbl_h), .tm_allbl_l(tm_allbl_l),
     .ngate_25(ngate_25), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol), .bgr(bgr),
     .fsm_blkadd(fsm_blkadd[3:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_coladd(fsm_coladd[9:0]), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi(vblinhi), .s_rd(s_rd[3:0]), .srdsup_hv(srdsup_hv),
     .ysup_25(ysup_25), .vpxa(vpxa));
ml_chip_nvcm_hvsw_8f Ihvsw ( .bgr(bgr),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .vpp_int(vpp_int), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd), .fsm_wpen(fsm_wpen),
     .s_rdin_hv(s_rdin_hv[3:0]), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .srdsup_hv(srdsup_hv), .s_rd(s_rd[3:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .tm_allbl_l(tm_allbl_l),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_pumpen(fsm_pumpen), .sb25sup_25(sb25sup_25),
     .fsm_lshven(fsm_lshven), .sbhvsup_hv(sbhvsup_hv), .vpxa(vpxa),
     .ysup_25(ysup_25), .ngate_25(ngate_25), .fsm_wgnden(fsm_wgnden),
     .vblinhi(vblinhi), .tm_wleqbl(tm_wleqbl), .vpp(vpp),
     .fsm_vrdwl(fsm_vrdwl[2:0]), .fsm_bgr_dis(fsm_bgr_dis),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_vpgmwl(fsm_vpgmwl[2:0]), .fsm_tm_testdec(fsm_tm_testdec));
nmoscap_25  C0 ( .MINUS(GND_), .PLUS(vddp_));
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(vddp_));

endmodule
// Library - ice8chip, Cell - sg_bufx10_ice8p, View - schematic
// LAST TIME SAVED: Sep  1 14:14:18 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module sg_bufx10_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - misc, Cell - nvcm_top_ice8p, View - schematic
// LAST TIME SAVED: Nov 17 16:51:37 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module nvcm_top_ice8p ( bp0, fsm_blkadd, fsm_blkadd_b, fsm_coladd,
     fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_redrow,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_recall,
     fsm_rowadd, fsm_sample, fsm_tm_allbank_sel, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_bgr_dis,
     fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_ref,
     fsm_tm_rprd, fsm_tm_tcol, fsm_tm_testdec, fsm_tm_testdec_wr,
     fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvpp, fsm_tm_xvpxa_int, fsm_trim_ipp,
     fsm_trim_multibl_read, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_trim_vbg, fsm_trim_vpgmwl, fsm_trim_vrdwl, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b, status_wip, clk,
     nv_dataout, nvcm_ce_b, nvcm_max_coladd, nvcm_max_rowadd, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_redrow, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_recall, fsm_sample, fsm_tm_allbank_sel,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_bgr_dis, fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode,
     fsm_tm_rprd, fsm_tm_tcol, fsm_tm_testdec, fsm_tm_testdec_wr,
     fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvpp, fsm_tm_xvpxa_int, fsm_trim_multibl_read, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b, status_wip;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

output [3:0]  fsm_blkadd_b;
output [8:0]  fsm_rowadd;
output [1:0]  fsm_tm_ref;
output [11:0]  fsm_coladd;
output [2:0]  fsm_trim_vrdwl;
output [3:0]  fsm_trim_vbg;
output [3:0]  fsm_blkadd;
output [3:0]  fsm_trim_ipp;
output [2:0]  fsm_trim_vpgmwl;
output [2:0]  fsm_trim_rrefrd;
output [2:0]  fsm_trim_rrefpgm;

input [11:0]  nvcm_max_coladd;
input [8:0]  nvcm_max_rowadd;
input [8:0]  nv_dataout;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - ice1chip, Cell - nvcm_ml_block_ice1f, View - schematic
// LAST TIME SAVED: Mar  2 18:16:48 2011
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module nvcm_ml_block_ice1f ( bp0, fsm_recall, fsm_tm_margin0_read,
     nvcm_boot, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b, vpp,
     clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b;

inout  vpp;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  fsm_blkadd;

wire  [2:0]  fsm_trim_vrdwl;

wire  [2:0]  fsm_trim_vpgmwl;

wire  [3:0]  fsm_trim_vbg;

wire  [2:0]  fsm_trim_rrefrd;

wire  [2:0]  fsm_trim_rrefpgm;

wire  [3:0]  fsm_trim_ipp;

wire  [8:0]  nv_dataout;

wire  [3:0]  fsm_blkadd_b;

wire  [1:0]  fsm_tm_ref_buf;

wire  [11:0]  fsm_coladd;

wire  [8:0]  fsm_rowadd;



ml_chip_nvcm_1f I_ml_chip_nvcm ( .fsm_tm_ref(fsm_tm_ref_buf[1:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .fsm_bgr_dis(fsm_bgr_dis),
     .tm_allbank_sel(fsm_tm_allbank_sel), .fsm_coladd(fsm_coladd[9:0]),
     .tm_wleqbl(fsm_tm_vwleqbl), .tm_testdec_wr(fsm_tm_testdec_wr),
     .tm_tcol(fsm_tm_tcol), .tm_dma(fsm_tm_dma),
     .tm_allwl_l(fsm_tm_allwl_l), .tm_allwl_h(fsm_tm_allwl_h),
     .tm_allbl_l(fsm_tm_allbl_l), .tm_allbl_h(fsm_tm_allbl_h),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vrdwl(fsm_trim_vrdwl[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxaint(fsm_tm_xvpxa_int), .fsm_tm_xvppint(fsm_tm_xvpp),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(rst_bd), .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rrow(fsm_nv_redrow), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_multibl_read(fsm_trim_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .nv_dataout(nv_dataout[8:0]), .vpp(vpp));
tiehi I442 ( .tiehi(tvdd_fsm));
tielo I369 ( .tielo(tgnd_fsm));
sg_bufx10_ice8p I541 ( .in(rst_b), .out(rst_bd));
nvcm_top_ice8p I_nvcm_top_ice8p ( .fsm_tm_bgr_dis(fsm_bgr_dis),
     .fsm_tm_allbank_sel(fsm_tm_allbank_sel),
     .fsm_coladd(fsm_coladd[11:0]), .nvcm_max_coladd({tgnd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tgnd_fsm, tvdd_fsm, tgnd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm, tvdd_fsm}),
     .nvcm_max_rowadd({tgnd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm,
     tgnd_fsm, tgnd_fsm, tvdd_fsm, tvdd_fsm, tvdd_fsm}),
     .status_wip(net249), .fsm_tm_ref(fsm_tm_ref_buf[1:0]),
     .fsm_tm_rprd(fsm_tm_rprd), .nvcm_boot(nvcm_boot),
     .spi_ss_b(spi_ss_b), .spi_sdi(spi_sdi),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_ce_b(nvcm_ce_b), .nv_dataout(nv_dataout[8:0]), .clk(clk),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .nvcm_relextspi(nvcm_relextspi), .nvcm_rdy(nvcm_rdy),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_tm_xvbg(fsm_tm_xvbg),
     .fsm_trim_vrdwl(fsm_trim_vrdwl[2:0]),
     .fsm_trim_vpgmwl(fsm_trim_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_multibl_read(fsm_trim_multibl_read),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_xvpxa_int(fsm_tm_xvpxa_int), .fsm_tm_xvpp(fsm_tm_xvpp),
     .fsm_tm_xforce(fsm_tm_xforce), .fsm_tm_vwleqbl(fsm_tm_vwleqbl),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_testdec_wr(fsm_tm_testdec_wr),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_tcol(fsm_tm_tcol),
     .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_margin0_read(fsm_tm_margin0_read),
     .fsm_tm_dma(fsm_tm_dma), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_sample(fsm_sample),
     .fsm_rowadd(fsm_rowadd[8:0]), .fsm_recall(fsm_recall),
     .fsm_rd(fsm_rd), .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmien(fsm_pgmien), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_redrow(fsm_nv_redrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_din(fsm_din),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .bp0(bp0));

endmodule
// Library - leafcell, Cell - bram_bufferx16_2inv, View - schematic
// LAST TIME SAVED: May 13 10:13:11 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_bufferx16_2inv ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I4 ( .A(net6), .Y(out));
inv I3 ( .A(in), .Y(net6));

endmodule
// Library - xpmem, Cell - ml_dff_bl, View - schematic
// LAST TIME SAVED: May 11 18:38:30 2010
// NETLIST TIME: May  5 11:56:46 2011
`timescale 1ns / 1ns 

module ml_dff_bl ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_clk_buf, View - schematic
// LAST TIME SAVED: Aug  9 18:57:25 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_clk_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_powersurg_buf, View - schematic
// LAST TIME SAVED: Jun 18 17:30:09 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_powersurg_buf ( o, in );
output  o;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I404 ( .A(net016), .Y(net012));
inv_hvt I405 ( .A(net012), .Y(o));
inv_hvt I391 ( .A(net77), .Y(net016));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_sch, View - schematic
// LAST TIME SAVED: Nov  8 11:11:57 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_sch ( dataout, bl, prec_sup, cram_prec, cram_pullup_b,
     cram_write, data_muxsel, datain, latch_clock, latch_reset,
     prec_hold_b, smc_wdic_clk );
output  dataout;

inout  bl, prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, datain,
     latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff Idff ( .R(latch_reset), .D(dff_in), .CLK(latch_clock),
     .QN(write_data_b), .Q(dff_data));
pch_hvt  MP8 ( .D(net0148), .B(vdd_), .G(dataout), .S(vdd_));
pch_hvt  MP9 ( .D(bl), .B(vdd_), .G(net084), .S(net0148));
pch_hvt  M0 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  M3 ( .D(net0110), .B(vdd_), .G(cram_write), .S(prec_sup));
pch_hvt  MP12 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  M2 ( .D(bl), .B(vdd_), .G(prec_hold_b), .S(net0110));
pch_hvt  MP4 ( .D(net0143), .B(vdd_), .G(cram_pullup_b), .S(vdd_));
pch_hvt  MP5 ( .D(sa_out), .B(vdd_), .G(bl), .S(net0143));
nch_hvt  MN12 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN8 ( .D(sa_out), .B(gnd_), .G(cram_pullup_b), .S(gnd_));
nch_hvt  M1 ( .D(net0166), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN3 ( .D(sa_out), .B(gnd_), .G(bl), .S(gnd_));
nch_hvt  MN6 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
nor2_hvt I223 ( .A(net084), .B(write_data_b), .Y(n_gate));
inv_hvt I163 ( .A(write_data_b), .Y(dataout));
inv_hvt I159 ( .A(cram_prec), .Y(net0161));
inv_hvt I160 ( .A(cram_write), .Y(net084));
mux2_hvt I161 ( .in1(sa_out), .in0(datain), .out(latch_in),
     .sel(data_muxsel));
mux2_hvt I164 ( .in1(dff_data), .in0(latch_in), .out(dff_in),
     .sel(smc_wdic_clk));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_bram10k, View - schematic
// LAST TIME SAVED: Aug  4 18:43:48 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tile_bram10k ( cram_prec_out, cram_write_out, data_out,
     para_out, bl, prec_sup, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, datain, latch_clock, latch_reset,
     para_en, para_in, prec_hold_b, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out, para_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, para_en, para_in, prec_hold_b,
     smc_wdic_clk;

inout [41:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:0]  data_in;

wire  [4:1]  data_dummy_in;

wire  [14:0]  ck;

wire  [41:0]  dataout;



mux2_hvt I216 ( .in1(net119), .in0(dataout[6]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I208 ( .in1(data_dummy_in[2]), .in0(dataout[3]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I209 ( .in1(data_dummy_in[3]), .in0(dataout[4]),
     .out(data_in[3]), .sel(data_muxsel1));
mux2_hvt I196 ( .in1(data_dummy_in[1]), .in0(dataout[2]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I210 ( .in1(data_dummy_in[4]), .in0(dataout[5]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I217 ( .in1(para_in), .in0(dataout[1]), .out(data_out_mux),
     .sel(para_en));
inv_hvt I262 ( .A(data_out_mux), .Y(net151));
inv_hvt I261 ( .A(net151), .Y(data_in[0]));
inv_hvt I175 ( .A(dataout[1]), .Y(net154));
inv_hvt I176 ( .A(net154), .Y(para_out));
inv_hvt I172 ( .A(net160), .Y(data_out));
inv_hvt I171 ( .A(dataout[41]), .Y(net160));
inv_hvt I201 ( .A(latch_clock), .Y(net0133));
inv_hvt I207 ( .A(net0105), .Y(ck[14]));
inv_hvt I206 ( .A(net0107), .Y(net0105));
inv_hvt I205 ( .A(net0133), .Y(net0107));
ml_dff_bl I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net97), .Q(net119));
ml_dff_bl I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net92), .Q(data_dummy_in[4]));
ml_dff_bl I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net87), .Q(data_dummy_in[2]));
ml_dff_bl I179 ( .R(latch_reset), .D(data_in[0]), .CLK(ck[14]),
     .QN(net82), .Q(data_dummy_in[1]));
ml_dff_bl I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net77), .Q(data_dummy_in[3]));
ml_blsa_clk_buf I192_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I192_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I192_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I192_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I192_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I192_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I192_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I192_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I192_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I192_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I192_0_ ( .in(latch_clock), .o(ck[0]));
ml_powersurg_buf I165 ( .in(cram_prec), .o(net162));
ml_powersurg_buf I163 ( .in(net162), .o(net164));
ml_powersurg_buf I162 ( .in(net170), .o(net166));
ml_powersurg_buf I169 ( .in(net166), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(cram_write), .o(net170));
ml_powersurg_buf I168 ( .in(net164), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[14]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[15]),
     .dataout(dataout[15]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[13]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[14]),
     .dataout(dataout[14]), .cram_prec(net164));

endmodule
// Library - xpmem, Cell - ml_blsa_tile, View - schematic
// LAST TIME SAVED: Jan  7 13:26:29 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tile ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [53:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [53:0]  dataout;

wire  [13:0]  ck;



inv_hvt I172 ( .A(net48), .Y(data_out));
inv_hvt I171 ( .A(dataout[53]), .Y(net48));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_powersurg_buf I161 ( .in(cram_write), .o(net53));
ml_powersurg_buf I165 ( .in(net57), .o(net55));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net57));
ml_powersurg_buf I163 ( .in(net55), .o(net59));
ml_powersurg_buf I162 ( .in(net65), .o(net61));
ml_powersurg_buf I169 ( .in(net61), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net53), .o(net65));
ml_powersurg_buf I168 ( .in(net59), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_47_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[47]),
     .dataout(dataout[47]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_46_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[46]),
     .dataout(dataout[46]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_45_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[45]),
     .dataout(dataout[45]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_44_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[44]),
     .dataout(dataout[44]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_43_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[43]),
     .dataout(dataout[43]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_42_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[42]),
     .dataout(dataout[42]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net55));
ml_blsa_sch I170_53_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[53]), .dataout(dataout[53]),
     .cram_prec(net57));
ml_blsa_sch I170_52_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[52]), .dataout(dataout[52]),
     .cram_prec(net57));
ml_blsa_sch I170_51_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[51]), .dataout(dataout[51]),
     .cram_prec(net57));
ml_blsa_sch I170_50_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[50]), .dataout(dataout[50]),
     .cram_prec(net57));
ml_blsa_sch I170_49_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[49]), .dataout(dataout[49]),
     .cram_prec(net57));
ml_blsa_sch I170_48_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .data_muxsel(data_muxsel),
     .cram_write(net53), .bl(bl[48]), .dataout(dataout[48]),
     .cram_prec(net57));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net59));

endmodule
// Library - xpmem, Cell - ml_blprecwrt_en, View - schematic
// LAST TIME SAVED: Aug  5 16:47:07 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blprecwrt_en ( data_out, action, clkin, data_in, rst );
output  data_out;

input  action, clkin, data_in, rst;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor3_hvt I105 ( .B(net86), .Y(net94), .A(net98), .C(rst));
nor2_hvt I103 ( .A(net88), .B(net94), .Y(net98));
inv_hvt I66 ( .A(net89), .Y(net88));
inv_hvt I168 ( .A(action), .Y(net86));
inv_hvt I165 ( .A(net98), .Y(data_out));
nand3_hvt I160 ( .Y(net89), .B(data_in), .C(action), .A(clkin));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_bram10k, View - schematic
// LAST TIME SAVED: Oct 20 17:35:57 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex2_bram10k ( data_out, latch_clock_out, para_out,
     prec_out, wrt_out, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, datain, latch_clock_in, latch_reset,
     para_en, para_in, prec_in, smc_clk_dpr, smc_wdic_clk, smc_write,
     wrt_in );
output  data_out, latch_clock_out, para_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, para_en, para_in, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in;

inout [95:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



tiehi I284 ( .tiehi(prec_hold_b));
pch_hvt  M3 ( .D(prec_sup), .B(vdd_), .G(net095), .S(vdd_));
nor2_hvt I385 ( .A(latch_reset), .B(net092), .Y(net067));
inv_hvt I198 ( .A(prec_hold_b), .Y(net095));
inv_hvt I189 ( .A(net100), .Y(latch_clock_out));
inv_hvt I191 ( .A(latch_clock_in), .Y(net100));
inv_hvt I193 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I196 ( .A(net067), .Y(net068));
inv_hvt I197 ( .A(net0130), .Y(net0105));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));
inv_hvt I187 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I188 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I192 ( .A(latch_reset), .Y(net94));
inv_hvt I194 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I190 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I195 ( .A(smc_wdic_clk), .Y(net088));
ml_blsa_tile_bram10k tile0 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .para_en(para_en), .para_in(para_in),
     .para_out(para_out), .bl(bl[41:0]),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_out),
     .cram_prec_out(prec_en_last));
ml_blsa_tile tile1 ( .prec_sup(prec_sup), .prec_hold_b(prec_hold_b),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[95:42]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net092));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net068), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net0130));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));

endmodule
// Library - xpmem, Cell - ml_buf_ice5, View - schematic
// LAST TIME SAVED: Aug  4 15:14:20 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_buf_ice5 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_last, View - schematic
// LAST TIME SAVED: Aug  4 18:09:54 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tile_last ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [17:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:0]  ck;

wire  [17:0]  dataout;



ml_dff Idff ( .R(latch_reset), .D(dataout[16]), .CLK(ck[0]),
     .QN(net50), .Q(net45));
ml_dff I179 ( .R(latch_reset), .D(net58), .CLK(ck[0]), .QN(net49),
     .Q(net61));
mux2_hvt I174 ( .in1(net45), .in0(dataout[17]), .out(net58),
     .sel(data_muxsel));
tiehis I185 ( .tiehi(net040));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_buf_ice5 I205 ( .in(net61), .o(data_out), .sel(net040));
ml_powersurg_buf I169 ( .in(cram_write), .o(cram_write_out));
ml_powersurg_buf I168 ( .in(cram_prec), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[16]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[17]), .dataout(dataout[17]));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[15]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[16]), .dataout(dataout[16]));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));

endmodule
// Library - leafcell, Cell - bram_sdo_reg, View - schematic
// LAST TIME SAVED: Jul  8 11:50:49 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_sdo_reg ( do, tielo, clk, di );
output  do, tielo;

input  clk, di;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff I_bm_sdo_dff ( .R(tielo), .D(di), .CLK(clk), .QN(net11),
     .Q(net018));
bram_bufferx16_2inv I51 ( .in(net018), .out(do));
tielo I_tielo ( .tielo(tielo));

endmodule
// Library - leafcell, Cell - bram_bufferx4, View - schematic
// LAST TIME SAVED: Aug 12 09:08:27 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module bram_bufferx4 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex1_last_ice1f, View - schematic
// LAST TIME SAVED: Jan 20 18:04:52 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex1_last_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [71:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I385 ( .A(net0111), .B(latch_reset), .Y(net0121));
ml_blsa_tile_last Iml_blsa_tile_last ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .bl(bl[71:54]),
     .latch_reset(latch_reset_buf), .datain(datain_io),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_1st), .cram_prec_out(prec_en_1st),
     .latch_clock(latch_clock_out), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blsa_tile Iml_blsa_tile_0 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_dic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_1st), .cram_prec(prec_en_1st),
     .data_out(datain_io), .cram_write_out(wrt_out),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
tiehi I284 ( .tiehi(prec_hold_b));
pch_hvt  M0 ( .D(prec_sup), .B(vdd_), .G(vdd_), .S(vdd_));
inv_hvt I197 ( .A(prec_hold_b), .Y(vdd_));
inv_hvt I194 ( .A(smc_wdic_clk), .Y(net0125));
inv_hvt I196 ( .A(net0124), .Y(net066));
inv_hvt I187 ( .A(net0121), .Y(net068));
inv_hvt I193 ( .A(latch_reset), .Y(net0127));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net0133));
inv_hvt I204 ( .A(net0137), .Y(latch_clock_out));
inv_hvt I208 ( .A(net0125), .Y(smc_dic_clk_buf));
inv_hvt I192 ( .A(latch_clock_in), .Y(net0137));
inv_hvt I190 ( .A(net0139), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net0139));
inv_hvt I203 ( .A(net0133), .Y(cram_pullup_b_buf));
inv_hvt I207 ( .A(net0127), .Y(latch_reset_buf));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net068), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net0124));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net0111));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex1_ice1f, View - schematic
// LAST TIME SAVED: Jan 20 17:58:11 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex1_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [53:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_0 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_out), .cram_prec_out(prec_en_last),
     .bl(bl[53:0]));
tiehi I284 ( .tiehi(prec_hold_b));
pch_hvt  M3 ( .D(prec_sup), .B(vdd_), .G(net075), .S(vdd_));
nor2_hvt I385 ( .A(latch_reset), .B(net049), .Y(net051));
inv_hvt I186 ( .A(data_muxsel), .Y(net084));
inv_hvt I190 ( .A(net084), .Y(data_muxsel_buf));
inv_hvt I199 ( .A(latch_clock_in), .Y(net0100));
inv_hvt I200 ( .A(prec_hold_b), .Y(net075));
inv_hvt I221 ( .A(net096), .Y(net054));
inv_hvt I201 ( .A(net051), .Y(net052));
inv_hvt I198 ( .A(net0100), .Y(latch_clock_out));
inv_hvt I197 ( .A(net090), .Y(cram_pullup_b_buf));
inv_hvt I205 ( .A(smc_wdic_clk), .Y(net094));
inv_hvt I204 ( .A(net094), .Y(smc_wdic_clk_buf));
inv_hvt I196 ( .A(cram_pullup_b), .Y(net090));
inv_hvt I203 ( .A(net086), .Y(latch_reset_buf));
inv_hvt I202 ( .A(latch_reset), .Y(net086));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net052), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net096));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net049));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_1st, View - schematic
// LAST TIME SAVED: Aug  4 18:53:38 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tile_1st ( cram_prec_out, cram_write_out, data_out, bl,
     prec_sup, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, prec_hold_b,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;

inout  prec_sup;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, prec_hold_b, smc_wdic_clk;

inout [55:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:1]  data_dummy_in;

wire  [55:0]  dataout;

wire  [5:1]  data_in;

wire  [14:0]  ck;



ml_dff I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net132), .Q(net154));
ml_dff I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net137), .Q(data_dummy_in[4]));
ml_dff I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net142), .Q(data_dummy_in[2]));
ml_dff I179 ( .R(latch_reset), .D(datain), .CLK(ck[14]), .QN(net147),
     .Q(data_dummy_in[1]));
ml_dff I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net152), .Q(data_dummy_in[3]));
inv_hvt I171 ( .A(dataout[55]), .Y(net121));
inv_hvt I172 ( .A(net121), .Y(data_out));
inv_hvt I224 ( .A(net0130), .Y(ck[14]));
inv_hvt I225 ( .A(net0129), .Y(net0130));
inv_hvt I226 ( .A(net0126), .Y(net0129));
inv_hvt I229 ( .A(latch_clock), .Y(net0122));
inv_hvt I227 ( .A(net0124), .Y(net0126));
inv_hvt I228 ( .A(net0122), .Y(net0124));
mux2_hvt I197 ( .in1(net154), .in0(dataout[4]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I232 ( .in1(data_dummy_in[2]), .in0(dataout[1]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I230 ( .in1(data_dummy_in[4]), .in0(dataout[3]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I233 ( .in1(data_dummy_in[1]), .in0(dataout[0]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I231 ( .in1(data_dummy_in[3]), .in0(dataout[2]),
     .out(data_in[3]), .sel(data_muxsel1));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_blsa_sch Iml_blsa_sch_15_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[14]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_14_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[13]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_13_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[12]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_12_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[11]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_11_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[10]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_10_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[9]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_9_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[8]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_8_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[7]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_7_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[6]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_6_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_5_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_4_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[4]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_3_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[3]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_2_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[2]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_1_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[1]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_0_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(datain), .cram_prec(cram_prec_out),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_47_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[47]),
     .dataout(dataout[47]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_46_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[46]),
     .dataout(dataout[46]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_45_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[45]),
     .dataout(dataout[45]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_44_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[44]),
     .dataout(dataout[44]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_43_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[43]),
     .dataout(dataout[43]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_42_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[42]),
     .dataout(dataout[42]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_41_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[41]),
     .dataout(dataout[41]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_40_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[40]),
     .dataout(dataout[40]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_39_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[39]),
     .dataout(dataout[39]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_38_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[38]),
     .dataout(dataout[38]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_37_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[37]),
     .dataout(dataout[37]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_36_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[36]),
     .dataout(dataout[36]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_35_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[35]),
     .dataout(dataout[35]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_34_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[34]),
     .dataout(dataout[34]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_33_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[33]),
     .dataout(dataout[33]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_32_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[32]),
     .dataout(dataout[32]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_55_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[54]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[55]),
     .dataout(dataout[55]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_54_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[53]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[54]),
     .dataout(dataout[54]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_53_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[53]),
     .dataout(dataout[53]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_52_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[52]),
     .dataout(dataout[52]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_51_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[51]),
     .dataout(dataout[51]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_50_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[50]),
     .dataout(dataout[50]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_49_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[49]),
     .dataout(dataout[49]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_48_ ( .prec_hold_b(prec_hold_b), .prec_sup(prec_sup),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[48]),
     .dataout(dataout[48]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_31_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[31]),
     .dataout(dataout[31]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_30_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[30]),
     .dataout(dataout[30]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_29_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[29]),
     .dataout(dataout[29]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_28_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[28]),
     .dataout(dataout[28]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_27_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[27]),
     .dataout(dataout[27]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_26_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[26]),
     .dataout(dataout[26]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_25_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[25]),
     .dataout(dataout[25]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_24_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[24]),
     .dataout(dataout[24]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_23_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[23]),
     .dataout(dataout[23]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_22_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[22]),
     .dataout(dataout[22]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_21_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[21]),
     .dataout(dataout[21]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_20_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[20]),
     .dataout(dataout[20]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_19_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[19]),
     .dataout(dataout[19]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_18_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[18]),
     .dataout(dataout[18]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_17_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[17]),
     .dataout(dataout[17]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_16_ ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[16]),
     .dataout(dataout[16]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_powersurg_buf I161 ( .in(cram_write), .o(net104));
ml_powersurg_buf I165 ( .in(net108), .o(net106));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net108));
ml_powersurg_buf I163 ( .in(net106), .o(net110));
ml_powersurg_buf I162 ( .in(net116), .o(net112));
ml_powersurg_buf I169 ( .in(net112), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net104), .o(net116));
ml_powersurg_buf I168 ( .in(net110), .o(cram_prec_out));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_1st_ice1f, View - schematic
// LAST TIME SAVED: Jan 20 17:52:04 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_tilex2_1st_ice1f ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, smc_write, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, smc_write, wrt_in;

inout [109:0]  bl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_1 ( .prec_hold_b(prec_hold_b),
     .prec_sup(prec_sup), .cram_pullup_b(cram_pullup_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_wdic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_in), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[109:56]));
ml_blsa_tile_1st Iml_blsa_tile_1st_0 ( .prec_sup(prec_sup),
     .prec_hold_b(prec_hold_b), .bl(bl[55:0]),
     .cram_pullup_b(cram_pullup_buf), .latch_clock(latch_clock_out),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .datain(datain), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_mid),
     .cram_prec(prec_en_mid), .data_out(data_tile),
     .cram_write_out(wrt_out), .cram_prec_out(prec_en_last));
nor2_hvt I385 ( .A(latch_reset), .B(net86), .Y(net117));
pch_hvt  M3 ( .D(prec_sup), .B(vdd_), .G(net106), .S(vdd_));
tiehi I284 ( .tiehi(prec_hold_b));
inv_hvt I190 ( .A(net095), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net095));
inv_hvt I202 ( .A(latch_reset), .Y(net0113));
inv_hvt I203 ( .A(net0113), .Y(latch_reset_buf));
inv_hvt I196 ( .A(cram_pullup_b), .Y(net0109));
inv_hvt I204 ( .A(net0105), .Y(smc_wdic_clk_buf));
inv_hvt I200 ( .A(prec_hold_b), .Y(net106));
inv_hvt I205 ( .A(smc_wdic_clk), .Y(net0105));
inv_hvt I221 ( .A(net138), .Y(net110));
inv_hvt I197 ( .A(net0109), .Y(cram_pullup_buf));
inv_hvt I198 ( .A(net099), .Y(latch_clock_out));
inv_hvt I199 ( .A(latch_clock_in), .Y(net099));
inv_hvt I201 ( .A(net117), .Y(net118));
ml_blprecwrt_en Iprec_hd_wrt ( .rst(net118), .data_in(prec_out),
     .clkin(prec_out), .action(smc_write), .data_out(net138));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(net86));

endmodule
// Library - xpmem, Cell - ml_buf_ice1f, View - schematic
// LAST TIME SAVED: Jan  7 14:21:36 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_buf_ice1f ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_bank_ice1f, View - schematic
// LAST TIME SAVED: Mar  8 09:38:22 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_blsa_bank_ice1f ( cm_sdo_u, bl, banksel, cm_sdi_u,
     cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk,
     smc_write );


input  banksel, cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk,
     smc_write;

output [1:0]  cm_sdo_u;

inout [331:0]  bl;

input [1:0]  cm_sdi_u;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tilex2_bram10k I_lt_34 ( .smc_write(smc_write_buf),
     .para_en(cor_en_8bpcfg_buf), .para_in(sdi1_buf),
     .para_out(para_out), .bl(bl[259:164]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net0137),
     .latch_clock_out(net0171), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret), .wrt_in(wrt_out_5),
     .prec_in(prec_out_5), .latch_reset(latch_reset_buf),
     .datain(data_out_2), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_34),
     .prec_out(prec_out_34), .data_out(data_out_34));
ml_blsa_tilex1_last_ice1f I_lt_5 ( .smc_write(smc_write_buf),
     .bl(bl[331:260]), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(smc_clk), .latch_clock_out(net0137),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf),
     .wrt_in(cram_write_buf), .prec_in(net377),
     .latch_reset(latch_reset_buf), .datain(data_out_34),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_5), .prec_out(prec_out_5),
     .data_out(cm_sdo_u[1]));
ml_blsa_tilex1_ice1f I_lt_2 ( .smc_write(smc_write_buf),
     .bl(bl[163:110]), .cram_pullup_b(net0161),
     .latch_clock_in(net0171), .latch_clock_out(net393),
     .smc_wdic_clk(net0158), .smc_clk_dpr(net0165),
     .wrt_in(wrt_out_34), .prec_in(prec_out_34),
     .latch_reset(latch_reset_buf), .datain(data_out_01),
     .data_muxsel1(net0152), .data_muxsel(net0149),
     .cram_write(net0146), .cram_prec(net0155), .wrt_out(wrt_out_2),
     .prec_out(prec_out_2), .data_out(data_out_2));
ml_blsa_tilex2_1st_ice1f I_lt_01 ( .smc_write(smc_write_buf),
     .wrt_in(wrt_out_2), .prec_in(prec_out_2),
     .latch_reset(latch_reset_buf), .datain(net0140),
     .data_muxsel1(net0152), .data_muxsel(net0149),
     .cram_write(net0146), .bl(bl[109:0]), .cram_prec(net0155),
     .wrt_out(wrt_out_01), .prec_out(prec_out_01),
     .data_out(data_out_01), .latch_clock_in(net393),
     .cram_pullup_b(net0161), .latch_clock_out(net440),
     .smc_wdic_clk(net0158), .smc_clk_dpr(net0354));
ml_buf_ice1f I291 ( .in(net0160), .o(net0165),
     .sel(smc_clk_buf_b_ret));
ml_buf_ice1f I292 ( .in(net0160), .o(net0354), .sel(smc_clk_buf));
ml_buf_ice1f I284 ( .in(net0160), .o(net0140), .sel(sdi0_buf));
ml_buf_ice1f I247 ( .in(cm_sdi_u[1]), .o(sdi1_buf), .sel(net527));
ml_buf_ice1f I249 ( .in(net519), .o(cor_en_8bpcfg_buf), .sel(net527));
ml_buf_ice1f I285 ( .in(net0160), .o(net0146), .sel(cram_write_buf));
ml_buf_ice1f I265 ( .in(net527), .o(cm_sdo_u[0]), .sel(net451));
ml_buf_ice1f I257 ( .in(smc_wdic_clk), .o(smc_wdic_clk_buf),
     .sel(banksel));
ml_buf_ice1f I203 ( .in(data_muxsel1), .o(data_muxsel1_buf),
     .sel(banksel));
ml_buf_ice1f I205 ( .in(latch_reset), .o(latch_reset_buf),
     .sel(net529));
ml_buf_ice1f I207 ( .in(cram_write), .o(cram_write_buf),
     .sel(banksel));
ml_buf_ice1f I208 ( .in(cram_pullup_logic_b), .o(cram_pullup_b_buf),
     .sel(cram_pullup_logic_b));
ml_buf_ice1f I288 ( .in(net0160), .o(net0149), .sel(data_muxsel_buf));
ml_buf_ice1f I201 ( .in(cram_prec), .o(cram_prec_buf), .sel(banksel));
ml_buf_ice1f I289 ( .in(net0160), .o(net0152), .sel(data_muxsel1_buf));
ml_buf_ice1f I294b ( .in(banksel), .o(smc_write_buf), .sel(smc_write));
ml_buf_ice1f I216 ( .in(net528), .o(net474), .sel(net528));
ml_buf_ice1f I286 ( .in(net0160), .o(net0155), .sel(cram_prec_buf));
ml_buf_ice1f I8 ( .in(net0160), .o(net0158), .sel(smc_wdic_clk_buf));
ml_buf_ice1f I290 ( .in(net0160), .o(net0161),
     .sel(cram_pullup_b_buf));
ml_buf_ice1f I245 ( .in(cm_sdi_u[0]), .o(sdi0_buf), .sel(net527));
ml_buf_ice1f I187 ( .in(smc_clk), .o(smc_clk_buf), .sel(smc_clk));
ml_buf_ice1f I188 ( .in(net525), .o(smc_clk_buf_b_ret), .sel(net525));
ml_buf_ice1f I204 ( .in(data_muxsel), .o(data_muxsel_buf),
     .sel(banksel));
ml_buf_ice1f I227 ( .in(net532), .o(net489), .sel(net532));
nor3_hvt I217 ( .B(net531), .Y(net492), .A(net531), .C(net531));
nor3_hvt I220 ( .B(net500), .Y(net496), .A(net500), .C(net500));
nor3_hvt I218 ( .B(net492), .Y(net500), .A(net492), .C(net492));
nand3_hvt I231 ( .Y(net503), .B(net507), .C(net507), .A(net507));
nand3_hvt I230 ( .Y(net507), .B(net511), .C(net511), .A(net511));
nand3_hvt I224 ( .Y(net511), .B(net526), .C(net526), .A(net526));
nor2_hvt I254 ( .B(net515), .Y(net522), .A(cram_pullup_b));
inv_hvt I253 ( .A(cor_en_8bpcfg_b), .Y(net519));
inv_hvt I256 ( .A(banksel), .Y(net515));
inv_hvt I255 ( .A(net522), .Y(cram_pullup_logic_b));
inv_hvt I189 ( .A(smc_clk), .Y(net525));
tiehi I268 ( .tiehi(net526));
tiehi I272 ( .tiehi(net527));
tiehi I287 ( .tiehi(net0160));
tiehi I271 ( .tiehi(net528));
tiehi I273 ( .tiehi(net529));
tiehi I267 ( .tiehi(net377));
tiehi I270 ( .tiehi(net531));
tiehi I269 ( .tiehi(net532));
ml_dff_bl I_ml_dff_bl ( .R(latch_reset_buf), .D(para_out),
     .CLK(smc_clk), .QN(net536), .Q(net451));

endmodule
// Library - ice1chip, Cell - CHIP_route_top_ice1f, View - schematic
// LAST TIME SAVED: Mar  7 16:46:33 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module CHIP_route_top_ice1f ( cm_sdo_u1, cm_sdo_u3, bl_top,
     cm_banksel_bltld3, cm_banksel_bltrd1, cm_clk_bltld3,
     cm_clk_bltrd1, cm_prec_bltld3, cm_sdi_u1d3, cm_sdi_u3d2,
     core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1r,
     smc_write_bltl1d1, smc_write_bltld3 );


input  cm_clk_bltld3, cm_clk_bltrd1, cm_prec_bltld3, core_por_b_rowu1,
     core_por_b_rowu3, cram_prec_bltrd1, cram_pullup_b_bltrd1,
     cram_pullup_bltld3, cram_write_bltld3, cram_write_bltrd1,
     data_muxsel1_bltld3, data_muxsel1_bltrd1, data_muxsel_bltld3,
     data_muxsel_bltrd1, en_8bconfig_b_bltld3, en_8bconfig_b_bltrd1,
     smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1r, smc_write_bltl1d1,
     smc_write_bltld3;

output [1:0]  cm_sdo_u1;
output [1:0]  cm_sdo_u3;

inout [663:0]  bl_top;

input [3:3]  cm_banksel_bltrd1;
input [1:0]  cm_sdi_u1d3;
input [1:0]  cm_sdi_u3d2;
input [1:1]  cm_banksel_bltld3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_blsa_bank_ice1f I_bltr ( .smc_write(smc_write_bltl1d1),
     .bl(bl_top[663:332]), .smc_wdic_clk(smc_wdis_dclk_bltrd1r),
     .smc_clk(cm_clk_bltrd1), .cm_sdi_u(cm_sdi_u3d2[1:0]),
     .latch_reset(core_por_b_rowu3), .cm_sdo_u(cm_sdo_u3[1:0]),
     .data_muxsel1(data_muxsel1_bltrd1),
     .data_muxsel(data_muxsel_bltrd1), .cram_write(cram_write_bltrd1),
     .cram_prec(cram_prec_bltrd1),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltrd1),
     .cram_pullup_b(cram_pullup_b_bltrd1),
     .banksel(cm_banksel_bltrd1[3]));
ml_blsa_bank_ice1f I_bltlu1 ( .smc_write(smc_write_bltld3),
     .bl({bl_top[0], bl_top[1], bl_top[2], bl_top[3], bl_top[4],
     bl_top[5], bl_top[6], bl_top[7], bl_top[8], bl_top[9], bl_top[10],
     bl_top[11], bl_top[12], bl_top[13], bl_top[14], bl_top[15],
     bl_top[16], bl_top[17], bl_top[18], bl_top[19], bl_top[20],
     bl_top[21], bl_top[22], bl_top[23], bl_top[24], bl_top[25],
     bl_top[26], bl_top[27], bl_top[28], bl_top[29], bl_top[30],
     bl_top[31], bl_top[32], bl_top[33], bl_top[34], bl_top[35],
     bl_top[36], bl_top[37], bl_top[38], bl_top[39], bl_top[40],
     bl_top[41], bl_top[42], bl_top[43], bl_top[44], bl_top[45],
     bl_top[46], bl_top[47], bl_top[48], bl_top[49], bl_top[50],
     bl_top[51], bl_top[52], bl_top[53], bl_top[54], bl_top[55],
     bl_top[56], bl_top[57], bl_top[58], bl_top[59], bl_top[60],
     bl_top[61], bl_top[62], bl_top[63], bl_top[64], bl_top[65],
     bl_top[66], bl_top[67], bl_top[68], bl_top[69], bl_top[70],
     bl_top[71], bl_top[72], bl_top[73], bl_top[74], bl_top[75],
     bl_top[76], bl_top[77], bl_top[78], bl_top[79], bl_top[80],
     bl_top[81], bl_top[82], bl_top[83], bl_top[84], bl_top[85],
     bl_top[86], bl_top[87], bl_top[88], bl_top[89], bl_top[90],
     bl_top[91], bl_top[92], bl_top[93], bl_top[94], bl_top[95],
     bl_top[96], bl_top[97], bl_top[98], bl_top[99], bl_top[100],
     bl_top[101], bl_top[102], bl_top[103], bl_top[104], bl_top[105],
     bl_top[106], bl_top[107], bl_top[108], bl_top[109], bl_top[110],
     bl_top[111], bl_top[112], bl_top[113], bl_top[114], bl_top[115],
     bl_top[116], bl_top[117], bl_top[118], bl_top[119], bl_top[120],
     bl_top[121], bl_top[122], bl_top[123], bl_top[124], bl_top[125],
     bl_top[126], bl_top[127], bl_top[128], bl_top[129], bl_top[130],
     bl_top[131], bl_top[132], bl_top[133], bl_top[134], bl_top[135],
     bl_top[136], bl_top[137], bl_top[138], bl_top[139], bl_top[140],
     bl_top[141], bl_top[142], bl_top[143], bl_top[144], bl_top[145],
     bl_top[146], bl_top[147], bl_top[148], bl_top[149], bl_top[150],
     bl_top[151], bl_top[152], bl_top[153], bl_top[154], bl_top[155],
     bl_top[156], bl_top[157], bl_top[158], bl_top[159], bl_top[160],
     bl_top[161], bl_top[162], bl_top[163], bl_top[164], bl_top[165],
     bl_top[166], bl_top[167], bl_top[168], bl_top[169], bl_top[170],
     bl_top[171], bl_top[172], bl_top[173], bl_top[174], bl_top[175],
     bl_top[176], bl_top[177], bl_top[178], bl_top[179], bl_top[180],
     bl_top[181], bl_top[182], bl_top[183], bl_top[184], bl_top[185],
     bl_top[186], bl_top[187], bl_top[188], bl_top[189], bl_top[190],
     bl_top[191], bl_top[192], bl_top[193], bl_top[194], bl_top[195],
     bl_top[196], bl_top[197], bl_top[198], bl_top[199], bl_top[200],
     bl_top[201], bl_top[202], bl_top[203], bl_top[204], bl_top[205],
     bl_top[206], bl_top[207], bl_top[208], bl_top[209], bl_top[210],
     bl_top[211], bl_top[212], bl_top[213], bl_top[214], bl_top[215],
     bl_top[216], bl_top[217], bl_top[218], bl_top[219], bl_top[220],
     bl_top[221], bl_top[222], bl_top[223], bl_top[224], bl_top[225],
     bl_top[226], bl_top[227], bl_top[228], bl_top[229], bl_top[230],
     bl_top[231], bl_top[232], bl_top[233], bl_top[234], bl_top[235],
     bl_top[236], bl_top[237], bl_top[238], bl_top[239], bl_top[240],
     bl_top[241], bl_top[242], bl_top[243], bl_top[244], bl_top[245],
     bl_top[246], bl_top[247], bl_top[248], bl_top[249], bl_top[250],
     bl_top[251], bl_top[252], bl_top[253], bl_top[254], bl_top[255],
     bl_top[256], bl_top[257], bl_top[258], bl_top[259], bl_top[260],
     bl_top[261], bl_top[262], bl_top[263], bl_top[264], bl_top[265],
     bl_top[266], bl_top[267], bl_top[268], bl_top[269], bl_top[270],
     bl_top[271], bl_top[272], bl_top[273], bl_top[274], bl_top[275],
     bl_top[276], bl_top[277], bl_top[278], bl_top[279], bl_top[280],
     bl_top[281], bl_top[282], bl_top[283], bl_top[284], bl_top[285],
     bl_top[286], bl_top[287], bl_top[288], bl_top[289], bl_top[290],
     bl_top[291], bl_top[292], bl_top[293], bl_top[294], bl_top[295],
     bl_top[296], bl_top[297], bl_top[298], bl_top[299], bl_top[300],
     bl_top[301], bl_top[302], bl_top[303], bl_top[304], bl_top[305],
     bl_top[306], bl_top[307], bl_top[308], bl_top[309], bl_top[310],
     bl_top[311], bl_top[312], bl_top[313], bl_top[314], bl_top[315],
     bl_top[316], bl_top[317], bl_top[318], bl_top[319], bl_top[320],
     bl_top[321], bl_top[322], bl_top[323], bl_top[324], bl_top[325],
     bl_top[326], bl_top[327], bl_top[328], bl_top[329], bl_top[330],
     bl_top[331]}), .smc_wdic_clk(smc_wdis_dclk_bltld3),
     .smc_clk(cm_clk_bltld3), .cm_sdi_u(cm_sdi_u1d3[1:0]),
     .latch_reset(core_por_b_rowu1), .cm_sdo_u(cm_sdo_u1[1:0]),
     .data_muxsel1(data_muxsel1_bltld3),
     .data_muxsel(data_muxsel_bltld3), .cram_write(cram_write_bltld3),
     .cram_prec(cm_prec_bltld3),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltld3),
     .cram_pullup_b(cram_pullup_bltld3),
     .banksel(cm_banksel_bltld3[1]));

endmodule
// Library - xpmem, Cell - ml_buf_ice5_2, View - schematic
// LAST TIME SAVED: Jun 14 11:22:45 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_buf_ice5_2 ( o, in, sel );
output  o;

input  in, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_rowdrv2_last, View - schematic
// LAST TIME SAVED: Aug 18 15:57:39 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_rowdrv2_last ( pgate, reset, smc_rsr_out, vddctrl, wl,
     wl_rd_sup, wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write
     );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
ml_dff I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));

endmodule
// Library - xpmem, Cell - ml_rowdrvsup2, View - schematic
// LAST TIME SAVED: Jul 23 17:04:42 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_rowdrvsup2 ( wl_rd_sup, wl_rden_b );
inout  wl_rd_sup, wl_rden_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R2 ( .MINUS(net089), .PLUS(net095), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net0104), .PLUS(net0110), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net095), .PLUS(net0158), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(wl_rd_sup), .PLUS(net0104), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(net080), .PLUS(net092), .BULK(gnd_));
rppolywo_m  R3 ( .MINUS(net092), .PLUS(net089), .BULK(gnd_));
rppolywo_m  R9 ( .MINUS(net083), .PLUS(net086), .BULK(gnd_));
rppolywo_m  R8 ( .MINUS(net086), .PLUS(net080), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(net077), .PLUS(net083), .BULK(gnd_));
rppolywo_m  R13 ( .MINUS(net0108), .PLUS(net0107), .BULK(gnd_));
rppolywo_m  R11 ( .MINUS(net071), .PLUS(net077), .BULK(gnd_));
rppolywo_m  R12 ( .MINUS(net0108), .PLUS(net071), .BULK(gnd_));
rppolywo_m  R15 ( .MINUS(net0113), .PLUS(wl_rd_sup), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net0110), .PLUS(net045), .BULK(gnd_));
rppolywo_m  R14 ( .MINUS(net0107), .PLUS(net0113), .BULK(gnd_));
nch_hvt  MN16 ( .D(wl_rd_sup), .B(gnd_), .G(act_rd_b), .S(gnd_));
nch_hvt  MN14 ( .D(net0158), .B(gnd_), .G(act_rd), .S(gnd_));
pch_hvt  MP13 ( .D(wl_rden_b), .B(vdd_), .G(net059), .S(vdd_));
pch_hvt  MP15 ( .D(net045), .B(vdd_), .G(act_rd_b), .S(vdd_));
inv_hvt I217 ( .A(wl_rden_b), .Y(net0142));
inv_hvt I220 ( .A(net0142), .Y(act_rd_b));
inv_hvt I180 ( .A(act_rd_b), .Y(act_rd));
tielo I223 ( .tielo(net059));

endmodule
// Library - ice8chip, Cell - clk_mux_2to1_ice8p, View - schematic
// LAST TIME SAVED: Nov  5 16:41:18 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module clk_mux_2to1_ice8p ( clk, cbit, cbitb, min, prog );
output  clk;

input  cbit, cbitb, prog;

input [1:0]  min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I_inv0 ( .A(prog), .Y(net030));
nand2_lvt I_nand2_1 ( .A(st2), .Y(clkb), .B(net030));
inv_lvt I_inv2 ( .A(clkb), .Y(clk));
txgate_lvt I_txgate_hvt0 ( .in(min[0]), .out(st2), .pp(cbit),
     .nn(cbitb));
txgate_lvt I_txgate_hvt1 ( .in(min[1]), .out(st2), .pp(cbitb),
     .nn(cbit));

endmodule
// Library - xpmem, Cell - ml_rowdrv2, View - schematic
// LAST TIME SAVED: Jul 14 10:46:41 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_rowdrv2 ( pgate, reset, smc_rsr_out, vddctrl, wl, wl_rd_sup,
     wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
ml_dff I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile_last, View - schematic
// LAST TIME SAVED: Jan 24 11:25:01 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_rowdrv_tile_last ( pgate, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  reset;
output [15:0]  wl;
output [15:0]  vddctrl;
output [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



nor2_hvt I211 ( .A(smc_rsr_out[15]), .Y(net049), .B(smc_rsr_inc_out));
inv_hvt I215 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I216 ( .A(net041), .Y(por_rst_buf));
inv_hvt I217 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I391 ( .A(net049), .Y(smc_rsr_inc_last));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I213 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net079));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I214 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I212 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I190 ( .A(net079), .Y(smc_rsr_1st_out));
ml_rowdrv2_last Iml_rowdrv2_last ( .smc_rsr_inc(smc_rsr_inc_last),
     .smc_rsr_in(smc_rsr_out[14]), .rsr_rst(rsr_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_rst(cram_rst_buf),
     .smc_rsr_out(smc_rsr_out[15]), .reset(reset[15]), .wl(wl[15]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile, View - schematic
// LAST TIME SAVED: Jul 23 16:59:38 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_rowdrv_tile ( pgate, por_rst_out, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  por_rst_out, smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  vddctrl;
output [15:0]  pgate;
output [15:0]  wl;
output [15:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



inv_hvt I223 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I216 ( .A(cram_rst), .Y(net057));
inv_hvt I218 ( .A(net069), .Y(smc_write_buf));
inv_hvt I215 ( .A(cram_vddoff), .Y(net061));
inv_hvt I219 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I220 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I214 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I213 ( .A(smc_write), .Y(net069));
inv_hvt I221 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I212 ( .A(cram_wl_en), .Y(net055));
inv_hvt I217 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I190 ( .A(net037), .Y(smc_rsr_1st_out));
inv_hvt I211 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net037));
inv_hvt I210 ( .A(rsr_rst), .Y(net047));
inv_hvt I192 ( .A(por_rst), .Y(net041));
inv_hvt I222 ( .A(net041), .Y(por_rst_out));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I224 ( .A(net055), .Y(cram_wl_en_buf));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_15_ ( .reset(reset[15]), .wl(wl[15]),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[14]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[15]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_rowdrv_bank_ice1f, View - schematic
// LAST TIME SAVED: Mar  8 10:01:50 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_rowdrv_bank_ice1f ( jtag_rowtest_mode_b, last_rsr, pgate,
     reset, vddctrl, wl, banksel, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst,
     smc_rsr_inc, smc_write, trst_b );
output  jtag_rowtest_mode_b, last_rsr;

input  banksel, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst, smc_rsr_inc,
     smc_write, trst_b;

output [143:0]  reset;
output [143:0]  vddctrl;
output [143:0]  wl;
output [143:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  smc_rsr_1st_out_buf;

wire  [8:0]  smc_rsr_out;

wire  [7:0]  por_rst_out;

wire  [7:0]  smc_rsr_inc_out;

wire  [8:0]  smc_rsr_1st_out;



tielo I252 ( .tielo(net0130));
nand3_hvt I231 ( .Y(net186), .B(net190), .C(net190), .A(net190));
nand3_hvt I230 ( .Y(net190), .B(net195), .C(net195), .A(net195));
nand3_hvt I224 ( .B(net131), .Y(net195), .A(net131), .C(net131));
nand2_hvt I233 ( .A(smc_rsr_inc), .B(banksel), .Y(net181));
mux2_hvt I161 ( .in1(jtag_clk), .in0(net263), .out(net184),
     .sel(net256));
nor3_hvt I238 ( .B(por_rst), .Y(net248), .A(net208), .C(trst));
nor3_hvt I232 ( .C(rsr_rst), .A(jtag_rowtest_rst), .B(net0130),
     .Y(net213));
nor3_hvt I218 ( .B(net225), .Y(net215), .A(net225), .C(net225));
nor3_hvt I220 ( .B(net215), .Y(net219), .A(net215), .C(net215));
nor3_hvt I217 ( .C(net131), .A(net131), .B(net131), .Y(net225));
nor3_hvt I244 ( .B(por_rst), .Y(net227), .A(net276),
     .C(smc_rsr_1st_out_buf[0]));
nor2_hvt I239 ( .A(jtag_rowtest_rst), .B(net248), .Y(net208));
nor2_hvt I193 ( .A(por_rst), .B(rsr_set_1st), .Y(net252));
nor2_hvt I245 ( .A(rsr_set_1st), .B(net227), .Y(net276));
inv_hvt I247 ( .A(net256), .Y(jtag_rowtest_mode_b));
inv_hvt I241 ( .A(net208), .Y(net256));
inv_hvt I192 ( .A(net213), .Y(rsr_set_1st));
inv_hvt I234 ( .A(net181), .Y(net263));
inv_hvt I35 ( .A(net264), .Y(smc_rsr_1st_out_buf[0]));
inv_hvt I240 ( .A(trst_b), .Y(trst));
inv_hvt I210 ( .A(net268), .Y(last_rsr));
inv_hvt I391 ( .A(net252), .Y(rst_row_reg));
inv_hvt I36 ( .A(smc_rsr_1st_out[0]), .Y(net264));
inv_hvt I209 ( .A(smc_rsr_out[8]), .Y(net268));
inv_hvt I205 ( .A(net276), .Y(smc_rsr_in_1st));
tiehi I269 ( .tiehi(net162));
tiehi I249 ( .tiehi(net131));
tiehi I250 ( .tiehi(net132));
ml_buf_ice5_2 I227 ( .in(net131), .o(net134), .sel(net131));
ml_buf_ice5_2 I216 ( .in(net131), .o(net137), .sel(net131));
ml_buf_ice5_2 I198 ( .sel(banksel), .in(cram_wl_en),
     .o(cram_wl_en_buf));
ml_buf_ice5_2 I196 ( .sel(banksel), .in(cram_rst), .o(cram_rst_buf));
ml_buf_ice5_2 I199 ( .sel(net132), .in(por_rst), .o(por_rst_buf));
ml_buf_ice5_2 I197 ( .sel(banksel), .in(cram_vddoff),
     .o(cram_vddoff_buf));
ml_buf_ice5_2 I195 ( .sel(banksel), .in(cram_pgateoff),
     .o(cram_pgateoff_buf));
ml_buf_ice5_2 I201 ( .sel(banksel), .in(smc_write), .o(smc_write_buf));
ml_buf_ice5_2 I203 ( .sel(net184), .in(net184), .o(smc_rsr_inc_buf));
ml_buf_ice5_2 I213 ( .in(net162), .o(net161), .sel(net162));
ml_rowdrv_tile_last I_ml_rowdrv_tile_last (
     .smc_rsr_inc_out(smc_rsr_inc_out_last), .pgate(pgate[143:128]),
     .wl(wl[143:128]), .vddctrl(vddctrl[143:128]),
     .reset(reset[143:128]), .smc_rsr_1st_out(smc_rsr_1st_out[8]),
     .smcc_rsr_out(smc_rsr_out[8]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_buf), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[7]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf));
ml_rowdrv_tile I_ml_rowdrv_tile_7_ ( .por_rst_out(por_rst_out[7]),
     .smc_rsr_inc_out(smc_rsr_inc_out[7]),
     .smcc_rsr_out(smc_rsr_out[7]),
     .smc_rsr_1st_out(smc_rsr_1st_out[7]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out_last), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[6]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[127:112]), .vddctrl(vddctrl[127:112]),
     .reset(reset[127:112]), .pgate(pgate[127:112]));
ml_rowdrv_tile I_ml_rowdrv_tile_6_ ( .por_rst_out(por_rst_out[6]),
     .smc_rsr_inc_out(smc_rsr_inc_out[6]),
     .smcc_rsr_out(smc_rsr_out[6]),
     .smc_rsr_1st_out(smc_rsr_1st_out[6]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[7]), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[5]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[111:96]), .vddctrl(vddctrl[111:96]), .reset(reset[111:96]),
     .pgate(pgate[111:96]));
ml_rowdrv_tile I_ml_rowdrv_tile_5_ ( .por_rst_out(por_rst_out[5]),
     .smc_rsr_inc_out(smc_rsr_inc_out[5]),
     .smcc_rsr_out(smc_rsr_out[5]),
     .smc_rsr_1st_out(smc_rsr_1st_out[5]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[6]), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[4]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[95:80]), .vddctrl(vddctrl[95:80]), .reset(reset[95:80]),
     .pgate(pgate[95:80]));
ml_rowdrv_tile I_ml_rowdrv_tile_4_ ( .por_rst_out(por_rst_out[4]),
     .smc_rsr_inc_out(smc_rsr_inc_out[4]),
     .smcc_rsr_out(smc_rsr_out[4]),
     .smc_rsr_1st_out(smc_rsr_1st_out[4]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[5]), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[3]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[79:64]), .vddctrl(vddctrl[79:64]), .reset(reset[79:64]),
     .pgate(pgate[79:64]));
ml_rowdrv_tile I_ml_rowdrv_tile_3_ ( .por_rst_out(por_rst_out[3]),
     .smc_rsr_inc_out(smc_rsr_inc_out[3]),
     .smcc_rsr_out(smc_rsr_out[3]),
     .smc_rsr_1st_out(smc_rsr_1st_out[3]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[4]), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[2]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[63:48]), .vddctrl(vddctrl[63:48]), .reset(reset[63:48]),
     .pgate(pgate[63:48]));
ml_rowdrv_tile I_ml_rowdrv_tile_2_ ( .por_rst_out(por_rst_out[2]),
     .smc_rsr_inc_out(smc_rsr_inc_out[2]),
     .smcc_rsr_out(smc_rsr_out[2]),
     .smc_rsr_1st_out(smc_rsr_1st_out[2]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[3]), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[1]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[47:32]), .vddctrl(vddctrl[47:32]), .reset(reset[47:32]),
     .pgate(pgate[47:32]));
ml_rowdrv_tile I_ml_rowdrv_tile_1_ ( .por_rst_out(por_rst_out[1]),
     .smc_rsr_inc_out(smc_rsr_inc_out[1]),
     .smcc_rsr_out(smc_rsr_out[1]),
     .smc_rsr_1st_out(smc_rsr_1st_out[1]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[2]), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[0]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[31:16]), .vddctrl(vddctrl[31:16]), .reset(reset[31:16]),
     .pgate(pgate[31:16]));
ml_rowdrv_tile I_ml_rowdrv_tile_0_ ( .por_rst_out(por_rst_out[0]),
     .smc_rsr_inc_out(smc_rsr_inc_out[0]),
     .smcc_rsr_out(smc_rsr_out[0]),
     .smc_rsr_1st_out(smc_rsr_1st_out[0]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[1]), .smc_rsr_in(smc_rsr_in_1st),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[15:0]), .vddctrl(vddctrl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]));

endmodule
// Library - ice8chip, Cell - sg_dffbuf_modified, View - schematic
// LAST TIME SAVED: Aug 19 09:09:59 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module sg_dffbuf_modified ( dffout, clk, d, r );
output  dffout;

input  clk, d, r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff I0 ( .R(r), .D(d), .CLK(clk), .QN(net9), .Q(net10));
sg_bufx10_ice8p I5 ( .in(net10), .out(dffout));

endmodule
// Library - ice1chip, Cell - CHIP_route_lft_ice1f, View - schematic
// LAST TIME SAVED: Apr 22 10:30:29 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module CHIP_route_lft_ice1f ( cm_banksel_bltld3_1_, cm_clk_bltld3,
     cm_sdi_u1d3, cm_sdo_u1d1, core_por_b_rowu1, cram_prec_bltld3,
     cram_pullup_bltld3, cram_write_bltld3, data_muxsel1_bltld3,
     data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     last_rsr, pgate_l, reset_l, smc_wdis_dclk_bltld3,
     smc_write_bltld3, vdd_cntl_l, wl_l, cm_banksel_blbld1,
     cm_banksel_blbld, cm_clk_blbld, cm_sdi_u1d, cm_sdo_u1,
     core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0 );
output  cm_banksel_bltld3_1_, cm_clk_bltld3, core_por_b_rowu1,
     cram_prec_bltld3, cram_pullup_bltld3, cram_write_bltld3,
     data_muxsel1_bltld3, data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     smc_wdis_dclk_bltld3, smc_write_bltld3;

input  cm_clk_blbld, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;

output [1:0]  cm_sdo_u1d1;
output [287:0]  reset_l;
output [287:0]  wl_l;
output [1:0]  cm_sdi_u1d3;
output [287:0]  vdd_cntl_l;
output [1:0]  last_rsr;
output [287:0]  pgate_l;

input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdi_u1d;
input [1:1]  cm_banksel_blbld;
input [0:0]  cm_banksel_blbld1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdi_u1d0;

wire  [1:0]  net299;

wire  [1:1]  cm_banksel_bltld;

wire  [1:0]  cm_sdo_u1d0;

wire  [1:0]  dff_out;



ml_rowdrv_bank_ice1f I_ml_rowdrv_bank1f_bot ( .wl(wl_l[143:0]),
     .pgate(pgate_l[143:0]), .reset(reset_l[143:0]),
     .vddctrl(vdd_cntl_l[143:0]), .trst_b(j_rst_bl0),
     .smc_write(smc_writel0),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu0_b),
     .last_rsr(last_rsr[0]), .banksel(cm_banksel_blbld1[0]),
     .cram_pgateoff(cram_pgateoffl0), .cram_rst(cram_rstl0),
     .cram_vddoff(cram_vddoffl0), .cram_wl_en(cram_wl_enl0),
     .jtag_clk(tck_padl0), .jtag_rowtest_rst(row_testl1),
     .por_rst(core_por_bbl0), .rsr_rst(smc_rsr_rstl0),
     .smc_rsr_inc(smc_row_incl0));
ml_rowdrv_bank_ice1f I_ml_rowdrv_bank1f_top ( .wl({wl_l[144],
     wl_l[145], wl_l[146], wl_l[147], wl_l[148], wl_l[149], wl_l[150],
     wl_l[151], wl_l[152], wl_l[153], wl_l[154], wl_l[155], wl_l[156],
     wl_l[157], wl_l[158], wl_l[159], wl_l[160], wl_l[161], wl_l[162],
     wl_l[163], wl_l[164], wl_l[165], wl_l[166], wl_l[167], wl_l[168],
     wl_l[169], wl_l[170], wl_l[171], wl_l[172], wl_l[173], wl_l[174],
     wl_l[175], wl_l[176], wl_l[177], wl_l[178], wl_l[179], wl_l[180],
     wl_l[181], wl_l[182], wl_l[183], wl_l[184], wl_l[185], wl_l[186],
     wl_l[187], wl_l[188], wl_l[189], wl_l[190], wl_l[191], wl_l[192],
     wl_l[193], wl_l[194], wl_l[195], wl_l[196], wl_l[197], wl_l[198],
     wl_l[199], wl_l[200], wl_l[201], wl_l[202], wl_l[203], wl_l[204],
     wl_l[205], wl_l[206], wl_l[207], wl_l[208], wl_l[209], wl_l[210],
     wl_l[211], wl_l[212], wl_l[213], wl_l[214], wl_l[215], wl_l[216],
     wl_l[217], wl_l[218], wl_l[219], wl_l[220], wl_l[221], wl_l[222],
     wl_l[223], wl_l[224], wl_l[225], wl_l[226], wl_l[227], wl_l[228],
     wl_l[229], wl_l[230], wl_l[231], wl_l[232], wl_l[233], wl_l[234],
     wl_l[235], wl_l[236], wl_l[237], wl_l[238], wl_l[239], wl_l[240],
     wl_l[241], wl_l[242], wl_l[243], wl_l[244], wl_l[245], wl_l[246],
     wl_l[247], wl_l[248], wl_l[249], wl_l[250], wl_l[251], wl_l[252],
     wl_l[253], wl_l[254], wl_l[255], wl_l[256], wl_l[257], wl_l[258],
     wl_l[259], wl_l[260], wl_l[261], wl_l[262], wl_l[263], wl_l[264],
     wl_l[265], wl_l[266], wl_l[267], wl_l[268], wl_l[269], wl_l[270],
     wl_l[271], wl_l[272], wl_l[273], wl_l[274], wl_l[275], wl_l[276],
     wl_l[277], wl_l[278], wl_l[279], wl_l[280], wl_l[281], wl_l[282],
     wl_l[283], wl_l[284], wl_l[285], wl_l[286], wl_l[287]}),
     .pgate({pgate_l[144], pgate_l[145], pgate_l[146], pgate_l[147],
     pgate_l[148], pgate_l[149], pgate_l[150], pgate_l[151],
     pgate_l[152], pgate_l[153], pgate_l[154], pgate_l[155],
     pgate_l[156], pgate_l[157], pgate_l[158], pgate_l[159],
     pgate_l[160], pgate_l[161], pgate_l[162], pgate_l[163],
     pgate_l[164], pgate_l[165], pgate_l[166], pgate_l[167],
     pgate_l[168], pgate_l[169], pgate_l[170], pgate_l[171],
     pgate_l[172], pgate_l[173], pgate_l[174], pgate_l[175],
     pgate_l[176], pgate_l[177], pgate_l[178], pgate_l[179],
     pgate_l[180], pgate_l[181], pgate_l[182], pgate_l[183],
     pgate_l[184], pgate_l[185], pgate_l[186], pgate_l[187],
     pgate_l[188], pgate_l[189], pgate_l[190], pgate_l[191],
     pgate_l[192], pgate_l[193], pgate_l[194], pgate_l[195],
     pgate_l[196], pgate_l[197], pgate_l[198], pgate_l[199],
     pgate_l[200], pgate_l[201], pgate_l[202], pgate_l[203],
     pgate_l[204], pgate_l[205], pgate_l[206], pgate_l[207],
     pgate_l[208], pgate_l[209], pgate_l[210], pgate_l[211],
     pgate_l[212], pgate_l[213], pgate_l[214], pgate_l[215],
     pgate_l[216], pgate_l[217], pgate_l[218], pgate_l[219],
     pgate_l[220], pgate_l[221], pgate_l[222], pgate_l[223],
     pgate_l[224], pgate_l[225], pgate_l[226], pgate_l[227],
     pgate_l[228], pgate_l[229], pgate_l[230], pgate_l[231],
     pgate_l[232], pgate_l[233], pgate_l[234], pgate_l[235],
     pgate_l[236], pgate_l[237], pgate_l[238], pgate_l[239],
     pgate_l[240], pgate_l[241], pgate_l[242], pgate_l[243],
     pgate_l[244], pgate_l[245], pgate_l[246], pgate_l[247],
     pgate_l[248], pgate_l[249], pgate_l[250], pgate_l[251],
     pgate_l[252], pgate_l[253], pgate_l[254], pgate_l[255],
     pgate_l[256], pgate_l[257], pgate_l[258], pgate_l[259],
     pgate_l[260], pgate_l[261], pgate_l[262], pgate_l[263],
     pgate_l[264], pgate_l[265], pgate_l[266], pgate_l[267],
     pgate_l[268], pgate_l[269], pgate_l[270], pgate_l[271],
     pgate_l[272], pgate_l[273], pgate_l[274], pgate_l[275],
     pgate_l[276], pgate_l[277], pgate_l[278], pgate_l[279],
     pgate_l[280], pgate_l[281], pgate_l[282], pgate_l[283],
     pgate_l[284], pgate_l[285], pgate_l[286], pgate_l[287]}),
     .reset({reset_l[144], reset_l[145], reset_l[146], reset_l[147],
     reset_l[148], reset_l[149], reset_l[150], reset_l[151],
     reset_l[152], reset_l[153], reset_l[154], reset_l[155],
     reset_l[156], reset_l[157], reset_l[158], reset_l[159],
     reset_l[160], reset_l[161], reset_l[162], reset_l[163],
     reset_l[164], reset_l[165], reset_l[166], reset_l[167],
     reset_l[168], reset_l[169], reset_l[170], reset_l[171],
     reset_l[172], reset_l[173], reset_l[174], reset_l[175],
     reset_l[176], reset_l[177], reset_l[178], reset_l[179],
     reset_l[180], reset_l[181], reset_l[182], reset_l[183],
     reset_l[184], reset_l[185], reset_l[186], reset_l[187],
     reset_l[188], reset_l[189], reset_l[190], reset_l[191],
     reset_l[192], reset_l[193], reset_l[194], reset_l[195],
     reset_l[196], reset_l[197], reset_l[198], reset_l[199],
     reset_l[200], reset_l[201], reset_l[202], reset_l[203],
     reset_l[204], reset_l[205], reset_l[206], reset_l[207],
     reset_l[208], reset_l[209], reset_l[210], reset_l[211],
     reset_l[212], reset_l[213], reset_l[214], reset_l[215],
     reset_l[216], reset_l[217], reset_l[218], reset_l[219],
     reset_l[220], reset_l[221], reset_l[222], reset_l[223],
     reset_l[224], reset_l[225], reset_l[226], reset_l[227],
     reset_l[228], reset_l[229], reset_l[230], reset_l[231],
     reset_l[232], reset_l[233], reset_l[234], reset_l[235],
     reset_l[236], reset_l[237], reset_l[238], reset_l[239],
     reset_l[240], reset_l[241], reset_l[242], reset_l[243],
     reset_l[244], reset_l[245], reset_l[246], reset_l[247],
     reset_l[248], reset_l[249], reset_l[250], reset_l[251],
     reset_l[252], reset_l[253], reset_l[254], reset_l[255],
     reset_l[256], reset_l[257], reset_l[258], reset_l[259],
     reset_l[260], reset_l[261], reset_l[262], reset_l[263],
     reset_l[264], reset_l[265], reset_l[266], reset_l[267],
     reset_l[268], reset_l[269], reset_l[270], reset_l[271],
     reset_l[272], reset_l[273], reset_l[274], reset_l[275],
     reset_l[276], reset_l[277], reset_l[278], reset_l[279],
     reset_l[280], reset_l[281], reset_l[282], reset_l[283],
     reset_l[284], reset_l[285], reset_l[286], reset_l[287]}),
     .vddctrl({vdd_cntl_l[144], vdd_cntl_l[145], vdd_cntl_l[146],
     vdd_cntl_l[147], vdd_cntl_l[148], vdd_cntl_l[149],
     vdd_cntl_l[150], vdd_cntl_l[151], vdd_cntl_l[152],
     vdd_cntl_l[153], vdd_cntl_l[154], vdd_cntl_l[155],
     vdd_cntl_l[156], vdd_cntl_l[157], vdd_cntl_l[158],
     vdd_cntl_l[159], vdd_cntl_l[160], vdd_cntl_l[161],
     vdd_cntl_l[162], vdd_cntl_l[163], vdd_cntl_l[164],
     vdd_cntl_l[165], vdd_cntl_l[166], vdd_cntl_l[167],
     vdd_cntl_l[168], vdd_cntl_l[169], vdd_cntl_l[170],
     vdd_cntl_l[171], vdd_cntl_l[172], vdd_cntl_l[173],
     vdd_cntl_l[174], vdd_cntl_l[175], vdd_cntl_l[176],
     vdd_cntl_l[177], vdd_cntl_l[178], vdd_cntl_l[179],
     vdd_cntl_l[180], vdd_cntl_l[181], vdd_cntl_l[182],
     vdd_cntl_l[183], vdd_cntl_l[184], vdd_cntl_l[185],
     vdd_cntl_l[186], vdd_cntl_l[187], vdd_cntl_l[188],
     vdd_cntl_l[189], vdd_cntl_l[190], vdd_cntl_l[191],
     vdd_cntl_l[192], vdd_cntl_l[193], vdd_cntl_l[194],
     vdd_cntl_l[195], vdd_cntl_l[196], vdd_cntl_l[197],
     vdd_cntl_l[198], vdd_cntl_l[199], vdd_cntl_l[200],
     vdd_cntl_l[201], vdd_cntl_l[202], vdd_cntl_l[203],
     vdd_cntl_l[204], vdd_cntl_l[205], vdd_cntl_l[206],
     vdd_cntl_l[207], vdd_cntl_l[208], vdd_cntl_l[209],
     vdd_cntl_l[210], vdd_cntl_l[211], vdd_cntl_l[212],
     vdd_cntl_l[213], vdd_cntl_l[214], vdd_cntl_l[215],
     vdd_cntl_l[216], vdd_cntl_l[217], vdd_cntl_l[218],
     vdd_cntl_l[219], vdd_cntl_l[220], vdd_cntl_l[221],
     vdd_cntl_l[222], vdd_cntl_l[223], vdd_cntl_l[224],
     vdd_cntl_l[225], vdd_cntl_l[226], vdd_cntl_l[227],
     vdd_cntl_l[228], vdd_cntl_l[229], vdd_cntl_l[230],
     vdd_cntl_l[231], vdd_cntl_l[232], vdd_cntl_l[233],
     vdd_cntl_l[234], vdd_cntl_l[235], vdd_cntl_l[236],
     vdd_cntl_l[237], vdd_cntl_l[238], vdd_cntl_l[239],
     vdd_cntl_l[240], vdd_cntl_l[241], vdd_cntl_l[242],
     vdd_cntl_l[243], vdd_cntl_l[244], vdd_cntl_l[245],
     vdd_cntl_l[246], vdd_cntl_l[247], vdd_cntl_l[248],
     vdd_cntl_l[249], vdd_cntl_l[250], vdd_cntl_l[251],
     vdd_cntl_l[252], vdd_cntl_l[253], vdd_cntl_l[254],
     vdd_cntl_l[255], vdd_cntl_l[256], vdd_cntl_l[257],
     vdd_cntl_l[258], vdd_cntl_l[259], vdd_cntl_l[260],
     vdd_cntl_l[261], vdd_cntl_l[262], vdd_cntl_l[263],
     vdd_cntl_l[264], vdd_cntl_l[265], vdd_cntl_l[266],
     vdd_cntl_l[267], vdd_cntl_l[268], vdd_cntl_l[269],
     vdd_cntl_l[270], vdd_cntl_l[271], vdd_cntl_l[272],
     vdd_cntl_l[273], vdd_cntl_l[274], vdd_cntl_l[275],
     vdd_cntl_l[276], vdd_cntl_l[277], vdd_cntl_l[278],
     vdd_cntl_l[279], vdd_cntl_l[280], vdd_cntl_l[281],
     vdd_cntl_l[282], vdd_cntl_l[283], vdd_cntl_l[284],
     vdd_cntl_l[285], vdd_cntl_l[286], vdd_cntl_l[287]}),
     .smc_write(smc_write_bltld3), .smc_rsr_inc(net303),
     .rsr_rst(net289), .por_rst(core_por_b_rowu1),
     .jtag_rowtest_rst(net345), .jtag_clk(net305), .cram_wl_en(net273),
     .cram_vddoff(net335), .cram_rst(net319), .cram_pgateoff(net295),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu1_b),
     .last_rsr(last_rsr[1]), .banksel(net231), .trst_b(net311));
tielo I74 ( .tielo(net219));
sg_bufx10_ice8p I28 ( .in(smc_writel0), .out(net221));
sg_bufx10_ice8p I35 ( .in(net291), .out(net223));
sg_bufx10_ice8p I45 ( .in(row_testl1), .out(net225));
sg_bufx10_ice8p I44 ( .in(net225), .out(net227));
sg_bufx10_ice8p I2 ( .in(cram_write_bltld), .out(net229));
sg_bufx10_ice8p I67 ( .in(cm_banksel_bltld[1]), .out(net231));
sg_bufx10_ice8p I39 ( .in(net237), .out(net233));
sg_bufx10_ice8p I4 ( .in(data_muxsel1_blbld),
     .out(data_muxsel1_bltld));
sg_bufx10_ice8p I40 ( .in(cram_wl_enl0), .out(net237));
sg_bufx10_ice8p I37 ( .in(cram_vddoffl0), .out(net239));
sg_bufx10_ice8p I22 ( .in(core_por_bbl0), .out(net241));
sg_bufx10_ice8p I5 ( .in(data_muxsel1_bltld), .out(net243));
sg_bufx10_ice8p I527 ( .in(net327), .out(en_8bconfig_b_bltld3));
sg_bufx10_ice8p I523 ( .in(net283), .out(data_muxsel_bltld3));
sg_bufx10_ice8p I524 ( .in(net243), .out(data_muxsel1_bltld3));
sg_bufx10_ice8p I526 ( .in(net343), .out(cram_prec_bltld3));
sg_bufx10_ice8p I33 ( .in(cram_rstl0), .out(net253));
sg_bufx10_ice8p I70_1_ ( .in(cm_sdo_u1[1]), .out(cm_sdo_u1d0[1]));
sg_bufx10_ice8p I70_0_ ( .in(cm_sdo_u1[0]), .out(cm_sdo_u1d0[0]));
sg_bufx10_ice8p I528 ( .in(net337), .out(smc_wdis_dclk_bltld3));
sg_bufx10_ice8p I18 ( .in(smc_rsr_rstl0), .out(net259));
sg_bufx10_ice8p I529 ( .in(net293), .out(cram_pullup_bltld3));
sg_bufx10_ice8p I3 ( .in(cram_write_blbld), .out(cram_write_bltld));
sg_bufx10_ice8p I532 ( .in(net363), .out(cm_clk_bltld3));
sg_bufx10_ice8p I79 ( .in(cm_clk_blbld), .out(cm_clk_bltld));
sg_bufx10_ice8p I8 ( .in(cram_pullup_blbld), .out(cram_pullup_bltld));
sg_bufx10_ice8p I7 ( .in(data_muxsel_blbld), .out(data_muxsel_bltld));
sg_bufx10_ice8p I554 ( .in(net233), .out(net273));
sg_bufx10_ice8p I27 ( .in(net221), .out(net275));
sg_bufx10_ice8p I25 ( .in(smc_row_incl0), .out(net277));
sg_bufx10_ice8p I47 ( .in(net357), .out(net279));
sg_bufx10_ice8p I68_1_ ( .in(cm_sdi_u1d[1]), .out(cm_sdi_u1d0[1]));
sg_bufx10_ice8p I68_0_ ( .in(cm_sdi_u1d[0]), .out(cm_sdi_u1d0[0]));
sg_bufx10_ice8p I6 ( .in(data_muxsel_bltld), .out(net283));
sg_bufx10_ice8p I38 ( .in(net239), .out(net285));
sg_bufx10_ice8p I19 ( .in(net259), .out(net287));
sg_bufx10_ice8p I546 ( .in(net287), .out(net289));
sg_bufx10_ice8p I36 ( .in(cram_pgateoffl0), .out(net291));
sg_bufx10_ice8p I9 ( .in(cram_pullup_bltld), .out(net293));
sg_bufx10_ice8p I547 ( .in(net223), .out(net295));
sg_bufx10_ice8p I552 ( .in(net275), .out(smc_write_bltld3));
sg_bufx10_ice8p I69_1_ ( .in(cm_sdi_u1d0[1]), .out(net299[0]));
sg_bufx10_ice8p I69_0_ ( .in(cm_sdi_u1d0[0]), .out(net299[1]));
sg_bufx10_ice8p I549 ( .in(net349), .out(net303));
sg_bufx10_ice8p I544 ( .in(net279), .out(net305));
sg_bufx10_ice8p I530_1_ ( .in(net299[0]), .out(cm_sdi_u1d3[1]));
sg_bufx10_ice8p I530_0_ ( .in(net299[1]), .out(cm_sdi_u1d3[0]));
sg_bufx10_ice8p I545 ( .in(net353), .out(net311));
sg_bufx10_ice8p I531 ( .in(net231), .out(cm_banksel_bltld3_1_));
sg_bufx10_ice8p I551 ( .in(net331), .out(net319));
sg_bufx10_ice8p I553 ( .in(net355), .out(core_por_b_rowu1));
sg_bufx10_ice8p I81 ( .in(cm_clk_bltld), .out(net363));
sg_bufx10_ice8p I15 ( .in(en_8bconfig_b_blbld),
     .out(en_8bconfig_b_bltld));
sg_bufx10_ice8p I14 ( .in(en_8bconfig_b_bltld), .out(net327));
sg_bufx10_ice8p I0 ( .in(cram_prec_blbld), .out(cram_prec_bltld));
sg_bufx10_ice8p I34 ( .in(net253), .out(net331));
sg_bufx10_ice8p I49 ( .in(j_rst_bl0), .out(net333));
sg_bufx10_ice8p I550 ( .in(net285), .out(net335));
sg_bufx10_ice8p I13 ( .in(smc_wdis_dclk_bltld), .out(net337));
sg_bufx10_ice8p I66 ( .in(cm_banksel_blbld[1]),
     .out(cm_banksel_bltld[1]));
sg_bufx10_ice8p I80_1_ ( .in(dff_out[1]), .out(cm_sdo_u1d1[1]));
sg_bufx10_ice8p I80_0_ ( .in(dff_out[0]), .out(cm_sdo_u1d1[0]));
sg_bufx10_ice8p I1 ( .in(cram_prec_bltld), .out(net343));
sg_bufx10_ice8p I548 ( .in(net227), .out(net345));
sg_bufx10_ice8p I525 ( .in(net229), .out(cram_write_bltld3));
sg_bufx10_ice8p I26 ( .in(net277), .out(net349));
sg_bufx10_ice8p I12 ( .in(smc_wdis_dclk_blbld),
     .out(smc_wdis_dclk_bltld));
sg_bufx10_ice8p I48 ( .in(net333), .out(net353));
sg_bufx10_ice8p I21 ( .in(net241), .out(net355));
sg_bufx10_ice8p I46 ( .in(tck_padl0), .out(net357));
sg_dffbuf_modified I73_1_ ( .d(cm_sdo_u1d0[1]), .clk(net363),
     .dffout(dff_out[1]), .r(net219));
sg_dffbuf_modified I73_0_ ( .d(cm_sdo_u1d0[0]), .clk(net363),
     .dffout(dff_out[0]), .r(net219));
sg_dffbuf_modified I77 ( .d(last_rsr[0]), .clk(net363),
     .dffout(last_rsr0), .r(net219));

endmodule
// Library - leafcell, Cell - creset_filter, View - schematic
// LAST TIME SAVED: Sep 30 15:04:05 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module creset_filter ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I11 ( .in(net042), .out(out));
nch_hvt  M0 ( .D(net13), .B(gnd_), .G(in), .S(gnd_));
nch_hvt  MN31 ( .D(net17), .B(gnd_), .G(net9), .S(gnd_));
rppolywo_m  R0 ( .MINUS(net17), .PLUS(pbias), .BULK(gnd_));
pch_hvt  M3 ( .D(net13), .B(vdd_), .G(net042), .S(vdd_));
pch_hvt  M2 ( .D(net13), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  M1 ( .D(vdd_), .B(vdd_), .G(net13), .S(vdd_));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(net9), .S(vdd_));
inv_hvt I6 ( .A(net13), .Y(net042));
inv_hvt I4 ( .A(in), .Y(net9));

endmodule
// Library - ice8chip, Cell - bram_bufferx16_ice8p, View - schematic
// LAST TIME SAVED: Aug  6 14:53:07 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module bram_bufferx16_ice8p ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I5 ( .A(net07), .Y(net09));
inv_hvt I2 ( .A(in), .Y(net07));
inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(net09), .Y(net6));

endmodule
// Library - ice8chip, Cell - eh_io_pup_2_new_ice8p, View - schematic
// LAST TIME SAVED: Aug 25 11:50:10 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module eh_io_pup_2_new_ice8p ( por_b, core_por_b, vdd_io );
output  por_b;

input  core_por_b, vdd_io;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M8 ( .D(net104), .B(gnd_), .G(v_in), .S(net104));
nch_lvt  M23 ( .D(net104), .B(gnd_), .G(v_in), .S(net0196));
sg_bufx10_ice8p I_clkbuf ( .in(net84), .out(por_b));
nch_na25  M27 ( .D(net0224), .B(gnd_), .G(net0224), .S(net0132));
nch_na25  M24 ( .D(net0132), .B(gnd_), .G(net0132), .S(net0220));
nch_na25  M25 ( .D(net0220), .B(gnd_), .G(net0220), .S(net0216));
nch_na25  M9 ( .D(net158), .B(gnd_), .G(net158), .S(net154));
nch_na25  M13 ( .D(net150), .B(gnd_), .G(net150), .S(net162));
nch_na25  M16 ( .D(v_in), .B(gnd_), .G(net147), .S(net0195));
nch_na25  M20 ( .D(net162), .B(gnd_), .G(net162), .S(net0112));
nch_na25  M12 ( .D(net154), .B(gnd_), .G(net154), .S(net150));
nch_na25  M26 ( .D(net0216), .B(gnd_), .G(net0216), .S(gnd_));
nch_na25  M21 ( .D(net0112), .B(gnd_), .G(net0112), .S(gnd_));
rppolywo_m  R66 ( .MINUS(gnd_), .PLUS(net145), .BULK(gnd_));
nch_25  MN6 ( .D(net0195), .B(gnd_), .G(net145), .S(gnd_));
nch_25  M10 ( .D(net0195), .B(gnd_), .G(net147), .S(net158));
nch_25  M14 ( .D(v_in), .B(gnd_), .G(net147), .S(net0224));
nch_hvt  M22 ( .D(net104), .B(gnd_), .G(v_in), .S(net104));
nch_hvt  MN1 ( .D(net0196), .B(gnd_), .G(core_por_b), .S(gnd_));
nch_hvt  M2 ( .D(net84), .B(gnd_), .G(net104), .S(gnd_));
pch_hvt  M17 ( .D(net104), .B(vdd_), .G(v_in), .S(vdd_));
pch_hvt  MP8 ( .D(net104), .B(vdd_), .G(core_por_b), .S(vdd_));
pch_hvt  M0 ( .D(net84), .B(vdd_), .G(net104), .S(vdd_));
pch_25  M1 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
pch_25  M5 ( .D(net0195), .B(vdd_io), .G(net0195), .S(vdd_io));
pch_25  M3 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
pch_25  M7 ( .D(net0195), .B(vdd_io), .G(net145), .S(net0195));
pch_25  M6 ( .D(net0195), .B(vdd_io), .G(net0195), .S(vdd_io));
pch_25  M4 ( .D(net0195), .B(vdd_io), .G(net0195), .S(vdd_io));
vdd_tiehigh I96 ( .vdd_tieh(net147));

endmodule
// Library - ice8chip, Cell - eh_core_pup_2, View - schematic
// LAST TIME SAVED: Sep  7 10:17:18 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module eh_core_pup_2 ( por_b );
output  por_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I7 ( .A(out_1), .Y(out_2));
inv_hvt I9 ( .A(out_2), .Y(out_3));
inv_hvt I11 ( .A(out_3), .Y(por_b));
nch_hvt  M3 ( .D(gnd_), .B(gnd_), .G(out_2), .S(gnd_));
nch_hvt  M4 ( .D(gnd_), .B(gnd_), .G(net148), .S(gnd_));
nch_hvt  M0 ( .D(out_1), .B(gnd_), .G(net148), .S(gnd_));
nch_hvt  M5 ( .D(gnd_), .B(gnd_), .G(net148), .S(gnd_));
nch_hvt  M1 ( .D(out_1), .B(gnd_), .G(out_2), .S(gnd_));
rppolywo  R10 ( .MINUS(net130), .PLUS(net109));
rppolywo  R12 ( .MINUS(net154), .PLUS(net157));
rppolywo  R6 ( .MINUS(out_1), .PLUS(net124));
rppolywo  R9 ( .MINUS(net118), .PLUS(net130));
rppolywo  R15 ( .MINUS(net166), .PLUS(div_1));
rppolywo  R13 ( .MINUS(net157), .PLUS(net145));
rppolywo  R1 ( .MINUS(net068), .PLUS(net048));
rppolywo  R2 ( .MINUS(net067), .PLUS(net068));
rppolywo  R4 ( .MINUS(net142), .PLUS(net148));
rppolywo  R5 ( .MINUS(div_1), .PLUS(net142));
rppolywo  R41 ( .MINUS(net039), .PLUS(net042));
rppolywo  R40 ( .MINUS(net042), .PLUS(vdd_));
rppolywo  R11 ( .MINUS(net109), .PLUS(net154));
rppolywo  R0 ( .MINUS(net048), .PLUS(net039));
rppolywo  R8 ( .MINUS(net127), .PLUS(net118));
rppolywo  R14 ( .MINUS(net145), .PLUS(net166));
rppolywo  R3 ( .MINUS(net148), .PLUS(net067));
rppolywo  R7 ( .MINUS(net124), .PLUS(net127));

endmodule
// Library - ice8chip, Cell - clk_mux2to1_ice8p, View - schematic
// LAST TIME SAVED: Nov  9 10:58:23 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module clk_mux2to1_ice8p ( gnet, bl, min0, min1, min2, min3, pgate_l,
     pgate_r, prog, reset_l, reset_r, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r );


input  prog;

output [3:0]  gnet;

inout [3:0]  bl;

input [1:0]  min2;
input [1:0]  pgate_l;
input [1:0]  reset_l;
input [1:0]  min0;
input [1:0]  reset_r;
input [1:0]  min1;
input [1:0]  min3;
input [1:0]  vdd_cntl_r;
input [1:0]  wl_l;
input [1:0]  vdd_cntl_l;
input [1:0]  pgate_r;
input [1:0]  wl_r;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [7:0]  cbitb;

wire  [7:0]  cbit;

wire  [1:0]  l_vdd;



clk_mux_2to1_ice8p I_clkmux3 ( .prog(prog), .cbit(cbit[3]),
     .cbitb(cbitb[3]), .min(min3[1:0]), .clk(gnet[3]));
clk_mux_2to1_ice8p I_clkmux1 ( .prog(prog), .cbit(cbit[1]),
     .cbitb(cbitb[1]), .min(min1[1:0]), .clk(gnet[1]));
clk_mux_2to1_ice8p I_clkmux2 ( .prog(prog), .cbit(cbit[2]),
     .cbitb(cbitb[2]), .min(min2[1:0]), .clk(gnet[2]));
clk_mux_2to1_ice8p I_clkmux0 ( .prog(prog), .cbit(cbit[0]),
     .cbitb(cbitb[0]), .min(min0[1:0]), .clk(gnet[0]));
pch_hvt  I_pch_hvt_l_1_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(l_vdd[0]));
pch_hvt  I_pch_hvt_l_0_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(l_vdd[1]));
pch_hvt  M0_1_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_r[1]), .S(r_vdd[1]));
pch_hvt  M0_0_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl_r[0]), .S(r_vdd[0]));
cram2x2 I_cram2x2_lft ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset_l[1:0]), .q(cbit[3:0]), .wl(wl_l[1:0]),
     .r_vdd({l_vdd[0], l_vdd[1]}), .pgate(pgate_l[1:0]));
cram2x2 I_cram2x2_rgt ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset_r[1:0]), .q(cbit[7:4]), .wl(wl_r[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate_r[1:0]));

endmodule
// Library - ice8chip, Cell - SMC_CORE_POR_right_ice8p, View -
//schematic
// LAST TIME SAVED: Sep 29 09:25:02 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module SMC_CORE_POR_right_ice8p ( core_por_b0, core_por_bb, smc_por_b,
     creset_b, smc_core_por_bottom1, smc_core_por_bottom2,
     vddio_rightbank );
output  core_por_b0, core_por_bb, smc_por_b;

input  creset_b, smc_core_por_bottom1, smc_core_por_bottom2,
     vddio_rightbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



sg_bufx10_ice8p I500 ( .in(net032), .out(core_por_bb));
eh_io_pup_2_new_ice8p Ieh_io_pup_2_new_ice8p ( .core_por_b(net026),
     .vdd_io(vddio_rightbank), .por_b(net3));
eh_core_pup_2 Ieh_core_pup_2 ( .por_b(net026));
nand2_hvt I6 ( .A(net026), .Y(net021), .B(creset_b));
inv_hvt I11 ( .A(net04), .Y(smc_por_b));
inv_hvt I701 ( .A(core_por_b0), .Y(net032));
inv_hvt I7 ( .A(net021), .Y(core_por_b0));
nand4_hvt I2 ( .D(core_por_b0), .C(smc_core_por_bottom2), .A(net3),
     .Y(net04), .B(smc_core_por_bottom1));

endmodule
// Library - ice8chip, Cell - smc_and_jtag_ice8p, View - schematic
// LAST TIME SAVED: Sep 30 15:13:23 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module smc_and_jtag_ice8p ( bm_bank_sdi, bm_banksel, bm_clk, bm_init,
     bm_rcapmux_en, bm_sa, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_banksel, cm_clk, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2, cm_sdi_u3, data_muxsel, data_muxsel1,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0, j_hiz_b,
     j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck, j_tdi,
     j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, psdo, rst_b,
     smc_load_nvcm_bstream, smc_osc_fsel, smc_oscoff_b, smc_podt_off,
     smc_podt_rst, smc_read, smc_row_inc, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rsr_rst, smc_rwl_en, smc_seq_rst,
     smc_wcram_rst, smc_wdis_dclk, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, tdo_oe_pad, tdo_pad,
     bm_bank_sdo, boot, bp0, bschain_sdo, cdone_in, cm_last_rsr,
     cm_monitor_cell, cm_sdo_u0, cm_sdo_u1, cm_sdo_u2, cm_sdo_u3,
     cnt_podt_out, coldboot_sel, creset_b, idcode_msb20bits, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     osc_clk, por_b, psdi, spi_clk_in, spi_sdi, spi_ss_in_b, tck_pad,
     tdi_pad, tms_pad, trst_pad, warmboot_sel );
output  bm_clk, bm_init, bm_rcapmux_en, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_clk, data_muxsel,
     data_muxsel1, en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0,
     j_hiz_b, j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck,
     j_tdi, j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, rst_b,
     smc_load_nvcm_bstream, smc_oscoff_b, smc_podt_off, smc_podt_rst,
     smc_read, smc_row_inc, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rsr_rst, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_wdis_dclk, smc_write, smc_wset_prec, smc_wset_precgnd,
     smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_oe_pad, tdo_pad;

input  boot, bp0, bschain_sdo, cdone_in, cm_last_rsr, cnt_podt_out,
     creset_b, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, osc_clk, por_b, spi_clk_in, spi_sdi,
     spi_ss_in_b, tck_pad, tdi_pad, tms_pad, trst_pad;

output [10:0]  bm_sa;
output [1:0]  cm_sdi_u2;
output [1:0]  smc_osc_fsel;
output [3:0]  bm_banksel;
output [3:0]  cm_banksel;
output [7:1]  psdo;
output [1:0]  cm_sdi_u3;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_sdi_u0;
output [3:0]  bm_bank_sdi;

input [3:0]  cm_monitor_cell;
input [1:0]  cm_sdo_u0;
input [7:1]  psdi;
input [1:0]  coldboot_sel;
input [1:0]  warmboot_sel;
input [19:0]  idcode_msb20bits;
input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdo_u2;
input [3:0]  bm_bank_sdo;
input [1:0]  cm_sdo_u3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - ice8chip, Cell - ml_cram_logic_ice8p, View - schematic
// LAST TIME SAVED: Oct 22 15:51:24 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_cram_logic_ice8p ( cram_pgateoff, cram_prec, cram_pullup_b,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, smc_clk_out, por,
     smc_clk, smc_read, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rwl_en, smc_seq_rst, smc_wcram_rst, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en );
output  cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, smc_clk_out;

input  por, smc_clk, smc_read, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_write, smc_wset_prec, smc_wset_precgnd, smc_wwlwrt_dis,
     smc_wwlwrt_en;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C2 ( .MINUS(GND_), .PLUS(net326));
nmoscap_25  C1 ( .MINUS(GND_), .PLUS(net306));
nmoscap_25  C0 ( .MINUS(GND_), .PLUS(net314));
tielo I480 ( .tielo(net235));
sg_bufx10_ice8p I461 ( .in(net321), .out(cram_pullup_b));
sg_bufx10_ice8p I446 ( .in(net245), .out(cram_prec));
sg_bufx10_ice8p I457 ( .in(net234), .out(cram_wl_en));
sg_bufx10_ice8p I467 ( .in(net226), .out(cram_pgateoff));
sg_bufx10_ice8p I447 ( .in(cram_write_int), .out(cram_write));
sg_bufx10_ice8p I526 ( .in(net295), .out(cram_vddoff));
nand2_hvt I213 ( .A(net285), .Y(net222), .B(net311));
mux2_hvt I430 ( .in1(net407), .in0(net254), .out(net226),
     .sel(net235));
mux2_hvt I428 ( .in1(cram_write_int), .in0(net319), .out(net230),
     .sel(net285));
mux2_hvt I429 ( .in1(net254), .in0(net230), .out(net234),
     .sel(net235));
mux2_hvt I295 ( .in1(net255), .in0(net293), .out(net238),
     .sel(net285));
nor2_hvt I402 ( .A(net240), .B(smc_wset_precgnd), .Y(net242));
nor2_hvt I329 ( .A(net287), .B(smc_seq_rst), .Y(net245));
nor2_hvt I398 ( .A(smc_rpull_b), .B(net247), .Y(net248));
nor2_hvt I393 ( .A(set_wl_write), .B(reset_logic), .Y(net251));
nor2_hvt I364 ( .A(net426), .B(smc_seq_rst), .Y(net254));
nor2_hvt I400 ( .A(net255), .B(smc_wset_prec), .Y(net257));
nor2_hvt I366 ( .A(reset_logic), .B(net417), .Y(net260));
nor2_hvt I223 ( .A(net359), .B(por), .Y(net263));
nor2_hvt I390 ( .A(smc_write), .B(smc_seq_rst), .Y(net266));
nor2_hvt I392 ( .A(net240), .B(cram_rst), .Y(net269));
nor2_hvt I389 ( .A(net442), .B(reset_logic), .Y(net272));
nor2_hvt I385 ( .A(smc_rprec), .B(net274), .Y(net368));
nor2_hvt I414 ( .A(net276), .B(smc_wwlwrt_en), .Y(net278));
nor2_hvt I391 ( .A(cram_rst), .B(reset_logic), .Y(net281));
inv_hvt I458 ( .A(net272), .Y(rst_rpull_rwl));
inv_hvt I452 ( .A(net266), .Y(net285));
inv_hvt I451 ( .A(net238), .Y(net287));
inv_hvt I459 ( .A(smc_rwl_en), .Y(net289));
inv_hvt I373 ( .A(set_wl_write), .Y(net314));
inv_hvt I346 ( .A(net368), .Y(net293));
inv_hvt I464 ( .A(net222), .Y(net295));
inv_hvt I468 ( .A(net456), .Y(net297));
inv_hvt I454 ( .A(net260), .Y(dis_pgatewrt));
inv_hvt I403 ( .A(net242), .Y(net444));
inv_hvt I450 ( .A(net257), .Y(net303));
inv_hvt I448 ( .A(net281), .Y(net443));
inv_hvt I442 ( .A(net306), .Y(net307));
inv_hvt I444 ( .A(net315), .Y(net306));
inv_hvt I453 ( .A(net269), .Y(net311));
inv_hvt I445 ( .A(net307), .Y(net326));
inv_hvt I435 ( .A(net314), .Y(net315));
inv_hvt I4 ( .A(sm_clk_b), .Y(smc_clk_out));
inv_hvt I421 ( .A(net421), .Y(net319));
inv_hvt I462 ( .A(net247), .Y(net321));
inv_hvt I3 ( .A(smc_clk), .Y(sm_clk_b));
inv_hvt I449 ( .A(net251), .Y(net325));
inv_hvt I443 ( .A(net326), .Y(cram_write_int));
inv_hvt I465 ( .A(cram_rst_int_b), .Y(cram_rst));
inv_hvt I456 ( .A(net263), .Y(reset_logic));
inv_hvt I463 ( .A(net451), .Y(net247));
inv_hvt I460 ( .A(net248), .Y(net335));
inv_hvt I466 ( .A(net297), .Y(cram_rst_int_b));
inv_hvt I256 ( .A(net436), .Y(set_wl_write));
inv_hvt I455 ( .A(net278), .Y(net341));
nor3_hvt I472 ( .B(net347), .Y(net343), .A(net347), .C(net347));
nor3_hvt I471 ( .B(net351), .Y(net347), .A(net351), .C(net351));
nor3_hvt I470 ( .B(net363), .Y(net351), .A(net363), .C(net363));
nor3_hvt I217 ( .B(vdd_tieh), .Y(net355), .A(vdd_tieh), .C(vdd_tieh));
nor3_hvt I386 ( .B(smc_seq_rst), .Y(net359), .A(smc_write),
     .C(smc_read));
nor3_hvt I469 ( .B(net355), .Y(net363), .A(net355), .C(net355));
nor3_hvt I387 ( .B(smc_rwl_en), .Y(net274), .A(net368),
     .C(reset_logic));
nand3_hvt I476 ( .Y(net370), .B(net386), .C(net386), .A(net386));
nand3_hvt I477 ( .Y(net374), .B(net370), .C(net370), .A(net370));
nand3_hvt I478 ( .Y(net378), .B(net374), .C(net374), .A(net374));
nand3_hvt I479 ( .Y(net382), .B(net378), .C(net378), .A(net378));
nand3_hvt I426 ( .Y(net386), .B(vdd_tieh), .C(vdd_tieh), .A(vdd_tieh));
ml_dff I432 ( .R(dis_pgatewrt), .D(net412), .CLK(smc_clk_out),
     .QN(net406), .Q(net407));
ml_dff I431 ( .R(dis_pgatewrt), .D(net254), .CLK(sm_clk_b),
     .QN(net411), .Q(net412));
ml_dff I411 ( .R(reset_logic), .D(smc_wwlwrt_dis), .CLK(smc_clk),
     .QN(net416), .Q(net417));
ml_dff I408 ( .R(rst_rpull_rwl), .D(vdd_tieh), .CLK(net289),
     .QN(net421), .Q(net400));
ml_dff I405 ( .R(dis_pgatewrt), .D(vdd_tieh), .CLK(set_wl_write),
     .QN(net426), .Q(net399));
ml_dff I412 ( .R(net325), .D(net303), .CLK(smc_clk_out), .QN(net394),
     .Q(net255));
ml_dff I410 ( .R(dis_pgatewrt), .D(net341), .CLK(smc_clk_out),
     .QN(net436), .Q(net276));
ml_dff I108 ( .R(reset_logic), .D(smc_rrst_pullwlen),
     .CLK(smc_clk_out), .QN(net402), .Q(net442));
ml_dff I413 ( .R(net443), .D(net444), .CLK(smc_clk_out), .QN(net446),
     .Q(net240));
ml_dff I407 ( .R(rst_rpull_rwl), .D(net335), .CLK(smc_clk_out),
     .QN(net451), .Q(net397));
ml_dff I406 ( .R(reset_logic), .D(smc_wcram_rst), .CLK(smc_clk_out),
     .QN(net456), .Q(net457));
tiehi I427 ( .tiehi(vdd_tieh));

endmodule
// Library - xpmem, Cell - ml_dff_osc, View - schematic
// LAST TIME SAVED: Oct  7 11:47:56 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_dff_osc ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - misc, Cell - ml_mux3_hvt, View - schematic
// LAST TIME SAVED: May 13 15:14:37 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_mux3_hvt ( out, in0, in1, in2, sel );
output  out;

input  in0, in1, in2;

input [3:0]  sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I21 ( .A(sel[0]), .Y(net30));
inv_hvt I24 ( .A(sel[1]), .Y(net28));
inv_hvt I25 ( .A(sel[2]), .Y(net26));
txgate_hvt I23 ( .in(in1), .out(out), .pp(net28), .nn(sel[1]));
txgate_hvt I20 ( .in(in0), .out(out), .pp(net30), .nn(sel[0]));
txgate_hvt I26 ( .in(in2), .out(out), .pp(net26), .nn(sel[2]));
nch_hvt  MN19 ( .D(out), .B(gnd_), .G(sel[3]), .S(gnd_));

endmodule
// Library - misc, Cell - ml_osc_stage, View - schematic
// LAST TIME SAVED: Sep 30 16:59:25 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_osc_stage ( out, clkin, oscen_b, pbias, sel_trim );
output  out;

input  clkin, oscen_b, pbias;

input [3:0]  sel_trim;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C5 ( .MINUS(gnd_), .PLUS(loadbot_0));
nmoscap_25  C6 ( .MINUS(gnd_), .PLUS(loadbot_1));
nmoscap_25  C4 ( .MINUS(gnd_), .PLUS(loadbot_2));
nch_hvt  MN41 ( .D(loadbot_0), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN39 ( .D(loadbot_2), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN29 ( .D(out), .B(gnd_), .G(in_bot), .S(gnd_));
nch_hvt  MN42 ( .D(loadbot_1), .B(gnd_), .G(net419), .S(gnd_));
pch_hvt  M3 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net456));
pch_hvt  M2 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net452));
pch_hvt  MP30 ( .D(net452), .B(vdd_), .G(oscen_b), .S(vdd_));
pch_hvt  MP72 ( .D(net456), .B(vdd_), .G(sel_trim[2]), .S(net452));
pch_hvt  MP33 ( .D(out), .B(vdd_), .G(in_bot), .S(vdd_));
inv_hvt I229 ( .A(net403), .Y(net419));
nor2_hvt I228 ( .A(clkin), .B(oscen_b), .Y(net403));
ml_mux3_hvt Iml_mux3_hvt_bot ( .in1(loadbot_1), .in0(loadbot_0),
     .out(in_bot), .sel(sel_trim[3:0]), .in2(loadbot_2));

endmodule
// Library - misc, Cell - ml_osc_logic, View - schematic
// LAST TIME SAVED: Oct  7 11:48:52 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_osc_logic ( sel_trim, clkin, smc_osc_fsel, smc_oscen );

input  clkin, smc_oscen;

output [3:0]  sel_trim;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:1]  in_sel;



ml_dff_osc I174 ( .R(reset_ff), .D(net050), .CLK(clkin_buf_b),
     .QN(net150), .Q(net172));
ml_dff_osc I238 ( .R(reset_ff), .D(net050), .CLK(clkin_buf),
     .QN(net154), .Q(net177));
ml_dff_osc I244 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf),
     .QN(net155), .Q(net182));
ml_dff_osc I245 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf_b),
     .QN(net153), .Q(net187));
ml_dff_osc I242 ( .R(reset_ff), .D(net048), .CLK(clkin_buf_b),
     .QN(net191), .Q(net192));
ml_dff_osc I243 ( .R(reset_ff), .D(net048), .CLK(clkin_buf),
     .QN(net152), .Q(net197));
nor2_hvt I256 ( .A(smc_osc_fsel[1]), .B(smc_osc_fsel[0]),
     .Y(in_sel[2]));
inv_hvt I293 ( .A(net197), .Y(net052));
inv_hvt I263 ( .A(clkin_buf), .Y(net065));
inv_hvt I283 ( .A(clkin_buf_b), .Y(clkin_buf));
inv_hvt I284 ( .A(smc_oscen), .Y(reset_ff));
inv_hvt I282 ( .A(clkin), .Y(clkin_buf_b));
inv_hvt I255 ( .A(smc_osc_fsel[1]), .Y(in_sel[1]));
inv_hvt I294 ( .A(net192), .Y(net054));
inv_hvt I295 ( .A(net177), .Y(net057));
inv_hvt I296 ( .A(net172), .Y(net061));
inv_hvt I261 ( .A(in_sel[2]), .Y(net050));
inv_hvt I262 ( .A(in_sel[1]), .Y(net048));
inv_hvt I299 ( .A(net059), .Y(net0143));
inv_hvt I297 ( .A(net065), .Y(net063));
inv_hvt I302 ( .A(net094), .Y(net096));
inv_hvt I298 ( .A(net063), .Y(net059));
inv_hvt I304 ( .A(net0143), .Y(net092));
inv_hvt I303 ( .A(net092), .Y(net094));
inv_hvt I301 ( .A(net096), .Y(clkin_buf_delay));
inv_hvt I285 ( .A(net058), .Y(sel_trim[3]));
tiehis I281 ( .tiehi(net058));
ml_mux2_hvt I279 ( .in1(net182), .in0(net187), .out(sel_trim[0]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I277 ( .in1(net057), .in0(net061), .out(sel_trim[2]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I278 ( .in1(net052), .in0(net054), .out(sel_trim[1]),
     .sel(clkin_buf_delay));

endmodule
// Library - misc, Cell - ml_osc, View - schematic
// LAST TIME SAVED: Oct  7 11:48:19 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_osc ( clk_out, smc_osc_fsel, smc_oscen );
output  clk_out;

input  smc_oscen;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sel_trim;



ml_dff_osc I174 ( .R(oscen_b), .D(clkby2_b), .CLK(clk_dffin),
     .QN(clkby2_b), .Q(clkby2));
ml_dff_osc I279 ( .R(oscen_b), .D(net063), .CLK(net0115), .QN(net063),
     .Q(net066));
rppolywo_m  R18 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net437), .PLUS(net383), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R3 ( .MINUS(net366), .PLUS(net076), .BULK(gnd_));
rppolywo_m  R2 ( .MINUS(net383), .PLUS(net366), .BULK(gnd_));
rppolywo_m  R5 ( .MINUS(net070), .PLUS(pbias), .BULK(gnd_));
rppolywo_m  R4 ( .MINUS(net076), .PLUS(net070), .BULK(gnd_));
nch_hvt  MN31 ( .D(net437), .B(gnd_), .G(smc_oscen), .S(gnd_));
pch_hvt  M0 ( .D(net0101), .B(vdd_), .G(oscen_b), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(net0101));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(smc_oscen), .S(vdd_));
nand2_hvt I175 ( .A(out_bot), .Y(clk_dffin), .B(out_top));
inv_hvt I280 ( .A(clkby2), .Y(net0115));
inv_hvt I222 ( .A(clkby2), .Y(clkby2_b_buf));
inv_hvt I220 ( .A(clkby2_b), .Y(clkby2_buf));
inv_hvt I176 ( .A(net063), .Y(clk_out));
inv_hvt I198 ( .A(smc_oscen), .Y(oscen_b));
ml_osc_stage Istage_bot ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_b_buf), .out(out_bot), .sel_trim(sel_trim[3:0]));
ml_osc_stage Istage_top ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_buf), .out(out_top), .sel_trim(sel_trim[3:0]));
ml_osc_logic Iosc_logic ( .sel_trim(sel_trim[3:0]),
     .smc_oscen(smc_oscen), .smc_osc_fsel(smc_osc_fsel[1:0]),
     .clkin(clk_out));

endmodule
// Library - misc, Cell - ml_osc_top, View - schematic
// LAST TIME SAVED: Oct 13 10:43:19 2010
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ml_osc_top ( cnt_podt_out, smc_clk, crst_b, por_b, smc_osc_fsel,
     smc_oscoff_b, smc_podt_off, smc_podt_rst );
output  cnt_podt_out, smc_clk;

input  crst_b, por_b, smc_oscoff_b, smc_podt_off, smc_podt_rst;

input [1:0]  smc_osc_fsel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  q_b;

wire  [10:0]  q;



ml_dff_osc I230 ( .R(cnt_rst), .D(net076), .CLK(q_b[10]), .QN(net067),
     .Q(net063));
ml_dff_osc I243 ( .R(rst_off_latch), .D(net0174), .CLK(clk_out_b),
     .QN(smc_off_b), .Q(net0152));
ml_dff_osc I228_10_ ( .R(cnt_rst), .D(q_b[10]), .CLK(q[9]),
     .QN(q_b[10]), .Q(q[10]));
ml_dff_osc I228_9_ ( .R(cnt_rst), .D(q_b[9]), .CLK(q[8]), .QN(q_b[9]),
     .Q(q[9]));
ml_dff_osc I228_8_ ( .R(cnt_rst), .D(q_b[8]), .CLK(q[7]), .QN(q_b[8]),
     .Q(q[8]));
ml_dff_osc I228_7_ ( .R(cnt_rst), .D(q_b[7]), .CLK(q[6]), .QN(q_b[7]),
     .Q(q[7]));
ml_dff_osc I228_6_ ( .R(cnt_rst), .D(q_b[6]), .CLK(q[5]), .QN(q_b[6]),
     .Q(q[6]));
ml_dff_osc I228_5_ ( .R(cnt_rst), .D(q_b[5]), .CLK(q[4]), .QN(q_b[5]),
     .Q(q[5]));
ml_dff_osc I228_4_ ( .R(cnt_rst), .D(q_b[4]), .CLK(q[3]), .QN(q_b[4]),
     .Q(q[4]));
ml_dff_osc I228_3_ ( .R(cnt_rst), .D(q_b[3]), .CLK(q[2]), .QN(q_b[3]),
     .Q(q[3]));
ml_dff_osc I228_2_ ( .R(cnt_rst), .D(q_b[2]), .CLK(q[1]), .QN(q_b[2]),
     .Q(q[2]));
ml_dff_osc I228_1_ ( .R(cnt_rst), .D(q_b[1]), .CLK(q[0]), .QN(q_b[1]),
     .Q(q[1]));
ml_dff_osc I228_0_ ( .R(cnt_rst), .D(q_b[0]), .CLK(clk_in),
     .QN(q_b[0]), .Q(q[0]));
nand2_hvt I227 ( .A(smc_off_b), .B(rst_osc_b), .Y(disable_osc));
nand2_hvt I270 ( .A(crst_b), .Y(net064), .B(por_b));
inv_hvt I233 ( .A(clk_out), .Y(clk_out_b));
inv_hvt I271 ( .A(net064), .Y(rst_osc_b));
inv_hvt I267 ( .A(net078), .Y(clk_in));
inv_hvt I262 ( .A(net067), .Y(cnt_podt_out));
inv_hvt I275 ( .A(smc_oscoff_b), .Y(net0174));
inv_hvt I277 ( .A(net054), .Y(cnt_rst));
inv_hvt I229 ( .A(rst_osc_b), .Y(net090));
inv_hvt I253 ( .A(net0124), .Y(rst_off_latch));
inv_hvt I232 ( .A(clk_out_b), .Y(smc_clk));
nor2_hvt I272 ( .A(net066), .B(disable_osc), .Y(smc_oscen));
nor2_hvt I266 ( .A(clk_out), .B(smc_podt_off), .Y(net078));
nor2_hvt I273 ( .A(smc_oscoff_b), .B(rst_osc_b), .Y(net066));
nor2_hvt I276 ( .A(net090), .B(smc_podt_rst), .Y(net054));
nor2_hvt I274 ( .A(smc_oscoff_b), .B(cnt_rst), .Y(net0124));
tiehis I179 ( .tiehi(net076));
ml_osc Iml_osc ( .smc_osc_fsel(smc_osc_fsel[1:0]), .clk_out(clk_out),
     .smc_oscen(smc_oscen));

endmodule
// Library - ice1chip, Cell - CHIP_route_lft2rgt_ice1f, View -
//schematic
// LAST TIME SAVED: Apr 28 15:21:41 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module CHIP_route_lft2rgt_ice1f ( bm_banksel_i[3:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa[7:0], bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i[3:0], bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0,
     cdone_out, ceb0, cm_banksel_blbrd_2_, cm_banksel_bldld[1:0],
     cm_banksel_bltrd1_3_, cm_clk_blbrd, cm_clk_bltrd1, cm_sdi_u0[1:0],
     cm_sdi_u1[1:0], cm_sdi_u2d[1:0], cm_sdi_u3d2[1:0], core_por_b0,
     core_por_b1, core_por_b_rowu3, core_por_bb, cram_pgateoff,
     cram_prec, cram_prec_bltrd1, cram_pullup_b, cram_pullup_b_bltrd1,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, cram_write_bltrd1,
     data_muxsel1_blbrd, data_muxsel1_bltrd1, data_muxsel_blbrd,
     data_muxsel_bltrd1, en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1,
     end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     last_rsr[1:0], md_spi_b, mode0, mux_jtag_sel, nvcm_spi_sdi,
     nvcm_spi_ss_b, pgate_r[287:0], reset_b_r[287:0], row_test0, rst_b,
     sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1,
     smc_write0, smc_write_bltl1d1, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, update0, vdd_cntl_r[287:0], wl_r[287:0],
     bm_sdo_o[3:0], bp0, cdone_in, cm_sdo_u0d1[1:0], cm_sdo_u1d3[1:0],
     cm_sdo_u2d1[1:0], cm_sdo_u3[1:0], creset_b_int, fabric_out_12_00,
     fabric_out_13_01, fabric_out_13_02, fromsdo, last_rsr3, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, spi_ss_in_bbank[4:0],
     tck_pad, tdi_pad, tms_pad, trstb_pad, vddio_rightbank );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bltrd1_3_, cm_clk_blbrd,
     cm_clk_bltrd1, core_por_b0, core_por_b1, core_por_b_rowu3,
     core_por_bb, cram_pgateoff, cram_prec, cram_prec_bltrd1,
     cram_pullup_b, cram_pullup_b_bltrd1, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, cram_write_bltrd1, data_muxsel1_blbrd,
     data_muxsel1_bltrd1, data_muxsel_blbrd, data_muxsel_bltrd1,
     en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1, end_of_startup,
     gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, mux_jtag_sel, nvcm_spi_sdi, nvcm_spi_ss_b, row_test0,
     rst_b, sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1,
     smc_write0, smc_write_bltl1d1, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, update0;

input  bp0, cdone_in, creset_b_int, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fromsdo, last_rsr3, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, tck_pad, tdi_pad,
     tms_pad, trstb_pad, vddio_rightbank;

output [287:0]  reset_b_r;
output [3:0]  bm_sdi_i;
output [1:0]  cm_banksel_bldld;
output [1:0]  cm_sdi_u3d2;
output [287:0]  pgate_r;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_sdi_u2d;
output [10:0]  bm_sa;
output [1:0]  last_rsr;
output [287:0]  vdd_cntl_r;
output [1:0]  cm_sdi_u0;
output [287:0]  wl_r;
output [3:0]  bm_banksel_i;

input [1:0]  cm_sdo_u0d1;
input [1:0]  cm_sdo_u3;
input [1:0]  cm_sdo_u2d1;
input [1:0]  cm_sdo_u1d3;
input [3:0]  bm_sdo_o;
input [4:0]  spi_ss_in_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net447;

wire  [1:0]  net350;

wire  [1:0]  cdsbus0;

wire  [3:0]  cm_banksel;

wire  [1:0]  net334;

wire  [1:0]  net446;

wire  [1:0]  net332;

wire  [1:0]  smc_osco_fsel;

wire  [1:0]  dff_out_top;

wire  [1:0]  net354;

wire  [6:0]  net0409;

wire  [1:0]  net336;

wire  [1:0]  net448;

wire  [1:0]  net346;



tiehi I_tiehi ( .tiehi(tvdd_idcode));
CHIP_route_lft_ice1f I_chip_route_lft2rgt_ice1f (
     .pgate_l(pgate_r[287:0]), .reset_l(reset_b_r[287:0]),
     .vdd_cntl_l(vdd_cntl_r[287:0]), .wl_l(wl_r[287:0]),
     .tck_padl0(j_tck), .smc_writel0(smc_write0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbrd),
     .smc_rsr_rstl0(smc_rsr_rst), .smc_row_incl0(smc_row_inc),
     .row_testl1(row_test0), .j_rst_bl0(j_rst_b),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbrd),
     .data_muxsel_blbld(data_muxsel_blbrd),
     .data_muxsel1_blbld(data_muxsel1_blbrd),
     .cram_write_blbld(cram_write), .cram_wl_enl0(cram_wl_en),
     .cram_vddoffl0(cram_vddoff), .cram_rstl0(cram_rst),
     .cram_pullup_blbld(cram_pullup_b), .cram_prec_blbld(cram_prec),
     .cram_pgateoffl0(cram_pgateoff), .core_por_bbl0(core_por_bb),
     .cm_sdo_u1(cm_sdo_u3[1:0]), .cm_sdi_u1d(cdsbus0[1:0]),
     .cm_clk_blbld(cm_clk_blbrd), .cm_banksel_blbld(cm_banksel[3]),
     .cm_banksel_blbld1(cm_banksel_blbrd_2_),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltrd1),
     .last_rsr(last_rsr[1:0]), .last_rsr0(net485),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu2_b),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltrd1),
     .data_muxsel1_bltld3(data_muxsel1_bltrd1),
     .cram_write_bltld3(cram_write_bltrd1),
     .cram_pullup_bltld3(cram_pullup_b_bltrd1),
     .cram_prec_bltld3(cram_prec_bltrd1),
     .core_por_b_rowu1(core_por_b_rowu3),
     .smc_write_bltld3(smc_write_bltl1d1),
     .cm_sdo_u1d1(dff_out_top[1:0]), .cm_sdi_u1d3(cm_sdi_u3d2[1:0]),
     .cm_clk_bltld3(cm_clk_bltrd1),
     .cm_banksel_bltld3_1_(cm_banksel_bltrd1_3_));
creset_filter I561 ( .in(creset_b_int), .out(crst_filterout));
bram_bufferx16_ice8p I702 ( .in(core_por_b0), .out(core_por_b1));
sg_bufx10_ice8p I558 ( .in(net441), .out(end_of_startup));
sg_bufx10_ice8p I559 ( .in(net439), .out(gsr));
sg_bufx10_ice8p I560 ( .in(net440), .out(gint_hz));
sg_bufx10_ice8p I550_1_ ( .in(net346[0]), .out(net332[0]));
sg_bufx10_ice8p I550_0_ ( .in(net346[1]), .out(net332[1]));
sg_bufx10_ice8p I476_1_ ( .in(net350[0]), .out(net334[0]));
sg_bufx10_ice8p I476_0_ ( .in(net350[1]), .out(net334[1]));
sg_bufx10_ice8p I478_1_ ( .in(net354[0]), .out(net336[0]));
sg_bufx10_ice8p I478_0_ ( .in(net354[1]), .out(net336[1]));
sg_bufx10_ice8p I479_1_ ( .in(net334[0]), .out(cm_sdi_u0[1]));
sg_bufx10_ice8p I479_0_ ( .in(net334[1]), .out(cm_sdi_u0[0]));
sg_bufx10_ice8p I480_1_ ( .in(net336[0]), .out(cm_sdi_u2d[1]));
sg_bufx10_ice8p I480_0_ ( .in(net336[1]), .out(cm_sdi_u2d[0]));
sg_bufx10_ice8p I481_1_ ( .in(net332[0]), .out(cm_sdi_u1[1]));
sg_bufx10_ice8p I481_0_ ( .in(net332[1]), .out(cm_sdi_u1[0]));
sg_bufx10_ice8p I551 ( .in(en_8bconfig_b_blbrd), .out(net0327));
sg_bufx10_ice8p I722_1_ ( .in(net447[0]), .out(net346[0]));
sg_bufx10_ice8p I722_0_ ( .in(net447[1]), .out(net346[1]));
sg_bufx10_ice8p I683_1_ ( .in(cm_banksel[1]),
     .out(cm_banksel_bldld[1]));
sg_bufx10_ice8p I683_0_ ( .in(cm_banksel[0]),
     .out(cm_banksel_bldld[0]));
sg_bufx10_ice8p I664_1_ ( .in(net448[0]), .out(net350[0]));
sg_bufx10_ice8p I664_0_ ( .in(net448[1]), .out(net350[1]));
sg_bufx10_ice8p I681 ( .in(cm_banksel[2]), .out(cm_banksel_blbrd_2_));
sg_bufx10_ice8p I723_1_ ( .in(net446[0]), .out(net354[0]));
sg_bufx10_ice8p I723_0_ ( .in(net446[1]), .out(net354[1]));
SMC_CORE_POR_right_ice8p I_SMC_CORE_POR_right (
     .core_por_b0(core_por_b0), .core_por_bb(core_por_bb),
     .vddio_rightbank(vddio_rightbank), .smc_por_b(smc_por_b0),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .creset_b(crst_filterout));
smc_and_jtag_ice8p I_smc_and_jtag_ice8p ( .bm_sa(bm_sa[10:0]),
     .warmboot_sel({fabric_out_13_02, fabric_out_13_01}),
     .trst_pad(trstb_pad), .tms_pad(tms_pad), .tdi_pad(tdi_pad),
     .tck_pad(tck_pad), .spi_ss_in_b(spi_ss_in_bbank[4]),
     .cdone_in(cdone_in), .spi_sdi(spi_ss_in_bbank[2]),
     .spi_clk_in(spi_ss_in_bbank[3]), .psdi({net497, net497, net497,
     net497, net497, net497, net497}), .por_b(smc_por_b0),
     .osc_clk(osc_clk), .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .idcode_msb20bits({tgnd_idcode, tgnd_idcode, tgnd_idcode,
     tvdd_idcode, tgnd_idcode, tgnd_idcode, tgnd_idcode, tvdd_idcode,
     tgnd_idcode, tgnd_idcode, tgnd_idcode, tgnd_idcode, tgnd_idcode,
     tgnd_idcode, tgnd_idcode, tgnd_idcode, tgnd_idcode, tgnd_idcode,
     tgnd_idcode, tvdd_idcode}), .creset_b(crst_filterout),
     .coldboot_sel(spi_ss_in_bbank[1:0]), .cnt_podt_out(cnt_podt_out),
     .cm_sdo_u3(dff_out_top[1:0]), .cm_sdo_u2(cm_sdo_u2d1[1:0]),
     .cm_sdo_u1(cm_sdo_u1d3[1:0]), .cm_sdo_u0(cm_sdo_u0d1[1:0]),
     .cm_monitor_cell({net497, net497, net497, net497}),
     .cm_last_rsr(last_rsr3), .bschain_sdo(fromsdo), .bp0(bp0),
     .boot(fabric_out_12_00), .bm_bank_sdo(bm_sdo_o[3:0]),
     .tdo_pad(totdopad), .tdo_oe_pad(sdo_enable),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out),
     .smc_wwlwrt_en(smc_wwlwrt_en), .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wdis_dclk(smc_wdis_dclk_blbrd),
     .smc_wcram_rst(smc_wcram_rst), .smc_seq_rst(smc_seq_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rsr_rst(smc_rsr_rst),
     .smc_rrst_pullwlen(smc_rrst_pullwlen), .smc_rpull_b(smc_rpull_b),
     .smc_rprec(smc_rprec), .smc_row_inc(smc_row_inc),
     .smc_read(smc_read), .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .psdo({net0409[0], net0409[1], net0409[2], net0409[3], net0409[4],
     net0409[5], net0409[6]}), .nvcm_spi_ss_b(nvcm_spi_ss_b),
     .nvcm_spi_sdi(nvcm_spi_sdi), .md_spi_b(md_spi_b),
     .j_upd_dr(update0), .j_tdi(j_tdi), .j_tck(j_tck),
     .j_shift0(shift0), .j_sft_dr(shiftromsmc), .j_rst_b(j_rst_b),
     .j_row_test(row_test0), .j_mode(mode0), .j_hiz_b(hiz_b0),
     .j_ceb0(ceb0), .gsr(net439), .gint_hz(net440),
     .end_of_startup(net441), .en_8bconfig_b(en_8bconfig_b_blbrd),
     .data_muxsel1(data_muxsel1_blbrd),
     .data_muxsel(data_muxsel_blbrd), .cm_sdi_u3(cdsbus0[1:0]),
     .cm_sdi_u2({net446[0], net446[1]}), .cm_sdi_u1({net447[0],
     net447[1]}), .cm_sdi_u0({net448[0], net448[1]}), .cm_clk(cm_clk),
     .cm_banksel(cm_banksel[3:0]), .cdone_out(cdone_out),
     .bs_en(bs_en0), .bm_wdummymux_en(bm_wdummymux_en_i),
     .bm_sweb(bm_sweb_i), .bm_sreb(bm_sreb_i), .bm_sclkrw(bm_sclkrw_i),
     .bm_rcapmux_en(bm_rcapmux_en_i), .bm_init(bm_init_i),
     .bm_clk(bm_sclk_i), .bm_banksel(bm_banksel_i[3:0]),
     .bm_bank_sdi(bm_sdi_i[3:0]));
ml_cram_logic_ice8p ml_cram_logic_ice8p_1f (
     .smc_wwlwrt_en(smc_wwlwrt_en), .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wcram_rst(smc_wcram_rst), .smc_seq_rst(smc_seq_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rrst_pullwlen(smc_rrst_pullwlen),
     .smc_rpull_b(smc_rpull_b), .smc_rprec(smc_rprec),
     .smc_read(smc_read), .smc_clk(cm_clk), .por(core_por_bb),
     .smc_clk_out(cm_clk_blbrd), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff));
inv_hvt Imux4jtag_sel ( .A(trstb_pad), .Y(mux_jtag_sel));
ml_osc_top I_ml_osc_top ( .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]), .por_b(core_por_b0),
     .crst_b(crst_filterout), .smc_clk(osc_clk),
     .cnt_podt_out(cnt_podt_out));
tielo I_tielo ( .tielo(tgnd_idcode));
tielo I553 ( .tielo(net497));

endmodule
// Library - xpmem, Cell - cram2x2x5, View - schematic
// LAST TIME SAVED: May 11 15:38:01 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module cram2x2x5 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [19:0]  q_b;
output [19:0]  q;

inout [9:0]  bl;

input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  r_gnd;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - ice1chip, Cell - CHIP_route_bot_ice1f_blbank, View -
//schematic
// LAST TIME SAVED: Mar  8 09:53:19 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module CHIP_route_bot_ice1f_blbank ( cm_sdo_u0, cm_sdo_u2, bl_bot,
     cm_banksel_blbld1_0_, cm_banksel_blbrd_2_, cm_clk_blbld,
     cm_clk_blbrd, cm_sdi_u0d1, cm_sdi_u2d, core_por_bb, core_por_bbl0,
     cram_prec, cram_prec_blbld, cram_pullup_b, cram_pullup_blbld,
     cram_write, cram_write_blbld, data_muxsel1_blbld,
     data_muxsel1_blbrd, data_muxsel_blbld, data_muxsel_blbrd,
     en_8bconfig_b_blbld, en_8bconfig_b_blbrd, smc_wdis_dclk_blbld,
     smc_wdis_dclk_blbrd, smc_write, smc_writel0 );


input  cm_banksel_blbld1_0_, cm_banksel_blbrd_2_, cm_clk_blbld,
     cm_clk_blbrd, core_por_bb, core_por_bbl0, cram_prec,
     cram_prec_blbld, cram_pullup_b, cram_pullup_blbld, cram_write,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel1_blbrd,
     data_muxsel_blbld, data_muxsel_blbrd, en_8bconfig_b_blbld,
     en_8bconfig_b_blbrd, smc_wdis_dclk_blbld, smc_wdis_dclk_blbrd,
     smc_write, smc_writel0;

output [1:0]  cm_sdo_u2;
output [1:0]  cm_sdo_u0;

inout [663:0]  bl_bot;

input [1:0]  cm_sdi_u2d;
input [1:0]  cm_sdi_u0d1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



CHIP_route_top_ice1f I_CHIP_route_top_ice1f ( .bl_top(bl_bot[663:0]),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_blbld),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_blbrd),
     .en_8bconfig_b_bltld3(en_8bconfig_b_blbld),
     .data_muxsel_bltrd1(data_muxsel_blbrd),
     .data_muxsel_bltld3(data_muxsel_blbld),
     .data_muxsel1_bltrd1(data_muxsel1_blbrd),
     .data_muxsel1_bltld3(data_muxsel1_blbld),
     .cram_write_bltrd1(cram_write),
     .cram_write_bltld3(cram_write_blbld),
     .cram_pullup_bltld3(cram_pullup_blbld),
     .cram_pullup_b_bltrd1(cram_pullup_b),
     .cram_prec_bltrd1(cram_prec), .core_por_b_rowu3(core_por_bb),
     .core_por_b_rowu1(core_por_bbl0), .cm_sdi_u3d2(cm_sdi_u2d[1:0]),
     .cm_sdi_u1d3(cm_sdi_u0d1[1:0]), .cm_prec_bltld3(cram_prec_blbld),
     .cm_clk_bltrd1(cm_clk_blbrd), .cm_clk_bltld3(cm_clk_blbld),
     .cm_banksel_bltrd1(cm_banksel_blbrd_2_),
     .cm_banksel_bltld3(cm_banksel_blbld1_0_),
     .cm_sdo_u3(cm_sdo_u2[1:0]), .cm_sdo_u1(cm_sdo_u0[1:0]),
     .smc_write_bltld3(smc_writel0), .smc_write_bltl1d1(smc_write));

endmodule
// Library - ice1chip, Cell - CHIP_route_bot_ice1f, View - schematic
// LAST TIME SAVED: Apr 22 10:25:51 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module CHIP_route_bot_ice1f ( cm_banksel_blbld1_0_,
     cm_banksel_blbld_1_, cm_clk_blbld, cm_sdi_u1d, cm_sdo_u0d1,
     cm_sdo_u1d3, cm_sdo_u2d1, core_por_b2, core_por_bbl0,
     cram_pgateoffl0, cram_prec_blbld, cram_pullup_blbld, cram_rstl0,
     cram_vddoffl0, cram_wl_enl0, cram_write_blbld, data_muxsel1_blbld,
     data_muxsel_blbld, en_8bconfig_b_blbld, j_rst_bl0, last_rsr3,
     row_testl1, smc_core_por_bottom1, smc_core_por_bottom2,
     smc_row_incl0, smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0,
     spi_ss_in_bbankd, tck_padl0, bl_bot, cm_banksel,
     cm_banksel_blbrd_2_, cm_clk_blbrd, cm_sdi_u0, cm_sdi_u1,
     cm_sdi_u2d, cm_sdo_u1d1, core_por_b0, core_por_bb, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     spi_ss_in_bbank, vddio_botbank, vddio_spi );
output  cm_banksel_blbld1_0_, cm_banksel_blbld_1_, cm_clk_blbld,
     core_por_b2, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, last_rsr3, row_testl1,
     smc_core_por_bottom1, smc_core_por_bottom2, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;


input  cm_banksel_blbrd_2_, cm_clk_blbrd, core_por_b0, core_por_bb,
     cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     vddio_botbank, vddio_spi;

output [1:0]  cm_sdo_u2d1;
output [4:0]  spi_ss_in_bbankd;
output [1:0]  cm_sdo_u0d1;
output [1:0]  cm_sdi_u1d;
output [1:0]  cm_sdo_u1d3;

inout [663:0]  bl_bot;

input [1:0]  cm_sdi_u0;
input [4:0]  spi_ss_in_bbank;
input [1:0]  cm_sdi_u2d;
input [1:0]  cm_sdi_u1;
input [1:0]  cm_sdo_u1d1;
input [1:0]  cm_banksel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1_buf;

wire  [1:0]  net233;

wire  [1:0]  cm_sdo_u0_buf;

wire  [1:0]  net297;

wire  [1:0]  dff_u2_d0;

wire  [1:0]  cm_sdi_u2d_buf;

wire  [1:0]  net321;

wire  [1:0]  net229;

wire  [1:0]  net317;

wire  [1:0]  net235;

wire  [1:0]  net234;

wire  [1:0]  cm_sdi_u0d1;

wire  [1:0]  cm_sdo_u2;

wire  [1:0]  dff_u0_d1;

wire  [1:0]  dff_u1_d1;

wire  [1:0]  cm_sdo_u0;



CHIP_route_bot_ice1f_blbank I_CHIP_route_bot_ice1f_blbank (
     .bl_bot(bl_bot[663:0]), .smc_writel0(smc_writel0),
     .smc_write(smc_write), .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_write(cram_write),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_pullup_b(cram_pullup_b), .cram_prec_blbld(cram_prec_blbld),
     .cram_prec(cram_prec), .core_por_bbl0(core_por_bbl0),
     .core_por_bb(core_por_bb), .cm_sdi_u2d(cm_sdi_u2d_buf[1:0]),
     .cm_sdi_u0d1(cm_sdi_u0d1[1:0]), .cm_clk_blbrd(cm_clk_blbrd),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1_0_),
     .cm_sdo_u0(cm_sdo_u0[1:0]), .cm_sdo_u2(cm_sdo_u2[1:0]));
tielo I561_1_ ( .tielo(net229[0]));
tielo I561_0_ ( .tielo(net229[1]));
tielo I562 ( .tielo(net230));
tielo I563 ( .tielo(net231));
tielo I564 ( .tielo(net232));
tielo I559_1_ ( .tielo(net233[0]));
tielo I559_0_ ( .tielo(net233[1]));
tielo I560_1_ ( .tielo(net234[0]));
tielo I560_0_ ( .tielo(net234[1]));
sg_bufx10_ice8p I532_1_ ( .in(net235[0]), .out(cm_sdi_u1d[1]));
sg_bufx10_ice8p I532_0_ ( .in(net235[1]), .out(cm_sdi_u1d[0]));
sg_bufx10_ice8p I484 ( .in(cram_pgateoff), .out(net327));
sg_bufx10_ice8p I482 ( .in(net239), .out(cram_pgateoffl0));
sg_bufx10_ice8p I516 ( .in(net241), .out(cm_banksel_blbld_1_));
sg_bufx10_ice8p I474 ( .in(net243), .out(net245));
sg_bufx10_ice8p I475 ( .in(net245), .out(smc_writel0));
sg_bufx10_ice8p I480 ( .in(net247), .out(net283));
sg_bufx10_ice8p I333 ( .in(j_rst_b), .out(j_rst_bl0));
sg_bufx10_ice8p I336 ( .in(core_por_bb), .out(net361));
sg_bufx10_ice8p I523 ( .in(smc_clk_mid), .out(cm_clk_blbld));
sg_bufx10_ice8p I478 ( .in(cram_vddoff), .out(net363));
sg_bufx10_ice8p I488 ( .in(predata_cram_pullup_b), .out(net295));
sg_bufx10_ice8p I473 ( .in(smc_write), .out(net243));
sg_bufx10_ice8p I496 ( .in(en_8bconfig_b_blbrd),
     .out(predata_en_8bconfig_b));
sg_bufx10_ice8p I527_1_ ( .in(cm_sdi_u0[1]), .out(net321[0]));
sg_bufx10_ice8p I527_0_ ( .in(cm_sdi_u0[0]), .out(net321[1]));
sg_bufx10_ice8p I459 ( .in(smc_row_inc), .out(net377));
sg_bufx10_ice8p I491 ( .in(cram_write), .out(predata_cram_write));
sg_bufx10_ice8p I568_4_ ( .in(spi_ss_in_bbank[4]),
     .out(spi_ss_in_bbankd[4]));
sg_bufx10_ice8p I568_3_ ( .in(spi_ss_in_bbank[3]),
     .out(spi_ss_in_bbankd[3]));
sg_bufx10_ice8p I568_2_ ( .in(spi_ss_in_bbank[2]),
     .out(spi_ss_in_bbankd[2]));
sg_bufx10_ice8p I568_1_ ( .in(spi_ss_in_bbank[1]),
     .out(spi_ss_in_bbankd[1]));
sg_bufx10_ice8p I568_0_ ( .in(spi_ss_in_bbank[0]),
     .out(spi_ss_in_bbankd[0]));
sg_bufx10_ice8p I467 ( .in(predata_muxsel1), .out(net291));
sg_bufx10_ice8p I505 ( .in(net273), .out(smc_rsr_rstl0));
sg_bufx10_ice8p I567 ( .in(core_por_b0), .out(core_por_b2));
sg_bufx10_ice8p I521 ( .in(net277), .out(cm_banksel_blbld1_0_));
sg_bufx10_ice8p I175 ( .in(net279), .out(data_muxsel_blbld));
sg_bufx10_ice8p I492 ( .in(net281), .out(cram_write_blbld));
sg_bufx10_ice8p I481 ( .in(net283), .out(cram_rstl0));
sg_bufx10_ice8p I439 ( .in(j_tck), .out(tck_padl0));
sg_bufx10_ice8p I495 ( .in(net287), .out(en_8bconfig_b_blbld));
sg_bufx10_ice8p I570 ( .in(net289), .out(core_por_bbl0));
sg_bufx10_ice8p I466 ( .in(net291), .out(data_muxsel1_blbld));
sg_bufx10_ice8p I486 ( .in(net293), .out(cram_prec_blbld));
sg_bufx10_ice8p I489 ( .in(net295), .out(cram_pullup_blbld));
sg_bufx10_ice8p I531_1_ ( .in(net297[0]), .out(net235[0]));
sg_bufx10_ice8p I531_0_ ( .in(net297[1]), .out(net235[1]));
sg_bufx10_ice8p I485 ( .in(cram_prec), .out(predata_cram_prec));
sg_bufx10_ice8p I533_1_ ( .in(cm_sdi_u1[1]), .out(net297[0]));
sg_bufx10_ice8p I533_0_ ( .in(cm_sdi_u1[0]), .out(net297[1]));
sg_bufx10_ice8p I520 ( .in(net303), .out(net277));
sg_bufx10_ice8p I517 ( .in(net305), .out(net241));
sg_bufx10_ice8p I493 ( .in(predata_cram_write), .out(net281));
sg_bufx10_ice8p I519 ( .in(cm_banksel[0]), .out(net303));
sg_bufx10_ice8p I509 ( .in(net311), .out(row_testl1));
sg_bufx10_ice8p I469 ( .in(net313), .out(smc_row_incl0));
sg_bufx10_ice8p I504 ( .in(smc_rsr_rst), .out(net331));
sg_bufx10_ice8p I529_1_ ( .in(net317[0]), .out(cm_sdi_u0d1[1]));
sg_bufx10_ice8p I529_0_ ( .in(net317[1]), .out(cm_sdi_u0d1[0]));
sg_bufx10_ice8p I476 ( .in(net319), .out(cram_vddoffl0));
sg_bufx10_ice8p I530_1_ ( .in(net321[0]), .out(net317[0]));
sg_bufx10_ice8p I530_0_ ( .in(net321[1]), .out(net317[1]));
sg_bufx10_ice8p I471 ( .in(net323), .out(net347));
sg_bufx10_ice8p I510 ( .in(net325), .out(net311));
sg_bufx10_ice8p I483 ( .in(net327), .out(net239));
sg_bufx10_ice8p I464 ( .in(predata_muxsel), .out(net279));
sg_bufx10_ice8p I503 ( .in(net331), .out(net273));
sg_bufx10_ice8p I494 ( .in(predata_en_8bconfig_b), .out(net287));
sg_bufx10_ice8p I490 ( .in(cram_pullup_b),
     .out(predata_cram_pullup_b));
sg_bufx10_ice8p I479 ( .in(cram_rst), .out(net247));
sg_bufx10_ice8p I465 ( .in(data_muxsel1_blbrd), .out(predata_muxsel1));
sg_bufx10_ice8p I525 ( .in(cm_clk_blbrd), .out(predata_smc_clk_out));
sg_bufx10_ice8p I518 ( .in(cm_banksel[1]), .out(net305));
sg_bufx10_ice8p I524 ( .in(predata_smc_clk_out), .out(smc_clk_mid));
sg_bufx10_ice8p I470 ( .in(net347), .out(cram_wl_enl0));
sg_bufx10_ice8p I511 ( .in(row_test0), .out(net325));
sg_bufx10_ice8p I293 ( .in(last_rsr1), .out(last_rsr2));
sg_bufx10_ice8p I541_1_ ( .in(dff_u0_d1[1]), .out(cm_sdo_u0d1[1]));
sg_bufx10_ice8p I541_0_ ( .in(dff_u0_d1[0]), .out(cm_sdo_u0d1[0]));
sg_bufx10_ice8p I539_1_ ( .in(cm_sdo_u1d1[1]), .out(cm_sdo_u1_buf[1]));
sg_bufx10_ice8p I539_0_ ( .in(cm_sdo_u1d1[0]), .out(cm_sdo_u1_buf[0]));
sg_bufx10_ice8p I455 ( .in(data_muxsel_blbrd), .out(predata_muxsel));
sg_bufx10_ice8p I526_1_ ( .in(cm_sdi_u2d[1]), .out(cm_sdi_u2d_buf[1]));
sg_bufx10_ice8p I526_0_ ( .in(cm_sdi_u2d[0]), .out(cm_sdi_u2d_buf[0]));
sg_bufx10_ice8p I569 ( .in(net361), .out(net289));
sg_bufx10_ice8p I477 ( .in(net363), .out(net319));
sg_bufx10_ice8p I566 ( .in(net387), .out(last_rsr3));
sg_bufx10_ice8p I540_1_ ( .in(dff_u1_d1[1]), .out(cm_sdo_u1d3[1]));
sg_bufx10_ice8p I540_0_ ( .in(dff_u1_d1[0]), .out(cm_sdo_u1d3[0]));
sg_bufx10_ice8p I497 ( .in(smc_wdis_dclk_blbrd),
     .out(predata_smc_wdis_dclk));
sg_bufx10_ice8p I487 ( .in(predata_cram_prec), .out(net293));
sg_bufx10_ice8p I498 ( .in(net373), .out(smc_wdis_dclk_blbld));
sg_bufx10_ice8p I499 ( .in(predata_smc_wdis_dclk), .out(net373));
sg_bufx10_ice8p I330 ( .in(net377), .out(net313));
sg_bufx10_ice8p I472 ( .in(cram_wl_en), .out(net323));
sg_dffbuf_modified I462_1_ ( .d(cm_sdo_u0_buf[1]), .clk(smc_clk_mid),
     .dffout(dff_u0_d1[1]), .r(net229[0]));
sg_dffbuf_modified I462_0_ ( .d(cm_sdo_u0_buf[0]), .clk(smc_clk_mid),
     .dffout(dff_u0_d1[0]), .r(net229[1]));
sg_dffbuf_modified I565 ( .d(last_rsr2), .clk(smc_clk_mid),
     .dffout(net387), .r(net232));
sg_dffbuf_modified I537_1_ ( .d(cm_sdo_u1_buf[1]), .clk(smc_clk_mid),
     .dffout(dff_u1_d1[1]), .r(net234[0]));
sg_dffbuf_modified I537_0_ ( .d(cm_sdo_u1_buf[0]), .clk(smc_clk_mid),
     .dffout(dff_u1_d1[0]), .r(net234[1]));
sg_dffbuf_modified I545_1_ ( .d(dff_u2_d0[1]),
     .clk(predata_smc_clk_out), .dffout(cm_sdo_u2d1[1]), .r(net231));
sg_dffbuf_modified I545_0_ ( .d(dff_u2_d0[0]),
     .clk(predata_smc_clk_out), .dffout(cm_sdo_u2d1[0]), .r(net231));
sg_dffbuf_modified I546_1_ ( .d(cm_sdo_u2[1]),
     .clk(predata_smc_clk_out), .dffout(dff_u2_d0[1]), .r(net230));
sg_dffbuf_modified I546_0_ ( .d(cm_sdo_u2[0]),
     .clk(predata_smc_clk_out), .dffout(dff_u2_d0[0]), .r(net230));
sg_dffbuf_modified I535_1_ ( .d(cm_sdo_u0[1]), .clk(cm_clk_blbld),
     .dffout(cm_sdo_u0_buf[1]), .r(net233[0]));
sg_dffbuf_modified I535_0_ ( .d(cm_sdo_u0[0]), .clk(cm_clk_blbld),
     .dffout(cm_sdo_u0_buf[0]), .r(net233[1]));
eh_io_pup_2_new_ice8p Ipor_spi ( .core_por_b(core_por_b0),
     .vdd_io(vddio_spi), .por_b(smc_core_por_bottom2));
eh_io_pup_2_new_ice8p Ipor_iob ( .core_por_b(core_por_b0),
     .vdd_io(vddio_botbank), .por_b(smc_core_por_bottom1));

endmodule
// Library - ice1chip, Cell - ring_route00_ice1f, View - schematic
// LAST TIME SAVED: Apr 22 10:57:27 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ring_route00_ice1f ( bm_banksel_i, bm_init_i, bm_rcapmux_en_i,
     bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bs_en0, cdone_out, ceb0, end_of_startup,
     gint_hz, gsr, hiz_b0, j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr, md_spi_b, mode0,
     mux_jtag_sel_b, pgate_l, pgate_r, reset_b_l, reset_b_r,
     sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_pad, update0, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r, bl_bot, bl_top, vppin, bm_sdo_o, cdone_in, creset_b_int,
     fabric_out_12_00, fabric_out_13_01, fabric_out_13_02, fromsdo,
     spi_ss_in_bbank, tck_pad, tdi_pad, tms_pad, trstb_pad,
     vddio_bottombank, vddio_spi );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     end_of_startup, gint_hz, gsr, hiz_b0, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, mux_jtag_sel_b, sdo_enable, shift0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, tdo_pad, update0;

inout  vppin;

input  cdone_in, creset_b_int, fabric_out_12_00, fabric_out_13_01,
     fabric_out_13_02, fromsdo, tck_pad, tdi_pad, tms_pad, trstb_pad,
     vddio_bottombank, vddio_spi;

output [287:0]  vdd_cntl_l;
output [287:0]  reset_b_r;
output [7:0]  bm_sa_i;
output [287:0]  vdd_cntl_r;
output [3:0]  last_rsr;
output [287:0]  wl_l;
output [287:0]  pgate_l;
output [287:0]  reset_b_l;
output [3:0]  bm_sdi_i;
output [287:0]  pgate_r;
output [3:0]  bm_banksel_i;
output [287:0]  wl_r;

inout [663:0]  bl_top;
inout [663:0]  bl_bot;

input [3:0]  bm_sdo_o;
input [4:0]  spi_ss_in_bbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1d1;

wire  [1:0]  cm_banksel;

wire  [1:0]  cm_sdi_u1d3;

wire  [1:0]  cm_sdi_u1;

wire  [1:1]  cm_banksel_bltld3;

wire  [1:0]  cm_sdi_u3d2;

wire  [1:0]  cm_sdi_u2d;

wire  [1:0]  cm_sdo_u2d1;

wire  [1:0]  cm_sdi_u1d;

wire  [1:0]  cm_sdo_u0d1;

wire  [1:0]  cm_sdo_u3;

wire  [4:0]  spi_ss_in_bbankd;

wire  [1:0]  cm_sdi_u0;

wire  [3:3]  cm_banksel_bltrd1;

wire  [1:0]  cm_sdo_u1d3;

wire  [1:0]  cm_sdo_u1;



nvcm_ml_block_ice1f I_nvcm_ml_block_ice1f ( .spi_ss_b(nvcm_spi_ss_b),
     .spi_sdi(nvcm_spi_sdi), .rst_b(rst_b), .nvcm_ce_b(cdone_in),
     .clk(spi_clk_out2fsm), .spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .spi_sdo(nvcm_spi_sdo), .nvcm_rdy(nvcm_rdy),
     .nvcm_boot(nvcm_boot),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream),
     .fsm_tm_margin0_read(net398), .fsm_recall(net399), .bp0(bp0),
     .vpp(vppin), .nvcm_relextspi(nvcm_relextspi));
CHIP_route_top_ice1f I_CHIP_route_top_ice1f ( .bl_top(bl_top[663:0]),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltld1),
     .data_muxsel1_bltrd1(data_muxsel1_bltld3),
     .data_muxsel1_bltld3(data_muxsel1_bltld1),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_bltld3),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1),
     .core_por_b_rowu3(core_por_b_rowu3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .cm_prec_bltld3(cm_prec_bltld3), .cm_clk_bltrd1(cm_clk_bltrd1),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cm_banksel_bltrd1(cm_banksel_bltrd1[3]),
     .cm_banksel_bltld3(cm_banksel_bltld3[1]),
     .cm_sdo_u3(cm_sdo_u3[1:0]), .cm_sdo_u1(cm_sdo_u1[1:0]),
     .smc_write_bltld3(smc_write_bltld3),
     .smc_write_bltl1d1(smc_write_bltl1d1r));
CHIP_route_lft2rgt_ice1f I_CHIP_route_rgt_ice1f ( bm_banksel_i[3:0],
     bm_init_i, bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i[3:0], bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0,
     cdone_out, ceb0, cm_banksel_blbrd_2_, cm_banksel[1:0],
     cm_banksel_bltrd1[3], cm_clk_blbrd, cm_clk_bltrd1, cm_sdi_u0[1:0],
     cm_sdi_u1[1:0], cm_sdi_u2d[1:0], cm_sdi_u3d2[1:0], core_por_b0,
     net228, core_por_b_rowu3, core_por_bb, cram_pgateoff, cram_prec,
     cram_prec_bltrd1, cram_pullup_b, cram_pullup_b_bltrd1, cram_rst,
     cram_vddoff, cram_wl_en, cram_write, cram_write_bltrd1,
     data_muxsel1_blbrd, data_muxsel1_bltld3, data_muxsel_blbrd,
     data_muxsel_bltrd1, en_8bconfig_b_blbrd, en_8bconfig_b_bltrd1,
     end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     last_rsr[3:2], md_spi_b, mode0, mux_jtag_sel_b, nvcm_spi_sdi,
     nvcm_spi_ss_b, pgate_r[287:0], reset_b_r[287:0], row_test0, rst_b,
     sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rsr, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1, smc_write,
     smc_write_bltl1d1r, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_pad, update0, vdd_cntl_r[287:0], wl_r[287:0],
     bm_sdo_o[3:0], bp0, cdone_in, cm_sdo_u0d1[1:0], cm_sdo_u1d3[1:0],
     cm_sdo_u2d1[1:0], cm_sdo_u3[1:0], creset_b_int, fabric_out_12_00,
     fabric_out_13_01, fabric_out_13_02, fromsdo, last_rsr3, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, spi_ss_in_bbankd[4:0],
     tck_pad, tdi_pad, tms_pad, trstb_pad, vddp_);
CHIP_route_lft_ice1f I_CHIP_route_lft_ice1f ( .pgate_l(pgate_l[287:0]),
     .reset_l(reset_b_l[287:0]), .vdd_cntl_l(vdd_cntl_l[287:0]),
     .wl_l(wl_l[287:0]), .smc_write_bltld3(smc_write_bltld3),
     .tck_padl0(tck_padl0), .smc_writel0(smc_writel0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .smc_rsr_rstl0(smc_rsr_rstl0), .smc_row_incl0(smc_row_incl0),
     .row_testl1(row_testl1), .j_rst_bl0(j_rst_bl0),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_wl_enl0(cram_wl_enl0),
     .cram_vddoffl0(cram_vddoffl0), .cram_rstl0(cram_rstl0),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld),
     .cram_pgateoffl0(cram_pgateoffl0), .core_por_bbl0(core_por_bbl0),
     .cm_sdo_u1(cm_sdo_u1[1:0]), .cm_sdi_u1d(cm_sdi_u1d[1:0]),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbld(cm_banksel_blbld_1_),
     .cm_banksel_blbld1(cm_banksel_blbld1_0_),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3),
     .last_rsr(last_rsr[1:0]), .last_rsr0(last_rsr0),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel_bltld3(data_muxsel_bltld1),
     .data_muxsel1_bltld3(data_muxsel1_bltld1),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_bltld3),
     .cram_prec_bltld3(cm_prec_bltld3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdo_u1d1(cm_sdo_u1d1[1:0]), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cm_banksel_bltld3_1_(cm_banksel_bltld3[1]));
CHIP_route_bot_ice1f I_CHIP_route_bot_ice1f ( .bl_bot(bl_bot[663:0]),
     .core_por_b2(core_por_b2),
     .spi_ss_in_bbankd(spi_ss_in_bbankd[4:0]),
     .spi_ss_in_bbank(spi_ss_in_bbank[4:0]), .vddio_spi(vddio_spi),
     .vddio_botbank(vddio_bottombank), .smc_write(smc_write),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_rsr_rst(smc_rsr_rsr), .smc_row_inc(smc_row_inc),
     .row_test0(row_test0), .last_rsr1(last_rsr0), .j_tck(j_tck),
     .j_rst_b(j_rst_b), .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_blbrd(data_muxsel1_blbrd), .cram_write(cram_write),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff),
     .core_por_bb(core_por_bb), .core_por_b0(core_por_b0),
     .cm_sdo_u1d1(cm_sdo_u1d1[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .cm_clk_blbrd(cm_clk_blbrd),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .cm_banksel(cm_banksel[1:0]), .tck_padl0(tck_padl0),
     .smc_writel0(smc_writel0),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .smc_rsr_rstl0(smc_rsr_rstl0), .smc_row_incl0(smc_row_incl0),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .row_testl1(row_testl1), .last_rsr3(last_rsr3),
     .j_rst_bl0(j_rst_bl0), .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .cram_write_blbld(cram_write_blbld), .cram_wl_enl0(cram_wl_enl0),
     .cram_vddoffl0(cram_vddoffl0), .cram_rstl0(cram_rstl0),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld),
     .cram_pgateoffl0(cram_pgateoffl0), .core_por_bbl0(core_por_bbl0),
     .cm_sdo_u2d1(cm_sdo_u2d1[1:0]), .cm_sdo_u1d3(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0d1(cm_sdo_u0d1[1:0]), .cm_sdi_u1d(cm_sdi_u1d[1:0]),
     .cm_clk_blbld(cm_clk_blbld),
     .cm_banksel_blbld_1_(cm_banksel_blbld_1_),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1_0_));
sg_bufx10_ice8p I_clkbuf ( .in(spi_clk_out), .out(spi_clk_out2fsm));

endmodule
// Library - ice1chip, Cell - LVDS_INBUFFER_ice1f, View - schematic
// LAST TIME SAVED: Apr 20 16:11:20 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module LVDS_INBUFFER_ice1f ( indiff, in_padn, in_padp, vddio, cbit[2],
     cbit[3], cbit[4] );
output  indiff;

inout  in_padn, in_padp, vddio;


input [4:2]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor3_hvt I56 ( .B(net0113), .Y(net0161), .A(cbit[3]), .C(cbit[2]));
nch_25od33  M10 ( .D(net1132), .B(gnd_), .G(net1138), .S(gnd_));
nch_25od33  M8 ( .D(net1138), .B(gnd_), .G(comp_out_25), .S(gnd_));
nch_25od33  M1 ( .D(lvdsen_b_25), .B(gnd_), .G(lvdsen_25), .S(gnd_));
pch_25od33  M9 ( .D(net1138), .B(vddio), .G(comp_out_25), .S(vddio));
pch_25od33  M0 ( .D(comp_out_25), .B(vddio), .G(lvdsen_25), .S(vddio));
pch_25od33  M11 ( .D(net1132), .B(vddio), .G(net1138), .S(vddio));
pch_25od33  M18 ( .D(comp_out_25), .B(vddio), .G(in_padp),
     .S(net1180));
pch_25od33  M13 ( .D(net1180), .B(vddio), .G(net1203), .S(net1184));
pch_25od33  M12 ( .D(net1184), .B(vddio), .G(lvdsen_b_25), .S(vddio));
pch_25od33  M19 ( .D(net1203), .B(vddio), .G(in_padn), .S(net1180));
pch_25od33  M2 ( .D(lvdsen_b_25), .B(vddio), .G(lvdsen_25), .S(vddio));
inv_hvt I129 ( .A(net0161), .Y(net1191));
inv_hvt I131 ( .A(indiff_b), .Y(indiff));
inv_hvt I55 ( .A(cbit[4]), .Y(net0113));
nch_25  x8 ( .D(indiff_b), .B(GND_), .G(net1138), .S(gnd_));
nch_25  M17 ( .D(net1204), .B(gnd_), .G(lvdsen_25), .S(gnd_));
nch_25  M16 ( .D(net1212), .B(gnd_), .G(net1203), .S(net1204));
nch_25  M23 ( .D(net0153), .B(GND_), .G(net1132), .S(gnd_));
nch_25  M21 ( .D(net1203), .B(GND_), .G(in_padn), .S(net1212));
nch_25  M20 ( .D(comp_out_25), .B(GND_), .G(in_padp), .S(net1212));
nch_25  x20 ( .D(lvdsen_25), .B(GND_), .G(net1191), .S(gnd_));
nch_25  x19 ( .D(net1149), .B(GND_), .G(net0161), .S(gnd_));
pch_25  x18 ( .D(net1149), .B(vddio), .G(lvdsen_25), .S(vddio));
pch_25  M5 ( .D(lvdsen_25), .B(vddio), .G(net1149), .S(vddio));
pch_hvt  x12 ( .D(indiff_b), .B(vdd_), .G(net0153), .S(vdd_));
pch_hvt  x13 ( .D(net0153), .B(vdd_), .G(indiff_b), .S(vdd_));

endmodule
// Library - ice1chip, Cell - PLVDS_pair, View - schematic
// LAST TIME SAVED: Apr 20 16:11:22 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module PLVDS_pair ( c_n, c_p, PAD_n, PAD_p, POC, cbit, i_n, i_p, oen_n,
     oen_p, tiegnd, vddio );
output  c_n, c_p;

inout  PAD_n, PAD_p;

input  POC, i_n, i_p, oen_n, oen_p, tiegnd, vddio;

input [4:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



LVDS_INBUFFER_ice1f I_LVDS_INBUFFER ( indiff, in_padn_1, in_padp_0,
     vddio, cbit[3], cbit[2], cbit[4]);
PDUW08SDGZ_G_NOR I_ppart_0 ( .IE(cbit[3]), .POC(POC), .indiff(indiff),
     .PAD4LVDS(in_padp_0), .VDDIO(vddio), .REN(cbit[1]), .PAD(PAD_p),
     .C(c_p), .OEN(oen_p), .I(i_p));
PDUW08SDGZ_G_NOR I_npart_1 ( .IE(cbit[2]), .POC(POC), .indiff(tiegnd),
     .PAD4LVDS(in_padn_1), .VDDIO(vddio), .REN(cbit[0]), .PAD(PAD_n),
     .C(c_n), .OEN(oen_n), .I(i_n));

endmodule
// Library - kplibn40lp, Cell - diodN, View - schematic
// LAST TIME SAVED: May  3 17:09:20 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module diodN ( n1, n2 );
input  n1, n2;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_mac  M2 ( .D(n2), .B(gnd_), .G(n2), .S(n1));

endmodule
// Library - kplibn40lp, Cell - oneNodeN, View - schematic
// LAST TIME SAVED: May  3 17:11:45 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module oneNodeN ( n1 );
input  n1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M2 ( .D(n1), .B(n1), .G(n1), .S(n1));

endmodule
// Library - kplibn40lp, Cell - oneNodeP, View - schematic
// LAST TIME SAVED: May  3 17:12:12 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module oneNodeP ( n1 );
input  n1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch  M2 ( .D(n1), .B(n1), .G(n1), .S(n1));

endmodule
// Library - kplibn40lp, Cell - twoNodeP, View - schematic
// LAST TIME SAVED: May  3 17:13:23 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module twoNodeP ( n1, n2 );
input  n1, n2;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch  M2 ( .D(n2), .B(n2), .G(n1), .S(n2));

endmodule
// Library - kplibn40lp, Cell - twoNodeN, View - schematic
// LAST TIME SAVED: May  3 17:13:01 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module twoNodeN ( n1, n2 );
input  n1, n2;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M2 ( .D(n1), .B(n1), .G(n2), .S(n1));

endmodule
// Library - leafcell, Cell - sbox11to9_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:53:05 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox11to9_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  b;
inout [9:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_l10 ( .prog(prog), .in6(t[4]), .in5(t[10]), .in4(r[2]),
     .in3(r[10]), .in2(r[7]), .in1(b[10]), .in0(b[5]), .out(l[10]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t10 ( .prog(prog), .in6(r[4]), .in5(r[10]), .in4(b[2]),
     .in3(b[10]), .in2(b[7]), .in1(l[10]), .in0(l[5]), .out(t[10]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t11 ( .prog(prog), .in6(r[5]), .in5(r[11]), .in4(b[3]),
     .in3(b[11]), .in2(b[8]), .in1(l[11]), .in0(l[6]), .out(t[11]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t9 ( .prog(prog), .in6(r[3]), .in5(r[9]), .in4(b[1]),
     .in3(b[9]), .in2(b[6]), .in1(l[9]), .in0(l[4]), .out(t[9]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l11 ( .prog(prog), .in6(t[5]), .in5(t[11]), .in4(r[3]),
     .in3(r[11]), .in2(r[8]), .in1(b[11]), .in0(b[6]), .out(l[11]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l9 ( .prog(prog), .in6(t[3]), .in5(t[9]), .in4(r[1]),
     .in3(r[9]), .in2(r[6]), .in1(b[9]), .in0(b[4]), .out(l[9]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - kplibn40lp, Cell - dcapP, View - schematic
// LAST TIME SAVED: Apr 15 15:28:46 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module dcapP ( n1, n2 );
input  n1, n2;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_mac  M2 ( .D(n2), .B(n1), .G(n1), .S(n1));

endmodule
// Library - kplibn40lp, Cell - dcapN, View - schematic
// LAST TIME SAVED: Apr 15 15:27:32 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module dcapN ( n1, n2 );
input  n1, n2;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_mac  M2 ( .D(n2), .B(n1), .G(n1), .S(n1));

endmodule
// Library - misc, Cell - ABIWTCZ4, View - schematic
// LAST TIME SAVED: Apr 18 15:12:04 2011
// NETLIST TIME: May  5 11:56:47 2011
`timescale 1ns / 1ns 

module ABIWTCZ4 ( LOCK, PLLOUT, BYPASS, DIVF0, DIVF1, DIVF2, DIVF3,
     DIVF4, DIVF5, DIVF6, DIVQ0, DIVQ1, DIVQ2, DIVR0, DIVR1, DIVR2,
     DIVR3, FB, FSE, RANGE0, RANGE1, RANGE2, REF, RESET, VDDA );
output  LOCK, PLLOUT;

input  BYPASS, DIVF0, DIVF1, DIVF2, DIVF3, DIVF4, DIVF5, DIVF6, DIVQ0,
     DIVQ1, DIVQ2, DIVR0, DIVR1, DIVR2, DIVR3, FB, FSE, RANGE0, RANGE1,
     RANGE2, REF, RESET, VDDA;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_tri_2 Itrinv_mahvc_d_o_r ( .Tb(N00AESU), .T(N00AETM), .A(N00AEQU),
     .Y(N00AETQ));
inv_tri_2 I_trinv_mahqc_d_o_r ( .Tb(N00AEQN), .T(N00AERD), .A(N00AEQW),
     .Y(N00AERH));
inv_tri_2 Itinv_mahwk_l_w_z ( .Tb(N00AESV), .T(N00AEUC), .A(N00AEQV),
     .Y(N00AEUG));
inv_tri_2 Itrinv_mahrk_l_u_x ( .Tb(N00AEQO), .T(N00AERT), .A(N00AEQX),
     .Y(N00AERY));
nor4_hvt Inor4_xmafnf_g_h_i_oi_j_k_l ( .B(N00ADWK), .Y(N00ADWN),
     .D(N00ADWV), .A(N00ADWL), .C(N00ADWW));
nor3 nor3_XMAHOH_XMAHOI_XMAHOJ_XMAHOM_XMAHOK_XMAHOL ( .B(RANGE2),
     .Y(N00AEQE), .A(RANGE1), .C(RANGE0));
nor3 nor3_XMAHJN_XMAHJO_XMAHJP_XMAHJS_XMAHJQ_XMAHJR ( .B(DIVQ0),
     .Y(N00AEOY), .A(DIVQ1), .C(DIVQ2));
nor3 nor3_XMAFOC_XMAFOD_XMAFOE_XMAFOH_XMAFOG_XMAFOF ( .B(N00ADWV),
     .Y(N00ADWX), .A(N00ADRR), .C(N00ADWN));
nor3 nor3_XMAFMZ_XMAFNA_XMAFNB_XMAFNE_XMAFND_XMAFNC ( .B(N00ADWK),
     .Y(N00ADWM), .A(N00ADRR), .C(N00ADWN));
txgate xfer_XMAHWH_XMAHWS ( .in(N00AEUF), .out(N00AEUG), .pp(N00AEUC),
     .nn(N00AESV));
txgate xfer_XMAHUZ_XMAHVK ( .in(N00AETP), .out(N00AETQ), .pp(N00AETM),
     .nn(N00AESU));
txgate xfer_XMAHTR_XMAHUC ( .in(N00AESZ), .out(N00AETA), .pp(N00AEQL),
     .nn(N00AESW));
txgate xfer_XMAHSV_XMAHTF ( .in(N00AESR), .out(N00AESN), .pp(N00AEQL),
     .nn(N00AERB));
txgate xfer_XMAHSS_XMAHSZ ( .in(N00AESQ), .out(N00AEQQ), .pp(N00AEQP),
     .nn(N00AEQL));
txgate xfer_XMAHRO_XMAHSB ( .in(N00AERX), .out(N00AERY), .pp(N00AERT),
     .nn(N00AEQO));
txgate xfer_XMAHPZ_XMAHQK ( .in(N00AERG), .out(N00AERH), .pp(N00AERD),
     .nn(N00AEQN));
txgate xfer_XMAHPO_XMAHPP ( .in(DIVR3), .out(DIVR3), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAHPM_XMAHPN ( .in(DIVR2), .out(DIVR2), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAHPK_XMAHPL ( .in(DIVR1), .out(DIVR1), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAHPI_XMAHPJ ( .in(DIVR0), .out(DIVR0), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAHGW_XMAHHH ( .in(N00AEOC), .out(N00AEOD), .pp(N00AEJV),
     .nn(N00AEJU));
txgate xfer_XMAHFT_XMAHGQ ( .in(N00AENO), .out(N00AEJY), .pp(N00AENS),
     .nn(N00AENV));
txgate xfer_XMAHFR_XMAHGO ( .in(N00AENQ), .out(N00AENR), .pp(N00AEJV),
     .nn(N00AEJU));
txgate xfer_XMAHFH_XMAHGE ( .in(N00AENO), .out(N00AEJX), .pp(N00AENV),
     .nn(N00AENS));
txgate xfer_XMAHEF_XMAHFC ( .in(N00AENC), .out(N00AEJZ), .pp(N00AENG),
     .nn(N00AEMZ));
txgate xfer_XMAHED_XMAHFA ( .in(N00AENE), .out(N00AENF), .pp(N00AEJV),
     .nn(N00AEJU));
txgate xfer_XMAHDT_XMAHEQ ( .in(N00AENC), .out(N00AEJX), .pp(N00AEMZ),
     .nn(N00AENG));
txgate xfer_XMAHDB_XMAHDC ( .in(DIVQ0), .out(DIVQ0), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAHCZ_XMAHDA ( .in(DIVQ1), .out(DIVQ1), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAHCX_XMAHCY ( .in(DIVQ2), .out(DIVQ2), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAHAV_XMAHBS ( .in(N00AEMI), .out(N00AEMH), .pp(N00AEMM),
     .nn(N00AEMG));
txgate xfer_XMAHAT_XMAHBQ ( .in(N00AEMK), .out(N00AEML), .pp(N00AEKA),
     .nn(N00AEKB));
txgate xfer_XMAHAJ_XMAHBG ( .in(N00AEMI), .out(N00AEJZ), .pp(N00AEMG),
     .nn(N00AEMM));
txgate xfer_XMAGYP_XMAGZM ( .in(N00AELR), .out(N00AELQ), .pp(N00AELV),
     .nn(N00AELP));
txgate xfer_XMAGYN_XMAGZK ( .in(N00AELT), .out(N00AELU), .pp(N00AEKA),
     .nn(N00AEKB));
txgate xfer_XMAGYD_XMAGZA ( .in(N00AELR), .out(N00AEKE), .pp(N00AELP),
     .nn(N00AELV));
txgate xfer_XMAGWJ_XMAGXG ( .in(N00AELB), .out(N00AELA), .pp(N00AELF),
     .nn(N00AEKZ));
txgate xfer_XMAGWH_XMAGXE ( .in(N00AELD), .out(N00AELE), .pp(N00AEKA),
     .nn(N00AEKB));
txgate xfer_XMAGVX_XMAGWU ( .in(N00AELB), .out(N00AEKD), .pp(N00AEKZ),
     .nn(N00AELF));
txgate xfer_XMAGUD_XMAGVA ( .in(N00AEKL), .out(N00AEKK), .pp(N00AEKP),
     .nn(N00AEKJ));
txgate xfer_XMAGUB_XMAGUY ( .in(N00AEKN), .out(N00AEKO), .pp(N00AEKA),
     .nn(N00AEKB));
txgate xfer_XMAGTR_XMAGUO ( .in(N00AEKL), .out(N00AEKC), .pp(N00AEKJ),
     .nn(N00AEKP));
txgate xfer_XMAGSI_XMAGSJ ( .in(BYPASS), .out(BYPASS), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAGSG_XMAGSH ( .in(RESET), .out(RESET), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAGKY_XMAGLJ ( .in(N00AEGZ), .out(N00AEHA), .pp(N00AEGW),
     .nn(N00AEFP));
txgate xfer_XMAGJQ_XMAGKB ( .in(N00AEGJ), .out(N00AEGK), .pp(N00AEGG),
     .nn(N00AEFO));
txgate xfer_XMAGII_XMAGIT ( .in(N00AEFT), .out(N00AEFU), .pp(N00ADZO),
     .nn(N00AEFQ));
txgate xfer_XMAGHM_XMAGHW ( .in(N00AEFL), .out(N00AEFH), .pp(N00ADZO),
     .nn(N00AEAF));
txgate xfer_XMAGHJ_XMAGHQ ( .in(N00AEFK), .out(N00ADZV), .pp(N00ADZU),
     .nn(N00ADZO));
txgate xfer_XMAGGF_XMAGGS ( .in(N00AEER), .out(N00AEES), .pp(N00AEEN),
     .nn(N00ADZT));
txgate xfer_XMAGEQ_XMAGFB ( .in(N00AEEA), .out(N00AEEB), .pp(N00AEDX),
     .nn(N00ADZS));
txgate xfer_XMAGAZ_XMAGBK ( .in(N00AECS), .out(N00AECT), .pp(N00AECP),
     .nn(N00AEBI));
txgate xfer_XMAFZR_XMAGAC ( .in(N00AECC), .out(N00AECD), .pp(N00AEBZ),
     .nn(N00AEBH));
txgate xfer_XMAFYJ_XMAFYU ( .in(N00AEBM), .out(N00AEBN), .pp(N00AEAX),
     .nn(N00AEBJ));
txgate xfer_XMAFWD_XMAFWE ( .in(DIVF6), .out(DIVF6), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFWB_XMAFWC ( .in(DIVF5), .out(DIVF5), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFVZ_XMAFWA ( .in(DIVF4), .out(DIVF4), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFVX_XMAFVY ( .in(DIVF3), .out(DIVF3), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFVV_XMAFVW ( .in(DIVF2), .out(DIVF2), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFVT_XMAFVU ( .in(DIVF1), .out(DIVF1), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFVR_XMAFVS ( .in(DIVF0), .out(DIVF0), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFOQ_XMAFOR ( .in(RANGE0), .out(RANGE0), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFOO_XMAFOP ( .in(RANGE1), .out(RANGE1), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFOM_XMAFON ( .in(RANGE2), .out(RANGE2), .pp(vdd_),
     .nn(gnd_));
txgate xfer_XMAFJK_XMAFJU ( .in(N00ADUT), .out(N00ADUS), .pp(gnd_),
     .nn(vdd_));
txgate xfer_XMAFHR_XMAFIA ( .in(N00ADUI), .out(N00ADUF), .pp(N00ADUB),
     .nn(N00ADTZ));
txgate xfer_XMAFHM_XMAFHX ( .in(N00ADUE), .out(N00ADUH), .pp(N00ADTZ),
     .nn(N00ADUB));
txgate xfer_XMAFGP_XMAFGY ( .in(N00ADUB), .out(N00ADTX), .pp(N00ADTT),
     .nn(N00ADTR));
txgate xfer_XMAFGK_XMAFGV ( .in(N00ADTW), .out(N00ADUA), .pp(N00ADTR),
     .nn(N00ADTT));
txgate xfer_XMAFFN_XMAFFW ( .in(N00ADTT), .out(N00ADTP), .pp(N00ADTL),
     .nn(N00ADTJ));
txgate xfer_XMAFFI_XMAFFT ( .in(N00ADTO), .out(N00ADTS), .pp(N00ADTJ),
     .nn(N00ADTL));
txgate xfer_XMAFEL_XMAFEU ( .in(N00ADTL), .out(N00ADTH), .pp(N00ADTD),
     .nn(N00ADTB));
txgate xfer_XMAFEG_XMAFER ( .in(N00ADTG), .out(N00ADTK), .pp(N00ADTB),
     .nn(N00ADTD));
txgate xfer_XMAFDJ_XMAFDS ( .in(N00ADTD), .out(N00ADSZ), .pp(N00ADSV),
     .nn(N00ADST));
txgate xfer_XMAFDE_XMAFDP ( .in(N00ADSY), .out(N00ADTC), .pp(N00ADST),
     .nn(N00ADSV));
txgate xfer_XMAFCH_XMAFCQ ( .in(N00ADSV), .out(N00ADSR), .pp(N00ADSK),
     .nn(N00ADSI));
txgate xfer_XMAFCC_XMAFCN ( .in(N00ADSQ), .out(N00ADSU), .pp(N00ADSI),
     .nn(N00ADSK));
txgate xfer_XMAFBF_XMAFBO ( .in(N00ADSK), .out(N00ADSG), .pp(N00ADSM),
     .nn(N00ADSP));
txgate xfer_XMAFBA_XMAFBL ( .in(N00ADSF), .out(N00ADSJ), .pp(N00ADSP),
     .nn(N00ADSM));
txgate xfer_XMAEXL_XMAEXM ( .in(REF), .out(REF), .pp(vdd_), .nn(gnd_));
txgate xfer_XMAEXJ_XMAEXK ( .in(FB), .out(FB), .pp(vdd_), .nn(gnd_));
txgate xfer_XMAEXH_XMAEXI ( .in(FSE), .out(FSE), .pp(vdd_), .nn(gnd_));
nand2 nand2_XMAIAW_XMAIAX_XMAIAV_XMAIAU ( .A(N00AEQM), .Y(N00AERS),
     .B(DIVR3));
nand2 nand2_XMAIAS_XMAIAT_XMAIAR_XMAIAQ ( .A(N00AEQU), .Y(N00AEQS),
     .B(N00AEQV));
nand2 nand2_XMAIAO_XMAIAP_XMAIAN_XMAIAM ( .A(N00AERC), .Y(N00AERB),
     .B(N00AEVW));
nand2 nand2_XMAIAK_XMAIAL_XMAIAJ_XMAIAI ( .A(N00AEQR), .Y(N00AEVT),
     .B(N00AEVS));
nand2 nand2_XMAHYM_XMAHYN_XMAHYL_XMAHYK ( .A(N00AEQU), .Y(N00AEQY),
     .B(N00AEVC));
nand2 nand2_XMAHXW_XMAHXX_XMAHXV_XMAHXU ( .A(N00AEQM), .Y(N00AETL),
     .B(DIVR0));
nand2 nand2_XMAHXS_XMAHXT_XMAHXR_XMAHXQ ( .A(N00AEQM), .Y(N00AEUB),
     .B(DIVR1));
nand2 nand2_XMAHXO_XMAHXP_XMAHXN_XMAHXM ( .A(N00AEQM), .Y(N00AEUR),
     .B(DIVR2));
nand2 nand2_XMAHXK_XMAHXL_XMAHXJ_XMAHXI ( .A(N00AEQT), .Y(N00AESU),
     .B(N00AEQL));
nand2 nand2_XMAHMT_XMAHMU_XMAHMN_XMAHMO ( .A(N00AEPO), .Y(N00AEPS),
     .B(N00AEPP));
nand2 nand2_XMAHLN_XMAHLO_XMAHLM_XMAHLL ( .A(N00AEPM), .Y(N00AEPO),
     .B(N00AEJP));
nand2 nand2_XMAHLJ_XMAHLK_XMAHLI_XMAHLH ( .A(N00AEPN), .Y(N00AEPP),
     .B(N00AEJS));
nand2 nand2_XMAHKX_XMAHKY_XMAHKT_XMAHKU ( .A(N00AEPE), .Y(N00AEJP),
     .B(N00AEPD));
nand2 nand2_XMAHKR_XMAHKS_XMAHKQ_XMAHKP ( .A(REF), .Y(N00AEPE),
     .B(N00AEPH));
nand2 nand2_XMAHKN_XMAHKO_XMAHKM_XMAHKL ( .A(N00AEJR), .Y(N00AEPD),
     .B(N00AEPF));
nand2 nand2_XMAHIT_XMAHIU_XMAHIS_XMAHIR ( .A(N00AEOM), .Y(N00AEOR),
     .B(DIVQ0));
nand2 nand2_XMAHIP_XMAHIQ_XMAHIO_XMAHIN ( .A(DIVQ0), .Y(N00AEOT),
     .B(DIVQ1));
nand2 nand2_XMAHIL_XMAHIM_XMAHIK_XMAHIJ ( .A(N00AEJX), .Y(N00AENB),
     .B(N00AEOR));
nand2 nand2_XMAHIH_XMAHII_XMAHIC_XMAHHZ ( .A(N00AEJS), .Y(N00AEJU),
     .B(N00AEOO));
nand2 nand2_XMAHCV_XMAHCW_XMAHCQ_XMAHCN ( .A(N00AEJX), .Y(N00AEKA),
     .B(N00AEMZ));
nand2 nand2_XMAGQT_XMAGQU_XMAGQS_XMAGQR ( .A(N00AEIH), .Y(N00AEDQ),
     .B(N00ADZR));
nand2 nand2_XMAGQP_XMAGQQ_XMAGQO_XMAGQN ( .A(N00ADZR), .Y(N00AEFE),
     .B(DIVF4));
nand2 nand2_XMAGQL_XMAGQM_XMAGQK_XMAGQJ ( .A(N00ADZR), .Y(N00AEEM),
     .B(DIVF3));
nand2 nand2_XMAGQH_XMAGQI_XMAGQG_XMAGQF ( .A(N00ADZZ), .Y(N00AEIV),
     .B(N00AEAA));
nand2 nand2_XMAGQD_XMAGQE_XMAGQC_XMAGQB ( .A(N00AEAG), .Y(N00AEAF),
     .B(N00AEJB));
nand2 nand2_XMAGPZ_XMAGQA_XMAGPY_XMAGPX ( .A(N00ADZW), .Y(N00AEIY),
     .B(N00AEIX));
nand2 nand2_XMAGND_XMAGNE_XMAGNC_XMAGNB ( .A(N00ADZZ), .Y(N00AEHW),
     .B(N00AEAD));
nand2 nand2_XMAGMN_XMAGMO_XMAGMM_XMAGML ( .A(N00ADZR), .Y(N00AEGF),
     .B(DIVF0));
nand2 nand2_XMAGMJ_XMAGMK_XMAGMI_XMAGMH ( .A(N00ADZR), .Y(N00AEGV),
     .B(DIVF1));
nand2 nand2_XMAGMF_XMAGMG_XMAGME_XMAGMD ( .A(N00ADZR), .Y(N00AEHL),
     .B(DIVF2));
nand2 nand2_XMAGMB_XMAGMC_XMAGMA_XMAGLZ ( .A(N00ADZY), .Y(N00AEFO),
     .B(N00ADZO));
nand2 nand2_XMAGDY_XMAGDZ_XMAGDX_XMAGDW ( .A(N00AEAT), .Y(N00AEAY),
     .B(N00AEBD));
nand2 nand2_XMAGDU_XMAGDV_XMAGDT_XMAGDS ( .A(N00AEAO), .Y(N00AEAS),
     .B(N00AEBD));
nand2 nand2_XMAGDQ_XMAGDR_XMAGDP_XMAGDO ( .A(N00AEDQ), .Y(N00AEAN),
     .B(N00ADZQ));
nand2 nand2_XMAGCO_XMAGCP_XMAGCN_XMAGCM ( .A(N00AEBD), .Y(N00AEBY),
     .B(DIVF5));
nand2 nand2_XMAGCK_XMAGCL_XMAGCJ_XMAGCI ( .A(N00AEBD), .Y(N00AECO),
     .B(DIVF6));
nand2 nand2_XMAGCC_XMAGCD_XMAGCB_XMAGCA ( .A(N00AEAU), .Y(N00AEBH),
     .B(N00AEAX));
nand2 nand2_XMAFXX_XMAFXY_XMAFXO_XMAFXP ( .A(N00AEBA), .Y(N00AEAX),
     .B(N00AEAS));
nand2 nand2_XMAFQF_XMAFQG_XMAFQE_XMAFQD ( .A(N00ADXW), .Y(N00ADXZ),
     .B(RANGE1));
nand2 nand2_XMAFQB_XMAFQC_XMAFQA_XMAFPZ ( .A(RANGE2), .Y(N00ADYB),
     .B(RANGE0));
nand2 nand2_XMAFPX_XMAFPY_XMAFPW_XMAFPV ( .A(N00ADYB), .Y(N00ADYA),
     .B(N00ADXZ));
nand2 nand2_XMAFPT_XMAFPU_XMAFPS_XMAFPR ( .A(RANGE2), .Y(N00ADXT),
     .B(RANGE1));
nand2 nand2_XMAFIR_XMAFIS_XMAFIQ_XMAFIP ( .A(N00ADUL), .Y(N00ADSN),
     .B(N00ADUO));
nand2 nand2_XMAFIN_XMAFIO_XMAFIM_XMAFIL ( .A(N00ADUO), .Y(N00ADUN),
     .B(N00ADUI));
nand2 nand2_XMAFAR_XMAFAS_XMAFAQ_XMAFAP ( .A(N00ADRP), .Y(N00ADRM),
     .B(N00ADSE));
nand2 nand2_XMAEZD_XMAEZE_XMAEZC_XMAEZB ( .A(N00ADQU), .Y(N00ADQR),
     .B(N00ADRJ));
nand3 Inand3_mahsh_i_j_k_l_m ( .Y(N00AERU), .B(N00AEQR), .C(N00AESK),
     .A(vdd_));
nand3 nand3_XMAIBV_XMAIBW_XMAIBX_XMAIBS_XMAIBT_XMAIBU ( .Y(N00AEVN),
     .B(N00AEVK), .C(N00AEQW), .A(N00AEQV));
nand3 nand3_XMAHYH_XMAHYI_XMAHYJ_XMAHYE_XMAHYF_XMAHYG ( .Y(N00AEUY),
     .B(N00AEQW), .C(N00AEQV), .A(N00AEQU));
nand3 nand3_XMAHYB_XMAHYC_XMAHYD_XMAHXY_XMAHXZ_XMAHYA ( .Y(N00AESV),
     .B(N00AEQT), .C(N00AEQL), .A(N00AEQU));
nand3 nand3_XMAHIY_XMAHIZ_XMAHJA_XMAHIV_XMAHIW_XMAHIX ( .Y(N00AEMZ),
     .B(N00AEJT), .C(N00AEMW), .A(N00AEOT));
nand3 nand3_XMAGRO_XMAGRP_XMAGRQ_XMAGRL_XMAGRM_XMAGRN ( .Y(N00AEIR),
     .B(N00AEIO), .C(N00AEAB), .A(N00AEAA));
nand3 nand3_XMAGMY_XMAGMZ_XMAGNA_XMAGMV_XMAGMW_XMAGMX ( .Y(N00AEHS),
     .B(N00AEAB), .C(N00AEAA), .A(N00ADZZ));
nand3 nand3_XMAGMS_XMAGMT_XMAGMU_XMAGMP_XMAGMQ_XMAGMR ( .Y(N00AEFP),
     .B(N00ADZY), .C(N00ADZO), .A(N00ADZZ));
nand3 nand3_XMAGLW_XMAGLX_XMAGLY_XMAGLT_XMAGLU_XMAGLV ( .Y(N00AEGX),
     .B(N00ADZP), .C(N00ADZQ), .A(N00AEHL));
nand3 nand3_XMAGKO_XMAGKP_XMAGKQ_XMAGKL_XMAGKM_XMAGKN ( .Y(N00AEGH),
     .B(N00ADZP), .C(N00ADZQ), .A(N00AEGV));
nand3 nand3_XMAGJG_XMAGJH_XMAGJI_XMAGJD_XMAGJE_XMAGJF ( .Y(N00AEFR),
     .B(N00ADZP), .C(N00ADZQ), .A(N00AEGF));
nand3 nand3_XMAGHB_XMAGHC_XMAGHD_XMAGGY_XMAGGZ_XMAGHA ( .Y(N00AEEO),
     .B(N00ADZP), .C(N00ADZQ), .A(N00AEFE));
nand3 nand3_XMAGFO_XMAGFP_XMAGFQ_XMAGFL_XMAGFM_XMAGFN ( .Y(N00AEDY),
     .B(N00ADZP), .C(N00ADZQ), .A(N00AEEM));
nand3 nand3_XMAGEG_XMAGEH_XMAGEI_XMAGEA_XMAGEC_XMAGEE ( .Y(N00AEAT),
     .B(N00AEAU), .C(N00AEAV), .A(N00AEAW));
nand3 nand3_XMAGCT_XMAGCU_XMAGCV_XMAGCQ_XMAGCR_XMAGCS ( .Y(N00AEBI),
     .B(N00AEAU), .C(N00AEAX), .A(N00AEAV));
nand3 i_nand3_mahxc_d_e_f_g_h ( .Y(N00AEUD), .B(N00AEQR), .C(N00AEUR),
     .A(vdd_));
nand3 I_nand3_mahqu_v_w_x_y_z ( .Y(N00AERE), .B(vdd_), .C(N00AERS),
     .A(N00AEQR));
inv inv_XMAIAG_XMAIAH ( .A(N00AEVT), .Y(N00AEQZ));
inv inv_XMAIAE_XMAIAF ( .A(N00ADRR), .Y(N00AEQM));
inv inv_XMAIAC_XMAIAD ( .A(N00AEVD), .Y(N00AEVS));
inv inv_XMAIAA_XMAIAB ( .A(N00AEQL), .Y(N00AEQP));
inv inv_XMAHZY_XMAHZZ ( .A(N00AERA), .Y(N00ADSE));
inv inv_XMAHZW_XMAHZX ( .A(N00AERB), .Y(N00AEQL));
inv inv_XMAHZU_XMAHZV ( .A(N00ADQL), .Y(N00AERC));
inv inv_XMAHZS_XMAHZT ( .A(N00AEUY), .Y(N00AEVR));
inv inv_XMAHZQ_XMAHZR ( .A(N00AEQS), .Y(N00AEVQ));
inv inv_XMAHXA_XMAHXB ( .A(N00AESV), .Y(N00AEUC));
inv inv_XMAHWM_XMAHWR ( .A(N00AEUG), .Y(N00AEQV));
inv inv_XMAHWF_XMAHWQ ( .A(N00AEUE), .Y(N00AEUF));
inv inv_XMAHVS_XMAHVT ( .A(N00AESU), .Y(N00AETM));
inv inv_XMAHVE_XMAHVJ ( .A(N00AETQ), .Y(N00AEQU));
inv inv_XMAHUX_XMAHVI ( .A(N00AETO), .Y(N00AETP));
inv inv_XMAHUK_XMAHUL ( .A(N00AEQL), .Y(N00AESW));
inv inv_XMAHTW_XMAHUB ( .A(N00AETA), .Y(N00AEQT));
inv inv_XMAHTP_XMAHUA ( .A(N00AESY), .Y(N00AESZ));
inv inv_XMAHSX_XMAHTH ( .A(N00AESQ), .Y(N00AESR));
inv inv_XMAHST_XMAHTG ( .A(N00AESN), .Y(N00AEQR));
inv inv_XMAHSP_XMAHSY ( .A(N00AEQM), .Y(N00AESO));
inv inv_XMAHSF_XMAHSG ( .A(N00AEQO), .Y(N00AERT));
inv inv_XMAHRS_XMAHRT ( .A(N00AEQX), .Y(N00AESD));
inv inv_XMAHRR_XMAHSE ( .A(N00AERW), .Y(N00AERX));
inv inv_XMAHRQ_XMAHSD ( .A(N00AERV), .Y(N00AERW));
inv inv_XMAHRJ_XMAHSC ( .A(N00AERY), .Y(N00AEQX));
inv inv_XMAHQS_XMAHQT ( .A(N00AEQN), .Y(N00AERD));
inv inv_XMAHQE_XMAHQJ ( .A(N00AERH), .Y(N00AEQW));
inv inv_XMAHPX_XMAHQI ( .A(N00AERF), .Y(N00AERG));
inv inv_XMAHNP_XMAHNQ ( .A(RESET), .Y(N00AEQD));
inv inv_XMAHNN_XMAHNO ( .A(N00AEJS), .Y(N00AEJQ));
inv inv_XMAHNL_XMAHNM ( .A(N00AEOY), .Y(N00AEQC));
inv inv_XMAHNJ_XMAHNK ( .A(N00AEQB), .Y(N00AEPG));
inv inv_XMAHNH_XMAHNI ( .A(N00AEJQ), .Y(N00ADRD));
inv inv_XMAHNF_XMAHNG ( .A(N00AEQA), .Y(N00ADRR));
inv inv_XMAHMS_XMAHMW ( .A(N00AEPT), .Y(PLLOUT));
inv inv_XMAHMR_XMAHMV ( .A(N00AEPS), .Y(N00AEPT));
inv inv_XMAHJX_XMAHJY ( .A(N00AEPF), .Y(N00AEPH));
inv inv_XMAHJV_XMAHJW ( .A(N00AEPG), .Y(N00AEPF));
inv inv_XMAHHX_XMAHHY ( .A(N00AEOM), .Y(N00AENV));
inv inv_XMAHHV_XMAHHW ( .A(DIVQ2), .Y(N00AEMW));
inv inv_XMAHHT_XMAHHU ( .A(RESET), .Y(N00AEJT));
inv inv_XMAHHR_XMAHHS ( .A(N00AEJT), .Y(N00AEJW));
inv inv_XMAHHP_XMAHHQ ( .A(N00AEJU), .Y(N00AEJV));
inv inv_XMAHHB_XMAHHG ( .A(N00AEOD), .Y(N00AEJY));
inv inv_XMAHGU_XMAHHF ( .A(N00AEOB), .Y(N00AEOC));
inv inv_XMAHFS_XMAHGP ( .A(N00AENP), .Y(N00AENQ));
inv inv_XMAHFN_XMAHGF ( .A(N00AENR), .Y(N00AEJX));
inv inv_XMAHFJ_XMAHGG ( .A(N00AENV), .Y(N00AENS));
inv inv_XMAHEE_XMAHFB ( .A(N00AEND), .Y(N00AENE));
inv inv_XMAHDZ_XMAHER ( .A(N00AENF), .Y(N00AEJR));
inv inv_XMAHDV_XMAHET ( .A(N00AEMZ), .Y(N00AENG));
inv inv_XMAHCL_XMAHCM ( .A(N00AEKA), .Y(N00AEKB));
inv inv_XMAHCJ_XMAHCK ( .A(N00AEJW), .Y(N00AEKI));
inv inv_XMAHCF_XMAHCG ( .A(N00AEJZ), .Y(N00AEMH));
inv inv_XMAHCD_XMAHCE ( .A(N00AEMG), .Y(N00AEMU));
inv inv_XMAHAU_XMAHBR ( .A(N00AEMJ), .Y(N00AEMK));
inv inv_XMAHAP_XMAHBH ( .A(N00AEML), .Y(N00AEJZ));
inv inv_XMAHAL_XMAHBI ( .A(N00AEMG), .Y(N00AEMM));
inv inv_XMAGZZ_XMAHAA ( .A(N00AEKE), .Y(N00AELQ));
inv inv_XMAGZX_XMAGZY ( .A(N00AELP), .Y(N00AEKG));
inv inv_XMAGYO_XMAGZL ( .A(N00AELS), .Y(N00AELT));
inv inv_XMAGYJ_XMAGZB ( .A(N00AELU), .Y(N00AEKE));
inv inv_XMAGYF_XMAGZC ( .A(N00AELP), .Y(N00AELV));
inv inv_XMAGXT_XMAGXU ( .A(N00AEKD), .Y(N00AELA));
inv inv_XMAGXR_XMAGXS ( .A(N00AEKZ), .Y(N00AEKF));
inv inv_XMAGWI_XMAGXF ( .A(N00AELC), .Y(N00AELD));
inv inv_XMAGWD_XMAGWV ( .A(N00AELE), .Y(N00AEKD));
inv inv_XMAGVZ_XMAGWW ( .A(N00AEKZ), .Y(N00AELF));
inv inv_XMAGVN_XMAGVO ( .A(N00AEKC), .Y(N00AEKK));
inv inv_XMAGVL_XMAGVM ( .A(N00AEKJ), .Y(N00AEKH));
inv inv_XMAGUC_XMAGUZ ( .A(N00AEKM), .Y(N00AEKN));
inv inv_XMAGTX_XMAGUP ( .A(N00AEKO), .Y(N00AEKC));
inv inv_XMAGTT_XMAGUQ ( .A(N00AEKJ), .Y(N00AEKP));
inv inv_XMAGPV_XMAGPW ( .A(N00AEIY), .Y(N00AEAE));
inv inv_XMAGPT_XMAGPU ( .A(N00ADRR), .Y(N00ADZR));
inv inv_XMAGPR_XMAGPS ( .A(N00AEHX), .Y(N00AEIH));
inv inv_XMAGPP_XMAGPQ ( .A(N00AEIC), .Y(N00AEIX));
inv inv_XMAGPN_XMAGPO ( .A(N00ADZW), .Y(N00AEAH));
inv inv_XMAGPL_XMAGPM ( .A(N00AEAH), .Y(N00ADZP));
inv inv_XMAGPJ_XMAGPK ( .A(N00ADZO), .Y(N00ADZU));
inv inv_XMAGPH_XMAGPI ( .A(N00AEAF), .Y(N00ADZO));
inv inv_XMAGPF_XMAGPG ( .A(N00ADQN), .Y(N00AEAG));
inv inv_XMAGPD_XMAGPE ( .A(N00AEHS), .Y(N00AEIW));
inv inv_XMAGPB_XMAGPC ( .A(N00AEIV), .Y(N00AEIU));
inv inv_XMAGLR_XMAGLS ( .A(N00AEFP), .Y(N00AEGW));
inv inv_XMAGLD_XMAGLI ( .A(N00AEHA), .Y(N00AEAA));
inv inv_XMAGKW_XMAGLH ( .A(N00AEGY), .Y(N00AEGZ));
inv inv_XMAGKJ_XMAGKK ( .A(N00AEFO), .Y(N00AEGG));
inv inv_XMAGJV_XMAGKA ( .A(N00AEGK), .Y(N00ADZZ));
inv inv_XMAGJO_XMAGJZ ( .A(N00AEGI), .Y(N00AEGJ));
inv inv_XMAGJB_XMAGJC ( .A(N00ADZO), .Y(N00AEFQ));
inv inv_XMAGIN_XMAGIS ( .A(N00AEFU), .Y(N00ADZY));
inv inv_XMAGIG_XMAGIR ( .A(N00AEFS), .Y(N00AEFT));
inv inv_XMAGHO_XMAGHY ( .A(N00AEFK), .Y(N00AEFL));
inv inv_XMAGHK_XMAGHX ( .A(N00AEFH), .Y(N00ADZW));
inv inv_XMAGHG_XMAGHP ( .A(N00ADZR), .Y(N00AEFI));
inv inv_XMAGGW_XMAGGX ( .A(N00ADZT), .Y(N00AEEN));
inv inv_XMAGGJ_XMAGGK ( .A(N00AEAC), .Y(N00AEEX));
inv inv_XMAGGI_XMAGGV ( .A(N00AEEQ), .Y(N00AEER));
inv inv_XMAGGH_XMAGGU ( .A(N00AEEP), .Y(N00AEEQ));
inv inv_XMAGGA_XMAGGT ( .A(N00AEES), .Y(N00AEAC));
inv inv_XMAGFJ_XMAGFK ( .A(N00ADZS), .Y(N00AEDX));
inv inv_XMAGEV_XMAGFA ( .A(N00AEEB), .Y(N00AEAB));
inv inv_XMAGEO_XMAGEZ ( .A(N00AEDZ), .Y(N00AEEA));
inv inv_XMAGDM_XMAGDN ( .A(N00ADRR), .Y(N00AEBD));
inv inv_XMAGDK_XMAGDL ( .A(N00AEAY), .Y(N00AEAZ));
inv inv_XMAGDI_XMAGDJ ( .A(N00AEDO), .Y(N00AEAL));
inv inv_XMAGDG_XMAGDH ( .A(N00AEAZ), .Y(N00ADZQ));
inv inv_XMAGDE_XMAGDF ( .A(N00AEAX), .Y(N00AEDO));
inv inv_XMAGBS_XMAGBT ( .A(N00AEBI), .Y(N00AECP));
inv inv_XMAGBE_XMAGBJ ( .A(N00AECT), .Y(N00AEAW));
inv inv_XMAGAX_XMAGBI ( .A(N00AECR), .Y(N00AECS));
inv inv_XMAGAK_XMAGAL ( .A(N00AEBH), .Y(N00AEBZ));
inv inv_XMAFZW_XMAGAB ( .A(N00AECD), .Y(N00AEAV));
inv inv_XMAFZP_XMAGAA ( .A(N00AECB), .Y(N00AECC));
inv inv_XMAFZC_XMAFZD ( .A(N00AEAX), .Y(N00AEBJ));
inv inv_XMAFYO_XMAFYT ( .A(N00AEBN), .Y(N00AEAU));
inv inv_XMAFYH_XMAFYS ( .A(N00AEBL), .Y(N00AEBM));
inv inv_XMAFWQ_XMAFWY ( .A(N00AEAI), .Y(N00AEAJ));
inv inv_XMAFWP_XMAFWV ( .A(N00AEAK), .Y(N00AEAO));
inv inv_XMAFWO_XMAFWU ( .A(N00AEAO), .Y(N00AEAK));
inv inv_XMAFWK_XMAFWW ( .A(N00AEAJ), .Y(N00AEAI));
inv inv_XMAFPP_XMAFPQ ( .A(RANGE2), .Y(N00ADXW));
inv inv_XMAFPN_XMAFPO ( .A(RANGE1), .Y(N00ADXV));
inv inv_XMAFPL_XMAFPM ( .A(RANGE2), .Y(N00ADXU));
inv inv_XMAFPJ_XMAFPK ( .A(N00ADXT), .Y(N00ADXS));
inv inv_XMAFPH_XMAFPI ( .A(N00ADXQ), .Y(N00ADXR));
inv inv_XMAFPF_XMAFPG ( .A(RANGE0), .Y(N00ADXQ));
inv inv_XMAFKV_XMAFLV ( .A(N00ADVL), .Y(N00ADVJ));
inv inv_XMAFKR_XMAFLS ( .A(N00ADVI), .Y(N00ADVH));
inv inv_XMAFKQ_XMAFLR ( .A(N00ADVK), .Y(N00ADVI));
inv inv_XMAFJN_XMAFJY ( .A(N00ADRR), .Y(N00ADVB));
inv inv_XMAFJJ_XMAFJT ( .A(N00ADVA), .Y(N00ADUO));
inv inv_XMAFJG_XMAFJR ( .A(N00ADUZ), .Y(N00ADVA));
inv inv_XMAFJF_XMAFJQ ( .A(N00ADUY), .Y(N00ADUZ));
inv inv_XMAFJE_XMAFJP ( .A(N00ADUW), .Y(N00ADUY));
inv inv_XMAFJC_XMAFJO ( .A(N00ADUT), .Y(N00ADUW));
inv inv_XMAFIJ_XMAFIK ( .A(N00ADSP), .Y(N00ADSM));
inv inv_XMAFIH_XMAFII ( .A(N00ADRR), .Y(N00ADUL));
inv inv_XMAFIB_XMAFIC ( .A(LOCK), .Y(N00ADUI));
inv inv_XMAFHH_XMAFHT ( .A(N00ADUH), .Y(LOCK));
inv inv_XMAFHF_XMAFHS ( .A(N00ADUF), .Y(N00ADUE));
inv inv_XMAFGZ_XMAFHA ( .A(N00ADTZ), .Y(N00ADUB));
inv inv_XMAFGF_XMAFGR ( .A(N00ADUA), .Y(N00ADTZ));
inv inv_XMAFGD_XMAFGQ ( .A(N00ADTX), .Y(N00ADTW));
inv inv_XMAFFX_XMAFFY ( .A(N00ADTR), .Y(N00ADTT));
inv inv_XMAFFD_XMAFFP ( .A(N00ADTS), .Y(N00ADTR));
inv inv_XMAFFB_XMAFFO ( .A(N00ADTP), .Y(N00ADTO));
inv inv_XMAFEV_XMAFEW ( .A(N00ADTJ), .Y(N00ADTL));
inv inv_XMAFEB_XMAFEN ( .A(N00ADTK), .Y(N00ADTJ));
inv inv_XMAFDZ_XMAFEM ( .A(N00ADTH), .Y(N00ADTG));
inv inv_XMAFDT_XMAFDU ( .A(N00ADTB), .Y(N00ADTD));
inv inv_XMAFCZ_XMAFDL ( .A(N00ADTC), .Y(N00ADTB));
inv inv_XMAFCX_XMAFDK ( .A(N00ADSZ), .Y(N00ADSY));
inv inv_XMAFCR_XMAFCS ( .A(N00ADST), .Y(N00ADSV));
inv inv_XMAFBX_XMAFCJ ( .A(N00ADSU), .Y(N00ADST));
inv inv_XMAFBV_XMAFCI ( .A(N00ADSR), .Y(N00ADSQ));
inv inv_XMAFBP_XMAFBQ ( .A(N00ADSI), .Y(N00ADSK));
inv inv_XMAFAV_XMAFBH ( .A(N00ADSJ), .Y(N00ADSI));
inv inv_XMAFAT_XMAFBG ( .A(N00ADSG), .Y(N00ADSF));
inv inv_XMAFAN_XMAFAO ( .A(N00ADRQ), .Y(N00ADRZ));
inv inv_XMAFAD_XMAFAE ( .A(N00ADRK), .Y(N00ADQL));
inv inv_XMAEZP_XMAEZQ ( .A(N00ADRR), .Y(N00ADRQ));
inv inv_XMAEZN_XMAEZO ( .A(N00ADRL), .Y(N00ADRK));
inv inv_XMAEZL_XMAEZM ( .A(N00ADRM), .Y(N00ADQO));
inv inv_XMAEYZ_XMAEZA ( .A(N00ADQV), .Y(N00ADRE));
inv inv_XMAEYP_XMAEYQ ( .A(N00ADQP), .Y(N00ADQN));
inv inv_XMAEYB_XMAEYC ( .A(FSE), .Y(N00ADQV));
inv inv_XMAEXZ_XMAEYA ( .A(N00ADQQ), .Y(N00ADQP));
inv inv_XMAEXX_XMAEXY ( .A(N00ADQR), .Y(N00ADQM));
nor2 nor2_XMAICC_XMAICD_XMAICF_XMAICE ( .A(N00AEQR), .B(N00AEWG),
     .Y(N00AERA));
nor2 nor2_XMAIBY_XMAIBZ_XMAICB_XMAICA ( .A(DIVR0), .B(N00AEVS),
     .Y(N00AEWG));
nor2 nor2_XMAHZK_XMAHZL_XMAHZN_XMAHZP ( .A(N00AEVN), .B(N00AEQR),
     .Y(N00AEVC));
nor2 nor2_XMAHZE_XMAHZF_XMAHZH_XMAHZJ ( .A(N00AEQX), .B(N00AEQZ),
     .Y(N00AEVK));
nor2 nor2_XMAHYY_XMAHYZ_XMAHZB_XMAHZD ( .A(N00AEQT), .B(N00AEQY),
     .Y(N00AEQQ));
nor2 nor2_XMAHOD_XMAHOE_XMAHOG_XMAHOF ( .A(N00AEQD), .B(N00AEPG),
     .Y(N00AEPW));
nor2 nor2_XMAHNZ_XMAHOA_XMAHOC_XMAHOB ( .A(N00AEQC), .B(N00AEPG),
     .Y(N00AEPY));
nor2 nor2_XMAHNV_XMAHNW_XMAHNY_XMAHNX ( .A(N00AEPG), .B(RESET),
     .Y(N00AEQA));
nor2 nor2_XMAHNR_XMAHNS_XMAHNU_XMAHNT ( .A(BYPASS), .B(N00AEQE),
     .Y(N00AEQB));
nor2 nor2_XMAHNB_XMAHNC_XMAHNE_XMAHND ( .A(N00AEPY), .B(N00AEPW),
     .Y(N00AEPM));
nor2 nor2_XMAHMX_XMAHMY_XMAHNA_XMAHMZ ( .A(N00AEPM), .B(N00AEPW),
     .Y(N00AEPN));
nor2 nor2_XMAHJJ_XMAHJK_XMAHJM_XMAHJL ( .A(DIVQ2), .B(DIVQ1),
     .Y(N00AEOM));
nor2 nor2_XMAHJF_XMAHJG_XMAHJI_XMAHJH ( .A(RESET), .B(N00AEOY),
     .Y(N00AEOO));
nor2 nor2_XMAHJB_XMAHJC_XMAHJE_XMAHJD ( .A(DIVQ0), .B(DIVQ1),
     .Y(N00AEME));
nor2 nor2_XMAGOV_XMAGOW_XMAGOY_XMAGPA ( .A(N00AEIR), .B(N00ADZW),
     .Y(N00AEAD));
nor2 nor2_XMAGOP_XMAGOQ_XMAGOS_XMAGOU ( .A(N00AEAC), .B(N00AEAE),
     .Y(N00AEIO));
nor2 nor2_XMAGOJ_XMAGOK_XMAGOM_XMAGOO ( .A(N00ADZY), .B(N00AEHW),
     .Y(N00ADZV));
nor2 nor2_XMAFQL_XMAFQM_XMAFQO_XMAFQN ( .A(RANGE0), .B(N00ADXV),
     .Y(N00ADYF));
nor2 nor2_XMAFQH_XMAFQI_XMAFQK_XMAFQJ ( .A(N00ADYF), .B(N00ADXU),
     .Y(N00ADYE));
nor2 nor2_XMAFNW_XMAFNV_XMAFNY_XMAFNZ ( .A(N00ADWW), .B(N00ADWV),
     .Y(N00ADVK));
nor2 nor2_XMAFNR_XMAFNS_XMAFNU_XMAFNT ( .A(N00ADWW), .B(N00ADWX),
     .Y(N00ADWV));
nor2 nor2_XMAFNN_XMAFNO_XMAFNQ_XMAFNP ( .A(N00ADQO), .B(N00ADVK),
     .Y(N00ADWW));
nor2 nor2_XMAFMT_XMAFMS_XMAFMV_XMAFMW ( .A(N00ADWL), .B(N00ADWK),
     .Y(N00ADVL));
nor2 nor2_XMAFMO_XMAFMP_XMAFMR_XMAFMQ ( .A(N00ADWL), .B(N00ADWM),
     .Y(N00ADWK));
nor2 nor2_XMAFMK_XMAFML_XMAFMN_XMAFMM ( .A(N00ADQM), .B(N00ADVL),
     .Y(N00ADWL));
nor2 nor2_XMAFIT_XMAFIU_XMAFIW_XMAFIY ( .A(N00ADUN), .B(N00ADQO),
     .Y(N00ADSP));
diodN diod_XMAFJL ( .n2(gnd_), .n1(N00ADUV));
oneNodeN oneNodeXMAHPQ ( .n1(gnd_));
oneNodeN oneNodeXMAHLZ ( .n1(gnd_));
oneNodeN oneNodeXMAHLY ( .n1(gnd_));
oneNodeN oneNodeXMAHLX ( .n1(gnd_));
oneNodeN oneNodeXMAHLW ( .n1(gnd_));
oneNodeN oneNodeXMAHLU ( .n1(gnd_));
oneNodeN oneNodeXMAHLS ( .n1(gnd_));
oneNodeN oneNodeXMAHLR ( .n1(gnd_));
oneNodeN oneNodeXMAHLQ ( .n1(gnd_));
oneNodeN oneNodeXMAHLP ( .n1(gnd_));
oneNodeN oneNodeXMAHKZ ( .n1(gnd_));
oneNodeN oneNodeXMAHFY ( .n1(gnd_));
oneNodeN oneNodeXMAHFU ( .n1(gnd_));
oneNodeN oneNodeXMAHEK ( .n1(gnd_));
oneNodeN oneNodeXMAHDH ( .n1(gnd_));
oneNodeN oneNodeXMAHDG ( .n1(gnd_));
oneNodeN oneNodeXMAHDF ( .n1(gnd_));
oneNodeN oneNodeXMAHDE ( .n1(gnd_));
oneNodeN oneNodeXMAHBY ( .n1(gnd_));
oneNodeN oneNodeXMAHBA ( .n1(gnd_));
oneNodeN oneNodeXMAHAW ( .n1(gnd_));
oneNodeN oneNodeXMAGZS ( .n1(gnd_));
oneNodeN oneNodeXMAGYU ( .n1(gnd_));
oneNodeN oneNodeXMAGYQ ( .n1(gnd_));
oneNodeN oneNodeXMAGXM ( .n1(gnd_));
oneNodeN oneNodeXMAGWO ( .n1(gnd_));
oneNodeN oneNodeXMAGWK ( .n1(gnd_));
oneNodeN oneNodeXMAGVG ( .n1(gnd_));
oneNodeN oneNodeXMAGUI ( .n1(gnd_));
oneNodeN oneNodeXMAGUE ( .n1(gnd_));
oneNodeN oneNodeXMAGTH ( .n1(gnd_));
oneNodeN oneNodeXMAGTG ( .n1(gnd_));
oneNodeN oneNodeXMAGTF ( .n1(gnd_));
oneNodeN oneNodeXMAFWF ( .n1(gnd_));
oneNodeP oneNodeXMAHON ( .n1(vdd_));
oneNodeP oneNodeXMAHMK ( .n1(vdd_));
oneNodeP oneNodeXMAHMJ ( .n1(vdd_));
oneNodeP oneNodeXMAHMI ( .n1(vdd_));
oneNodeP oneNodeXMAHMH ( .n1(vdd_));
oneNodeP oneNodeXMAHMG ( .n1(vdd_));
oneNodeP oneNodeXMAHMF ( .n1(vdd_));
oneNodeP oneNodeXMAHME ( .n1(vdd_));
oneNodeP oneNodeXMAHMD ( .n1(vdd_));
oneNodeP oneNodeXMAHMB ( .n1(vdd_));
oneNodeP oneNodeXMAHKK ( .n1(vdd_));
oneNodeP oneNodeXMAHKI ( .n1(vdd_));
oneNodeP oneNodeXMAHKH ( .n1(vdd_));
oneNodeP oneNodeXMAHKF ( .n1(vdd_));
oneNodeP oneNodeXMAHKE ( .n1(vdd_));
oneNodeP oneNodeXMAHKD ( .n1(vdd_));
oneNodeP oneNodeXMAHGD ( .n1(vdd_));
oneNodeP oneNodeXMAHEP ( .n1(vdd_));
oneNodeP oneNodeXMAHEL ( .n1(vdd_));
oneNodeP oneNodeXMAHDO ( .n1(vdd_));
oneNodeP oneNodeXMAHDN ( .n1(vdd_));
oneNodeP oneNodeXMAHDM ( .n1(vdd_));
oneNodeP oneNodeXMAHDL ( .n1(vdd_));
oneNodeP oneNodeXMAHDK ( .n1(vdd_));
oneNodeP oneNodeXMAHBF ( .n1(vdd_));
oneNodeP oneNodeXMAGYZ ( .n1(vdd_));
oneNodeP oneNodeXMAGWT ( .n1(vdd_));
oneNodeP oneNodeXMAGUN ( .n1(vdd_));
oneNodeP oneNodeXMAGTK ( .n1(vdd_));
oneNodeP oneNodeXMAGTJ ( .n1(vdd_));
oneNodeP oneNodeXMAGTI ( .n1(vdd_));
oneNodeP oneNodeXMAFIG ( .n1(vdd_));
oneNodeP oneNodeXMAFIF ( .n1(vdd_));
oneNodeP oneNodeXMAFHY ( .n1(vdd_));
oneNodeP oneNodeXMAFHW ( .n1(vdd_));
oneNodeP oneNodeXMAFHE ( .n1(vdd_));
oneNodeP oneNodeXMAFHD ( .n1(vdd_));
oneNodeP oneNodeXMAFGW ( .n1(vdd_));
oneNodeP oneNodeXMAFGU ( .n1(vdd_));
oneNodeP oneNodeXMAFGC ( .n1(vdd_));
oneNodeP oneNodeXMAFGB ( .n1(vdd_));
oneNodeP oneNodeXMAFFU ( .n1(vdd_));
oneNodeP oneNodeXMAFFS ( .n1(vdd_));
oneNodeP oneNodeXMAFFA ( .n1(vdd_));
oneNodeP oneNodeXMAFEZ ( .n1(vdd_));
oneNodeP oneNodeXMAFES ( .n1(vdd_));
oneNodeP oneNodeXMAFEQ ( .n1(vdd_));
oneNodeP oneNodeXMAFDY ( .n1(vdd_));
oneNodeP oneNodeXMAFDX ( .n1(vdd_));
oneNodeP oneNodeXMAFDQ ( .n1(vdd_));
oneNodeP oneNodeXMAFDO ( .n1(vdd_));
oneNodeP oneNodeXMAFCW ( .n1(vdd_));
oneNodeP oneNodeXMAFCV ( .n1(vdd_));
oneNodeP oneNodeXMAFCO ( .n1(vdd_));
oneNodeP oneNodeXMAFCM ( .n1(vdd_));
oneNodeP oneNodeXMAFBU ( .n1(vdd_));
oneNodeP oneNodeXMAFBT ( .n1(vdd_));
oneNodeP oneNodeXMAFBM ( .n1(vdd_));
oneNodeP oneNodeXMAFBK ( .n1(vdd_));
twoNodeP twoNodeXMAFJW ( .n2(N00ADUT), .n1(vdd_));
twoNodeP twoNodeXMAFJV ( .n2(N00ADUS), .n1(vdd_));
twoNodeN twoNodeXMAFTW ( .n2(N00ADZB), .n1(gnd_));
twoNodeN twoNodeXMAFSZ ( .n2(N00ADZE), .n1(gnd_));
twoNodeN twoNodeXMAFJA ( .n2(N00ADUT), .n1(gnd_));
twoNodeN twoNodeXMAFIZ ( .n2(N00ADUS), .n1(gnd_));
dcapP dcap_XMAIBJ ( .n2(N00AEQN), .n1(vdd_));
dcapP dcap_XMAHVX ( .n2(N00AETN), .n1(vdd_));
dcapP dcap_XMAHUP ( .n2(N00AESX), .n1(vdd_));
dcapP dcap_XMAHOO ( .n2(N00AEJQ), .n1(vdd_));
dcapP dcap_XMAHMC ( .n2(N00AEPN), .n1(vdd_));
dcapP dcap_XMAHMA ( .n2(N00AEPM), .n1(vdd_));
dcapP dcap_XMAHKJ ( .n2(N00AEPH), .n1(vdd_));
dcapP dcap_XMAHKG ( .n2(N00AEPF), .n1(vdd_));
dcapP dcap_XMAHGC ( .n2(N00AENS), .n1(vdd_));
dcapP dcap_XMAHGB ( .n2(N00AEJX), .n1(vdd_));
dcapP dcap_XMAHGA ( .n2(N00AEJY), .n1(vdd_));
dcapP dcap_XMAHFZ ( .n2(N00AENP), .n1(vdd_));
dcapP dcap_XMAHEO ( .n2(N00AENG), .n1(vdd_));
dcapP dcap_XMAHEN ( .n2(N00AEJX), .n1(vdd_));
dcapP dcap_XMAHEM ( .n2(N00AEJZ), .n1(vdd_));
dcapP dcap_XMAHDJ ( .n2(N00AEJW), .n1(vdd_));
dcapP dcap_XMAHCI ( .n2(N00AEMH), .n1(vdd_));
dcapP dcap_XMAHCH ( .n2(N00AEMU), .n1(vdd_));
dcapP dcap_XMAHCC ( .n2(N00AEMX), .n1(vdd_));
dcapP dcap_XMAHBE ( .n2(N00AEMM), .n1(vdd_));
dcapP dcap_XMAHBD ( .n2(N00AEJZ), .n1(vdd_));
dcapP dcap_XMAHBC ( .n2(N00AEMH), .n1(vdd_));
dcapP dcap_XMAHBB ( .n2(N00AEMJ), .n1(vdd_));
dcapP dcap_XMAHAC ( .n2(N00AELQ), .n1(vdd_));
dcapP dcap_XMAHAB ( .n2(N00AEKG), .n1(vdd_));
dcapP dcap_XMAGZW ( .n2(N00AEMF), .n1(vdd_));
dcapP dcap_XMAGYY ( .n2(N00AELV), .n1(vdd_));
dcapP dcap_XMAGYX ( .n2(N00AEKE), .n1(vdd_));
dcapP dcap_XMAGYW ( .n2(N00AELQ), .n1(vdd_));
dcapP dcap_XMAGYV ( .n2(N00AELS), .n1(vdd_));
dcapP dcap_XMAGXW ( .n2(N00AELA), .n1(vdd_));
dcapP dcap_XMAGXV ( .n2(N00AEKF), .n1(vdd_));
dcapP dcap_XMAGXQ ( .n2(N00AELO), .n1(vdd_));
dcapP dcap_XMAGWS ( .n2(N00AELF), .n1(vdd_));
dcapP dcap_XMAGWR ( .n2(N00AEKD), .n1(vdd_));
dcapP dcap_XMAGWQ ( .n2(N00AELA), .n1(vdd_));
dcapP dcap_XMAGWP ( .n2(N00AELC), .n1(vdd_));
dcapP dcap_XMAGVQ ( .n2(N00AEKK), .n1(vdd_));
dcapP dcap_XMAGVP ( .n2(N00AEKH), .n1(vdd_));
dcapP dcap_XMAGVK ( .n2(N00AEKY), .n1(vdd_));
dcapP dcap_XMAGUM ( .n2(N00AEKP), .n1(vdd_));
dcapP dcap_XMAGUL ( .n2(N00AEKC), .n1(vdd_));
dcapP dcap_XMAGUK ( .n2(N00AEKK), .n1(vdd_));
dcapP dcap_XMAGUJ ( .n2(N00AEKM), .n1(vdd_));
dcapP dcap_XMAGRU ( .n2(N00ADRJ), .n1(vdd_));
dcapP dcap_XMAGRC ( .n2(N00ADZS), .n1(vdd_));
dcapP dcap_XMAGBY ( .n2(N00AECQ), .n1(vdd_));
dcapP dcap_XMAGAQ ( .n2(N00AECA), .n1(vdd_));
dcapP dcap_XMAFZI ( .n2(N00AEBK), .n1(vdd_));
dcapP dcap_XMAFIE ( .n2(N00ADUI), .n1(vdd_));
dcapP dcap_XMAFHZ ( .n2(N00ADUI), .n1(vdd_));
dcapP dcap_XMAFHC ( .n2(N00ADUB), .n1(vdd_));
dcapP dcap_XMAFGX ( .n2(N00ADUB), .n1(vdd_));
dcapP dcap_XMAFGA ( .n2(N00ADTT), .n1(vdd_));
dcapP dcap_XMAFFV ( .n2(N00ADTT), .n1(vdd_));
dcapP dcap_XMAFEY ( .n2(N00ADTL), .n1(vdd_));
dcapP dcap_XMAFET ( .n2(N00ADTL), .n1(vdd_));
dcapP dcap_XMAFDW ( .n2(N00ADTD), .n1(vdd_));
dcapP dcap_XMAFDR ( .n2(N00ADTD), .n1(vdd_));
dcapP dcap_XMAFCU ( .n2(N00ADSV), .n1(vdd_));
dcapP dcap_XMAFCP ( .n2(N00ADSV), .n1(vdd_));
dcapP dcap_XMAFBS ( .n2(N00ADSK), .n1(vdd_));
dcapP dcap_XMAFBN ( .n2(N00ADSK), .n1(vdd_));
dcapN dcap_XMAICH ( .n2(N00AEVW), .n1(gnd_));
dcapN dcap_XMAIAY ( .n2(N00AEVZ), .n1(gnd_));
dcapN dcap_XMAHYS ( .n2(N00AEVD), .n1(gnd_));
dcapN dcap_XMAHYO ( .n2(N00AEVD), .n1(gnd_));
dcapN dcap_XMAHLV ( .n2(N00AEPP), .n1(gnd_));
dcapN dcap_XMAHLT ( .n2(N00AEPO), .n1(gnd_));
dcapN dcap_XMAHLA ( .n2(N00AEJQ), .n1(gnd_));
dcapN dcap_XMAHKC ( .n2(N00AEPE), .n1(gnd_));
dcapN dcap_XMAHKB ( .n2(N00AEPH), .n1(gnd_));
dcapN dcap_XMAHKA ( .n2(N00AEPF), .n1(gnd_));
dcapN dcap_XMAHJZ ( .n2(N00AEPD), .n1(gnd_));
dcapN dcap_XMAHFX ( .n2(N00AENS), .n1(gnd_));
dcapN dcap_XMAHFW ( .n2(N00AEJX), .n1(gnd_));
dcapN dcap_XMAHFV ( .n2(N00AEJY), .n1(gnd_));
dcapN dcap_XMAHEJ ( .n2(N00AENG), .n1(gnd_));
dcapN dcap_XMAHEI ( .n2(N00AEJX), .n1(gnd_));
dcapN dcap_XMAHEH ( .n2(N00AEJZ), .n1(gnd_));
dcapN dcap_XMAHEG ( .n2(N00AEND), .n1(gnd_));
dcapN dcap_XMAHDI ( .n2(N00AENB), .n1(gnd_));
dcapN dcap_XMAHDD ( .n2(N00AEJW), .n1(gnd_));
dcapN dcap_XMAHBU ( .n2(N00AEMH), .n1(gnd_));
dcapN dcap_XMAHBT ( .n2(N00AEMU), .n1(gnd_));
dcapN dcap_XMAHAZ ( .n2(N00AEMM), .n1(gnd_));
dcapN dcap_XMAHAY ( .n2(N00AEJZ), .n1(gnd_));
dcapN dcap_XMAHAX ( .n2(N00AEMH), .n1(gnd_));
dcapN dcap_XMAGZO ( .n2(N00AELQ), .n1(gnd_));
dcapN dcap_XMAGZN ( .n2(N00AEKG), .n1(gnd_));
dcapN dcap_XMAGYT ( .n2(N00AELV), .n1(gnd_));
dcapN dcap_XMAGYS ( .n2(N00AEKE), .n1(gnd_));
dcapN dcap_XMAGYR ( .n2(N00AELQ), .n1(gnd_));
dcapN dcap_XMAGXI ( .n2(N00AELA), .n1(gnd_));
dcapN dcap_XMAGXH ( .n2(N00AEKF), .n1(gnd_));
dcapN dcap_XMAGWN ( .n2(N00AELF), .n1(gnd_));
dcapN dcap_XMAGWM ( .n2(N00AEKD), .n1(gnd_));
dcapN dcap_XMAGWL ( .n2(N00AELA), .n1(gnd_));
dcapN dcap_XMAGVD ( .n2(N00AEKX), .n1(gnd_));
dcapN dcap_XMAGVC ( .n2(N00AEKK), .n1(gnd_));
dcapN dcap_XMAGVB ( .n2(N00AEKH), .n1(gnd_));
dcapN dcap_XMAGUH ( .n2(N00AEKP), .n1(gnd_));
dcapN dcap_XMAGUG ( .n2(N00AEKC), .n1(gnd_));
dcapN dcap_XMAGUF ( .n2(N00AEKK), .n1(gnd_));
dcapN dcap_XMAGRW ( .n2(N00AEJB), .n1(gnd_));
dcapN dcap_XMAGOD ( .n2(N00AEDM), .n1(gnd_));
dcapN dcap_XMAGOC ( .n2(N00AEDM), .n1(gnd_));
dcapN dcap_XMAGNP ( .n2(N00AEIC), .n1(gnd_));
dcapN dcap_XMAGCE ( .n2(N00AEDG), .n1(gnd_));
dcapN dcap_XMAFJM ( .n2(N00ADUU), .n1(gnd_));
dcapN dcap_XMAFID ( .n2(N00ADUI), .n1(gnd_));
dcapN dcap_XMAFHO ( .n2(N00ADUF), .n1(gnd_));
dcapN dcap_XMAFHJ ( .n2(N00ADUI), .n1(gnd_));
dcapN dcap_XMAFHB ( .n2(N00ADUB), .n1(gnd_));
dcapN dcap_XMAFGM ( .n2(N00ADTX), .n1(gnd_));
dcapN dcap_XMAFGH ( .n2(N00ADUB), .n1(gnd_));
dcapN dcap_XMAFFZ ( .n2(N00ADTT), .n1(gnd_));
dcapN dcap_XMAFFK ( .n2(N00ADTP), .n1(gnd_));
dcapN dcap_XMAFFF ( .n2(N00ADTT), .n1(gnd_));
dcapN dcap_XMAFEX ( .n2(N00ADTL), .n1(gnd_));
dcapN dcap_XMAFEI ( .n2(N00ADTH), .n1(gnd_));
dcapN dcap_XMAFED ( .n2(N00ADTL), .n1(gnd_));
dcapN dcap_XMAFDV ( .n2(N00ADTD), .n1(gnd_));
dcapN dcap_XMAFDG ( .n2(N00ADSZ), .n1(gnd_));
dcapN dcap_XMAFDB ( .n2(N00ADTD), .n1(gnd_));
dcapN dcap_XMAFCT ( .n2(N00ADSV), .n1(gnd_));
dcapN dcap_XMAFCE ( .n2(N00ADSR), .n1(gnd_));
dcapN dcap_XMAFBZ ( .n2(N00ADSV), .n1(gnd_));
dcapN dcap_XMAFBR ( .n2(N00ADSK), .n1(gnd_));
dcapN dcap_XMAFBC ( .n2(N00ADSG), .n1(gnd_));
dcapN dcap_XMAFAX ( .n2(N00ADSK), .n1(gnd_));
dcapN dcap_XMAFAF ( .n2(N00ADRY), .n1(gnd_));
pch_mac  XMAICL ( .D(N00AEVW), .B(vdd_), .G(N00ADRR), .S(N00AEWJ));
pch_mac  XMAICK ( .D(N00AEWK), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAICJ ( .D(N00AEWJ), .B(vdd_), .G(N00AEWG), .S(N00AEWK));
pch_mac  XMAIBR ( .D(N00AEQO), .B(vdd_), .G(N00AEQW), .S(vdd_));
pch_mac  XMAIBQ ( .D(N00AEQO), .B(vdd_), .G(N00AEQV), .S(vdd_));
pch_mac  XMAIBP ( .D(N00AEQO), .B(vdd_), .G(N00AEQU), .S(vdd_));
pch_mac  XMAIBO ( .D(N00AEQO), .B(vdd_), .G(N00AEQT), .S(vdd_));
pch_mac  XMAIBN ( .D(N00AEQO), .B(vdd_), .G(N00AEQL), .S(vdd_));
pch_mac  XMAIBI ( .D(N00AEQN), .B(vdd_), .G(N00AEQV), .S(vdd_));
pch_mac  XMAIBH ( .D(N00AEQN), .B(vdd_), .G(N00AEQU), .S(vdd_));
pch_mac  XMAIBG ( .D(N00AEQN), .B(vdd_), .G(N00AEQT), .S(vdd_));
pch_mac  XMAIBF ( .D(N00AEQN), .B(vdd_), .G(N00AEQL), .S(vdd_));
pch_mac  XMAIBB ( .D(N00AESK), .B(vdd_), .G(N00AEQM), .S(vdd_));
pch_mac  XMAIBA ( .D(N00AESK), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAHZO ( .D(N00AEVC), .B(vdd_), .G(N00AEQR), .S(N00AEVO));
pch_mac  XMAHZM ( .D(N00AEVO), .B(vdd_), .G(N00AEVN), .S(vdd_));
pch_mac  XMAHZI ( .D(N00AEVK), .B(vdd_), .G(N00AEQZ), .S(N00AEVL));
pch_mac  XMAHZG ( .D(N00AEVL), .B(vdd_), .G(N00AEQX), .S(vdd_));
pch_mac  XMAHZC ( .D(N00AEQQ), .B(vdd_), .G(N00AEQY), .S(N00AEVI));
pch_mac  XMAHZA ( .D(N00AEVI), .B(vdd_), .G(N00AEQT), .S(vdd_));
pch_mac  XMAHYX ( .D(N00AEVH), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAHYW ( .D(N00AEVG), .B(vdd_), .G(DIVR3), .S(N00AEVH));
pch_mac  XMAHYV ( .D(N00AEVD), .B(vdd_), .G(gnd_), .S(N00AEVE));
pch_mac  XMAHYU ( .D(N00AEVF), .B(vdd_), .G(DIVR2), .S(N00AEVG));
pch_mac  XMAHYT ( .D(N00AEVE), .B(vdd_), .G(DIVR1), .S(N00AEVF));
pch_mac  XMAHWY ( .D(N00AEUM), .B(vdd_), .G(N00AEUF), .S(vdd_));
pch_mac  XMAHWX ( .D(N00AEUN), .B(vdd_), .G(N00AEQV), .S(vdd_));
pch_mac  XMAHWV ( .D(N00AEUE), .B(vdd_), .G(N00AEUD), .S(vdd_));
pch_mac  XMAHWU ( .D(N00AEUE), .B(vdd_), .G(N00AESV), .S(N00AEUN));
pch_mac  XMAHWT ( .D(N00AEUE), .B(vdd_), .G(N00AEUC), .S(N00AEUM));
pch_mac  XMAHVZ ( .D(N00AETN), .B(vdd_), .G(N00AEUB), .S(vdd_));
pch_mac  XMAHVY ( .D(N00AETN), .B(vdd_), .G(N00AEQR), .S(vdd_));
pch_mac  XMAHVQ ( .D(N00AETW), .B(vdd_), .G(N00AETP), .S(vdd_));
pch_mac  XMAHVP ( .D(N00AETX), .B(vdd_), .G(N00AEQU), .S(vdd_));
pch_mac  XMAHVN ( .D(N00AETO), .B(vdd_), .G(N00AETN), .S(vdd_));
pch_mac  XMAHVM ( .D(N00AETO), .B(vdd_), .G(N00AESU), .S(N00AETX));
pch_mac  XMAHVL ( .D(N00AETO), .B(vdd_), .G(N00AETM), .S(N00AETW));
pch_mac  XMAHUR ( .D(N00AESX), .B(vdd_), .G(N00AETL), .S(vdd_));
pch_mac  XMAHUQ ( .D(N00AESX), .B(vdd_), .G(N00AEQR), .S(vdd_));
pch_mac  XMAHUJ ( .D(N00AETI), .B(vdd_), .G(N00AEQT), .S(vdd_));
pch_mac  XMAHUI ( .D(N00AETG), .B(vdd_), .G(N00AESZ), .S(vdd_));
pch_mac  XMAHUH ( .D(N00AETH), .B(vdd_), .G(N00AEQT), .S(vdd_));
pch_mac  XMAHUG ( .D(N00AETA), .B(vdd_), .G(N00AESW), .S(N00AETI));
pch_mac  XMAHUF ( .D(N00AESY), .B(vdd_), .G(N00AESX), .S(vdd_));
pch_mac  XMAHUE ( .D(N00AESY), .B(vdd_), .G(N00AESW), .S(N00AETH));
pch_mac  XMAHUD ( .D(N00AESY), .B(vdd_), .G(N00AEQL), .S(N00AETG));
pch_mac  XMAHTE ( .D(N00AESQ), .B(vdd_), .G(N00AEQL), .S(N00AEST));
pch_mac  XMAHTD ( .D(N00AESS), .B(vdd_), .G(N00AEQR), .S(vdd_));
pch_mac  XMAHTC ( .D(N00AEST), .B(vdd_), .G(N00AESR), .S(vdd_));
pch_mac  XMAHTB ( .D(N00AESN), .B(vdd_), .G(N00AERB), .S(N00AESS));
pch_mac  XMAHTA ( .D(N00AESQ), .B(vdd_), .G(N00AEQM), .S(vdd_));
pch_mac  XMAHSA ( .D(N00AERV), .B(vdd_), .G(N00AERT), .S(N00AESG));
pch_mac  XMAHRZ ( .D(N00AERV), .B(vdd_), .G(N00AEQO), .S(N00AESH));
pch_mac  XMAHRY ( .D(N00AERV), .B(vdd_), .G(N00AERU), .S(vdd_));
pch_mac  XMAHRW ( .D(N00AESH), .B(vdd_), .G(N00AESD), .S(vdd_));
pch_mac  XMAHRV ( .D(N00AESG), .B(vdd_), .G(N00AERW), .S(vdd_));
pch_mac  XMAHQQ ( .D(N00AERN), .B(vdd_), .G(N00AERG), .S(vdd_));
pch_mac  XMAHQP ( .D(N00AERO), .B(vdd_), .G(N00AEQW), .S(vdd_));
pch_mac  XMAHQN ( .D(N00AERF), .B(vdd_), .G(N00AERE), .S(vdd_));
pch_mac  XMAHQM ( .D(N00AERF), .B(vdd_), .G(N00AEQN), .S(N00AERO));
pch_mac  XMAHQL ( .D(N00AERF), .B(vdd_), .G(N00AERD), .S(N00AERN));
pch_mac  XMAHPR ( .D(gnd_), .B(vdd_), .G(vdd_), .S(gnd_));
pch_mac  XMAHHO ( .D(N00AEOL), .B(vdd_), .G(N00AEJY), .S(vdd_));
pch_mac  XMAHHN ( .D(N00AEOJ), .B(vdd_), .G(N00AEOC), .S(vdd_));
pch_mac  XMAHHM ( .D(N00AEOK), .B(vdd_), .G(N00AENB), .S(vdd_));
pch_mac  XMAHHL ( .D(N00AEOD), .B(vdd_), .G(N00AEJU), .S(N00AEOL));
pch_mac  XMAHHK ( .D(N00AEOB), .B(vdd_), .G(N00AEJT), .S(vdd_));
pch_mac  XMAHHJ ( .D(N00AEOB), .B(vdd_), .G(N00AEJU), .S(N00AEOK));
pch_mac  XMAHHI ( .D(N00AEOB), .B(vdd_), .G(N00AEJV), .S(N00AEOJ));
pch_mac  XMAHGN ( .D(N00AENP), .B(vdd_), .G(N00AEJV), .S(N00AEOA));
pch_mac  XMAHGM ( .D(N00AENP), .B(vdd_), .G(N00AEJT), .S(vdd_));
pch_mac  XMAHGL ( .D(N00AENR), .B(vdd_), .G(N00AEJU), .S(N00AENZ));
pch_mac  XMAHGK ( .D(N00AEOA), .B(vdd_), .G(N00AENQ), .S(vdd_));
pch_mac  XMAHGJ ( .D(N00AENZ), .B(vdd_), .G(N00AEJX), .S(vdd_));
pch_mac  XMAHGI ( .D(N00AENY), .B(vdd_), .G(N00AENO), .S(vdd_));
pch_mac  XMAHGH ( .D(N00AENP), .B(vdd_), .G(N00AEJU), .S(N00AENY));
pch_mac  XMAHEZ ( .D(N00AEND), .B(vdd_), .G(N00AEJV), .S(N00AENK));
pch_mac  XMAHEY ( .D(N00AENF), .B(vdd_), .G(N00AEJU), .S(N00AENN));
pch_mac  XMAHEX ( .D(N00AENL), .B(vdd_), .G(N00AENE), .S(vdd_));
pch_mac  XMAHEW ( .D(N00AENN), .B(vdd_), .G(N00AEJR), .S(vdd_));
pch_mac  XMAHEV ( .D(N00AENM), .B(vdd_), .G(N00AENC), .S(vdd_));
pch_mac  XMAHEU ( .D(N00AEND), .B(vdd_), .G(N00AEJU), .S(N00AENM));
pch_mac  XMAHES ( .D(N00AENK), .B(vdd_), .G(N00AEJW), .S(N00AENL));
pch_mac  XMAHCB ( .D(N00AEMX), .B(vdd_), .G(N00AEMW), .S(vdd_));
pch_mac  XMAHCA ( .D(N00AEMG), .B(vdd_), .G(N00AEKE), .S(N00AEMX));
pch_mac  XMAHBZ ( .D(N00AEMG), .B(vdd_), .G(N00AEKG), .S(N00AEMX));
pch_mac  XMAHBP ( .D(N00AEMJ), .B(vdd_), .G(N00AEKA), .S(N00AEMT));
pch_mac  XMAHBO ( .D(N00AEMJ), .B(vdd_), .G(N00AEKI), .S(vdd_));
pch_mac  XMAHBN ( .D(N00AEML), .B(vdd_), .G(N00AEKB), .S(N00AEMS));
pch_mac  XMAHBM ( .D(N00AEMT), .B(vdd_), .G(N00AEMK), .S(vdd_));
pch_mac  XMAHBL ( .D(N00AEMS), .B(vdd_), .G(N00AEJZ), .S(vdd_));
pch_mac  XMAHBK ( .D(N00AEMR), .B(vdd_), .G(N00AEMI), .S(vdd_));
pch_mac  XMAHBJ ( .D(N00AEMJ), .B(vdd_), .G(N00AEKB), .S(N00AEMR));
pch_mac  XMAGZV ( .D(N00AEMF), .B(vdd_), .G(N00AEME), .S(vdd_));
pch_mac  XMAGZU ( .D(N00AELP), .B(vdd_), .G(N00AEKD), .S(N00AEMF));
pch_mac  XMAGZT ( .D(N00AELP), .B(vdd_), .G(N00AEKF), .S(N00AEMF));
pch_mac  XMAGZJ ( .D(N00AELS), .B(vdd_), .G(N00AEKA), .S(N00AEMC));
pch_mac  XMAGZI ( .D(N00AELS), .B(vdd_), .G(N00AEKI), .S(vdd_));
pch_mac  XMAGZH ( .D(N00AELU), .B(vdd_), .G(N00AEKB), .S(N00AEMB));
pch_mac  XMAGZG ( .D(N00AEMC), .B(vdd_), .G(N00AELT), .S(vdd_));
pch_mac  XMAGZF ( .D(N00AEMB), .B(vdd_), .G(N00AEKE), .S(vdd_));
pch_mac  XMAGZE ( .D(N00AEMA), .B(vdd_), .G(N00AELR), .S(vdd_));
pch_mac  XMAGZD ( .D(N00AELS), .B(vdd_), .G(N00AEKB), .S(N00AEMA));
pch_mac  XMAGXP ( .D(N00AELO), .B(vdd_), .G(DIVQ0), .S(vdd_));
pch_mac  XMAGXO ( .D(N00AEKZ), .B(vdd_), .G(N00AEKC), .S(N00AELO));
pch_mac  XMAGXN ( .D(N00AEKZ), .B(vdd_), .G(N00AEKH), .S(N00AELO));
pch_mac  XMAGXD ( .D(N00AELC), .B(vdd_), .G(N00AEKA), .S(N00AELM));
pch_mac  XMAGXC ( .D(N00AELC), .B(vdd_), .G(N00AEKI), .S(vdd_));
pch_mac  XMAGXB ( .D(N00AELE), .B(vdd_), .G(N00AEKB), .S(N00AELL));
pch_mac  XMAGXA ( .D(N00AELM), .B(vdd_), .G(N00AELD), .S(vdd_));
pch_mac  XMAGWZ ( .D(N00AELL), .B(vdd_), .G(N00AEKD), .S(vdd_));
pch_mac  XMAGWY ( .D(N00AELK), .B(vdd_), .G(N00AELB), .S(vdd_));
pch_mac  XMAGWX ( .D(N00AELC), .B(vdd_), .G(N00AEKB), .S(N00AELK));
pch_mac  XMAGVJ ( .D(N00AEKY), .B(vdd_), .G(DIVQ1), .S(vdd_));
pch_mac  XMAGVI ( .D(N00AEKJ), .B(vdd_), .G(gnd_), .S(N00AEKY));
pch_mac  XMAGVH ( .D(N00AEKJ), .B(vdd_), .G(gnd_), .S(N00AEKY));
pch_mac  XMAGUX ( .D(N00AEKM), .B(vdd_), .G(N00AEKA), .S(N00AEKW));
pch_mac  XMAGUW ( .D(N00AEKM), .B(vdd_), .G(N00AEKI), .S(vdd_));
pch_mac  XMAGUV ( .D(N00AEKO), .B(vdd_), .G(N00AEKB), .S(N00AEKV));
pch_mac  XMAGUU ( .D(N00AEKW), .B(vdd_), .G(N00AEKN), .S(vdd_));
pch_mac  XMAGUT ( .D(N00AEKV), .B(vdd_), .G(N00AEKC), .S(vdd_));
pch_mac  XMAGUS ( .D(N00AEKU), .B(vdd_), .G(N00AEKL), .S(vdd_));
pch_mac  XMAGUR ( .D(N00AEKM), .B(vdd_), .G(N00AEKB), .S(N00AEKU));
pch_mac  XMAGSA ( .D(N00AEJB), .B(vdd_), .G(N00ADRR), .S(N00AEJN));
pch_mac  XMAGRZ ( .D(N00AEJO), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAGRY ( .D(N00AEJN), .B(vdd_), .G(N00AEDM), .S(N00AEJO));
pch_mac  XMAGRT ( .D(N00ADRJ), .B(vdd_), .G(N00ADZX), .S(vdd_));
pch_mac  XMAGRK ( .D(N00ADZT), .B(vdd_), .G(N00AEAB), .S(vdd_));
pch_mac  XMAGRJ ( .D(N00ADZT), .B(vdd_), .G(N00AEAA), .S(vdd_));
pch_mac  XMAGRI ( .D(N00ADZT), .B(vdd_), .G(N00ADZZ), .S(vdd_));
pch_mac  XMAGRH ( .D(N00ADZT), .B(vdd_), .G(N00ADZY), .S(vdd_));
pch_mac  XMAGRG ( .D(N00ADZT), .B(vdd_), .G(N00ADZO), .S(vdd_));
pch_mac  XMAGRB ( .D(N00ADZS), .B(vdd_), .G(N00AEAA), .S(vdd_));
pch_mac  XMAGRA ( .D(N00ADZS), .B(vdd_), .G(N00ADZZ), .S(vdd_));
pch_mac  XMAGQZ ( .D(N00ADZS), .B(vdd_), .G(N00ADZY), .S(vdd_));
pch_mac  XMAGQY ( .D(N00ADZS), .B(vdd_), .G(N00ADZO), .S(vdd_));
pch_mac  XMAGOZ ( .D(N00AEAD), .B(vdd_), .G(N00ADZW), .S(N00AEIS));
pch_mac  XMAGOX ( .D(N00AEIS), .B(vdd_), .G(N00AEIR), .S(vdd_));
pch_mac  XMAGOT ( .D(N00AEIO), .B(vdd_), .G(N00AEAE), .S(N00AEIP));
pch_mac  XMAGOR ( .D(N00AEIP), .B(vdd_), .G(N00AEAC), .S(vdd_));
pch_mac  XMAGON ( .D(N00ADZV), .B(vdd_), .G(N00AEHW), .S(N00AEIM));
pch_mac  XMAGOL ( .D(N00AEIM), .B(vdd_), .G(N00ADZY), .S(vdd_));
pch_mac  XMAGOI ( .D(N00AEIL), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAGOH ( .D(N00AEIK), .B(vdd_), .G(gnd_), .S(N00AEIL));
pch_mac  XMAGOG ( .D(N00AEDM), .B(vdd_), .G(N00AEIH), .S(N00AEII));
pch_mac  XMAGOF ( .D(N00AEIJ), .B(vdd_), .G(DIVF6), .S(N00AEIK));
pch_mac  XMAGOE ( .D(N00AEII), .B(vdd_), .G(DIVF5), .S(N00AEIJ));
pch_mac  XMAGNY ( .D(N00AEIG), .B(vdd_), .G(DIVF4), .S(vdd_));
pch_mac  XMAGNX ( .D(N00AEIF), .B(vdd_), .G(DIVF3), .S(N00AEIG));
pch_mac  XMAGNW ( .D(N00AEIC), .B(vdd_), .G(gnd_), .S(N00AEID));
pch_mac  XMAGNV ( .D(N00AEIE), .B(vdd_), .G(DIVF2), .S(N00AEIF));
pch_mac  XMAGNU ( .D(N00AEID), .B(vdd_), .G(DIVF1), .S(N00AEIE));
pch_mac  XMAGNO ( .D(N00AEIB), .B(vdd_), .G(DIVF4), .S(vdd_));
pch_mac  XMAGNN ( .D(N00AEIA), .B(vdd_), .G(DIVF3), .S(N00AEIB));
pch_mac  XMAGNM ( .D(N00AEHX), .B(vdd_), .G(DIVF0), .S(N00AEHY));
pch_mac  XMAGNL ( .D(N00AEHZ), .B(vdd_), .G(DIVF2), .S(N00AEIA));
pch_mac  XMAGNK ( .D(N00AEHY), .B(vdd_), .G(DIVF1), .S(N00AEHZ));
pch_mac  XMAGLQ ( .D(N00AEHI), .B(vdd_), .G(N00AEAA), .S(vdd_));
pch_mac  XMAGLP ( .D(N00AEHG), .B(vdd_), .G(N00AEGZ), .S(vdd_));
pch_mac  XMAGLO ( .D(N00AEHH), .B(vdd_), .G(N00AEAA), .S(vdd_));
pch_mac  XMAGLN ( .D(N00AEHA), .B(vdd_), .G(N00AEFP), .S(N00AEHI));
pch_mac  XMAGLM ( .D(N00AEGY), .B(vdd_), .G(N00AEGX), .S(vdd_));
pch_mac  XMAGLL ( .D(N00AEGY), .B(vdd_), .G(N00AEFP), .S(N00AEHH));
pch_mac  XMAGLK ( .D(N00AEGY), .B(vdd_), .G(N00AEGW), .S(N00AEHG));
pch_mac  XMAGKI ( .D(N00AEGS), .B(vdd_), .G(N00ADZZ), .S(vdd_));
pch_mac  XMAGKH ( .D(N00AEGQ), .B(vdd_), .G(N00AEGJ), .S(vdd_));
pch_mac  XMAGKG ( .D(N00AEGR), .B(vdd_), .G(N00ADZZ), .S(vdd_));
pch_mac  XMAGKF ( .D(N00AEGK), .B(vdd_), .G(N00AEFO), .S(N00AEGS));
pch_mac  XMAGKE ( .D(N00AEGI), .B(vdd_), .G(N00AEGH), .S(vdd_));
pch_mac  XMAGKD ( .D(N00AEGI), .B(vdd_), .G(N00AEFO), .S(N00AEGR));
pch_mac  XMAGKC ( .D(N00AEGI), .B(vdd_), .G(N00AEGG), .S(N00AEGQ));
pch_mac  XMAGJA ( .D(N00AEGC), .B(vdd_), .G(N00ADZY), .S(vdd_));
pch_mac  XMAGIZ ( .D(N00AEGA), .B(vdd_), .G(N00AEFT), .S(vdd_));
pch_mac  XMAGIY ( .D(N00AEGB), .B(vdd_), .G(N00ADZY), .S(vdd_));
pch_mac  XMAGIX ( .D(N00AEFU), .B(vdd_), .G(N00AEFQ), .S(N00AEGC));
pch_mac  XMAGIW ( .D(N00AEFS), .B(vdd_), .G(N00AEFR), .S(vdd_));
pch_mac  XMAGIV ( .D(N00AEFS), .B(vdd_), .G(N00AEFQ), .S(N00AEGB));
pch_mac  XMAGIU ( .D(N00AEFS), .B(vdd_), .G(N00ADZO), .S(N00AEGA));
pch_mac  XMAGHV ( .D(N00AEFK), .B(vdd_), .G(N00ADZO), .S(N00AEFN));
pch_mac  XMAGHU ( .D(N00AEFM), .B(vdd_), .G(N00ADZW), .S(vdd_));
pch_mac  XMAGHT ( .D(N00AEFN), .B(vdd_), .G(N00AEFL), .S(vdd_));
pch_mac  XMAGHS ( .D(N00AEFH), .B(vdd_), .G(N00AEAF), .S(N00AEFM));
pch_mac  XMAGHR ( .D(N00AEFK), .B(vdd_), .G(N00ADZR), .S(vdd_));
pch_mac  XMAGGR ( .D(N00AEEP), .B(vdd_), .G(N00AEEN), .S(N00AEFA));
pch_mac  XMAGGQ ( .D(N00AEEP), .B(vdd_), .G(N00ADZT), .S(N00AEFB));
pch_mac  XMAGGP ( .D(N00AEEP), .B(vdd_), .G(N00AEEO), .S(vdd_));
pch_mac  XMAGGO ( .D(N00AEES), .B(vdd_), .G(N00ADZT), .S(N00AEEZ));
pch_mac  XMAGGN ( .D(N00AEFB), .B(vdd_), .G(N00AEEX), .S(vdd_));
pch_mac  XMAGGM ( .D(N00AEFA), .B(vdd_), .G(N00AEEQ), .S(vdd_));
pch_mac  XMAGGL ( .D(N00AEEZ), .B(vdd_), .G(N00AEAC), .S(vdd_));
pch_mac  XMAGFI ( .D(N00AEEJ), .B(vdd_), .G(N00AEAB), .S(vdd_));
pch_mac  XMAGFH ( .D(N00AEEH), .B(vdd_), .G(N00AEEA), .S(vdd_));
pch_mac  XMAGFG ( .D(N00AEEI), .B(vdd_), .G(N00AEAB), .S(vdd_));
pch_mac  XMAGFF ( .D(N00AEEB), .B(vdd_), .G(N00ADZS), .S(N00AEEJ));
pch_mac  XMAGFE ( .D(N00AEDZ), .B(vdd_), .G(N00AEDY), .S(vdd_));
pch_mac  XMAGFD ( .D(N00AEDZ), .B(vdd_), .G(N00ADZS), .S(N00AEEI));
pch_mac  XMAGFC ( .D(N00AEDZ), .B(vdd_), .G(N00AEDX), .S(N00AEEH));
pch_mac  XMAGDD ( .D(N00AEDL), .B(vdd_), .G(N00AEDM), .S(vdd_));
pch_mac  XMAGDC ( .D(N00AEDL), .B(vdd_), .G(N00AEDM), .S(vdd_));
pch_mac  XMAGDB ( .D(N00ADZX), .B(vdd_), .G(N00ADZW), .S(N00AEDL));
pch_mac  XMAGDA ( .D(N00ADZX), .B(vdd_), .G(N00AEAY), .S(N00AEDL));
pch_mac  XMAGCP ( .D(N00AEBY), .B(vdd_), .G(N00AEBD), .S(vdd_));
pch_mac  XMAGCO ( .D(N00AEBY), .B(vdd_), .G(DIVF5), .S(vdd_));
pch_mac  XMAGCL ( .D(N00AECO), .B(vdd_), .G(N00AEBD), .S(vdd_));
pch_mac  XMAGCK ( .D(N00AECO), .B(vdd_), .G(DIVF6), .S(vdd_));
pch_mac  XMAGCH ( .D(N00AEDE), .B(vdd_), .G(N00AEBD), .S(vdd_));
pch_mac  XMAGCG ( .D(N00AEDE), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAGCD ( .D(N00AEBH), .B(vdd_), .G(N00AEAU), .S(vdd_));
pch_mac  XMAGCC ( .D(N00AEBH), .B(vdd_), .G(N00AEAX), .S(vdd_));
pch_mac  XMAGBZ ( .D(N00AECQ), .B(vdd_), .G(N00AEDE), .S(vdd_));
pch_mac  XMAGBX ( .D(N00AECQ), .B(vdd_), .G(N00ADZQ), .S(vdd_));
pch_mac  XMAGBR ( .D(N00AEDB), .B(vdd_), .G(N00AEAW), .S(vdd_));
pch_mac  XMAGBQ ( .D(N00AECZ), .B(vdd_), .G(N00AECS), .S(vdd_));
pch_mac  XMAGBP ( .D(N00AEDA), .B(vdd_), .G(N00AEAW), .S(vdd_));
pch_mac  XMAGBO ( .D(N00AECT), .B(vdd_), .G(N00AEBI), .S(N00AEDB));
pch_mac  XMAGBN ( .D(N00AECR), .B(vdd_), .G(N00AECQ), .S(vdd_));
pch_mac  XMAGBM ( .D(N00AECR), .B(vdd_), .G(N00AEBI), .S(N00AEDA));
pch_mac  XMAGBL ( .D(N00AECR), .B(vdd_), .G(N00AECP), .S(N00AECZ));
pch_mac  XMAGAR ( .D(N00AECA), .B(vdd_), .G(N00AECO), .S(vdd_));
pch_mac  XMAGAP ( .D(N00AECA), .B(vdd_), .G(N00ADZQ), .S(vdd_));
pch_mac  XMAGAJ ( .D(N00AECL), .B(vdd_), .G(N00AEAV), .S(vdd_));
pch_mac  XMAGAI ( .D(N00AECJ), .B(vdd_), .G(N00AECC), .S(vdd_));
pch_mac  XMAGAH ( .D(N00AECK), .B(vdd_), .G(N00AEAV), .S(vdd_));
pch_mac  XMAGAG ( .D(N00AECD), .B(vdd_), .G(N00AEBH), .S(N00AECL));
pch_mac  XMAGAF ( .D(N00AECB), .B(vdd_), .G(N00AECA), .S(vdd_));
pch_mac  XMAGAE ( .D(N00AECB), .B(vdd_), .G(N00AEBH), .S(N00AECK));
pch_mac  XMAGAD ( .D(N00AECB), .B(vdd_), .G(N00AEBZ), .S(N00AECJ));
pch_mac  XMAFZJ ( .D(N00AEBK), .B(vdd_), .G(N00AEBY), .S(vdd_));
pch_mac  XMAFZH ( .D(N00AEBK), .B(vdd_), .G(N00ADZQ), .S(vdd_));
pch_mac  XMAFZB ( .D(N00AEBV), .B(vdd_), .G(N00AEAU), .S(vdd_));
pch_mac  XMAFZA ( .D(N00AEBT), .B(vdd_), .G(N00AEBM), .S(vdd_));
pch_mac  XMAFYZ ( .D(N00AEBU), .B(vdd_), .G(N00AEAU), .S(vdd_));
pch_mac  XMAFYY ( .D(N00AEBN), .B(vdd_), .G(N00AEBJ), .S(N00AEBV));
pch_mac  XMAFYX ( .D(N00AEBL), .B(vdd_), .G(N00AEBK), .S(vdd_));
pch_mac  XMAFYW ( .D(N00AEBL), .B(vdd_), .G(N00AEBJ), .S(N00AEBU));
pch_mac  XMAFYV ( .D(N00AEBL), .B(vdd_), .G(N00AEAX), .S(N00AEBT));
pch_mac  XMAFXZ ( .D(N00AEBA), .B(vdd_), .G(N00AEBD), .S(vdd_));
pch_mac  XMAFXY ( .D(N00AEAX), .B(vdd_), .G(N00AEBA), .S(vdd_));
pch_mac  XMAFXX ( .D(N00AEAX), .B(vdd_), .G(N00AEAS), .S(vdd_));
pch_mac  XMAFXW ( .D(N00AEBG), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAFXV ( .D(N00AEBA), .B(vdd_), .G(N00ADZW), .S(N00AEBF));
pch_mac  XMAFXU ( .D(N00AEBA), .B(vdd_), .G(N00ADZW), .S(N00AEBG));
pch_mac  XMAFXT ( .D(N00AEBF), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAFXC ( .D(N00AEAI), .B(vdd_), .G(N00AEAN), .S(N00AEAR));
pch_mac  XMAFXB ( .D(N00AEAQ), .B(vdd_), .G(N00AEAL), .S(vdd_));
pch_mac  XMAFXA ( .D(N00AEAR), .B(vdd_), .G(N00AEAL), .S(vdd_));
pch_mac  XMAFWZ ( .D(N00AEAI), .B(vdd_), .G(N00AEAN), .S(N00AEAQ));
pch_mac  XMAFWX ( .D(N00AEAK), .B(vdd_), .G(N00AEAI), .S(vdd_));
pch_mac  XMAFWG ( .D(gnd_), .B(vdd_), .G(vdd_), .S(gnd_));
pch_mac  XMAFQG ( .D(N00ADXZ), .B(vdd_), .G(N00ADXW), .S(vdd_));
pch_mac  XMAFQF ( .D(N00ADXZ), .B(vdd_), .G(RANGE1), .S(vdd_));
pch_mac  XMAFQC ( .D(N00ADYB), .B(vdd_), .G(RANGE2), .S(vdd_));
pch_mac  XMAFQB ( .D(N00ADYB), .B(vdd_), .G(RANGE0), .S(vdd_));
pch_mac  XMAFPY ( .D(N00ADYA), .B(vdd_), .G(N00ADYB), .S(vdd_));
pch_mac  XMAFPX ( .D(N00ADYA), .B(vdd_), .G(N00ADXZ), .S(vdd_));
pch_mac  XMAFPU ( .D(N00ADXT), .B(vdd_), .G(RANGE2), .S(vdd_));
pch_mac  XMAFPT ( .D(N00ADXT), .B(vdd_), .G(RANGE1), .S(vdd_));
pch_mac  XMAFOB ( .D(N00ADXB), .B(vdd_), .G(N00ADWV), .S(vdd_));
pch_mac  XMAFOA ( .D(N00ADVK), .B(vdd_), .G(N00ADWW), .S(N00ADXB));
pch_mac  XMAFMY ( .D(N00ADWR), .B(vdd_), .G(N00ADWK), .S(vdd_));
pch_mac  XMAFMX ( .D(N00ADVL), .B(vdd_), .G(N00ADWL), .S(N00ADWR));
pch_mac  XMAFMW ( .D(N00ADWQ), .B(vdd_), .G(N00ADWL), .S(vdd_));
pch_mac  XMAFMV ( .D(N00ADVL), .B(vdd_), .G(N00ADWK), .S(N00ADWQ));
pch_mac  XMAFMR ( .D(N00ADWK), .B(vdd_), .G(N00ADWM), .S(N00ADWP));
pch_mac  XMAFMQ ( .D(N00ADWP), .B(vdd_), .G(N00ADWL), .S(vdd_));
pch_mac  XMAFMF ( .D(N00ADWH), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAFME ( .D(N00ADUS), .B(vdd_), .G(N00ADVI), .S(vdd_));
pch_mac  XMAFMD ( .D(N00ADWJ), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAFMC ( .D(N00ADWI), .B(vdd_), .G(gnd_), .S(N00ADWJ));
pch_mac  XMAFMB ( .D(N00ADVC), .B(vdd_), .G(N00ADVJ), .S(N00ADWI));
pch_mac  XMAFMA ( .D(N00ADWG), .B(vdd_), .G(gnd_), .S(N00ADWH));
pch_mac  XMAFLZ ( .D(N00ADWF), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAFLY ( .D(N00ADWE), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAFLX ( .D(N00ADVD), .B(vdd_), .G(N00ADVJ), .S(N00ADWG));
pch_mac  XMAFLW ( .D(N00ADVE), .B(vdd_), .G(N00ADVJ), .S(N00ADWF));
pch_mac  XMAFLU ( .D(N00ADVF), .B(vdd_), .G(N00ADVJ), .S(N00ADWE));
pch_mac  XMAFLT ( .D(N00ADUS), .B(vdd_), .G(N00ADVJ), .S(vdd_));
pch_mac  XMAFLQ ( .D(N00ADVG), .B(vdd_), .G(N00ADVB), .S(vdd_));
pch_mac  XMAFJX ( .D(N00ADUV), .B(vdd_), .G(N00ADRR), .S(vdd_));
pch_mac  XMAFJS ( .D(N00ADUS), .B(vdd_), .G(N00ADVB), .S(vdd_));
pch_mac  XMAFIY ( .D(N00ADUR), .B(vdd_), .G(N00ADUN), .S(vdd_));
pch_mac  XMAFIX ( .D(N00ADSP), .B(vdd_), .G(N00ADQO), .S(N00ADUQ));
pch_mac  XMAFIW ( .D(N00ADSP), .B(vdd_), .G(N00ADQO), .S(N00ADUR));
pch_mac  XMAFIV ( .D(N00ADUQ), .B(vdd_), .G(N00ADUN), .S(vdd_));
pch_mac  XMAFHV ( .D(N00ADUF), .B(vdd_), .G(N00ADUE), .S(vdd_));
pch_mac  XMAFHU ( .D(N00ADUH), .B(vdd_), .G(LOCK), .S(vdd_));
pch_mac  XMAFGT ( .D(N00ADTX), .B(vdd_), .G(N00ADTW), .S(vdd_));
pch_mac  XMAFGS ( .D(N00ADUA), .B(vdd_), .G(N00ADTZ), .S(vdd_));
pch_mac  XMAFFR ( .D(N00ADTP), .B(vdd_), .G(N00ADTO), .S(vdd_));
pch_mac  XMAFFQ ( .D(N00ADTS), .B(vdd_), .G(N00ADTR), .S(vdd_));
pch_mac  XMAFEP ( .D(N00ADTH), .B(vdd_), .G(N00ADTG), .S(vdd_));
pch_mac  XMAFEO ( .D(N00ADTK), .B(vdd_), .G(N00ADTJ), .S(vdd_));
pch_mac  XMAFDN ( .D(N00ADSZ), .B(vdd_), .G(N00ADSY), .S(vdd_));
pch_mac  XMAFDM ( .D(N00ADTC), .B(vdd_), .G(N00ADTB), .S(vdd_));
pch_mac  XMAFCL ( .D(N00ADSR), .B(vdd_), .G(N00ADSQ), .S(vdd_));
pch_mac  XMAFCK ( .D(N00ADSU), .B(vdd_), .G(N00ADST), .S(vdd_));
pch_mac  XMAFBJ ( .D(N00ADSG), .B(vdd_), .G(N00ADSF), .S(vdd_));
pch_mac  XMAFBI ( .D(N00ADSJ), .B(vdd_), .G(N00ADSI), .S(vdd_));
pch_mac  XMAFAS ( .D(N00ADRM), .B(vdd_), .G(N00ADRP), .S(vdd_));
pch_mac  XMAFAR ( .D(N00ADRM), .B(vdd_), .G(N00ADSE), .S(vdd_));
pch_mac  XMAFAM ( .D(N00ADSC), .B(vdd_), .G(REF), .S(vdd_));
pch_mac  XMAFAL ( .D(N00ADRL), .B(vdd_), .G(N00ADRZ), .S(N00ADSC));
pch_mac  XMAFAK ( .D(N00ADSB), .B(vdd_), .G(gnd_), .S(vdd_));
pch_mac  XMAFAJ ( .D(N00ADRL), .B(vdd_), .G(N00ADRQ), .S(N00ADSB));
pch_mac  XMAFAC ( .D(N00ADRX), .B(vdd_), .G(N00ADRL), .S(vdd_));
pch_mac  XMAFAB ( .D(N00ADRN), .B(vdd_), .G(N00ADRL), .S(N00ADRX));
pch_mac  XMAEZY ( .D(N00ADRV), .B(vdd_), .G(N00ADRO), .S(vdd_));
pch_mac  XMAEZX ( .D(N00ADRP), .B(vdd_), .G(N00ADRO), .S(N00ADRV));
pch_mac  XMAEZU ( .D(N00ADRT), .B(vdd_), .G(N00ADRN), .S(vdd_));
pch_mac  XMAEZT ( .D(N00ADRO), .B(vdd_), .G(N00ADRN), .S(N00ADRT));
pch_mac  XMAEZE ( .D(N00ADQR), .B(vdd_), .G(N00ADQU), .S(vdd_));
pch_mac  XMAEZD ( .D(N00ADQR), .B(vdd_), .G(N00ADRJ), .S(vdd_));
pch_mac  XMAEYY ( .D(N00ADRH), .B(vdd_), .G(FB), .S(vdd_));
pch_mac  XMAEYX ( .D(N00ADQQ), .B(vdd_), .G(N00ADRE), .S(N00ADRH));
pch_mac  XMAEYW ( .D(N00ADRG), .B(vdd_), .G(N00ADRD), .S(vdd_));
pch_mac  XMAEYV ( .D(N00ADQQ), .B(vdd_), .G(N00ADQV), .S(N00ADRG));
pch_mac  XMAEYO ( .D(N00ADRB), .B(vdd_), .G(N00ADQQ), .S(vdd_));
pch_mac  XMAEYN ( .D(N00ADQS), .B(vdd_), .G(N00ADQQ), .S(N00ADRB));
pch_mac  XMAEYK ( .D(N00ADQZ), .B(vdd_), .G(N00ADQT), .S(vdd_));
pch_mac  XMAEYJ ( .D(N00ADQU), .B(vdd_), .G(N00ADQT), .S(N00ADQZ));
pch_mac  XMAEYG ( .D(N00ADQX), .B(vdd_), .G(N00ADQS), .S(vdd_));
pch_mac  XMAEYF ( .D(N00ADQT), .B(vdd_), .G(N00ADQS), .S(N00ADQX));
nch_mac  M0 ( .D(N00AERI), .B(gnd_), .G(N00AEQN), .S(N00AERF));
nch_mac  XMAICI ( .D(gnd_), .B(gnd_), .G(N00AEWG), .S(N00AEVW));
nch_mac  XMAICG ( .D(gnd_), .B(gnd_), .G(N00ADRR), .S(N00AEVW));
nch_mac  XMAIBM ( .D(gnd_), .B(gnd_), .G(N00AEQT), .S(N00AEWD));
nch_mac  XMAIBL ( .D(N00AEWD), .B(gnd_), .G(N00AEVR), .S(N00AEWC));
nch_mac  XMAIBK ( .D(N00AEWC), .B(gnd_), .G(N00AEQL), .S(N00AEQO));
nch_mac  XMAIBE ( .D(gnd_), .B(gnd_), .G(N00AEQT), .S(N00AEWB));
nch_mac  XMAIBD ( .D(N00AEWB), .B(gnd_), .G(N00AEVQ), .S(N00AEWA));
nch_mac  XMAIBC ( .D(N00AEWA), .B(gnd_), .G(N00AEQL), .S(N00AEQN));
nch_mac  XMAIAZ ( .D(N00AEVZ), .B(gnd_), .G(N00AEQM), .S(N00AESK));
nch_mac  XMAHYR ( .D(gnd_), .B(gnd_), .G(DIVR3), .S(N00AEVD));
nch_mac  XMAHYQ ( .D(gnd_), .B(gnd_), .G(DIVR2), .S(N00AEVD));
nch_mac  XMAHYP ( .D(gnd_), .B(gnd_), .G(DIVR1), .S(N00AEVD));
nch_mac  XMAHWP ( .D(gnd_), .B(gnd_), .G(N00AEUF), .S(N00AEUI));
nch_mac  XMAHWO ( .D(gnd_), .B(gnd_), .G(N00AEUD), .S(N00AEUK));
nch_mac  XMAHWN ( .D(N00AEUJ), .B(gnd_), .G(N00AEUC), .S(N00AEUE));
nch_mac  XMAHWJ ( .D(N00AEUK), .B(gnd_), .G(N00AEQV), .S(N00AEUJ));
nch_mac  XMAHWI ( .D(N00AEUH), .B(gnd_), .G(N00AESV), .S(N00AEUE));
nch_mac  XMAHWG ( .D(N00AEUI), .B(gnd_), .G(N00AEUD), .S(N00AEUH));
nch_mac  XMAHVW ( .D(gnd_), .B(gnd_), .G(N00AEUB), .S(N00AEUA));
nch_mac  XMAHVV ( .D(N00AEUA), .B(gnd_), .G(vdd_), .S(N00AETZ));
nch_mac  XMAHVU ( .D(N00AETZ), .B(gnd_), .G(N00AEQR), .S(N00AETN));
nch_mac  XMAHVH ( .D(gnd_), .B(gnd_), .G(N00AETP), .S(N00AETS));
nch_mac  XMAHVG ( .D(gnd_), .B(gnd_), .G(N00AETN), .S(N00AETU));
nch_mac  XMAHVF ( .D(N00AETT), .B(gnd_), .G(N00AETM), .S(N00AETO));
nch_mac  XMAHVB ( .D(N00AETU), .B(gnd_), .G(N00AEQU), .S(N00AETT));
nch_mac  XMAHVA ( .D(N00AETR), .B(gnd_), .G(N00AESU), .S(N00AETO));
nch_mac  XMAHUY ( .D(N00AETS), .B(gnd_), .G(N00AETN), .S(N00AETR));
nch_mac  XMAHUO ( .D(gnd_), .B(gnd_), .G(N00AETL), .S(N00AETK));
nch_mac  XMAHUN ( .D(N00AETK), .B(gnd_), .G(vdd_), .S(N00AETJ));
nch_mac  XMAHUM ( .D(N00AETJ), .B(gnd_), .G(N00AEQR), .S(N00AESX));
nch_mac  XMAHTZ ( .D(gnd_), .B(gnd_), .G(N00AESZ), .S(N00AETC));
nch_mac  XMAHTY ( .D(gnd_), .B(gnd_), .G(N00AESX), .S(N00AETE));
nch_mac  XMAHTX ( .D(N00AETD), .B(gnd_), .G(N00AEQL), .S(N00AESY));
nch_mac  XMAHTV ( .D(gnd_), .B(gnd_), .G(N00AEQT), .S(N00AETF));
nch_mac  XMAHTU ( .D(N00AETF), .B(gnd_), .G(N00AEQL), .S(N00AETA));
nch_mac  XMAHTT ( .D(N00AETE), .B(gnd_), .G(N00AEQT), .S(N00AETD));
nch_mac  XMAHTS ( .D(N00AETB), .B(gnd_), .G(N00AESW), .S(N00AESY));
nch_mac  XMAHTQ ( .D(N00AETC), .B(gnd_), .G(N00AESX), .S(N00AETB));
nch_mac  XMAHSW ( .D(gnd_), .B(gnd_), .G(N00AESR), .S(N00AESM));
nch_mac  XMAHSU ( .D(N00AESL), .B(gnd_), .G(N00AEQP), .S(N00AESQ));
nch_mac  XMAHSR ( .D(gnd_), .B(gnd_), .G(N00AEQR), .S(N00AESP));
nch_mac  XMAHSQ ( .D(N00AESP), .B(gnd_), .G(N00AEQL), .S(N00AESN));
nch_mac  XMAHSO ( .D(gnd_), .B(gnd_), .G(N00AESO), .S(N00AESN));
nch_mac  XMAHSN ( .D(N00AESM), .B(gnd_), .G(N00AEQM), .S(N00AESL));
nch_mac  XMAHRP ( .D(N00AESA), .B(gnd_), .G(N00AERU), .S(N00AESE));
nch_mac  XMAHRN ( .D(N00AESE), .B(gnd_), .G(N00AEQO), .S(N00AERV));
nch_mac  XMAHRM ( .D(N00AESB), .B(gnd_), .G(N00AESD), .S(N00AERZ));
nch_mac  XMAHRI ( .D(gnd_), .B(gnd_), .G(N00AERU), .S(N00AESB));
nch_mac  XMAHRH ( .D(gnd_), .B(gnd_), .G(N00AERW), .S(N00AESA));
nch_mac  XMAHRG ( .D(N00AERZ), .B(gnd_), .G(N00AERT), .S(N00AERV));
nch_mac  XMAHQH ( .D(gnd_), .B(gnd_), .G(N00AERG), .S(N00AERJ));
nch_mac  XMAHQG ( .D(gnd_), .B(gnd_), .G(N00AERE), .S(N00AERL));
nch_mac  XMAHQF ( .D(N00AERK), .B(gnd_), .G(N00AERD), .S(N00AERF));
nch_mac  XMAHQB ( .D(N00AERL), .B(gnd_), .G(N00AEQW), .S(N00AERK));
nch_mac  XMAHPY ( .D(N00AERJ), .B(gnd_), .G(N00AERE), .S(N00AERI));
nch_mac  XMAHMQ ( .D(gnd_), .B(gnd_), .G(N00AEPO), .S(N00AEPV));
nch_mac  XMAHMP ( .D(N00AEPV), .B(gnd_), .G(N00AEPP), .S(N00AEPS));
nch_mac  XMAHKW ( .D(gnd_), .B(gnd_), .G(N00AEPD), .S(N00AEPL));
nch_mac  XMAHKV ( .D(N00AEPL), .B(gnd_), .G(N00AEPE), .S(N00AEJP));
nch_mac  XMAHIG ( .D(gnd_), .B(gnd_), .G(N00AEOO), .S(N00AEOP));
nch_mac  XMAHIF ( .D(gnd_), .B(gnd_), .G(N00AEOO), .S(N00AEOP));
nch_mac  XMAHIE ( .D(gnd_), .B(gnd_), .G(N00AEOO), .S(N00AEOP));
nch_mac  XMAHID ( .D(N00AEOP), .B(gnd_), .G(N00AEJS), .S(N00AEJU));
nch_mac  XMAHIB ( .D(gnd_), .B(gnd_), .G(N00AEOO), .S(N00AEON));
nch_mac  XMAHIA ( .D(gnd_), .B(gnd_), .G(N00AEOO), .S(N00AEON));
nch_mac  XMAHHE ( .D(gnd_), .B(gnd_), .G(N00AEOC), .S(N00AEOF));
nch_mac  XMAHHD ( .D(gnd_), .B(gnd_), .G(N00AEJT), .S(N00AEOH));
nch_mac  XMAHHC ( .D(N00AEOG), .B(gnd_), .G(N00AEJV), .S(N00AEOB));
nch_mac  XMAHHA ( .D(gnd_), .B(gnd_), .G(N00AEJY), .S(N00AEOI));
nch_mac  XMAHGZ ( .D(N00AEOI), .B(gnd_), .G(N00AEJV), .S(N00AEOD));
nch_mac  XMAHGY ( .D(N00AEOH), .B(gnd_), .G(N00AENB), .S(N00AEOG));
nch_mac  XMAHGX ( .D(N00AEOE), .B(gnd_), .G(N00AEJU), .S(N00AEOB));
nch_mac  XMAHGV ( .D(N00AEOF), .B(gnd_), .G(N00AEJT), .S(N00AEOE));
nch_mac  XMAHFQ ( .D(N00AENT), .B(gnd_), .G(N00AEJU), .S(N00AENP));
nch_mac  XMAHFP ( .D(N00AENX), .B(gnd_), .G(N00AEJV), .S(N00AENR));
nch_mac  XMAHFO ( .D(gnd_), .B(gnd_), .G(N00AEJX), .S(N00AENX));
nch_mac  XMAHFM ( .D(gnd_), .B(gnd_), .G(N00AENQ), .S(N00AENU));
nch_mac  XMAHFL ( .D(N00AENW), .B(gnd_), .G(N00AEJV), .S(N00AENP));
nch_mac  XMAHFK ( .D(gnd_), .B(gnd_), .G(N00AENO), .S(N00AENW));
nch_mac  XMAHFI ( .D(N00AENU), .B(gnd_), .G(N00AEJT), .S(N00AENT));
nch_mac  XMAHEC ( .D(N00AENI), .B(gnd_), .G(N00AEJU), .S(N00AEND));
nch_mac  XMAHEB ( .D(N00AENJ), .B(gnd_), .G(N00AEJV), .S(N00AENF));
nch_mac  XMAHEA ( .D(gnd_), .B(gnd_), .G(N00AEJR), .S(N00AENJ));
nch_mac  XMAHDY ( .D(gnd_), .B(gnd_), .G(N00AENE), .S(N00AENI));
nch_mac  XMAHDX ( .D(N00AENH), .B(gnd_), .G(N00AEJV), .S(N00AEND));
nch_mac  XMAHDW ( .D(gnd_), .B(gnd_), .G(N00AENC), .S(N00AENH));
nch_mac  XMAHDU ( .D(gnd_), .B(gnd_), .G(N00AEJW), .S(N00AEND));
nch_mac  XMAHCU ( .D(gnd_), .B(gnd_), .G(N00AEMZ), .S(N00AENA));
nch_mac  XMAHCT ( .D(gnd_), .B(gnd_), .G(N00AEMZ), .S(N00AENA));
nch_mac  XMAHCS ( .D(gnd_), .B(gnd_), .G(N00AEMZ), .S(N00AENA));
nch_mac  XMAHCR ( .D(N00AENA), .B(gnd_), .G(N00AEJX), .S(N00AEKA));
nch_mac  XMAHCP ( .D(gnd_), .B(gnd_), .G(N00AEMZ), .S(N00AEMY));
nch_mac  XMAHCO ( .D(gnd_), .B(gnd_), .G(N00AEMZ), .S(N00AEMY));
nch_mac  XMAHBX ( .D(gnd_), .B(gnd_), .G(N00AEMW), .S(N00AEMG));
nch_mac  XMAHBW ( .D(N00AEMV), .B(gnd_), .G(N00AEKE), .S(N00AEMG));
nch_mac  XMAHBV ( .D(gnd_), .B(gnd_), .G(N00AEKG), .S(N00AEMV));
nch_mac  XMAHAS ( .D(N00AEMN), .B(gnd_), .G(N00AEKB), .S(N00AEMJ));
nch_mac  XMAHAR ( .D(N00AEMQ), .B(gnd_), .G(N00AEKA), .S(N00AEML));
nch_mac  XMAHAQ ( .D(gnd_), .B(gnd_), .G(N00AEJZ), .S(N00AEMQ));
nch_mac  XMAHAO ( .D(gnd_), .B(gnd_), .G(N00AEMK), .S(N00AEMO));
nch_mac  XMAHAN ( .D(N00AEMP), .B(gnd_), .G(N00AEKA), .S(N00AEMJ));
nch_mac  XMAHAM ( .D(gnd_), .B(gnd_), .G(N00AEMI), .S(N00AEMP));
nch_mac  XMAHAK ( .D(N00AEMO), .B(gnd_), .G(N00AEKI), .S(N00AEMN));
nch_mac  XMAGZR ( .D(gnd_), .B(gnd_), .G(N00AEME), .S(N00AELP));
nch_mac  XMAGZQ ( .D(N00AEMD), .B(gnd_), .G(N00AEKD), .S(N00AELP));
nch_mac  XMAGZP ( .D(gnd_), .B(gnd_), .G(N00AEKF), .S(N00AEMD));
nch_mac  XMAGYM ( .D(N00AELW), .B(gnd_), .G(N00AEKB), .S(N00AELS));
nch_mac  XMAGYL ( .D(N00AELZ), .B(gnd_), .G(N00AEKA), .S(N00AELU));
nch_mac  XMAGYK ( .D(gnd_), .B(gnd_), .G(N00AEKE), .S(N00AELZ));
nch_mac  XMAGYI ( .D(gnd_), .B(gnd_), .G(N00AELT), .S(N00AELX));
nch_mac  XMAGYH ( .D(N00AELY), .B(gnd_), .G(N00AEKA), .S(N00AELS));
nch_mac  XMAGYG ( .D(gnd_), .B(gnd_), .G(N00AELR), .S(N00AELY));
nch_mac  XMAGYE ( .D(N00AELX), .B(gnd_), .G(N00AEKI), .S(N00AELW));
nch_mac  XMAGXL ( .D(gnd_), .B(gnd_), .G(DIVQ0), .S(N00AEKZ));
nch_mac  XMAGXK ( .D(N00AELN), .B(gnd_), .G(N00AEKC), .S(N00AEKZ));
nch_mac  XMAGXJ ( .D(gnd_), .B(gnd_), .G(N00AEKH), .S(N00AELN));
nch_mac  XMAGWG ( .D(N00AELG), .B(gnd_), .G(N00AEKB), .S(N00AELC));
nch_mac  XMAGWF ( .D(N00AELJ), .B(gnd_), .G(N00AEKA), .S(N00AELE));
nch_mac  XMAGWE ( .D(gnd_), .B(gnd_), .G(N00AEKD), .S(N00AELJ));
nch_mac  XMAGWC ( .D(gnd_), .B(gnd_), .G(N00AELD), .S(N00AELH));
nch_mac  XMAGWB ( .D(N00AELI), .B(gnd_), .G(N00AEKA), .S(N00AELC));
nch_mac  XMAGWA ( .D(gnd_), .B(gnd_), .G(N00AELB), .S(N00AELI));
nch_mac  XMAGVY ( .D(N00AELH), .B(gnd_), .G(N00AEKI), .S(N00AELG));
nch_mac  XMAGVF ( .D(gnd_), .B(gnd_), .G(DIVQ1), .S(N00AEKJ));
nch_mac  XMAGVE ( .D(N00AEKX), .B(gnd_), .G(gnd_), .S(N00AEKJ));
nch_mac  XMAGUA ( .D(N00AEKQ), .B(gnd_), .G(N00AEKB), .S(N00AEKM));
nch_mac  XMAGTZ ( .D(N00AEKT), .B(gnd_), .G(N00AEKA), .S(N00AEKO));
nch_mac  XMAGTY ( .D(gnd_), .B(gnd_), .G(N00AEKC), .S(N00AEKT));
nch_mac  XMAGTW ( .D(gnd_), .B(gnd_), .G(N00AEKN), .S(N00AEKR));
nch_mac  XMAGTV ( .D(N00AEKS), .B(gnd_), .G(N00AEKA), .S(N00AEKM));
nch_mac  XMAGTU ( .D(gnd_), .B(gnd_), .G(N00AEKL), .S(N00AEKS));
nch_mac  XMAGTS ( .D(N00AEKR), .B(gnd_), .G(N00AEKI), .S(N00AEKQ));
nch_mac  XMAGRX ( .D(gnd_), .B(gnd_), .G(N00AEDM), .S(N00AEJB));
nch_mac  XMAGRV ( .D(gnd_), .B(gnd_), .G(N00ADRR), .S(N00AEJB));
nch_mac  XMAGRS ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00AEJM));
nch_mac  XMAGRR ( .D(N00AEJM), .B(gnd_), .G(N00ADZX), .S(N00ADRJ));
nch_mac  XMAGRF ( .D(gnd_), .B(gnd_), .G(N00ADZY), .S(N00AEJJ));
nch_mac  XMAGRE ( .D(N00AEJJ), .B(gnd_), .G(N00AEIW), .S(N00AEJI));
nch_mac  XMAGRD ( .D(N00AEJI), .B(gnd_), .G(N00ADZO), .S(N00ADZT));
nch_mac  XMAGQX ( .D(gnd_), .B(gnd_), .G(N00ADZY), .S(N00AEJH));
nch_mac  XMAGQW ( .D(N00AEJH), .B(gnd_), .G(N00AEIU), .S(N00AEJG));
nch_mac  XMAGQV ( .D(N00AEJG), .B(gnd_), .G(N00ADZO), .S(N00ADZS));
nch_mac  XMAGOB ( .D(gnd_), .B(gnd_), .G(DIVF6), .S(N00AEDM));
nch_mac  XMAGOA ( .D(gnd_), .B(gnd_), .G(DIVF5), .S(N00AEDM));
nch_mac  XMAGNZ ( .D(gnd_), .B(gnd_), .G(N00AEIH), .S(N00AEDM));
nch_mac  XMAGNT ( .D(gnd_), .B(gnd_), .G(DIVF4), .S(N00AEIC));
nch_mac  XMAGNS ( .D(gnd_), .B(gnd_), .G(DIVF3), .S(N00AEIC));
nch_mac  XMAGNR ( .D(gnd_), .B(gnd_), .G(DIVF2), .S(N00AEIC));
nch_mac  XMAGNQ ( .D(gnd_), .B(gnd_), .G(DIVF1), .S(N00AEIC));
nch_mac  XMAGNJ ( .D(gnd_), .B(gnd_), .G(DIVF4), .S(N00AEHX));
nch_mac  XMAGNI ( .D(gnd_), .B(gnd_), .G(DIVF3), .S(N00AEHX));
nch_mac  XMAGNH ( .D(gnd_), .B(gnd_), .G(DIVF2), .S(N00AEHX));
nch_mac  XMAGNG ( .D(gnd_), .B(gnd_), .G(DIVF1), .S(N00AEHX));
nch_mac  XMAGNF ( .D(gnd_), .B(gnd_), .G(DIVF0), .S(N00AEHX));
nch_mac  XMAGLG ( .D(gnd_), .B(gnd_), .G(N00AEGZ), .S(N00AEHC));
nch_mac  XMAGLF ( .D(gnd_), .B(gnd_), .G(N00AEGX), .S(N00AEHE));
nch_mac  XMAGLE ( .D(N00AEHD), .B(gnd_), .G(N00AEGW), .S(N00AEGY));
nch_mac  XMAGLC ( .D(gnd_), .B(gnd_), .G(N00AEAA), .S(N00AEHF));
nch_mac  XMAGLB ( .D(N00AEHF), .B(gnd_), .G(N00AEGW), .S(N00AEHA));
nch_mac  XMAGLA ( .D(N00AEHE), .B(gnd_), .G(N00AEAA), .S(N00AEHD));
nch_mac  XMAGKZ ( .D(N00AEHB), .B(gnd_), .G(N00AEFP), .S(N00AEGY));
nch_mac  XMAGKX ( .D(N00AEHC), .B(gnd_), .G(N00AEGX), .S(N00AEHB));
nch_mac  XMAGJY ( .D(gnd_), .B(gnd_), .G(N00AEGJ), .S(N00AEGM));
nch_mac  XMAGJX ( .D(gnd_), .B(gnd_), .G(N00AEGH), .S(N00AEGO));
nch_mac  XMAGJW ( .D(N00AEGN), .B(gnd_), .G(N00AEGG), .S(N00AEGI));
nch_mac  XMAGJU ( .D(gnd_), .B(gnd_), .G(N00ADZZ), .S(N00AEGP));
nch_mac  XMAGJT ( .D(N00AEGP), .B(gnd_), .G(N00AEGG), .S(N00AEGK));
nch_mac  XMAGJS ( .D(N00AEGO), .B(gnd_), .G(N00ADZZ), .S(N00AEGN));
nch_mac  XMAGJR ( .D(N00AEGL), .B(gnd_), .G(N00AEFO), .S(N00AEGI));
nch_mac  XMAGJP ( .D(N00AEGM), .B(gnd_), .G(N00AEGH), .S(N00AEGL));
nch_mac  XMAGIQ ( .D(gnd_), .B(gnd_), .G(N00AEFT), .S(N00AEFW));
nch_mac  XMAGIP ( .D(gnd_), .B(gnd_), .G(N00AEFR), .S(N00AEFY));
nch_mac  XMAGIO ( .D(N00AEFX), .B(gnd_), .G(N00ADZO), .S(N00AEFS));
nch_mac  XMAGIM ( .D(gnd_), .B(gnd_), .G(N00ADZY), .S(N00AEFZ));
nch_mac  XMAGIL ( .D(N00AEFZ), .B(gnd_), .G(N00ADZO), .S(N00AEFU));
nch_mac  XMAGIK ( .D(N00AEFY), .B(gnd_), .G(N00ADZY), .S(N00AEFX));
nch_mac  XMAGIJ ( .D(N00AEFV), .B(gnd_), .G(N00AEFQ), .S(N00AEFS));
nch_mac  XMAGIH ( .D(N00AEFW), .B(gnd_), .G(N00AEFR), .S(N00AEFV));
nch_mac  XMAGHN ( .D(gnd_), .B(gnd_), .G(N00AEFL), .S(N00AEFG));
nch_mac  XMAGHL ( .D(N00AEFF), .B(gnd_), .G(N00ADZU), .S(N00AEFK));
nch_mac  XMAGHI ( .D(gnd_), .B(gnd_), .G(N00ADZW), .S(N00AEFJ));
nch_mac  XMAGHH ( .D(N00AEFJ), .B(gnd_), .G(N00ADZO), .S(N00AEFH));
nch_mac  XMAGHF ( .D(gnd_), .B(gnd_), .G(N00AEFI), .S(N00AEFH));
nch_mac  XMAGHE ( .D(N00AEFG), .B(gnd_), .G(N00ADZR), .S(N00AEFF));
nch_mac  XMAGGG ( .D(N00AEEU), .B(gnd_), .G(N00AEEO), .S(N00AEEY));
nch_mac  XMAGGE ( .D(N00AEEY), .B(gnd_), .G(N00ADZT), .S(N00AEEP));
nch_mac  XMAGGD ( .D(N00AEEV), .B(gnd_), .G(N00AEEX), .S(N00AEET));
nch_mac  XMAGGC ( .D(N00AEEW), .B(gnd_), .G(N00AEEN), .S(N00AEES));
nch_mac  XMAGGB ( .D(gnd_), .B(gnd_), .G(N00AEAC), .S(N00AEEW));
nch_mac  XMAGFZ ( .D(gnd_), .B(gnd_), .G(N00AEEO), .S(N00AEEV));
nch_mac  XMAGFY ( .D(gnd_), .B(gnd_), .G(N00AEEQ), .S(N00AEEU));
nch_mac  XMAGFX ( .D(N00AEET), .B(gnd_), .G(N00AEEN), .S(N00AEEP));
nch_mac  XMAGEY ( .D(gnd_), .B(gnd_), .G(N00AEEA), .S(N00AEED));
nch_mac  XMAGEX ( .D(gnd_), .B(gnd_), .G(N00AEDY), .S(N00AEEF));
nch_mac  XMAGEW ( .D(N00AEEE), .B(gnd_), .G(N00AEDX), .S(N00AEDZ));
nch_mac  XMAGEU ( .D(gnd_), .B(gnd_), .G(N00AEAB), .S(N00AEEG));
nch_mac  XMAGET ( .D(N00AEEG), .B(gnd_), .G(N00AEDX), .S(N00AEEB));
nch_mac  XMAGES ( .D(N00AEEF), .B(gnd_), .G(N00AEAB), .S(N00AEEE));
nch_mac  XMAGER ( .D(N00AEEC), .B(gnd_), .G(N00ADZS), .S(N00AEDZ));
nch_mac  XMAGEP ( .D(N00AEED), .B(gnd_), .G(N00AEDY), .S(N00AEEC));
nch_mac  XMAGEF ( .D(gnd_), .B(gnd_), .G(N00AEAW), .S(N00AEDW));
nch_mac  XMAGED ( .D(N00AEDW), .B(gnd_), .G(N00AEAV), .S(N00AEDU));
nch_mac  XMAGEB ( .D(N00AEDU), .B(gnd_), .G(N00AEAU), .S(N00AEAT));
nch_mac  XMAGCZ ( .D(gnd_), .B(gnd_), .G(N00AEAY), .S(N00AEDN));
nch_mac  XMAGCY ( .D(N00AEDN), .B(gnd_), .G(N00ADZW), .S(N00ADZX));
nch_mac  XMAGCX ( .D(gnd_), .B(gnd_), .G(N00AEDM), .S(N00ADZX));
nch_mac  XMAGCN ( .D(N00AEDI), .B(gnd_), .G(N00AEBD), .S(N00AEBY));
nch_mac  XMAGCM ( .D(gnd_), .B(gnd_), .G(DIVF5), .S(N00AEDI));
nch_mac  XMAGCJ ( .D(N00AEDH), .B(gnd_), .G(N00AEBD), .S(N00AECO));
nch_mac  XMAGCI ( .D(gnd_), .B(gnd_), .G(DIVF6), .S(N00AEDH));
nch_mac  XMAGCF ( .D(N00AEDG), .B(gnd_), .G(N00AEBD), .S(N00AEDE));
nch_mac  XMAGCB ( .D(N00AEDF), .B(gnd_), .G(N00AEAX), .S(N00AEBH));
nch_mac  XMAGCA ( .D(gnd_), .B(gnd_), .G(N00AEAU), .S(N00AEDF));
nch_mac  XMAGBW ( .D(gnd_), .B(gnd_), .G(N00AEDE), .S(N00AEDD));
nch_mac  XMAGBV ( .D(N00AEDD), .B(gnd_), .G(N00ADZQ), .S(N00AEDC));
nch_mac  XMAGBU ( .D(N00AEDC), .B(gnd_), .G(vdd_), .S(N00AECQ));
nch_mac  XMAGBH ( .D(gnd_), .B(gnd_), .G(N00AECS), .S(N00AECV));
nch_mac  XMAGBG ( .D(gnd_), .B(gnd_), .G(N00AECQ), .S(N00AECX));
nch_mac  XMAGBF ( .D(N00AECW), .B(gnd_), .G(N00AECP), .S(N00AECR));
nch_mac  XMAGBD ( .D(gnd_), .B(gnd_), .G(N00AEAW), .S(N00AECY));
nch_mac  XMAGBC ( .D(N00AECY), .B(gnd_), .G(N00AECP), .S(N00AECT));
nch_mac  XMAGBB ( .D(N00AECX), .B(gnd_), .G(N00AEAW), .S(N00AECW));
nch_mac  XMAGBA ( .D(N00AECU), .B(gnd_), .G(N00AEBI), .S(N00AECR));
nch_mac  XMAGAY ( .D(N00AECV), .B(gnd_), .G(N00AECQ), .S(N00AECU));
nch_mac  XMAGAO ( .D(gnd_), .B(gnd_), .G(N00AECO), .S(N00AECN));
nch_mac  XMAGAN ( .D(N00AECN), .B(gnd_), .G(N00ADZQ), .S(N00AECM));
nch_mac  XMAGAM ( .D(N00AECM), .B(gnd_), .G(vdd_), .S(N00AECA));
nch_mac  XMAFZZ ( .D(gnd_), .B(gnd_), .G(N00AECC), .S(N00AECF));
nch_mac  XMAFZY ( .D(gnd_), .B(gnd_), .G(N00AECA), .S(N00AECH));
nch_mac  XMAFZX ( .D(N00AECG), .B(gnd_), .G(N00AEBZ), .S(N00AECB));
nch_mac  XMAFZV ( .D(gnd_), .B(gnd_), .G(N00AEAV), .S(N00AECI));
nch_mac  XMAFZU ( .D(N00AECI), .B(gnd_), .G(N00AEBZ), .S(N00AECD));
nch_mac  XMAFZT ( .D(N00AECH), .B(gnd_), .G(N00AEAV), .S(N00AECG));
nch_mac  XMAFZS ( .D(N00AECE), .B(gnd_), .G(N00AEBH), .S(N00AECB));
nch_mac  XMAFZQ ( .D(N00AECF), .B(gnd_), .G(N00AECA), .S(N00AECE));
nch_mac  XMAFZG ( .D(gnd_), .B(gnd_), .G(N00AEBY), .S(N00AEBX));
nch_mac  XMAFZF ( .D(N00AEBX), .B(gnd_), .G(N00ADZQ), .S(N00AEBW));
nch_mac  XMAFZE ( .D(N00AEBW), .B(gnd_), .G(vdd_), .S(N00AEBK));
nch_mac  XMAFYR ( .D(gnd_), .B(gnd_), .G(N00AEBM), .S(N00AEBP));
nch_mac  XMAFYQ ( .D(gnd_), .B(gnd_), .G(N00AEBK), .S(N00AEBR));
nch_mac  XMAFYP ( .D(N00AEBQ), .B(gnd_), .G(N00AEAX), .S(N00AEBL));
nch_mac  XMAFYN ( .D(gnd_), .B(gnd_), .G(N00AEAU), .S(N00AEBS));
nch_mac  XMAFYM ( .D(N00AEBS), .B(gnd_), .G(N00AEAX), .S(N00AEBN));
nch_mac  XMAFYL ( .D(N00AEBR), .B(gnd_), .G(N00AEAU), .S(N00AEBQ));
nch_mac  XMAFYK ( .D(N00AEBO), .B(gnd_), .G(N00AEBJ), .S(N00AEBL));
nch_mac  XMAFYI ( .D(N00AEBP), .B(gnd_), .G(N00AEBK), .S(N00AEBO));
nch_mac  XMAFXS ( .D(N00AEBE), .B(gnd_), .G(N00AEAX), .S(N00AEBA));
nch_mac  XMAFXR ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00AEBE));
nch_mac  XMAFXQ ( .D(gnd_), .B(gnd_), .G(N00AEBD), .S(N00AEBB));
nch_mac  XMAFXP ( .D(gnd_), .B(gnd_), .G(N00AEAS), .S(N00AEBC));
nch_mac  XMAFXO ( .D(N00AEBC), .B(gnd_), .G(N00AEBA), .S(N00AEAX));
nch_mac  XMAFXN ( .D(N00AEBB), .B(gnd_), .G(N00ADZW), .S(N00AEBA));
nch_mac  XMAFWT ( .D(N00AEAP), .B(gnd_), .G(N00AEAN), .S(N00AEAK));
nch_mac  XMAFWS ( .D(gnd_), .B(gnd_), .G(N00AEAL), .S(N00AEAI));
nch_mac  XMAFWR ( .D(gnd_), .B(gnd_), .G(N00AEAI), .S(N00AEAP));
nch_mac  XMAFWN ( .D(N00AEAM), .B(gnd_), .G(N00AEAN), .S(N00AEAK));
nch_mac  XMAFWM ( .D(gnd_), .B(gnd_), .G(N00AEAI), .S(N00AEAM));
nch_mac  XMAFWL ( .D(gnd_), .B(gnd_), .G(N00AEAL), .S(N00AEAI));
nch_mac  XMAFUN ( .D(gnd_), .B(gnd_), .G(N00ADYZ), .S(N00ADZI));
nch_mac  XMAFUM ( .D(gnd_), .B(gnd_), .G(N00ADZF), .S(N00ADZJ));
nch_mac  XMAFUL ( .D(gnd_), .B(gnd_), .G(N00ADRR), .S(N00ADZL));
nch_mac  XMAFUK ( .D(gnd_), .B(gnd_), .G(N00ADZL), .S(N00ADZK));
nch_mac  XMAFUJ ( .D(gnd_), .B(gnd_), .G(N00ADZK), .S(N00ADZJ));
nch_mac  XMAFUI ( .D(gnd_), .B(gnd_), .G(N00ADZJ), .S(N00ADZH));
nch_mac  XMAFUH ( .D(gnd_), .B(gnd_), .G(N00ADZH), .S(N00ADZG));
nch_mac  XMAFTU ( .D(gnd_), .B(gnd_), .G(N00ADZF), .S(N00ADZA));
nch_mac  XMAFTS ( .D(gnd_), .B(gnd_), .G(N00ADYZ), .S(N00ADZF));
nch_mac  XMAFTD ( .D(gnd_), .B(gnd_), .G(RANGE2), .S(N00ADZD));
nch_mac  XMAFTA ( .D(gnd_), .B(gnd_), .G(N00ADZC), .S(N00ADZE));
nch_mac  XMAFSY ( .D(gnd_), .B(gnd_), .G(N00ADZD), .S(N00ADZC));
nch_mac  XMAFSW ( .D(gnd_), .B(gnd_), .G(N00ADZA), .S(N00ADYZ));
nch_mac  XMAFSJ ( .D(N00ADXP), .B(gnd_), .G(N00ADYX), .S(N00ADVG));
nch_mac  XMAFSI ( .D(gnd_), .B(gnd_), .G(N00ADYY), .S(N00ADYX));
nch_mac  XMAFSH ( .D(gnd_), .B(gnd_), .G(N00ADXS), .S(N00ADYY));
nch_mac  XMAFSG ( .D(N00ADVF), .B(gnd_), .G(N00ADYX), .S(N00ADXP));
nch_mac  XMAFRZ ( .D(N00ADXN), .B(gnd_), .G(N00ADYV), .S(N00ADVG));
nch_mac  XMAFRY ( .D(gnd_), .B(gnd_), .G(N00ADYW), .S(N00ADYV));
nch_mac  XMAFRX ( .D(gnd_), .B(gnd_), .G(N00ADYE), .S(N00ADYW));
nch_mac  XMAFRW ( .D(N00ADVE), .B(gnd_), .G(N00ADYV), .S(N00ADXN));
nch_mac  XMAFRP ( .D(N00ADXL), .B(gnd_), .G(N00ADYT), .S(N00ADVG));
nch_mac  XMAFRO ( .D(gnd_), .B(gnd_), .G(N00ADYU), .S(N00ADYT));
nch_mac  XMAFRN ( .D(gnd_), .B(gnd_), .G(N00ADYA), .S(N00ADYU));
nch_mac  XMAFRM ( .D(N00ADVD), .B(gnd_), .G(N00ADYT), .S(N00ADXL));
nch_mac  XMAFRF ( .D(N00ADXJ), .B(gnd_), .G(N00ADYR), .S(N00ADVG));
nch_mac  XMAFRE ( .D(gnd_), .B(gnd_), .G(N00ADYS), .S(N00ADYR));
nch_mac  XMAFRD ( .D(gnd_), .B(gnd_), .G(N00ADXR), .S(N00ADYS));
nch_mac  XMAFRC ( .D(N00ADVC), .B(gnd_), .G(N00ADYR), .S(N00ADXJ));
nch_mac  XMAFQE ( .D(N00ADYD), .B(gnd_), .G(N00ADXW), .S(N00ADXZ));
nch_mac  XMAFQD ( .D(gnd_), .B(gnd_), .G(RANGE1), .S(N00ADYD));
nch_mac  XMAFQA ( .D(N00ADYC), .B(gnd_), .G(RANGE2), .S(N00ADYB));
nch_mac  XMAFPZ ( .D(gnd_), .B(gnd_), .G(RANGE0), .S(N00ADYC));
nch_mac  XMAFPW ( .D(N00ADXY), .B(gnd_), .G(N00ADYB), .S(N00ADYA));
nch_mac  XMAFPV ( .D(gnd_), .B(gnd_), .G(N00ADXZ), .S(N00ADXY));
nch_mac  XMAFPS ( .D(N00ADXX), .B(gnd_), .G(RANGE2), .S(N00ADXT));
nch_mac  XMAFPR ( .D(gnd_), .B(gnd_), .G(RANGE1), .S(N00ADXX));
nch_mac  XMAFNX ( .D(gnd_), .B(gnd_), .G(N00ADWN), .S(N00ADVK));
nch_mac  XMAFMU ( .D(gnd_), .B(gnd_), .G(N00ADWN), .S(N00ADVL));
nch_mac  XMAFMT ( .D(gnd_), .B(gnd_), .G(N00ADWK), .S(N00ADVL));
nch_mac  XMAFMS ( .D(gnd_), .B(gnd_), .G(N00ADWL), .S(N00ADVL));
nch_mac  XMAFMP ( .D(gnd_), .B(gnd_), .G(N00ADWL), .S(N00ADWK));
nch_mac  XMAFMO ( .D(gnd_), .B(gnd_), .G(N00ADWM), .S(N00ADWK));
nch_mac  XMAFLP ( .D(gnd_), .B(gnd_), .G(N00ADVB), .S(N00ADWD));
nch_mac  XMAFLO ( .D(N00ADWD), .B(gnd_), .G(N00ADVB), .S(N00ADWC));
nch_mac  XMAFLN ( .D(N00ADWC), .B(gnd_), .G(N00ADVB), .S(N00ADVZ));
nch_mac  XMAFLM ( .D(gnd_), .B(gnd_), .G(N00ADVB), .S(N00ADWB));
nch_mac  XMAFLL ( .D(N00ADWB), .B(gnd_), .G(N00ADVB), .S(N00ADVV));
nch_mac  XMAFLK ( .D(gnd_), .B(gnd_), .G(N00ADVB), .S(N00ADVR));
nch_mac  XMAFLJ ( .D(N00ADVY), .B(gnd_), .G(vdd_), .S(N00ADVC));
nch_mac  XMAFLI ( .D(N00ADWA), .B(gnd_), .G(N00ADVL), .S(N00ADUS));
nch_mac  XMAFLH ( .D(gnd_), .B(gnd_), .G(N00ADVK), .S(N00ADWA));
nch_mac  XMAFLG ( .D(N00ADVQ), .B(gnd_), .G(vdd_), .S(N00ADVE));
nch_mac  XMAFLF ( .D(N00ADVU), .B(gnd_), .G(vdd_), .S(N00ADVD));
nch_mac  XMAFLE ( .D(N00ADVZ), .B(gnd_), .G(N00ADVB), .S(N00ADVX));
nch_mac  XMAFLD ( .D(N00ADVW), .B(gnd_), .G(N00ADVH), .S(N00ADVY));
nch_mac  XMAFLC ( .D(N00ADVX), .B(gnd_), .G(vdd_), .S(N00ADVW));
nch_mac  XMAFLB ( .D(N00ADVV), .B(gnd_), .G(N00ADVB), .S(N00ADVT));
nch_mac  XMAFLA ( .D(N00ADVS), .B(gnd_), .G(N00ADVH), .S(N00ADVU));
nch_mac  XMAFKZ ( .D(N00ADVT), .B(gnd_), .G(vdd_), .S(N00ADVS));
nch_mac  XMAFKY ( .D(N00ADVR), .B(gnd_), .G(N00ADVB), .S(N00ADVP));
nch_mac  XMAFKX ( .D(N00ADVO), .B(gnd_), .G(N00ADVH), .S(N00ADVQ));
nch_mac  XMAFKW ( .D(N00ADVP), .B(gnd_), .G(vdd_), .S(N00ADVO));
nch_mac  XMAFKU ( .D(N00ADVM), .B(gnd_), .G(vdd_), .S(N00ADVN));
nch_mac  XMAFKT ( .D(N00ADVN), .B(gnd_), .G(N00ADVH), .S(N00ADVF));
nch_mac  XMAFKS ( .D(gnd_), .B(gnd_), .G(N00ADVB), .S(N00ADVM));
nch_mac  XMAFJI ( .D(N00ADUU), .B(gnd_), .G(N00ADVB), .S(N00ADUS));
nch_mac  XMAFJH ( .D(N00ADUX), .B(gnd_), .G(N00ADUY), .S(N00ADUW));
nch_mac  XMAFJD ( .D(gnd_), .B(gnd_), .G(N00ADUT), .S(N00ADUX));
nch_mac  XMAFJB ( .D(gnd_), .B(gnd_), .G(N00ADUV), .S(N00ADUU));
nch_mac  XMAFIU ( .D(gnd_), .B(gnd_), .G(N00ADUN), .S(N00ADSP));
nch_mac  XMAFIT ( .D(gnd_), .B(gnd_), .G(N00ADQO), .S(N00ADSP));
nch_mac  XMAFHQ ( .D(gnd_), .B(gnd_), .G(N00ADUB), .S(N00ADUK));
nch_mac  XMAFHP ( .D(N00ADUK), .B(gnd_), .G(N00ADSN), .S(N00ADUF));
nch_mac  XMAFHN ( .D(gnd_), .B(gnd_), .G(N00ADSN), .S(LOCK));
nch_mac  XMAFHL ( .D(N00ADUJ), .B(gnd_), .G(LOCK), .S(N00ADUH));
nch_mac  XMAFHK ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADUJ));
nch_mac  XMAFHI ( .D(N00ADUG), .B(gnd_), .G(N00ADUE), .S(N00ADUF));
nch_mac  XMAFHG ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADUG));
nch_mac  XMAFGO ( .D(gnd_), .B(gnd_), .G(N00ADTT), .S(N00ADUD));
nch_mac  XMAFGN ( .D(N00ADUD), .B(gnd_), .G(N00ADSN), .S(N00ADTX));
nch_mac  XMAFGL ( .D(gnd_), .B(gnd_), .G(N00ADSN), .S(N00ADTZ));
nch_mac  XMAFGJ ( .D(N00ADUC), .B(gnd_), .G(N00ADTZ), .S(N00ADUA));
nch_mac  XMAFGI ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADUC));
nch_mac  XMAFGG ( .D(N00ADTY), .B(gnd_), .G(N00ADTW), .S(N00ADTX));
nch_mac  XMAFGE ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADTY));
nch_mac  XMAFFM ( .D(gnd_), .B(gnd_), .G(N00ADTL), .S(N00ADTV));
nch_mac  XMAFFL ( .D(N00ADTV), .B(gnd_), .G(N00ADSN), .S(N00ADTP));
nch_mac  XMAFFJ ( .D(gnd_), .B(gnd_), .G(N00ADSN), .S(N00ADTR));
nch_mac  XMAFFH ( .D(N00ADTU), .B(gnd_), .G(N00ADTR), .S(N00ADTS));
nch_mac  XMAFFG ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADTU));
nch_mac  XMAFFE ( .D(N00ADTQ), .B(gnd_), .G(N00ADTO), .S(N00ADTP));
nch_mac  XMAFFC ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADTQ));
nch_mac  XMAFEK ( .D(gnd_), .B(gnd_), .G(N00ADTD), .S(N00ADTN));
nch_mac  XMAFEJ ( .D(N00ADTN), .B(gnd_), .G(N00ADSN), .S(N00ADTH));
nch_mac  XMAFEH ( .D(gnd_), .B(gnd_), .G(N00ADSN), .S(N00ADTJ));
nch_mac  XMAFEF ( .D(N00ADTM), .B(gnd_), .G(N00ADTJ), .S(N00ADTK));
nch_mac  XMAFEE ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADTM));
nch_mac  XMAFEC ( .D(N00ADTI), .B(gnd_), .G(N00ADTG), .S(N00ADTH));
nch_mac  XMAFEA ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADTI));
nch_mac  XMAFDI ( .D(gnd_), .B(gnd_), .G(N00ADSV), .S(N00ADTF));
nch_mac  XMAFDH ( .D(N00ADTF), .B(gnd_), .G(N00ADSN), .S(N00ADSZ));
nch_mac  XMAFDF ( .D(gnd_), .B(gnd_), .G(N00ADSN), .S(N00ADTB));
nch_mac  XMAFDD ( .D(N00ADTE), .B(gnd_), .G(N00ADTB), .S(N00ADTC));
nch_mac  XMAFDC ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADTE));
nch_mac  XMAFDA ( .D(N00ADTA), .B(gnd_), .G(N00ADSY), .S(N00ADSZ));
nch_mac  XMAFCY ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADTA));
nch_mac  XMAFCG ( .D(gnd_), .B(gnd_), .G(N00ADSK), .S(N00ADSX));
nch_mac  XMAFCF ( .D(N00ADSX), .B(gnd_), .G(N00ADSN), .S(N00ADSR));
nch_mac  XMAFCD ( .D(gnd_), .B(gnd_), .G(N00ADSN), .S(N00ADST));
nch_mac  XMAFCB ( .D(N00ADSW), .B(gnd_), .G(N00ADST), .S(N00ADSU));
nch_mac  XMAFCA ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADSW));
nch_mac  XMAFBY ( .D(N00ADSS), .B(gnd_), .G(N00ADSQ), .S(N00ADSR));
nch_mac  XMAFBW ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADSS));
nch_mac  XMAFBE ( .D(gnd_), .B(gnd_), .G(N00ADSM), .S(N00ADSO));
nch_mac  XMAFBD ( .D(N00ADSO), .B(gnd_), .G(N00ADSN), .S(N00ADSG));
nch_mac  XMAFBB ( .D(gnd_), .B(gnd_), .G(N00ADSN), .S(N00ADSI));
nch_mac  XMAFAZ ( .D(N00ADSL), .B(gnd_), .G(N00ADSI), .S(N00ADSJ));
nch_mac  XMAFAY ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADSL));
nch_mac  XMAFAW ( .D(N00ADSH), .B(gnd_), .G(N00ADSF), .S(N00ADSG));
nch_mac  XMAFAU ( .D(gnd_), .B(gnd_), .G(vdd_), .S(N00ADSH));
nch_mac  XMAFAQ ( .D(N00ADSD), .B(gnd_), .G(N00ADRP), .S(N00ADRM));
nch_mac  XMAFAP ( .D(gnd_), .B(gnd_), .G(N00ADSE), .S(N00ADSD));
nch_mac  XMAFAI ( .D(gnd_), .B(gnd_), .G(REF), .S(N00ADSA));
nch_mac  XMAFAH ( .D(N00ADSA), .B(gnd_), .G(N00ADRQ), .S(N00ADRL));
nch_mac  XMAFAG ( .D(N00ADRY), .B(gnd_), .G(N00ADRZ), .S(N00ADRL));
nch_mac  XMAFAA ( .D(gnd_), .B(gnd_), .G(N00ADRL), .S(N00ADRW));
nch_mac  XMAEZZ ( .D(N00ADRW), .B(gnd_), .G(N00ADRL), .S(N00ADRN));
nch_mac  XMAEZW ( .D(gnd_), .B(gnd_), .G(N00ADRO), .S(N00ADRU));
nch_mac  XMAEZV ( .D(N00ADRU), .B(gnd_), .G(N00ADRO), .S(N00ADRP));
nch_mac  XMAEZS ( .D(gnd_), .B(gnd_), .G(N00ADRN), .S(N00ADRS));
nch_mac  XMAEZR ( .D(N00ADRS), .B(gnd_), .G(N00ADRN), .S(N00ADRO));
nch_mac  XMAEZC ( .D(N00ADRI), .B(gnd_), .G(N00ADQU), .S(N00ADQR));
nch_mac  XMAEZB ( .D(gnd_), .B(gnd_), .G(N00ADRJ), .S(N00ADRI));
nch_mac  XMAEYU ( .D(gnd_), .B(gnd_), .G(FB), .S(N00ADRF));
nch_mac  XMAEYT ( .D(N00ADRF), .B(gnd_), .G(N00ADQV), .S(N00ADQQ));
nch_mac  XMAEYS ( .D(N00ADRC), .B(gnd_), .G(N00ADRE), .S(N00ADQQ));
nch_mac  XMAEYR ( .D(gnd_), .B(gnd_), .G(N00ADRD), .S(N00ADRC));
nch_mac  XMAEYM ( .D(gnd_), .B(gnd_), .G(N00ADQQ), .S(N00ADRA));
nch_mac  XMAEYL ( .D(N00ADRA), .B(gnd_), .G(N00ADQQ), .S(N00ADQS));
nch_mac  XMAEYI ( .D(gnd_), .B(gnd_), .G(N00ADQT), .S(N00ADQY));
nch_mac  XMAEYH ( .D(N00ADQY), .B(gnd_), .G(N00ADQT), .S(N00ADQU));
nch_mac  XMAEYE ( .D(gnd_), .B(gnd_), .G(N00ADQS), .S(N00ADQW));
nch_mac  XMAEYD ( .D(N00ADQW), .B(gnd_), .G(N00ADQS), .S(N00ADQT));
nch_mac  XMAEWV ( .D(gnd_), .B(gnd_), .G(N00AAAC), .S(N00AAAF));
nch_mac  XMAEWU ( .D(N00AAAE), .B(gnd_), .G(N00AAAC), .S(N00AAAB));
nch_mac  XMAEWR ( .D(gnd_), .B(gnd_), .G(N00AAAD), .S(N00AAAC));
nch_mac  XMAEWQ ( .D(gnd_), .B(gnd_), .G(N00AAAB), .S(VDDA));
nch_mac  XMAEWS ( .D(gnd_), .B(gnd_), .G(N00AAAA), .S(N00AAAD));
nch_mac  XMAEWT ( .D(N00AAAF), .B(gnd_), .G(N00AAAC), .S(N00AAAE));
rpodwo_m  XAGSM ( .MINUS(N00AEJS), .PLUS(N00ADZG), .BULK(vdd_));
pdio  DAGSK ( .PLUS(N00AEJS), .MINUS(vdd_));
pdio  DAFSP ( .PLUS(N00ADXS), .MINUS(VDDA));
pdio  DAFSF ( .PLUS(N00ADYE), .MINUS(VDDA));
pdio  DAFRV ( .PLUS(N00ADYA), .MINUS(VDDA));
pdio  DAFRL ( .PLUS(N00ADXR), .MINUS(VDDA));
pdio  DAGSL ( .PLUS(N00ADZG), .MINUS(vdd_));
rppolywo_m  XAFRB ( .MINUS(N00ADXF), .PLUS(N00ADXP), .BULK(VDDA));
rppolywo_m  XAFRA ( .MINUS(N00ADXF), .PLUS(N00ADYQ), .BULK(VDDA));
rppolywo_m  XAFQZ ( .MINUS(N00ADYQ), .PLUS(N00ADXN), .BULK(VDDA));
rppolywo_m  XAFQY ( .MINUS(N00ADXF), .PLUS(N00ADYP), .BULK(VDDA));
rppolywo_m  XAFQX ( .MINUS(N00ADYO), .PLUS(N00ADYN), .BULK(VDDA));
rppolywo_m  XAFQW ( .MINUS(N00ADYP), .PLUS(N00ADYO), .BULK(VDDA));
rppolywo_m  XAFQV ( .MINUS(N00ADYN), .PLUS(N00ADXL), .BULK(VDDA));
rppolywo_m  XAFQU ( .MINUS(N00ADXF), .PLUS(N00ADYK), .BULK(VDDA));
rppolywo_m  XAFQT ( .MINUS(N00ADYM), .PLUS(N00ADYI), .BULK(VDDA));
rppolywo_m  XAFQS ( .MINUS(N00ADYL), .PLUS(N00ADYM), .BULK(VDDA));
rppolywo_m  XAFQR ( .MINUS(N00ADYJ), .PLUS(N00ADYL), .BULK(VDDA));
rppolywo_m  XAFQQ ( .MINUS(N00ADYK), .PLUS(N00ADYJ), .BULK(VDDA));
rppolywo_m  XAFQP ( .MINUS(N00ADYI), .PLUS(N00ADXJ), .BULK(VDDA));
rppolywo_m  XAEXG ( .MINUS(N00AAAK), .PLUS(N00AAAJ), .BULK(gnd_));
rppolywo_m  XAEXD ( .MINUS(VDDA), .PLUS(N00AAAI), .BULK(gnd_));
rppolywo_m  XAEXE ( .MINUS(N00AAAJ), .PLUS(N00AAAA), .BULK(gnd_));
rppolywo_m  XAEXF ( .MINUS(N00AAAI), .PLUS(N00AAAK), .BULK(gnd_));

endmodule
// Library - io, Cell - PVDD1DGZ_G, View - schematic
// LAST TIME SAVED: Sep  3 14:17:09 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module PVDD1DGZ_G ( VDD );
inout  VDD;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD2DGZ_G, View - schematic
// LAST TIME SAVED: Sep  3 14:16:20 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module PVDD2DGZ_G ( VDDPST );
inout  VDDPST;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD2POC_G, View - schematic
// LAST TIME SAVED: Sep  3 14:39:22 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module PVDD2POC_G ( POC, VDDPST );
output  POC;

inout  VDDPST;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVSS3DGZ_G, View - schematic
// LAST TIME SAVED: Sep 17 14:47:58 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module PVSS3DGZ_G ( VDDPST, VSS );
inout  VDDPST, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - ice1chip, Cell - IO_lft_bank_ice1f_v2, View - schematic
// LAST TIME SAVED: Apr 20 16:04:40 2011
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module IO_lft_bank_ice1f_v2 ( in, pll_lock, pllout, pad, ien, lvds_en,
     oen, out, pll_bypass, pll_cbit, pll_fb, pll_fse, pll_ref,
     pll_reset, ren, vdda );
output  pll_lock, pllout;


input  pll_bypass, pll_fb, pll_fse, pll_ref, pll_reset, vdda;

output [23:0]  in;

inout [23:0]  pad;

input [23:0]  ien;
input [23:0]  oen;
input [23:0]  ren;
input [11:0]  lvds_en;
input [23:0]  out;
input [16:0]  pll_cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  ienb;



PLVDS_pair plvds_1_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[2]), .oen_n(oen[3]),
     .PAD_n(pad[3]), .c_p(in[2]), .c_n(in[3]), .PAD_p(pad[2]),
     .i_n(out[3]), .i_p(out[2]), .cbit({lvds_en[1], ienb[2], ienb[3],
     ren[2], ren[3]}));
PLVDS_pair plvds_0_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[0]), .oen_n(oen[1]),
     .PAD_n(pad[1]), .c_p(in[0]), .c_n(in[1]), .PAD_p(pad[0]),
     .i_n(out[1]), .i_p(out[0]), .cbit({lvds_en[0], ienb[0], ienb[1],
     ren[0], ren[1]}));
PLVDS_pair plvds2 ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[4]), .oen_n(oen[5]),
     .PAD_n(pad[5]), .c_p(in[4]), .c_n(in[5]), .PAD_p(pad[4]),
     .i_n(out[5]), .i_p(out[4]), .cbit({lvds_en[2], ienb[4], ienb[5],
     ren[4], ren[5]}));
PLVDS_pair plvds_5_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[10]), .oen_n(oen[11]),
     .PAD_n(pad[11]), .c_p(in[10]), .c_n(in[11]), .PAD_p(pad[10]),
     .i_n(out[11]), .i_p(out[10]), .cbit({lvds_en[5], ienb[10],
     ienb[11], ren[10], ren[11]}));
PLVDS_pair plvds_4_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[8]), .oen_n(oen[9]),
     .PAD_n(pad[9]), .c_p(in[8]), .c_n(in[9]), .PAD_p(pad[8]),
     .i_n(out[9]), .i_p(out[8]), .cbit({lvds_en[4], ienb[8], ienb[9],
     ren[8], ren[9]}));
PLVDS_pair plvds_3_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[6]), .oen_n(oen[7]),
     .PAD_n(pad[7]), .c_p(in[6]), .c_n(in[7]), .PAD_p(pad[6]),
     .i_n(out[7]), .i_p(out[6]), .cbit({lvds_en[3], ienb[6], ienb[7],
     ren[6], ren[7]}));
PLVDS_pair plvds6 ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[12]), .oen_n(oen[13]),
     .PAD_n(pad[13]), .c_p(in[12]), .c_n(in[13]), .PAD_p(pad[12]),
     .i_n(out[13]), .i_p(out[12]), .cbit({lvds_en[6], ienb[12],
     ienb[13], ren[12], ren[13]}));
PLVDS_pair plvds_9_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[18]), .oen_n(oen[19]),
     .PAD_n(pad[19]), .c_p(in[18]), .c_n(in[19]), .PAD_p(pad[18]),
     .i_n(out[19]), .i_p(out[18]), .cbit({lvds_en[9], ienb[18],
     ienb[19], ren[18], ren[19]}));
PLVDS_pair plvds_8_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[16]), .oen_n(oen[17]),
     .PAD_n(pad[17]), .c_p(in[16]), .c_n(in[17]), .PAD_p(pad[16]),
     .i_n(out[17]), .i_p(out[16]), .cbit({lvds_en[8], ienb[16],
     ienb[17], ren[16], ren[17]}));
PLVDS_pair plvds_7_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[14]), .oen_n(oen[15]),
     .PAD_n(pad[15]), .c_p(in[14]), .c_n(in[15]), .PAD_p(pad[14]),
     .i_n(out[15]), .i_p(out[14]), .cbit({lvds_en[7], ienb[14],
     ienb[15], ren[14], ren[15]}));
PLVDS_pair plvds_11_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[22]), .oen_n(oen[23]),
     .PAD_n(pad[23]), .c_p(in[22]), .c_n(in[23]), .PAD_p(pad[22]),
     .i_n(out[23]), .i_p(out[22]), .cbit({lvds_en[11], ienb[22],
     ienb[23], ren[22], ren[23]}));
PLVDS_pair plvds_10_ ( .tiegnd(tiegnd_lftpad), .POC(poc_lft),
     .vddio(vddio_leftbank), .oen_p(oen[20]), .oen_n(oen[21]),
     .PAD_n(pad[21]), .c_p(in[20]), .c_n(in[21]), .PAD_p(pad[20]),
     .i_n(out[21]), .i_p(out[20]), .cbit({lvds_en[10], ienb[20],
     ienb[21], ren[20], ren[21]}));
ABIWTCZ4 Ipll_bot ( .RESET(pll_reset), .REF(pll_ref),
     .RANGE2(pll_cbit[16]), .RANGE1(pll_cbit[15]),
     .RANGE0(pll_cbit[14]), .FSE(pll_fse), .FB(pll_fb),
     .DIVR3(pll_cbit[3]), .DIVR2(pll_cbit[2]), .DIVR1(pll_cbit[1]),
     .DIVR0(pll_cbit[0]), .DIVQ2(pll_cbit[13]), .DIVQ1(pll_cbit[12]),
     .DIVQ0(pll_cbit[11]), .DIVF5(pll_cbit[9]), .DIVF4(pll_cbit[8]),
     .DIVF3(pll_cbit[7]), .DIVF2(pll_cbit[6]), .DIVF1(pll_cbit[5]),
     .DIVF0(pll_cbit[4]), .BYPASS(pll_bypass), .PLLOUT(pllout),
     .LOCK(pll_lock), .VDDA(vdda), .DIVF6(pll_cbit[10]));
tielo4x I119 ( .tielo(tiegnd_lftpad));
inv_hvt I120_23_ ( .A(ien[23]), .Y(ienb[23]));
inv_hvt I120_22_ ( .A(ien[22]), .Y(ienb[22]));
inv_hvt I120_21_ ( .A(ien[21]), .Y(ienb[21]));
inv_hvt I120_20_ ( .A(ien[20]), .Y(ienb[20]));
inv_hvt I120_19_ ( .A(ien[19]), .Y(ienb[19]));
inv_hvt I120_18_ ( .A(ien[18]), .Y(ienb[18]));
inv_hvt I120_17_ ( .A(ien[17]), .Y(ienb[17]));
inv_hvt I120_16_ ( .A(ien[16]), .Y(ienb[16]));
inv_hvt I120_15_ ( .A(ien[15]), .Y(ienb[15]));
inv_hvt I120_14_ ( .A(ien[14]), .Y(ienb[14]));
inv_hvt I120_13_ ( .A(ien[13]), .Y(ienb[13]));
inv_hvt I120_12_ ( .A(ien[12]), .Y(ienb[12]));
inv_hvt I120_11_ ( .A(ien[11]), .Y(ienb[11]));
inv_hvt I120_10_ ( .A(ien[10]), .Y(ienb[10]));
inv_hvt I120_9_ ( .A(ien[9]), .Y(ienb[9]));
inv_hvt I120_8_ ( .A(ien[8]), .Y(ienb[8]));
inv_hvt I120_7_ ( .A(ien[7]), .Y(ienb[7]));
inv_hvt I120_6_ ( .A(ien[6]), .Y(ienb[6]));
inv_hvt I120_5_ ( .A(ien[5]), .Y(ienb[5]));
inv_hvt I120_4_ ( .A(ien[4]), .Y(ienb[4]));
inv_hvt I120_3_ ( .A(ien[3]), .Y(ienb[3]));
inv_hvt I120_2_ ( .A(ien[2]), .Y(ienb[2]));
inv_hvt I120_1_ ( .A(ien[1]), .Y(ienb[1]));
inv_hvt I120_0_ ( .A(ien[0]), .Y(ienb[0]));
PVDD1DGZ_G I129 ( .VDD(vdd_));
PVDD1DGZ_G I126_1_ ( .VDD(vdd_));
PVDD1DGZ_G I126_0_ ( .VDD(vdd_));
PVDD2DGZ_G I128 ( .VDDPST(vddio_leftbank));
PVDD2DGZ_G I121 ( .VDDPST(vddio_leftbank));
PVDD2DGZ_G I130 ( .VDDPST(vddio_leftbank));
PVDD2POC_G I122 ( .VDDPST(vddio_leftbank), .POC(poc_lft));
PVSS3DGZ_G gndummy12_1_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G gndummy12_0_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I123_1_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I123_0_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I127_1_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));
PVSS3DGZ_G I127_0_ ( .VSS(gnd_), .VDDPST(vddio_leftbank));

endmodule
// Library - misc, Cell - vpp_clamp_finger, View - schematic
// LAST TIME SAVED: Sep 17 15:01:43 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module vpp_clamp_finger ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .B(VSS), .D(net12), .G(VSS), .S(VSS));
nch_25  m1 ( .B(VSS), .D(VPP), .G(VDDIO), .S(net12));

endmodule
// Library - misc, Cell - vpp_clamp, View - schematic
// LAST TIME SAVED: Sep 17 14:58:48 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module vpp_clamp ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vpp_clamp_finger I0_3_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_2_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_1_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0_0_ ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));

endmodule
// Library - leafcell, Cell - sbox11to9_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:52:20 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox11to9_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  b;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r10 ( .prog(prog), .in6(b[4]), .in5(b[10]), .in4(l[2]),
     .in3(l[10]), .in2(l[7]), .in1(t[10]), .in0(t[5]), .out(r[10]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b10 ( .prog(prog), .in6(l[4]), .in5(l[10]), .in4(t[2]),
     .in3(t[10]), .in2(t[7]), .in1(r[10]), .in0(r[5]), .out(b[10]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b11 ( .prog(prog), .in6(l[5]), .in5(l[11]), .in4(t[3]),
     .in3(t[11]), .in2(t[8]), .in1(r[11]), .in0(r[6]), .out(b[11]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b9 ( .prog(prog), .in6(l[3]), .in5(l[9]), .in4(t[1]),
     .in3(t[9]), .in2(t[6]), .in1(r[9]), .in0(r[4]), .out(b[9]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r11 ( .prog(prog), .in6(b[5]), .in5(b[11]), .in4(l[3]),
     .in3(l[11]), .in2(l[8]), .in1(t[11]), .in0(t[6]), .out(r[11]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r9 ( .prog(prog), .in6(b[3]), .in5(b[9]), .in4(l[1]),
     .in3(l[9]), .in2(l[6]), .in1(t[9]), .in0(t[4]), .out(r[9]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - io, Cell - pvpp, View - schematic
// LAST TIME SAVED: Oct  4 15:01:12 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module pvpp ( vpp, vppin );
inout  vpp, vppin;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I60_15_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_14_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_13_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_12_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_11_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_10_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_9_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_8_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_7_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_6_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_5_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_4_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_3_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_2_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_1_ ( .vddp_tieh(vddio_in));
vddp_tiehigh I60_0_ ( .vddp_tieh(vddio_in));
rppolywo_m  R1 ( .MINUS(vpp), .PLUS(vppin), .BULK(gnd_));
vpp_clamp I59_15_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_14_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_13_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_12_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_11_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_10_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_9_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_8_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_7_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_6_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_5_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_4_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_3_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_2_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_1_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));
vpp_clamp I59_0_ ( .VSS(gnd_), .VDDIO(vddio_in), .VPP(vpp));

endmodule
// Library - ice1chip, Cell - IO_top_bank_ice1f, View - schematic
// LAST TIME SAVED: Apr 14 09:34:35 2011
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module IO_top_bank_ice1f ( in, pad, vpp, vppin, ien, oen, out, ren );

inout  vpp, vppin;


output [23:0]  in;

inout [23:0]  pad;

input [23:0]  out;
input [23:0]  ren;
input [23:0]  oen;
input [23:0]  ien;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net143;

wire  [10:0]  net217;

wire  [5:0]  net0166;

wire  [3:0]  net223;

wire  [23:0]  n_ienb;



tielo4x tielo4x_t ( .tielo(tiegnd_toppad));
pvpp vppfast_t ( .vppin(vppin), .vpp(vpp));
inv_hvt ien_inv_23_ ( .A(ien[23]), .Y(n_ienb[23]));
inv_hvt ien_inv_22_ ( .A(ien[22]), .Y(n_ienb[22]));
inv_hvt ien_inv_21_ ( .A(ien[21]), .Y(n_ienb[21]));
inv_hvt ien_inv_20_ ( .A(ien[20]), .Y(n_ienb[20]));
inv_hvt ien_inv_19_ ( .A(ien[19]), .Y(n_ienb[19]));
inv_hvt ien_inv_18_ ( .A(ien[18]), .Y(n_ienb[18]));
inv_hvt ien_inv_17_ ( .A(ien[17]), .Y(n_ienb[17]));
inv_hvt ien_inv_16_ ( .A(ien[16]), .Y(n_ienb[16]));
inv_hvt ien_inv_15_ ( .A(ien[15]), .Y(n_ienb[15]));
inv_hvt ien_inv_14_ ( .A(ien[14]), .Y(n_ienb[14]));
inv_hvt ien_inv_13_ ( .A(ien[13]), .Y(n_ienb[13]));
inv_hvt ien_inv_12_ ( .A(ien[12]), .Y(n_ienb[12]));
inv_hvt ien_inv_11_ ( .A(ien[11]), .Y(n_ienb[11]));
inv_hvt ien_inv_10_ ( .A(ien[10]), .Y(n_ienb[10]));
inv_hvt ien_inv_9_ ( .A(ien[9]), .Y(n_ienb[9]));
inv_hvt ien_inv_8_ ( .A(ien[8]), .Y(n_ienb[8]));
inv_hvt ien_inv_7_ ( .A(ien[7]), .Y(n_ienb[7]));
inv_hvt ien_inv_6_ ( .A(ien[6]), .Y(n_ienb[6]));
inv_hvt ien_inv_5_ ( .A(ien[5]), .Y(n_ienb[5]));
inv_hvt ien_inv_4_ ( .A(ien[4]), .Y(n_ienb[4]));
inv_hvt ien_inv_3_ ( .A(ien[3]), .Y(n_ienb[3]));
inv_hvt ien_inv_2_ ( .A(ien[2]), .Y(n_ienb[2]));
inv_hvt ien_inv_1_ ( .A(ien[1]), .Y(n_ienb[1]));
inv_hvt ien_inv_0_ ( .A(ien[0]), .Y(n_ienb[0]));
PVDD1DGZ_G vdd12_t_1_ ( .VDD(vdd_));
PVDD1DGZ_G vdd12_t_0_ ( .VDD(vdd_));
PVDD2POC_G vddio_poc2_t ( .VDDPST(vddio_topbank), .POC(poc_top));
PVDD2DGZ_G vcciodummy12_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vcciodummy12_0_ ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vddio1_t ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vddio34_t_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ_G vddio34_t_0_ ( .VDDPST(vddio_topbank));
PVSS3DGZ_G gnddummy12_1_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnddummy12_0_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnddummy34_1_ ( .VSS(gnd_), .VDDPST(vddp_));
PVSS3DGZ_G gnddummy34_0_ ( .VSS(gnd_), .VDDPST(vddp_));
PVSS3DGZ_G gnd23_t_1_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnd23_t_0_ ( .VSS(gnd_), .VDDPST(vddio_topbank));
PVSS3DGZ_G gnd1_t ( .VSS(gnd_), .VDDPST(vddio_topbank));
PDUW08SDGZ_G_NOR pad_t_10_ ( .REN(ren[10]), .C(in[10]), .OEN(oen[10]),
     .IE(n_ienb[10]), .I(out[10]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net173), .VDDIO(vddio_topbank), .PAD(pad[10]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_12_ ( .REN(ren[12]), .C(in[12]), .OEN(oen[12]),
     .IE(n_ienb[12]), .I(out[12]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net143[0]), .VDDIO(vddio_topbank), .PAD(pad[12]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_11_ ( .REN(ren[11]), .C(in[11]), .OEN(oen[11]),
     .IE(n_ienb[11]), .I(out[11]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net143[1]), .VDDIO(vddio_topbank), .PAD(pad[11]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_23_ ( .REN(ren[23]), .C(in[23]), .OEN(oen[23]),
     .IE(n_ienb[23]), .I(out[23]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[0]), .VDDIO(vddio_topbank), .PAD(pad[23]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_22_ ( .REN(ren[22]), .C(in[22]), .OEN(oen[22]),
     .IE(n_ienb[22]), .I(out[22]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[1]), .VDDIO(vddio_topbank), .PAD(pad[22]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_21_ ( .REN(ren[21]), .C(in[21]), .OEN(oen[21]),
     .IE(n_ienb[21]), .I(out[21]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[2]), .VDDIO(vddio_topbank), .PAD(pad[21]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_20_ ( .REN(ren[20]), .C(in[20]), .OEN(oen[20]),
     .IE(n_ienb[20]), .I(out[20]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[3]), .VDDIO(vddio_topbank), .PAD(pad[20]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_19_ ( .REN(ren[19]), .C(in[19]), .OEN(oen[19]),
     .IE(n_ienb[19]), .I(out[19]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[4]), .VDDIO(vddio_topbank), .PAD(pad[19]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_18_ ( .REN(ren[18]), .C(in[18]), .OEN(oen[18]),
     .IE(n_ienb[18]), .I(out[18]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[5]), .VDDIO(vddio_topbank), .PAD(pad[18]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_17_ ( .REN(ren[17]), .C(in[17]), .OEN(oen[17]),
     .IE(n_ienb[17]), .I(out[17]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[6]), .VDDIO(vddio_topbank), .PAD(pad[17]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_16_ ( .REN(ren[16]), .C(in[16]), .OEN(oen[16]),
     .IE(n_ienb[16]), .I(out[16]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[7]), .VDDIO(vddio_topbank), .PAD(pad[16]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_15_ ( .REN(ren[15]), .C(in[15]), .OEN(oen[15]),
     .IE(n_ienb[15]), .I(out[15]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[8]), .VDDIO(vddio_topbank), .PAD(pad[15]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_14_ ( .REN(ren[14]), .C(in[14]), .OEN(oen[14]),
     .IE(n_ienb[14]), .I(out[14]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[9]), .VDDIO(vddio_topbank), .PAD(pad[14]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_13_ ( .REN(ren[13]), .C(in[13]), .OEN(oen[13]),
     .IE(n_ienb[13]), .I(out[13]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net217[10]), .VDDIO(vddio_topbank), .PAD(pad[13]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_3_ ( .REN(ren[3]), .C(in[3]), .OEN(oen[3]),
     .IE(n_ienb[3]), .I(out[3]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[0]), .VDDIO(vddio_topbank), .PAD(pad[3]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_2_ ( .REN(ren[2]), .C(in[2]), .OEN(oen[2]),
     .IE(n_ienb[2]), .I(out[2]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[1]), .VDDIO(vddio_topbank), .PAD(pad[2]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_1_ ( .REN(ren[1]), .C(in[1]), .OEN(oen[1]),
     .IE(n_ienb[1]), .I(out[1]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[2]), .VDDIO(vddio_topbank), .PAD(pad[1]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_0_ ( .REN(ren[0]), .C(in[0]), .OEN(oen[0]),
     .IE(n_ienb[0]), .I(out[0]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net223[3]), .VDDIO(vddio_topbank), .PAD(pad[0]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_9_ ( .REN(ren[9]), .C(in[9]), .OEN(oen[9]),
     .IE(n_ienb[9]), .I(out[9]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[0]), .VDDIO(vddio_topbank), .PAD(pad[9]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_8_ ( .REN(ren[8]), .C(in[8]), .OEN(oen[8]),
     .IE(n_ienb[8]), .I(out[8]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[1]), .VDDIO(vddio_topbank), .PAD(pad[8]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_7_ ( .REN(ren[7]), .C(in[7]), .OEN(oen[7]),
     .IE(n_ienb[7]), .I(out[7]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[2]), .VDDIO(vddio_topbank), .PAD(pad[7]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_6_ ( .REN(ren[6]), .C(in[6]), .OEN(oen[6]),
     .IE(n_ienb[6]), .I(out[6]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[3]), .VDDIO(vddio_topbank), .PAD(pad[6]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_5_ ( .REN(ren[5]), .C(in[5]), .OEN(oen[5]),
     .IE(n_ienb[5]), .I(out[5]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[4]), .VDDIO(vddio_topbank), .PAD(pad[5]),
     .POC(poc_top));
PDUW08SDGZ_G_NOR pad_t_4_ ( .REN(ren[4]), .C(in[4]), .OEN(oen[4]),
     .IE(n_ienb[4]), .I(out[4]), .indiff(tiegnd_toppad),
     .PAD4LVDS(net0166[5]), .VDDIO(vddio_topbank), .PAD(pad[4]),
     .POC(poc_top));

endmodule
// Library - TSMC_IO, Cell - PDDW08SDGZ_G, View - schematic
// LAST TIME SAVED: Oct  4 08:25:43 2010
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module PDDW08SDGZ_G ( C, PAD, I, OEN, POC, REN, VDDIO );
output  C;

inout  PAD;

input  I, OEN, POC, REN, VDDIO;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - ice1chip, Cell - IO_rgt_bank_ice1f, View - schematic
// LAST TIME SAVED: Apr 14 09:34:07 2011
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module IO_rgt_bank_ice1f ( in, trstb_int, pad, TRSTb, ien, oen, out,
     ren );
output  trstb_int;


input  TRSTb;

output [24:0]  in;

inout [24:0]  pad;

input [24:0]  ien;
input [24:0]  oen;
input [25:0]  ren;
input [24:0]  out;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:0]  net144;

wire  [1:0]  net110;

wire  [1:0]  net154;

wire  [3:0]  net134;

wire  [3:0]  net115;

wire  [3:0]  net164;

wire  [1:0]  net117;

wire  [24:0]  n_ienb;

wire  [1:0]  net184;



tielo4x tielo4x_r ( .tielo(tiegnd_rgtpad));
tiehi4x tiehi4x_r ( .tiehi(tievdd_rgtpad));
inv_hvt I_ien_inv_24_ ( .A(ien[24]), .Y(n_ienb[24]));
inv_hvt I_ien_inv_23_ ( .A(ien[23]), .Y(n_ienb[23]));
inv_hvt I_ien_inv_22_ ( .A(ien[22]), .Y(n_ienb[22]));
inv_hvt I_ien_inv_21_ ( .A(ien[21]), .Y(n_ienb[21]));
inv_hvt I_ien_inv_20_ ( .A(ien[20]), .Y(n_ienb[20]));
inv_hvt I_ien_inv_19_ ( .A(ien[19]), .Y(n_ienb[19]));
inv_hvt I_ien_inv_18_ ( .A(ien[18]), .Y(n_ienb[18]));
inv_hvt I_ien_inv_17_ ( .A(ien[17]), .Y(n_ienb[17]));
inv_hvt I_ien_inv_16_ ( .A(ien[16]), .Y(n_ienb[16]));
inv_hvt I_ien_inv_15_ ( .A(ien[15]), .Y(n_ienb[15]));
inv_hvt I_ien_inv_14_ ( .A(ien[14]), .Y(n_ienb[14]));
inv_hvt I_ien_inv_13_ ( .A(ien[13]), .Y(n_ienb[13]));
inv_hvt I_ien_inv_12_ ( .A(ien[12]), .Y(n_ienb[12]));
inv_hvt I_ien_inv_11_ ( .A(ien[11]), .Y(n_ienb[11]));
inv_hvt I_ien_inv_10_ ( .A(ien[10]), .Y(n_ienb[10]));
inv_hvt I_ien_inv_9_ ( .A(ien[9]), .Y(n_ienb[9]));
inv_hvt I_ien_inv_8_ ( .A(ien[8]), .Y(n_ienb[8]));
inv_hvt I_ien_inv_7_ ( .A(ien[7]), .Y(n_ienb[7]));
inv_hvt I_ien_inv_6_ ( .A(ien[6]), .Y(n_ienb[6]));
inv_hvt I_ien_inv_5_ ( .A(ien[5]), .Y(n_ienb[5]));
inv_hvt I_ien_inv_4_ ( .A(ien[4]), .Y(n_ienb[4]));
inv_hvt I_ien_inv_3_ ( .A(ien[3]), .Y(n_ienb[3]));
inv_hvt I_ien_inv_2_ ( .A(ien[2]), .Y(n_ienb[2]));
inv_hvt I_ien_inv_1_ ( .A(ien[1]), .Y(n_ienb[1]));
inv_hvt I_ien_inv_0_ ( .A(ien[0]), .Y(n_ienb[0]));
PDDW08SDGZ_G trstb_r ( .REN(ren[25]), .C(trstb_int),
     .OEN(tievdd_rgtpad), .I(tiegnd_rgtpad), .VDDIO(vddio_rgtbank),
     .PAD(TRSTb), .POC(poc_rgt));
PVDD1DGZ_G vdd12_r_1_ ( .VDD(vdd_));
PVDD1DGZ_G vdd12_r_0_ ( .VDD(vdd_));
PDUW08SDGZ_G_NOR pad_r_13_ ( .REN(ren[13]), .C(in[13]), .OEN(oen[13]),
     .IE(n_ienb[13]), .I(out[13]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net154[0]), .VDDIO(vddio_rgtbank), .PAD(pad[13]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_12_ ( .REN(ren[12]), .C(in[12]), .OEN(oen[12]),
     .IE(n_ienb[12]), .I(out[12]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net154[1]), .VDDIO(vddio_rgtbank), .PAD(pad[12]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_7_ ( .REN(ren[7]), .C(in[7]), .OEN(oen[7]),
     .IE(n_ienb[7]), .I(out[7]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[0]), .VDDIO(vddio_rgtbank), .PAD(pad[7]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_6_ ( .REN(ren[6]), .C(in[6]), .OEN(oen[6]),
     .IE(n_ienb[6]), .I(out[6]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[1]), .VDDIO(vddio_rgtbank), .PAD(pad[6]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_5_ ( .REN(ren[5]), .C(in[5]), .OEN(oen[5]),
     .IE(n_ienb[5]), .I(out[5]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[2]), .VDDIO(vddio_rgtbank), .PAD(pad[5]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_4_ ( .REN(ren[4]), .C(in[4]), .OEN(oen[4]),
     .IE(n_ienb[4]), .I(out[4]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net164[3]), .VDDIO(vddio_rgtbank), .PAD(pad[4]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_3_ ( .REN(ren[3]), .C(in[3]), .OEN(oen[3]),
     .IE(n_ienb[3]), .I(out[3]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[0]), .VDDIO(vddio_rgtbank), .PAD(pad[3]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_2_ ( .REN(ren[2]), .C(in[2]), .OEN(oen[2]),
     .IE(n_ienb[2]), .I(out[2]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[1]), .VDDIO(vddio_rgtbank), .PAD(pad[2]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_1_ ( .REN(ren[1]), .C(in[1]), .OEN(oen[1]),
     .IE(n_ienb[1]), .I(out[1]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[2]), .VDDIO(vddio_rgtbank), .PAD(pad[1]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_0_ ( .REN(ren[0]), .C(in[0]), .OEN(oen[0]),
     .IE(n_ienb[0]), .I(out[0]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net115[3]), .VDDIO(vddio_rgtbank), .PAD(pad[0]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_9_ ( .REN(ren[9]), .C(in[9]), .OEN(oen[9]),
     .IE(n_ienb[9]), .I(out[9]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net184[0]), .VDDIO(vddio_rgtbank), .PAD(pad[9]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_8_ ( .REN(ren[8]), .C(in[8]), .OEN(oen[8]),
     .IE(n_ienb[8]), .I(out[8]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net184[1]), .VDDIO(vddio_rgtbank), .PAD(pad[8]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_11_ ( .REN(ren[11]), .C(in[11]), .OEN(oen[11]),
     .IE(n_ienb[11]), .I(out[11]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net117[0]), .VDDIO(vddio_rgtbank), .PAD(pad[11]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_10_ ( .REN(ren[10]), .C(in[10]), .OEN(oen[10]),
     .IE(n_ienb[10]), .I(out[10]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net117[1]), .VDDIO(vddio_rgtbank), .PAD(pad[10]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_24_ ( .REN(ren[24]), .C(in[24]), .OEN(oen[24]),
     .IE(n_ienb[24]), .I(out[24]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[0]), .VDDIO(vddio_rgtbank), .PAD(pad[24]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_23_ ( .REN(ren[23]), .C(in[23]), .OEN(oen[23]),
     .IE(n_ienb[23]), .I(out[23]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[1]), .VDDIO(vddio_rgtbank), .PAD(pad[23]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_22_ ( .REN(ren[22]), .C(in[22]), .OEN(oen[22]),
     .IE(n_ienb[22]), .I(out[22]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[2]), .VDDIO(vddio_rgtbank), .PAD(pad[22]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_21_ ( .REN(ren[21]), .C(in[21]), .OEN(oen[21]),
     .IE(n_ienb[21]), .I(out[21]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net134[3]), .VDDIO(vddio_rgtbank), .PAD(pad[21]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_18_ ( .REN(ren[18]), .C(in[18]), .OEN(oen[18]),
     .IE(n_ienb[18]), .I(out[18]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[0]), .VDDIO(vddio_rgtbank), .PAD(pad[18]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_17_ ( .REN(ren[17]), .C(in[17]), .OEN(oen[17]),
     .IE(n_ienb[17]), .I(out[17]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[1]), .VDDIO(vddio_rgtbank), .PAD(pad[17]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_16_ ( .REN(ren[16]), .C(in[16]), .OEN(oen[16]),
     .IE(n_ienb[16]), .I(out[16]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[2]), .VDDIO(vddio_rgtbank), .PAD(pad[16]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_15_ ( .REN(ren[15]), .C(in[15]), .OEN(oen[15]),
     .IE(n_ienb[15]), .I(out[15]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[3]), .VDDIO(vddio_rgtbank), .PAD(pad[15]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_14_ ( .REN(ren[14]), .C(in[14]), .OEN(oen[14]),
     .IE(n_ienb[14]), .I(out[14]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net144[4]), .VDDIO(vddio_rgtbank), .PAD(pad[14]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_20_ ( .REN(ren[20]), .C(in[20]), .OEN(oen[20]),
     .IE(n_ienb[20]), .I(out[20]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net110[0]), .VDDIO(vddio_rgtbank), .PAD(pad[20]),
     .POC(poc_rgt));
PDUW08SDGZ_G_NOR pad_r_19_ ( .REN(ren[19]), .C(in[19]), .OEN(oen[19]),
     .IE(n_ienb[19]), .I(out[19]), .indiff(tiegnd_rgtpad),
     .PAD4LVDS(net110[1]), .VDDIO(vddio_rgtbank), .PAD(pad[19]),
     .POC(poc_rgt));
PVDD2DGZ_G vcciodummy2 ( .VDDPST(vddp_));
PVDD2DGZ_G vddio12_r_1_ ( .VDDPST(vddio_rgtbank));
PVDD2DGZ_G vddio12_r_0_ ( .VDDPST(vddio_rgtbank));
PVDD2DGZ_G vddio2_r ( .VDDPST(vddio_rgtbank));
PVDD2DGZ_G vcciodummy1 ( .VDDPST(vddio_rgtbank));
PVDD2POC_G vddpoc_r ( .VDDPST(vddio_rgtbank), .POC(poc_rgt));
PVDD2POC_G vppv25_r ( .VDDPST(vddp_), .POC(net0123));
PVSS3DGZ_G gnd23_r_1_ ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnd23_r_0_ ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnddummy2 ( .VSS(gnd_), .VDDPST(vddp_));
PVSS3DGZ_G gnddummy1 ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnd3_r ( .VSS(gnd_), .VDDPST(vddio_rgtbank));
PVSS3DGZ_G gnd1_r ( .VSS(gnd_), .VDDPST(vddio_rgtbank));

endmodule
// Library - ice1chip, Cell - IO_bot_bank_ice1f, View - schematic
// LAST TIME SAVED: Apr 11 15:56:28 2011
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module IO_bot_bank_ice1f ( cdone_int, ctst_b_int, in, vddio_bottombank,
     vddio_spi, cdone, pad, cdone_out, ctst_b, ien, oen, out, ren );
output  cdone_int, ctst_b_int, vddio_bottombank, vddio_spi;

inout  cdone;

input  cdone_out, ctst_b;

output [23:0]  in;

inout [23:0]  pad;

input [23:0]  ien;
input [23:0]  out;
input [23:0]  oen;
input [23:0]  ren;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net188;

wire  [1:0]  net168;

wire  [7:0]  net241;

wire  [4:0]  net228;

wire  [1:0]  net237;

wire  [1:0]  net236;

wire  [1:0]  net234;

wire  [23:0]  n_ienb;



tiehi4x tiehi4x ( .tiehi(tievdd_botpad));
tielo4x tielo4x ( .tielo(tiegnd_botpad));
inv_hvt I_ien_inv_23_ ( .A(ien[23]), .Y(n_ienb[23]));
inv_hvt I_ien_inv_22_ ( .A(ien[22]), .Y(n_ienb[22]));
inv_hvt I_ien_inv_21_ ( .A(ien[21]), .Y(n_ienb[21]));
inv_hvt I_ien_inv_20_ ( .A(ien[20]), .Y(n_ienb[20]));
inv_hvt I_ien_inv_19_ ( .A(ien[19]), .Y(n_ienb[19]));
inv_hvt I_ien_inv_18_ ( .A(ien[18]), .Y(n_ienb[18]));
inv_hvt I_ien_inv_17_ ( .A(ien[17]), .Y(n_ienb[17]));
inv_hvt I_ien_inv_16_ ( .A(ien[16]), .Y(n_ienb[16]));
inv_hvt I_ien_inv_15_ ( .A(ien[15]), .Y(n_ienb[15]));
inv_hvt I_ien_inv_14_ ( .A(ien[14]), .Y(n_ienb[14]));
inv_hvt I_ien_inv_13_ ( .A(ien[13]), .Y(n_ienb[13]));
inv_hvt I_ien_inv_12_ ( .A(ien[12]), .Y(n_ienb[12]));
inv_hvt I_ien_inv_11_ ( .A(ien[11]), .Y(n_ienb[11]));
inv_hvt I_ien_inv_10_ ( .A(ien[10]), .Y(n_ienb[10]));
inv_hvt I_ien_inv_9_ ( .A(ien[9]), .Y(n_ienb[9]));
inv_hvt I_ien_inv_8_ ( .A(ien[8]), .Y(n_ienb[8]));
inv_hvt I_ien_inv_7_ ( .A(ien[7]), .Y(n_ienb[7]));
inv_hvt I_ien_inv_6_ ( .A(ien[6]), .Y(n_ienb[6]));
inv_hvt I_ien_inv_5_ ( .A(ien[5]), .Y(n_ienb[5]));
inv_hvt I_ien_inv_4_ ( .A(ien[4]), .Y(n_ienb[4]));
inv_hvt I_ien_inv_3_ ( .A(ien[3]), .Y(n_ienb[3]));
inv_hvt I_ien_inv_2_ ( .A(ien[2]), .Y(n_ienb[2]));
inv_hvt I_ien_inv_1_ ( .A(ien[1]), .Y(n_ienb[1]));
inv_hvt I_ien_inv_0_ ( .A(ien[0]), .Y(n_ienb[0]));
PVDD1DGZ_G vdd12_b_1_ ( .VDD(vdd_));
PVDD1DGZ_G vdd12_b_0_ ( .VDD(vdd_));
PVDD2POC_G vddiopoc2_b ( .VDDPST(vddio_bottombank), .POC(poc_bot));
PVDD2POC_G pvdd2poc_g_spivcc ( .VDDPST(vddio_spi), .POC(poc_spi));
PVDD2DGZ_G vddio3_b ( .VDDPST(vddio_bottombank));
PVDD2DGZ_G vcciodummy1 ( .VDDPST(vddio_bottombank));
PVDD2DGZ_G vddio1_b ( .VDDPST(vddio_bottombank));
PVDD2DGZ_G vcciodummy2 ( .VDDPST(vddio_spi));
PVSS3DGZ_G gnddummy1 ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd34_b_1_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd34_b_0_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd12_b_1_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnd12_b_0_ ( .VSS(gnd_), .VDDPST(vddio_bottombank));
PVSS3DGZ_G gnddummy2 ( .VSS(gnd_), .VDDPST(vddio_spi));
PVSS3DGZ_G gnd5 ( .VSS(gnd_), .VDDPST(vddio_spi));
PDUW08SDGZ_G_NOR pad_b_21_ ( .REN(ren[21]), .C(in[21]), .OEN(oen[21]),
     .IE(n_ienb[21]), .I(out[21]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net234[0]), .VDDIO(vddio_spi), .PAD(pad[21]),
     .POC(poc_spi));
PDUW08SDGZ_G_NOR pad_b_20_ ( .REN(ren[20]), .C(in[20]), .OEN(oen[20]),
     .IE(n_ienb[20]), .I(out[20]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net234[1]), .VDDIO(vddio_spi), .PAD(pad[20]),
     .POC(poc_spi));
PDUW08SDGZ_G_NOR pad_b_11_ ( .REN(ren[11]), .C(in[11]), .OEN(oen[11]),
     .IE(n_ienb[11]), .I(out[11]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net237[0]), .VDDIO(vddio_bottombank), .PAD(pad[11]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_10_ ( .REN(ren[10]), .C(in[10]), .OEN(oen[10]),
     .IE(n_ienb[10]), .I(out[10]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net237[1]), .VDDIO(vddio_bottombank), .PAD(pad[10]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_13_ ( .REN(ren[13]), .C(in[13]), .OEN(oen[13]),
     .IE(n_ienb[13]), .I(out[13]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net188[0]), .VDDIO(vddio_bottombank), .PAD(pad[13]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_12_ ( .REN(ren[12]), .C(in[12]), .OEN(oen[12]),
     .IE(n_ienb[12]), .I(out[12]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net188[1]), .VDDIO(vddio_bottombank), .PAD(pad[12]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_14_ ( .REN(ren[14]), .C(in[14]), .OEN(oen[14]),
     .IE(n_ienb[14]), .I(out[14]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net198), .VDDIO(vddio_bottombank), .PAD(pad[14]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_7_ ( .REN(ren[7]), .C(in[7]), .OEN(oen[7]),
     .IE(n_ienb[7]), .I(out[7]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[0]), .VDDIO(vddio_bottombank), .PAD(pad[7]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_6_ ( .REN(ren[6]), .C(in[6]), .OEN(oen[6]),
     .IE(n_ienb[6]), .I(out[6]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[1]), .VDDIO(vddio_bottombank), .PAD(pad[6]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_5_ ( .REN(ren[5]), .C(in[5]), .OEN(oen[5]),
     .IE(n_ienb[5]), .I(out[5]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[2]), .VDDIO(vddio_bottombank), .PAD(pad[5]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_4_ ( .REN(ren[4]), .C(in[4]), .OEN(oen[4]),
     .IE(n_ienb[4]), .I(out[4]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[3]), .VDDIO(vddio_bottombank), .PAD(pad[4]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_3_ ( .REN(ren[3]), .C(in[3]), .OEN(oen[3]),
     .IE(n_ienb[3]), .I(out[3]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[4]), .VDDIO(vddio_bottombank), .PAD(pad[3]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_2_ ( .REN(ren[2]), .C(in[2]), .OEN(oen[2]),
     .IE(n_ienb[2]), .I(out[2]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[5]), .VDDIO(vddio_bottombank), .PAD(pad[2]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_1_ ( .REN(ren[1]), .C(in[1]), .OEN(oen[1]),
     .IE(n_ienb[1]), .I(out[1]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[6]), .VDDIO(vddio_bottombank), .PAD(pad[1]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_0_ ( .REN(ren[0]), .C(in[0]), .OEN(oen[0]),
     .IE(n_ienb[0]), .I(out[0]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net241[7]), .VDDIO(vddio_bottombank), .PAD(pad[0]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_9_ ( .REN(ren[9]), .C(in[9]), .OEN(oen[9]),
     .IE(n_ienb[9]), .I(out[9]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net236[0]), .VDDIO(vddio_bottombank), .PAD(pad[9]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_8_ ( .REN(ren[8]), .C(in[8]), .OEN(oen[8]),
     .IE(n_ienb[8]), .I(out[8]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net236[1]), .VDDIO(vddio_bottombank), .PAD(pad[8]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_19_ ( .REN(ren[19]), .C(in[19]), .OEN(oen[19]),
     .IE(n_ienb[19]), .I(out[19]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[0]), .VDDIO(vddio_bottombank), .PAD(pad[19]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_18_ ( .REN(ren[18]), .C(in[18]), .OEN(oen[18]),
     .IE(n_ienb[18]), .I(out[18]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[1]), .VDDIO(vddio_bottombank), .PAD(pad[18]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_17_ ( .REN(ren[17]), .C(in[17]), .OEN(oen[17]),
     .IE(n_ienb[17]), .I(out[17]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[2]), .VDDIO(vddio_bottombank), .PAD(pad[17]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_16_ ( .REN(ren[16]), .C(in[16]), .OEN(oen[16]),
     .IE(n_ienb[16]), .I(out[16]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[3]), .VDDIO(vddio_bottombank), .PAD(pad[16]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_15_ ( .REN(ren[15]), .C(in[15]), .OEN(oen[15]),
     .IE(n_ienb[15]), .I(out[15]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net228[4]), .VDDIO(vddio_bottombank), .PAD(pad[15]),
     .POC(poc_bot));
PDUW08SDGZ_G_NOR ctst_b_b ( .REN(tiegnd_botpad), .C(ctst_b_int),
     .OEN(tievdd_botpad), .IE(tievdd_botpad), .I(tiegnd_botpad),
     .indiff(tiegnd_botpad), .PAD4LVDS(net233),
     .VDDIO(vddio_bottombank), .PAD(ctst_b), .POC(poc_bot));
PDUW08SDGZ_G_NOR cdone_b ( .REN(tiegnd_botpad), .C(cdone_int),
     .OEN(cdone_out), .IE(tievdd_botpad), .I(tiegnd_botpad),
     .indiff(tiegnd_botpad), .PAD4LVDS(net148),
     .VDDIO(vddio_bottombank), .PAD(cdone), .POC(poc_bot));
PDUW08SDGZ_G_NOR pad_b_23_ ( .REN(ren[23]), .C(in[23]), .OEN(oen[23]),
     .IE(n_ienb[23]), .I(out[23]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net168[0]), .VDDIO(vddio_spi), .PAD(pad[23]),
     .POC(poc_spi));
PDUW08SDGZ_G_NOR pad_b_22_ ( .REN(ren[22]), .C(in[22]), .OEN(oen[22]),
     .IE(n_ienb[22]), .I(out[22]), .indiff(tiegnd_botpad),
     .PAD4LVDS(net168[1]), .VDDIO(vddio_spi), .PAD(pad[22]),
     .POC(poc_spi));

endmodule
// Library - ice1chip, Cell - padring_ice1f, View - schematic
// LAST TIME SAVED: Apr 13 16:07:00 2011
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module padring_ice1f ( cdone_int, creset_b_int, in_bbank, in_lbank,
     in_rbank, in_tbank, pll_lock, pllout, trstb_int_pad,
     vddio_bottombank, vddio_spi, cdone, uio_bbank, uio_lbank,
     uio_rbank, uio_tbank, vpp, vppin, cdone_out, creset_b, ien,
     ien_bbank, ien_rbank, ien_tbank, lvds_en, oen_bbank, oen_lbank,
     oen_rbank, oen_tbank, out_bbank, out_lbank, out_rbank, out_tbank,
     pll_bypass, pll_cbit, pll_fb, pll_fse, pll_ref, pll_reset, ren,
     ren_bbank, ren_rbank, ren_tbank, trstb, vdda );
output  cdone_int, creset_b_int, pll_lock, pllout, trstb_int_pad,
     vddio_bottombank, vddio_spi;

inout  cdone, vpp, vppin;

input  cdone_out, creset_b, pll_bypass, pll_fb, pll_fse, pll_ref,
     pll_reset, trstb, vdda;

output [23:0]  in_tbank;
output [24:0]  in_rbank;
output [23:0]  in_bbank;
output [23:0]  in_lbank;

inout [24:0]  uio_rbank;
inout [23:0]  uio_bbank;
inout [23:0]  uio_tbank;
inout [23:0]  uio_lbank;

input [23:0]  ren_tbank;
input [23:0]  out_tbank;
input [16:0]  pll_cbit;
input [23:0]  ien_tbank;
input [25:0]  ren_rbank;
input [24:0]  ien_rbank;
input [23:0]  oen_tbank;
input [23:0]  ren_bbank;
input [23:0]  ien;
input [23:0]  ren;
input [23:0]  ien_bbank;
input [11:0]  lvds_en;
input [23:0]  out_lbank;
input [23:0]  oen_bbank;
input [23:0]  out_bbank;
input [24:0]  oen_rbank;
input [24:0]  out_rbank;
input [23:0]  oen_lbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



IO_lft_bank_ice1f_v2 iobank_l ( .ien(ien[23:0]),
     .lvds_en(lvds_en[11:0]), .ren(ren[23:0]), .pad(uio_lbank[23:0]),
     .in(in_lbank[23:0]), .oen(oen_lbank[23:0]), .out(out_lbank[23:0]),
     .vdda(vdda), .pll_ref(pll_ref), .pll_fse(pll_fse),
     .pll_cbit(pll_cbit[16:0]), .pll_fb(pll_fb),
     .pll_bypass(pll_bypass), .pll_lock(pll_lock), .pllout(pllout),
     .pll_reset(pll_reset));
IO_top_bank_ice1f iobank_t ( .vppin(vppin), .vpp(vpp),
     .ren(ren_tbank[23:0]), .out(out_tbank[23:0]),
     .oen(oen_tbank[23:0]), .ien(ien_tbank[23:0]), .in(in_tbank[23:0]),
     .pad(uio_tbank[23:0]));
IO_rgt_bank_ice1f iobank_r ( .ren(ren_rbank[25:0]),
     .ien(ien_rbank[24:0]), .oen(oen_rbank[24:0]), .in(in_rbank[24:0]),
     .pad(uio_rbank[24:0]), .out(out_rbank[24:0]), .TRSTb(trstb),
     .trstb_int(trstb_int_pad));
IO_bot_bank_ice1f iobank_b ( .vddio_bottombank(vddio_bottombank),
     .cdone_out(cdone_out), .ctst_b(creset_b), .ren(ren_bbank[23:0]),
     .out(out_bbank[23:0]), .oen(oen_bbank[23:0]),
     .ien(ien_bbank[23:0]), .in(in_bbank[23:0]), .pad(uio_bbank[23:0]),
     .vddio_spi(vddio_spi), .cdone(cdone), .cdone_int(cdone_int),
     .ctst_b_int(creset_b_int));

endmodule
// Library - ice1chip, Cell - ring_route_ice1f, View - schematic
// LAST TIME SAVED: Apr 13 16:08:16 2011
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module ring_route_ice1f ( bm_banksel_i, bm_init_i, bm_rcapmux_en_i,
     bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bs_en0, ceb0, end_of_startup, gint_hz, gsr,
     hiz_b0, in_bbank, in_lbank, in_rbank, in_tbank, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b,
     .cdsNet0(last_rsr[1]), .cdsNet0(last_rsr[0]),
     .cdsNet0(last_rsr[3]), .cdsNet0(last_rsr[2]), md_spi_b, mode0,
     mux_jtag_sel_b, pgate_l, pgate_r, pll_lock, pllout, reset_l,
     reset_r, sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, totdopad, trstb_pad, update0, vdd_cntl_l,
     vdd_cntl_r, wl_l, wl_r, bl_bot, bl_top, cdone, uio_bbank,
     uio_lbank, uio_rbank, uio_tbank, vpp, bm_sdo_o, creset_b,
     fabric_out_12_00, fabric_out_13_01, fabric_out_13_02, fromsdo,
     ien, ien_bbank, ien_rbank, ien_tbank, lvds_en, oen_bbank,
     oen_lbank, oen_rbank, oen_tbank, out_bbank, out_lbank, out_rbank,
     out_tbank, pll_bypass, pll_cbit, pll_fb, pll_fse, pll_ref,
     pll_reset, ren, ren_bbank, ren_rbank, ren_tbank, spi_ss_in_bbank,
     tck_pad, tdi_pad, tms_pad, trstb, vdda );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, ceb0, end_of_startup,
     gint_hz, gsr, hiz_b0, j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, md_spi_b, mode0, mux_jtag_sel_b,
     pll_lock, pllout, sdo_enable, shift0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, totdopad, trstb_pad, update0;

inout  cdone, vpp;

input  creset_b, fabric_out_12_00, fabric_out_13_01, fabric_out_13_02,
     fromsdo, pll_bypass, pll_fb, pll_fse, pll_ref, pll_reset, tck_pad,
     tdi_pad, tms_pad, trstb, vdda;

output [287:0]  reset_r;
output [287:0]  wl_l;
output [23:0]  in_lbank;
output [287:0]  reset_l;
output [3:0]  bm_banksel_i;
output [24:0]  in_rbank;
output [287:0]  vdd_cntl_l;
output [7:0]  bm_sa_i;
output [23:0]  in_tbank;
output [287:0]  wl_r;
output [3:0]  last_rsr;
output [287:0]  pgate_r;
output [3:0]  bm_sdi_i;
output [287:0]  vdd_cntl_r;
output [23:0]  in_bbank;
output [287:0]  pgate_l;

inout [24:0]  uio_rbank;
inout [663:0]  bl_bot;
inout [23:0]  uio_lbank;
inout [23:0]  uio_tbank;
inout [23:0]  uio_bbank;
inout [663:0]  bl_top;

input [23:0]  oen_bbank;
input [23:0]  out_bbank;
input [23:0]  ien_bbank;
input [3:0]  bm_sdo_o;
input [16:0]  pll_cbit;
input [11:0]  lvds_en;
input [23:0]  ien;
input [24:0]  oen_rbank;
input [23:0]  out_tbank;
input [23:0]  oen_tbank;
input [25:0]  ren_rbank;
input [23:0]  ren;
input [23:0]  out_lbank;
input [23:0]  ren_bbank;
input [24:0]  out_rbank;
input [23:0]  ien_tbank;
input [24:0]  ien_rbank;
input [23:0]  oen_lbank;
input [4:0]  spi_ss_in_bbank;
input [23:0]  ren_tbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ring_route00_ice1f I_ring_route00_ice1f (
     .spi_ss_in_bbank(spi_ss_in_bbank[4:0]),
     .fabric_out_12_00(fabric_out_12_00),
     .fabric_out_13_01(fabric_out_13_01),
     .fabric_out_13_02(fabric_out_13_02), .pgate_r(pgate_r[287:0]),
     .reset_b_r(reset_r[287:0]), .vdd_cntl_r(vdd_cntl_r[287:0]),
     .wl_r(wl_r[287:0]), .wl_l(wl_l[287:0]),
     .vdd_cntl_l(vdd_cntl_l[287:0]), .pgate_l(pgate_l[287:0]),
     .reset_b_l(reset_l[287:0]), .bl_top(bl_top[663:0]),
     .bl_bot(bl_bot[663:0]), .trstb_pad(trstb_pad), .tms_pad(tms_pad),
     .tdi_pad(tdi_pad), .tck_pad(tck_pad), .fromsdo(fromsdo),
     .creset_b_int(creset_b_int), .vddio_bottombank(vddio_bottombank),
     .vddio_spi(vddio_spi), .bm_sa_i(bm_sa_i[7:0]),
     .cdone_in(cdone_in), .bm_sdo_o(bm_sdo_o[3:0]), .vppin(vppin),
     .update0(update0), .tdo_pad(totdopad),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out), .shift0(shift0),
     .sdo_enable(sdo_enable), .mode0(mode0), .md_spi_b(md_spi_b),
     .last_rsr(last_rsr[3:0]),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .j_tdi(j_tdi), .j_tck(j_tck), .mux_jtag_sel_b(mux_jtag_sel_b),
     .hiz_b0(hiz_b0), .gsr(gsr), .gint_hz(gint_hz),
     .end_of_startup(end_of_startup), .ceb0(ceb0),
     .cdone_out(cdone_out), .bs_en0(bs_en0),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclk_i(bm_sclk_i),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bm_banksel_i(bm_banksel_i[3:0]));
padring_ice1f I_padring_ice1f ( .ien(ien[23:0]),
     .lvds_en(lvds_en[11:0]), .ren(ren[23:0]),
     .uio_lbank(uio_lbank[23:0]), .oen_lbank(oen_lbank[23:0]),
     .out_lbank(out_lbank[23:0]), .in_lbank(in_lbank[23:0]),
     .vdda(vdda), .pll_lock(pll_lock), .pllout(pllout),
     .pll_reset(pll_reset), .pll_bypass(pll_bypass), .pll_fb(pll_fb),
     .pll_cbit(pll_cbit[16:0]), .pll_fse(pll_fse), .pll_ref(pll_ref),
     .vddio_bottombank(vddio_bottombank), .uio_bbank(uio_bbank[23:0]),
     .uio_rbank(uio_rbank[24:0]), .uio_tbank(uio_tbank[23:0]),
     .in_bbank(in_bbank[23:0]), .in_rbank(in_rbank[24:0]),
     .in_tbank(in_tbank[23:0]), .ren_bbank(ren_bbank[23:0]),
     .oen_bbank(oen_bbank[23:0]), .oen_rbank(oen_rbank[24:0]),
     .oen_tbank(oen_tbank[23:0]), .out_bbank(out_bbank[23:0]),
     .out_rbank(out_rbank[24:0]), .out_tbank(out_tbank[23:0]),
     .ren_rbank(ren_rbank[25:0]), .ien_rbank(ien_rbank[24:0]),
     .ien_tbank(ien_tbank[23:0]), .ren_tbank(ren_tbank[23:0]),
     .ien_bbank(ien_bbank[23:0]), .vppin(vppin), .trstb(trstb),
     .creset_b(creset_b), .cdone_out(cdone_out),
     .creset_b_int(creset_b_int), .vpp(vpp), .cdone(cdone),
     .cdone_int(cdone_in), .trstb_int_pad(trstb_pad),
     .vddio_spi(vddio_spi));

endmodule
// Library - ice1chip, Cell - chip_ice1f, View - schematic
// LAST TIME SAVED: May  3 11:43:07 2011
// NETLIST TIME: May  5 11:56:48 2011
`timescale 1ns / 1ns 

module chip_ice1f ( cdone, uio_bbank, uio_lbank, uio_rbank, uio_tbank,
     vpp, creset_b, trstb, vdda );

inout  cdone, vpp;

input  creset_b, trstb, vdda;

inout [23:0]  uio_lbank;
inout [24:0]  uio_rbank;
inout [23:0]  uio_bbank;
inout [23:0]  uio_tbank;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [287:0]  vdd_cntl_l;

wire  [23:0]  in_lbank;

wire  [3:0]  bm_sdi_o;

wire  [3:0]  bm_banksel_i;

wire  [1:0]  gclk_r2clktv_b;

wire  [663:0]  bl_top;

wire  [23:0]  out_lbank;

wire  [23:0]  out_tbank;

wire  [1:0]  gclk_l2clktv_b;

wire  [287:0]  pgate_l;

wire  [3:0]  bm_sdo_o;

wire  [7:0]  fo_dlyadj;

wire  [287:0]  reset_l;

wire  [23:0]  oen_lbank;

wire  [24:0]  out_rbank;

wire  [23:0]  in_tbank;

wire  [287:0]  pgate_r;

wire  [23:0]  out_bbank;

wire  [23:0]  oen_bbank;

wire  [24:0]  oen_rbank;

wire  [287:0]  reset_r;

wire  [287:0]  wl_l;

wire  [24:0]  in_rbank;

wire  [287:0]  wl_r;

wire  [663:0]  bl_bot;

wire  [287:0]  vdd_cntl_r;

wire  [3:0]  last_rsr;

wire  [23:0]  oen_tbank;

wire  [11:10]  in_bbank_pll;

wire  [23:0]  in_bbank;

wire  [287:0]  cf_bbank;

wire  [7:0]  bm_sa_i;

wire  [287:0]  cf_tbank;

wire  [4:0]  spi_ss_in_bbank;

wire  [16:0]  pll_cbit;

wire  [383:0]  cf_lbank;

wire  [383:0]  cf_rbank;



pll_wrapbuf_ice1f pll_wrap ( gclk_l2clktv_b[1:0], gclk_r2clktv_b[1:0],
     in_bbank_pll[10], in_bbank_pll[11], pll_bypass, pll_cbit[16:0],
     pll_fb, pll_fse, pll_lock_out, pll_ref, pll_reset, pll_sdo,
     cf_bbank[159], cf_bbank[135], cf_lbank[9:1], cf_lbank[33:25],
     cf_lbank[57:49], cf_lbank[81:73], cf_lbank[97], cf_lbank[99],
     cf_lbank[101], fabric_out_06_00, fabric_out_07_00, fo_bypass,
     fo_dlyadj[7:0], fo_fb, fo_ref, fo_reset, fo_sck, fp_sdi, icegate,
     in_bbank[10], in_bbank[11], pll_lock, pllout, gint_hz);
quad_x4_ice1 iquad_x4 ( bm_sdo_o[3:0], cf_bbank[287:0],
     cf_lbank[383:0], cf_rbank[383:0], cf_tbank[287:0], icegate,
     fabric_out_06_00, fabric_out_07_00, fabric_out_12_00_wb,
     fabric_out_13_01, fabric_out_13_02, fo_bypass, fo_dlyadj[7:0],
     fo_fb, fo_ref, fo_reset, fo_sck, fp_sdi, oen_bbank[23:0],
     oen_lbank[23:0], oen_rbank[24:0], oen_tbank[23:0],
     out_bbank[23:0], out_lbank[23:0], out_rbank[24:0],
     out_tbank[23:0], fromsdo, spi_ss_in_bbank[4:0], tck_pad, tdi_pad,
     tms_pad, bl_bot[663:0], bl_top[663:0], bm_banksel_i[3:0],
     bm_init_i, bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i,
     bm_sdi_o[3:0], bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0,
     ceb, end_of_startup, gclk_l2clktv_b[1:0], gclk_r2clktv_b[1:0],
     hiz_b0, jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[0],
     last_rsr[1], last_rsr[2], last_rsr[3], md_spi_b, mode0,
     mux_jtag_sel_b, {in_bbank[23:12], in_bbank_pll[11],
     in_bbank_pll[10], in_bbank[9:0]}, in_lbank[23:0], in_rbank[24:0],
     in_tbank[23:0], pgate_l[287:0], pgate_r[287:0], pll_lock_out,
     pll_sdo, gint_hz, gsr, gsr, reset_l[287:0], reset_r[287:0], j_tdi,
     sdo_enable, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out, j_tck, totdopad, trstb_pad, update0,
     vdd_cntl_l[287:0], vdd_cntl_r[287:0], wl_l[287:0], wl_r[287:0]);
ring_route_ice1f I_ring_route1f ( bm_banksel_i[3:0], bm_init_i,
     bm_rcapmux_en_i, bm_sa_i[7:0], bm_sclk_i, bm_sclkrw_i,
     bm_sdi_o[3:0], bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0,
     ceb, end_of_startup, gint_hz, gsr, hiz_b0, in_bbank[23:0],
     in_lbank[23:0], in_rbank[24:0], in_tbank[23:0], j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr[1],
     last_rsr[0], last_rsr[3], last_rsr[2], md_spi_b, mode0,
     mux_jtag_sel_b, pgate_l[287:0], pgate_r[287:0], pll_lock, pllout,
     reset_l[287:0], reset_r[287:0], sdo_enable, shift0, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out, totdopad, trstb_pad, update0,
     vdd_cntl_l[287:0], vdd_cntl_r[287:0], wl_l[287:0], wl_r[287:0],
     bl_bot[663:0], bl_top[663:0], cdone, uio_bbank[23:0],
     uio_lbank[23:0], uio_rbank[24:0], uio_tbank[23:0], vpp,
     bm_sdo_o[3:0], creset_b, fabric_out_12_00_wb, fabric_out_13_01,
     fabric_out_13_02, fromsdo, {cf_lbank[324], cf_lbank[323],
     cf_lbank[300], cf_lbank[299], cf_lbank[276], cf_lbank[275],
     cf_lbank[252], cf_lbank[251], cf_lbank[228], cf_lbank[227],
     cf_lbank[204], cf_lbank[203], cf_lbank[180], cf_lbank[179],
     cf_lbank[132], cf_lbank[131], cf_lbank[108], cf_lbank[107],
     cf_lbank[84], cf_lbank[83], cf_lbank[60], cf_lbank[59],
     cf_lbank[36], cf_lbank[35]}, {cf_bbank[275], cf_bbank[276],
     cf_bbank[251], cf_bbank[252], cf_bbank[227], cf_bbank[228],
     cf_bbank[203], cf_bbank[204], cf_bbank[179], cf_bbank[180],
     cf_bbank[155], cf_bbank[156], cf_bbank[131], cf_bbank[132],
     cf_bbank[107], cf_bbank[108], cf_bbank[83], cf_bbank[84],
     cf_bbank[59], cf_bbank[60], cf_bbank[35], cf_bbank[36],
     cf_bbank[11], cf_bbank[12]}, {cf_rbank[347], cf_rbank[348],
     cf_rbank[323], cf_rbank[324], cf_rbank[299], cf_rbank[300],
     cf_rbank[251], cf_rbank[252], cf_rbank[227], cf_rbank[228],
     cf_rbank[203], cf_rbank[204], cf_rbank[179], cf_rbank[180],
     cf_rbank[155], cf_rbank[156], cf_rbank[131], cf_rbank[132],
     cf_rbank[83], cf_rbank[84], cf_rbank[59], cf_rbank[35],
     cf_rbank[36], cf_rbank[11], cf_rbank[12]}, {cf_tbank[275],
     cf_tbank[276], cf_tbank[251], cf_tbank[252], cf_tbank[227],
     cf_tbank[228], cf_tbank[203], cf_tbank[204], cf_tbank[179],
     cf_tbank[180], cf_tbank[155], cf_tbank[156], cf_tbank[131],
     cf_tbank[132], cf_tbank[107], cf_tbank[108], cf_tbank[83],
     cf_tbank[84], cf_tbank[59], cf_tbank[60], cf_tbank[35],
     cf_tbank[36], cf_tbank[11], cf_tbank[12]}, {cf_lbank[325],
     cf_lbank[301], cf_lbank[277], cf_lbank[253], cf_lbank[229],
     cf_lbank[205], cf_lbank[181], cf_lbank[133], cf_lbank[109],
     cf_lbank[85], cf_lbank[61], cf_lbank[37]}, oen_bbank[23:0],
     oen_lbank[23:0], oen_rbank[24:0], oen_tbank[23:0],
     out_bbank[23:0], out_lbank[23:0], out_rbank[24:0],
     out_tbank[23:0], pll_bypass, pll_cbit[16:0], pll_fb, pll_fse,
     pll_ref, pll_reset, {cf_lbank[322], cf_lbank[312], cf_lbank[298],
     cf_lbank[288], cf_lbank[274], cf_lbank[264], cf_lbank[250],
     cf_lbank[240], cf_lbank[226], cf_lbank[216], cf_lbank[202],
     cf_lbank[192], cf_lbank[178], cf_lbank[168], cf_lbank[130],
     cf_lbank[120], cf_lbank[106], cf_lbank[96], cf_lbank[82],
     cf_lbank[72], cf_lbank[58], cf_lbank[48], cf_lbank[34],
     cf_lbank[24]}, {cf_bbank[264], cf_bbank[274], cf_bbank[240],
     cf_bbank[250], cf_bbank[216], cf_bbank[226], cf_bbank[192],
     cf_bbank[202], cf_bbank[168], cf_bbank[178], cf_bbank[144],
     cf_bbank[154], cf_bbank[120], cf_bbank[130], cf_bbank[96],
     cf_bbank[106], cf_bbank[72], cf_bbank[82], cf_bbank[48],
     cf_bbank[58], cf_bbank[24], cf_bbank[34], cf_bbank[0],
     cf_bbank[10]}, {cf_rbank[38], cf_rbank[336], cf_rbank[346],
     cf_rbank[312], cf_rbank[322], cf_rbank[288], cf_rbank[298],
     cf_rbank[240], cf_rbank[250], cf_rbank[216], cf_rbank[226],
     cf_rbank[192], cf_rbank[202], cf_rbank[168], cf_rbank[178],
     cf_rbank[144], cf_rbank[154], cf_rbank[120], cf_rbank[130],
     cf_rbank[72], cf_rbank[82], cf_rbank[48], cf_rbank[24],
     cf_rbank[34], cf_rbank[0], cf_rbank[10]}, {cf_tbank[264],
     cf_tbank[274], cf_tbank[240], cf_tbank[250], cf_tbank[216],
     cf_tbank[226], cf_tbank[192], cf_tbank[202], cf_tbank[168],
     cf_tbank[178], cf_tbank[144], cf_tbank[154], cf_tbank[120],
     cf_tbank[130], cf_tbank[96], cf_tbank[106], cf_tbank[72],
     cf_tbank[82], cf_tbank[48], cf_tbank[58], cf_tbank[24],
     cf_tbank[34], cf_tbank[0], cf_tbank[10]}, spi_ss_in_bbank[4:0],
     tck_pad, tdi_pad, tms_pad, trstb, vdda);

endmodule
// Library - leafcell, Cell - sbox8to6_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:51:38 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox8to6_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  t;
inout [9:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  reset_b;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I554 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_l7 ( .prog(prog), .in6(t[1]), .in5(t[7]), .in4(r[11]),
     .in3(r[7]), .in2(r[4]), .in1(b[7]), .in0(b[2]), .out(l[7]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t7 ( .prog(prog), .in6(r[1]), .in5(r[7]), .in4(b[11]),
     .in3(b[7]), .in2(b[4]), .in1(l[7]), .in0(l[2]), .out(t[7]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t8 ( .prog(prog), .in6(r[2]), .in5(r[8]), .in4(b[0]),
     .in3(b[8]), .in2(b[5]), .in1(l[8]), .in0(l[3]), .out(t[8]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t6 ( .prog(prog), .in6(r[0]), .in5(r[6]), .in4(b[10]),
     .in3(b[6]), .in2(b[3]), .in1(l[6]), .in0(l[1]), .out(t[6]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l8 ( .prog(prog), .in6(t[2]), .in5(t[8]), .in4(r[0]),
     .in3(r[8]), .in2(r[5]), .in1(b[8]), .in0(b[3]), .out(l[8]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l6 ( .prog(prog), .in6(t[0]), .in5(t[6]), .in4(r[10]),
     .in3(r[6]), .in2(r[3]), .in1(b[6]), .in0(b[1]), .out(l[6]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox8to6_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:50:50 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox8to6_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r7 ( .prog(prog), .in6(b[1]), .in5(b[7]), .in4(l[11]),
     .in3(l[7]), .in2(l[4]), .in1(t[7]), .in0(t[2]), .out(r[7]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b7 ( .prog(prog), .in6(l[1]), .in5(l[7]), .in4(t[11]),
     .in3(t[7]), .in2(t[4]), .in1(r[7]), .in0(r[2]), .out(b[7]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b8 ( .prog(prog), .in6(l[2]), .in5(l[8]), .in4(t[0]),
     .in3(t[8]), .in2(t[5]), .in1(r[8]), .in0(r[3]), .out(b[8]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b6 ( .prog(prog), .in6(l[0]), .in5(l[6]), .in4(t[10]),
     .in3(t[6]), .in2(t[3]), .in1(r[6]), .in0(r[1]), .out(b[6]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r8 ( .prog(prog), .in6(b[2]), .in5(b[8]), .in4(l[0]),
     .in3(l[8]), .in2(l[5]), .in1(t[8]), .in0(t[3]), .out(r[8]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r6 ( .prog(prog), .in6(b[0]), .in5(b[6]), .in4(l[10]),
     .in3(l[6]), .in2(l[3]), .in1(t[6]), .in0(t[1]), .out(r[6]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox5to3_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:39:32 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox5to3_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [11:0]  l;
inout [11:0]  t;
inout [11:0]  b;
inout [11:0]  r;
inout [9:0]  bl;

input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_l4 ( .prog(prog), .in6(t[10]), .in5(t[4]), .in4(r[8]),
     .in3(r[4]), .in2(r[1]), .in1(b[4]), .in0(b[11]), .out(l[4]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_t4 ( .prog(prog), .in6(r[10]), .in5(r[4]), .in4(b[8]),
     .in3(b[4]), .in2(b[1]), .in1(l[4]), .in0(l[11]), .out(t[4]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_t5 ( .prog(prog), .in6(r[11]), .in5(r[5]), .in4(b[9]),
     .in3(b[5]), .in2(b[2]), .in1(l[5]), .in0(l[0]), .out(t[5]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t3 ( .prog(prog), .in6(r[9]), .in5(r[3]), .in4(b[7]),
     .in3(b[3]), .in2(b[0]), .in1(l[3]), .in0(l[10]), .out(t[3]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_l5 ( .prog(prog), .in6(t[11]), .in5(t[5]), .in4(r[9]),
     .in3(r[5]), .in2(r[2]), .in1(b[5]), .in0(b[0]), .out(l[5]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_l3 ( .prog(prog), .in6(t[9]), .in5(t[3]), .in4(r[7]),
     .in3(r[3]), .in2(r[0]), .in1(b[3]), .in0(b[10]), .out(l[3]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox5to3_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:38:42 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox5to3_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  b;

input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r4 ( .prog(prog), .in6(b[10]), .in5(b[4]), .in4(l[8]),
     .in3(l[4]), .in2(l[1]), .in1(t[4]), .in0(t[11]), .out(r[4]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_b4 ( .prog(prog), .in6(l[10]), .in5(l[4]), .in4(t[8]),
     .in3(t[4]), .in2(t[1]), .in1(r[4]), .in0(r[11]), .out(b[4]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_b5 ( .prog(prog), .in6(l[11]), .in5(l[5]), .in4(t[9]),
     .in3(t[5]), .in2(t[2]), .in1(r[5]), .in0(r[0]), .out(b[5]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b3 ( .prog(prog), .in6(l[9]), .in5(l[3]), .in4(t[7]),
     .in3(t[3]), .in2(t[0]), .in1(r[3]), .in0(r[10]), .out(b[3]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));
sbox7to1_220 I_r5 ( .prog(prog), .in6(b[11]), .in5(b[5]), .in4(l[9]),
     .in3(l[5]), .in2(l[2]), .in1(t[5]), .in0(t[0]), .out(r[5]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_r3 ( .prog(prog), .in6(b[9]), .in5(b[3]), .in4(l[7]),
     .in3(l[3]), .in2(l[0]), .in1(t[3]), .in0(t[10]), .out(r[3]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));

endmodule
// Library - leafcell, Cell - sbox2to0_p2_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:37:50 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox2to0_p2_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbitb;
output [19:0]  cbit;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  b;
inout [11:0]  l;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
sbox7to1_220 I_l1 ( .prog(prog), .in6(t[7]), .in5(t[1]), .in4(r[5]),
     .in3(r[1]), .in2(r[10]), .in1(b[1]), .in0(b[8]), .out(l[1]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_l0 ( .prog(prog), .in6(t[6]), .in5(t[0]), .in4(r[4]),
     .in3(r[0]), .in2(r[9]), .in1(b[0]), .in0(b[7]), .out(l[0]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));
sbox7to1_220 I_t1 ( .prog(prog), .in6(r[7]), .in5(r[1]), .in4(b[5]),
     .in3(b[1]), .in2(b[10]), .in1(l[1]), .in0(l[8]), .out(t[1]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_l2 ( .prog(prog), .in6(t[8]), .in5(t[2]), .in4(r[6]),
     .in3(r[2]), .in2(r[11]), .in1(b[2]), .in0(b[9]), .out(l[2]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_t2 ( .prog(prog), .in6(r[8]), .in5(r[2]), .in4(b[6]),
     .in3(b[2]), .in2(b[11]), .in1(l[2]), .in0(l[9]), .out(t[2]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_t0 ( .prog(prog), .in6(r[6]), .in5(r[0]), .in4(b[4]),
     .in3(b[0]), .in2(b[9]), .in1(l[0]), .in0(l[7]), .out(t[0]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));

endmodule
// Library - leafcell, Cell - pll_ml_dff, View - schematic
// LAST TIME SAVED: Jun  9 15:25:37 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pll_ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - leafcell, Cell - sbox2to0_p1_v2, View - schematic
// LAST TIME SAVED: Oct 18 10:53:10 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox2to0_p1_v2 ( cbit, cbitb, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [19:0]  cbit;
output [19:0]  cbitb;

inout [9:0]  bl;
inout [11:0]  b;
inout [11:0]  r;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



cram2x2x5 I_cram2x2x5 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
sbox7to1_220 I_r1 ( .prog(prog), .in6(b[7]), .in5(b[1]), .in4(l[5]),
     .in3(l[1]), .in2(l[10]), .in1(t[1]), .in0(t[8]), .out(r[1]),
     .cb({cbitb[10], cbitb[11], cbitb[14]}), .c({cbit[10], cbit[11],
     cbit[14]}));
sbox7to1_220 I_r0 ( .prog(prog), .in6(b[6]), .in5(b[0]), .in4(l[4]),
     .in3(l[0]), .in2(l[9]), .in1(t[0]), .in0(t[7]), .out(r[0]),
     .cb({cbitb[4], cbitb[3], cbitb[0]}), .c({cbit[4], cbit[3],
     cbit[0]}));
sbox7to1_220 I_b1 ( .prog(prog), .in6(l[7]), .in5(l[1]), .in4(t[5]),
     .in3(t[1]), .in2(t[10]), .in1(r[1]), .in0(r[8]), .out(b[1]),
     .cb({cbitb[9], cbitb[8], cbitb[12]}), .c({cbit[9], cbit[8],
     cbit[12]}));
sbox7to1_220 I_r2 ( .prog(prog), .in6(b[8]), .in5(b[2]), .in4(l[6]),
     .in3(l[2]), .in2(l[11]), .in1(t[2]), .in0(t[9]), .out(r[2]),
     .cb({cbitb[13], cbitb[18], cbitb[17]}), .c({cbit[13], cbit[18],
     cbit[17]}));
sbox7to1_220 I_b2 ( .prog(prog), .in6(l[8]), .in5(l[2]), .in4(t[6]),
     .in3(t[2]), .in2(t[11]), .in1(r[2]), .in0(r[9]), .out(b[2]),
     .cb({cbitb[19], cbitb[16], cbitb[15]}), .c({cbit[19], cbit[16],
     cbit[15]}));
sbox7to1_220 I_b0 ( .prog(prog), .in6(l[6]), .in5(l[0]), .in4(t[4]),
     .in3(t[0]), .in2(t[9]), .in1(r[0]), .in0(r[7]), .out(b[0]),
     .cb({cbitb[2], cbitb[1], cbitb[6]}), .c({cbit[2], cbit[1],
     cbit[6]}));

endmodule
// Library - leafcell, Cell - span4_switchandmem_v3, View - schematic
// LAST TIME SAVED: Oct 19 10:24:53 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module span4_switchandmem_v3 ( c, cc, b, bl, l, r, t, pgate, prog,
     reset_b, vdd_cntl, wl );


input  prog;

output [7:0]  c;
output [15:8]  cc;

inout [11:0]  r;
inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  b;

input [15:0]  reset_b;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  n2;

wire  [19:0]  net0236;

wire  [19:0]  n1;

wire  [19:0]  net0248;

wire  [19:0]  net0245;

wire  [19:0]  n3;

wire  [19:0]  net0177;

wire  [19:0]  net0241;

wire  [19:0]  n6;

wire  [19:0]  n5;

wire  [19:0]  n0;

wire  [19:0]  n4;

wire  [19:0]  net0201;

wire  [19:0]  n7;

wire  [19:0]  net0189;

wire  [19:0]  net0250;



sbox11to9_p2_v2 I_sbox11to9_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0241[0], net0241[1], net0241[2], net0241[3],
     net0241[4], net0241[5], net0241[6], net0241[7], net0241[8],
     net0241[9], net0241[10], net0241[11], net0241[12], net0241[13],
     net0241[14], net0241[15], net0241[16], net0241[17], net0241[18],
     net0241[19]}), .cbit({n7[19:8], cc[15], n7[6], cc[14], n7[4:0]}),
     .wl(wl[15:14]), .vdd_cntl(vdd_cntl[15:14]),
     .reset_b(reset_b[15:14]), .pgate(pgate[15:14]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox11to9_p1_v2 I_sbox11to9_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0236[0], net0236[1], net0236[2], net0236[3],
     net0236[4], net0236[5], net0236[6], net0236[7], net0236[8],
     net0236[9], net0236[10], net0236[11], net0236[12], net0236[13],
     net0236[14], net0236[15], net0236[16], net0236[17], net0236[18],
     net0236[19]}), .cbit({n6[19:8], cc[13], n6[6], cc[12], n6[4:0]}),
     .wl(wl[13:12]), .vdd_cntl(vdd_cntl[13:12]),
     .reset_b(reset_b[13:12]), .pgate(pgate[13:12]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox8to6_p2_v2 I_sbox8to6_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0248[0], net0248[1], net0248[2], net0248[3],
     net0248[4], net0248[5], net0248[6], net0248[7], net0248[8],
     net0248[9], net0248[10], net0248[11], net0248[12], net0248[13],
     net0248[14], net0248[15], net0248[16], net0248[17], net0248[18],
     net0248[19]}), .cbit({n5[19:8], cc[11], n5[6], cc[10], n5[4:0]}),
     .wl(wl[11:10]), .vdd_cntl(vdd_cntl[11:10]),
     .reset_b(reset_b[11:10]), .pgate(pgate[11:10]), .t(t[11:0]),
     .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]));
sbox8to6_p1_v2 I_sbox8to6_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0177[0], net0177[1], net0177[2], net0177[3],
     net0177[4], net0177[5], net0177[6], net0177[7], net0177[8],
     net0177[9], net0177[10], net0177[11], net0177[12], net0177[13],
     net0177[14], net0177[15], net0177[16], net0177[17], net0177[18],
     net0177[19]}), .cbit({n4[19:8], cc[9], n4[6], cc[8], n4[4:0]}),
     .wl(wl[9:8]), .vdd_cntl(vdd_cntl[9:8]), .reset_b(reset_b[9:8]),
     .pgate(pgate[9:8]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox5to3_p2_v2 I_sbox5to3_p2_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0189[0], net0189[1], net0189[2], net0189[3],
     net0189[4], net0189[5], net0189[6], net0189[7], net0189[8],
     net0189[9], net0189[10], net0189[11], net0189[12], net0189[13],
     net0189[14], net0189[15], net0189[16], net0189[17], net0189[18],
     net0189[19]}), .cbit({n3[19:8], c[7], n3[6], c[6], n3[4:0]}),
     .wl(wl[7:6]), .vdd_cntl(vdd_cntl[7:6]), .reset_b(reset_b[7:6]),
     .pgate(pgate[7:6]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox5to3_p1_v2 I_sbox5to3_p1_v2 ( .b(b[11:0]), .prog(prog),
     .cbitb({net0201[0], net0201[1], net0201[2], net0201[3],
     net0201[4], net0201[5], net0201[6], net0201[7], net0201[8],
     net0201[9], net0201[10], net0201[11], net0201[12], net0201[13],
     net0201[14], net0201[15], net0201[16], net0201[17], net0201[18],
     net0201[19]}), .cbit({n2[19:8], c[5], n2[6], c[4], n2[4:0]}),
     .wl(wl[5:4]), .vdd_cntl(vdd_cntl[5:4]), .reset_b(reset_b[5:4]),
     .pgate(pgate[5:4]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox2to0_p2_v2 I_sbox2to0_p2_v2 ( .b(b[11:0]), .cbitb({net0245[0],
     net0245[1], net0245[2], net0245[3], net0245[4], net0245[5],
     net0245[6], net0245[7], net0245[8], net0245[9], net0245[10],
     net0245[11], net0245[12], net0245[13], net0245[14], net0245[15],
     net0245[16], net0245[17], net0245[18], net0245[19]}),
     .cbit({n1[19:8], c[3], n1[6], c[2], n1[4:0]}), .wl(wl[3:2]),
     .vdd_cntl(vdd_cntl[3:2]), .reset_b(reset_b[3:2]), .prog(prog),
     .pgate(pgate[3:2]), .t(t[11:0]), .r(r[11:0]), .l(l[11:0]),
     .bl(bl[9:0]));
sbox2to0_p1_v2 I_sbox2to0_p1_v2 ( .cbitb({net0250[0], net0250[1],
     net0250[2], net0250[3], net0250[4], net0250[5], net0250[6],
     net0250[7], net0250[8], net0250[9], net0250[10], net0250[11],
     net0250[12], net0250[13], net0250[14], net0250[15], net0250[16],
     net0250[17], net0250[18], net0250[19]}), .cbit({n0[19:8], c[1],
     n0[6], c[0], n0[4:0]}), .wl(wl[1:0]), .vdd_cntl(vdd_cntl[1:0]),
     .reset_b(reset_b[1:0]), .prog(prog), .pgate(pgate[1:0]),
     .t(t[11:0]), .r(r[11:0]), .l(l[11:0]), .bl(bl[9:0]), .b(b[11:0]));

endmodule
// Library - leafcell, Cell - span4_ice8p, View - schematic
// LAST TIME SAVED: Jan 12 15:03:31 2011
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module span4_ice8p ( bram_cbit, ccntrl_cbit, bl, sp4_h_l, sp4_h_r,
     sp4_v_b, sp4_v_t, pgate, prog, reset_b, vdd_cntl, wl );


input  prog;

output [7:0]  bram_cbit;
output [7:0]  ccntrl_cbit;

inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_t;
inout [47:0]  sp4_h_r;
inout [9:0]  bl;

input [15:0]  vdd_cntl;
input [15:0]  reset_b;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  sp4_h_r_mid;

wire  [11:0]  sp4_v_b_mid;



rm7y  R0_47_ ( .MINUS(sp4_v_b[47]), .PLUS(sp4_v_t[34]));
rm7y  R0_46_ ( .MINUS(sp4_v_b[46]), .PLUS(sp4_v_t[35]));
rm7y  R0_45_ ( .MINUS(sp4_v_b[45]), .PLUS(sp4_v_t[32]));
rm7y  R0_44_ ( .MINUS(sp4_v_b[44]), .PLUS(sp4_v_t[33]));
rm7y  R0_43_ ( .MINUS(sp4_v_b[43]), .PLUS(sp4_v_t[30]));
rm7y  R0_42_ ( .MINUS(sp4_v_b[42]), .PLUS(sp4_v_t[31]));
rm7y  R0_41_ ( .MINUS(sp4_v_b[41]), .PLUS(sp4_v_t[28]));
rm7y  R0_40_ ( .MINUS(sp4_v_b[40]), .PLUS(sp4_v_t[29]));
rm7y  R0_39_ ( .MINUS(sp4_v_b[39]), .PLUS(sp4_v_t[26]));
rm7y  R0_38_ ( .MINUS(sp4_v_b[38]), .PLUS(sp4_v_t[27]));
rm7y  R0_37_ ( .MINUS(sp4_v_b[37]), .PLUS(sp4_v_t[24]));
rm7y  R0_36_ ( .MINUS(sp4_v_b[36]), .PLUS(sp4_v_t[25]));
rm7y  R0_35_ ( .MINUS(sp4_v_b[35]), .PLUS(sp4_v_t[22]));
rm7y  R0_34_ ( .MINUS(sp4_v_b[34]), .PLUS(sp4_v_t[23]));
rm7y  R0_33_ ( .MINUS(sp4_v_b[33]), .PLUS(sp4_v_t[20]));
rm7y  R0_32_ ( .MINUS(sp4_v_b[32]), .PLUS(sp4_v_t[21]));
rm7y  R0_31_ ( .MINUS(sp4_v_b[31]), .PLUS(sp4_v_t[18]));
rm7y  R0_30_ ( .MINUS(sp4_v_b[30]), .PLUS(sp4_v_t[19]));
rm7y  R0_29_ ( .MINUS(sp4_v_b[29]), .PLUS(sp4_v_t[16]));
rm7y  R0_28_ ( .MINUS(sp4_v_b[28]), .PLUS(sp4_v_t[17]));
rm7y  R0_27_ ( .MINUS(sp4_v_b[27]), .PLUS(sp4_v_t[14]));
rm7y  R0_26_ ( .MINUS(sp4_v_b[26]), .PLUS(sp4_v_t[15]));
rm7y  R0_25_ ( .MINUS(sp4_v_b[25]), .PLUS(sp4_v_t[12]));
rm7y  R0_24_ ( .MINUS(sp4_v_b[24]), .PLUS(sp4_v_t[13]));
rm7y  R0_23_ ( .MINUS(sp4_v_b[23]), .PLUS(sp4_v_t[10]));
rm7y  R0_22_ ( .MINUS(sp4_v_b[22]), .PLUS(sp4_v_t[11]));
rm7y  R0_21_ ( .MINUS(sp4_v_b[21]), .PLUS(sp4_v_t[8]));
rm7y  R0_20_ ( .MINUS(sp4_v_b[20]), .PLUS(sp4_v_t[9]));
rm7y  R0_19_ ( .MINUS(sp4_v_b[19]), .PLUS(sp4_v_t[6]));
rm7y  R0_18_ ( .MINUS(sp4_v_b[18]), .PLUS(sp4_v_t[7]));
rm7y  R0_17_ ( .MINUS(sp4_v_b[17]), .PLUS(sp4_v_t[4]));
rm7y  R0_16_ ( .MINUS(sp4_v_b[16]), .PLUS(sp4_v_t[5]));
rm7y  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[2]));
rm7y  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[3]));
rm7y  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[0]));
rm7y  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[1]));
rm7y  R0_11_ ( .MINUS(sp4_v_b_mid[11]), .PLUS(sp4_v_t[46]));
rm7y  R0_10_ ( .MINUS(sp4_v_b_mid[10]), .PLUS(sp4_v_t[47]));
rm7y  R0_9_ ( .MINUS(sp4_v_b_mid[9]), .PLUS(sp4_v_t[44]));
rm7y  R0_8_ ( .MINUS(sp4_v_b_mid[8]), .PLUS(sp4_v_t[45]));
rm7y  R0_7_ ( .MINUS(sp4_v_b_mid[7]), .PLUS(sp4_v_t[42]));
rm7y  R0_6_ ( .MINUS(sp4_v_b_mid[6]), .PLUS(sp4_v_t[43]));
rm7y  R0_5_ ( .MINUS(sp4_v_b_mid[5]), .PLUS(sp4_v_t[40]));
rm7y  R0_4_ ( .MINUS(sp4_v_b_mid[4]), .PLUS(sp4_v_t[41]));
rm7y  R0_3_ ( .MINUS(sp4_v_b_mid[3]), .PLUS(sp4_v_t[38]));
rm7y  R0_2_ ( .MINUS(sp4_v_b_mid[2]), .PLUS(sp4_v_t[39]));
rm7y  R0_1_ ( .MINUS(sp4_v_b_mid[1]), .PLUS(sp4_v_t[36]));
rm7y  R0_0_ ( .MINUS(sp4_v_b_mid[0]), .PLUS(sp4_v_t[37]));
span4_switchandmem_v3 I_span4_switchandmem_rev ( .cc(ccntrl_cbit[7:0]),
     .c(bram_cbit[7:0]), .wl(wl[15:0]), .vdd_cntl(vdd_cntl[15:0]),
     .reset_b(reset_b[15:0]), .prog(prog), .pgate(pgate[15:0]),
     .t(sp4_v_b_mid[11:0]), .r(sp4_h_r[11:0]), .l(sp4_h_r_mid[11:0]),
     .bl(bl[9:0]), .b(sp4_v_b[11:0]));
rm6w  R1_27_ ( .MINUS(sp4_h_r[47]), .PLUS(sp4_h_l[34]));
rm6w  R1_26_ ( .MINUS(sp4_h_r[46]), .PLUS(sp4_h_l[35]));
rm6w  R1_25_ ( .MINUS(sp4_h_r[45]), .PLUS(sp4_h_l[32]));
rm6w  R1_24_ ( .MINUS(sp4_h_r[44]), .PLUS(sp4_h_l[33]));
rm6w  R1_23_ ( .MINUS(sp4_h_r[43]), .PLUS(sp4_h_l[30]));
rm6w  R1_22_ ( .MINUS(sp4_h_r[42]), .PLUS(sp4_h_l[31]));
rm6w  R1_21_ ( .MINUS(sp4_h_r[41]), .PLUS(sp4_h_l[28]));
rm6w  R1_20_ ( .MINUS(sp4_h_r[40]), .PLUS(sp4_h_l[29]));
rm6w  R1_19_ ( .MINUS(sp4_h_r[39]), .PLUS(sp4_h_l[26]));
rm6w  R1_18_ ( .MINUS(sp4_h_r[38]), .PLUS(sp4_h_l[27]));
rm6w  R1_17_ ( .MINUS(sp4_h_r[37]), .PLUS(sp4_h_l[24]));
rm6w  R1_16_ ( .MINUS(sp4_h_r[36]), .PLUS(sp4_h_l[25]));
rm6w  R1_15_ ( .MINUS(sp4_h_r[35]), .PLUS(sp4_h_l[22]));
rm6w  R1_14_ ( .MINUS(sp4_h_r[34]), .PLUS(sp4_h_l[23]));
rm6w  R1_13_ ( .MINUS(sp4_h_r[23]), .PLUS(sp4_h_l[10]));
rm6w  R1_12_ ( .MINUS(sp4_h_r[22]), .PLUS(sp4_h_l[11]));
rm6w  R1_11_ ( .MINUS(sp4_h_r_mid[11]), .PLUS(sp4_h_l[46]));
rm6w  R1_10_ ( .MINUS(sp4_h_r_mid[10]), .PLUS(sp4_h_l[47]));
rm6w  R1_9_ ( .MINUS(sp4_h_r_mid[9]), .PLUS(sp4_h_l[44]));
rm6w  R1_8_ ( .MINUS(sp4_h_r_mid[8]), .PLUS(sp4_h_l[45]));
rm6w  R1_7_ ( .MINUS(sp4_h_r_mid[7]), .PLUS(sp4_h_l[42]));
rm6w  R1_6_ ( .MINUS(sp4_h_r_mid[6]), .PLUS(sp4_h_l[43]));
rm6w  R1_5_ ( .MINUS(sp4_h_r_mid[5]), .PLUS(sp4_h_l[40]));
rm6w  R1_4_ ( .MINUS(sp4_h_r_mid[4]), .PLUS(sp4_h_l[41]));
rm6w  R1_3_ ( .MINUS(sp4_h_r_mid[3]), .PLUS(sp4_h_l[38]));
rm6w  R1_2_ ( .MINUS(sp4_h_r_mid[2]), .PLUS(sp4_h_l[39]));
rm6w  R1_1_ ( .MINUS(sp4_h_r_mid[1]), .PLUS(sp4_h_l[36]));
rm6w  R1_0_ ( .MINUS(sp4_h_r_mid[0]), .PLUS(sp4_h_l[37]));
rm6w  R2_19_ ( .MINUS(sp4_h_r[33]), .PLUS(sp4_h_l[20]));
rm6w  R2_18_ ( .MINUS(sp4_h_r[32]), .PLUS(sp4_h_l[21]));
rm6w  R2_17_ ( .MINUS(sp4_h_r[31]), .PLUS(sp4_h_l[18]));
rm6w  R2_16_ ( .MINUS(sp4_h_r[30]), .PLUS(sp4_h_l[19]));
rm6w  R2_15_ ( .MINUS(sp4_h_r[29]), .PLUS(sp4_h_l[16]));
rm6w  R2_14_ ( .MINUS(sp4_h_r[28]), .PLUS(sp4_h_l[17]));
rm6w  R2_13_ ( .MINUS(sp4_h_r[27]), .PLUS(sp4_h_l[14]));
rm6w  R2_12_ ( .MINUS(sp4_h_r[26]), .PLUS(sp4_h_l[15]));
rm6w  R2_11_ ( .MINUS(sp4_h_r[25]), .PLUS(sp4_h_l[12]));
rm6w  R2_10_ ( .MINUS(sp4_h_r[24]), .PLUS(sp4_h_l[13]));
rm6w  R2_9_ ( .MINUS(sp4_h_r[21]), .PLUS(sp4_h_l[8]));
rm6w  R2_8_ ( .MINUS(sp4_h_r[20]), .PLUS(sp4_h_l[9]));
rm6w  R2_7_ ( .MINUS(sp4_h_r[19]), .PLUS(sp4_h_l[6]));
rm6w  R2_6_ ( .MINUS(sp4_h_r[18]), .PLUS(sp4_h_l[7]));
rm6w  R2_5_ ( .MINUS(sp4_h_r[17]), .PLUS(sp4_h_l[4]));
rm6w  R2_4_ ( .MINUS(sp4_h_r[16]), .PLUS(sp4_h_l[5]));
rm6w  R2_3_ ( .MINUS(sp4_h_r[15]), .PLUS(sp4_h_l[2]));
rm6w  R2_2_ ( .MINUS(sp4_h_r[14]), .PLUS(sp4_h_l[3]));
rm6w  R2_1_ ( .MINUS(sp4_h_r[13]), .PLUS(sp4_h_l[0]));
rm6w  R2_0_ ( .MINUS(sp4_h_r[12]), .PLUS(sp4_h_l[1]));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev0, View - schematic
// LAST TIME SAVED: Sep 17 15:03:29 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module clkmandcmuxrev0 ( clk, clkb, glb2local, s_r, cbit, cbitb,
     glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, min0, min1,
     min2, min3, prog );
output  clk, clkb, s_r;

input  prog;

output [3:0]  glb2local;

input [7:0]  min3;
input [7:0]  min2;
input [7:0]  min0;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g3;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g0;
input [5:0]  lc_trk_g1;
input [7:0]  min1;
input [31:0]  cbit;
input [31:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_mux8to1 I_clkmux8to1_0 ( .prog(prog), .inmuxo(glb2local[0]),
     .min(min3[7:0]), .cbit(cbit[16:13]), .cbitb(cbitb[16:13]));
clk_mux8to1 I_clkmux8to1_1 ( .prog(prog), .inmuxo(glb2local[1]),
     .min(min2[7:0]), .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I_clkmux8to1_3 ( .prog(prog), .inmuxo(glb2local[3]),
     .min(min0[7:0]), .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));
clk_mux8to1 I_clkmux8to1_2 ( .prog(prog), .inmuxo(glb2local[2]),
     .min(min1[7:0]), .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
clk_mux12to1 I_clkmux12to1 ( .prog(prog), .min({lc_trk_g3[1],
     lc_trk_g2[0], lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}),
     .clk(clk), .clkb(clkb), .cbitb({cbitb[31], cbitb[4], cbitb[3],
     cbitb[2], cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3],
     cbit[2], cbit[1], cbit[0]}), .cenb(ceb));
ce_clkm8to1 I_cemux8to1 ( .cbitb(cbitb[8:5]), .min({lc_trk_g3[3],
     lc_trk_g2[2], lc_trk_g1[3], lc_trk_g0[2], glb_netwk[7],
     glb_netwk[5], glb_netwk[3], glb_netwk[1]}), .cbit(cbit[8:5]),
     .moutb(ceb), .prog(prog));
sr_clkm8to1 I_srmux8to1 ( .cbitb(cbitb[12:9]), .min({lc_trk_g3[5],
     lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4], glb_netwk[6],
     glb_netwk[4], glb_netwk[2], glb_netwk[0]}), .cbit(cbit[12:9]),
     .mout(s_r), .prog(prog));

endmodule
// Library - leafcell, Cell - sbox1, View - schematic
// LAST TIME SAVED: Jun  8 15:19:03 2007
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module sbox1 ( b, l, r, t, c, cb, prog );
inout  b, l, r, t;

input  prog;

input [7:0]  cb;
input [7:0]  c;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



sbox1m3to1 I232 ( .in2(r), .cb(cb[7:6]), .op(t), .in0(l), .in1(b),
     .c(c[7:6]), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb(cb[3:2]), .op(l), .in0(b), .in1(t),
     .c(c[3:2]), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb(cb[1:0]), .op(b), .in0(l), .in1(t),
     .c(c[1:0]), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb(cb[5:4]), .op(r), .in0(l), .in1(t),
     .c(c[5:4]), .prog(prog));

endmodule
// Library - xpmem, Cell - cram16x4, View - schematic
// LAST TIME SAVED: Jun 24 17:57:57 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module cram16x4 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [63:0]  q_b;
output [63:0]  q;

inout [3:0]  bl;

input [15:0]  r_gnd;
input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 I16_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[1:0]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[15:14]));
cram2x2 I16_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[1:0]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[13:12]));
cram2x2 I16_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[1:0]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[11:10]));
cram2x2 I16_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[1:0]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[9:8]));
cram2x2 I16_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[1:0]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[7:6]));
cram2x2 I16_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[1:0]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[5:4]));
cram2x2 I16_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[1:0]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[3:2]));
cram2x2 I16_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[3:2]), .q_b(q_b[63:60]),
     .q(q[63:60]), .wl(wl[15:14]));
cram2x2 Imstake_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[3:2]), .q_b(q_b[59:56]),
     .q(q[59:56]), .wl(wl[13:12]));
cram2x2 Imstake_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[3:2]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[11:10]));
cram2x2 Imstake_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[3:2]), .q_b(q_b[51:48]), .q(q[51:48]),
     .wl(wl[9:8]));
cram2x2 Imstake_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[3:2]), .q_b(q_b[47:44]), .q(q[47:44]),
     .wl(wl[7:6]));
cram2x2 Imstake_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[3:2]), .q_b(q_b[43:40]), .q(q[43:40]),
     .wl(wl[5:4]));
cram2x2 Imstake_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[3:2]), .q_b(q_b[39:36]), .q(q[39:36]),
     .wl(wl[3:2]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[35:32]), .q(q[35:32]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - misc_module4_v3, View - schematic
// LAST TIME SAVED: Nov  5 15:38:16 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module misc_module4_v3 ( S_R, cbit, cbitb, clk, clkb, glb2local, sp4,
     bl, b, glb_netwk, l, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3,
     m, min0, min1, min2, min3, pgate, prog, r, reset_b, sp12,
     vdd_cntl, wl );
output  S_R, clk, clkb;


input  prog;

output [3:0]  glb2local;
output [7:0]  sp4;
output [63:0]  cbit;
output [63:0]  cbitb;

inout [3:0]  bl;

input [7:0]  sp12;
input [15:0]  pgate;
input [7:0]  min2;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [5:0]  lc_trk_g1;
input [1:0]  r;
input [7:0]  min1;
input [7:0]  glb_netwk;
input [1:0]  l;
input [5:0]  lc_trk_g0;
input [7:0]  min0;
input [1:0]  m;
input [5:0]  lc_trk_g2;
input [15:0]  reset_b;
input [5:0]  lc_trk_g3;
input [1:0]  b;
input [7:0]  min3;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  r_vdd;



inv_hvt I_inv2 ( .A(progb), .Y(progd));
inv_hvt I_inv1 ( .A(prog), .Y(progb));
pch_hvt  M0_15_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[15]), .S(r_vdd[15]));
pch_hvt  M0_14_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[14]), .S(r_vdd[14]));
pch_hvt  M0_13_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[13]), .S(r_vdd[13]));
pch_hvt  M0_12_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[12]), .S(r_vdd[12]));
pch_hvt  M0_11_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[11]), .S(r_vdd[11]));
pch_hvt  M0_10_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[10]), .S(r_vdd[10]));
pch_hvt  M0_9_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[9]), .S(r_vdd[9]));
pch_hvt  M0_8_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[8]), .S(r_vdd[8]));
pch_hvt  M0_7_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[7]), .S(r_vdd[7]));
pch_hvt  M0_6_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[6]), .S(r_vdd[6]));
pch_hvt  M0_5_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[5]), .S(r_vdd[5]));
pch_hvt  M0_4_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[4]), .S(r_vdd[4]));
pch_hvt  M0_3_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[3]), .S(r_vdd[3]));
pch_hvt  M0_2_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[2]), .S(r_vdd[2]));
pch_hvt  M0_1_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[1]), .S(r_vdd[1]));
pch_hvt  M0_0_ ( .D(vdd_), .B(vdd_), .G(vdd_cntl[0]), .S(r_vdd[0]));
clkmandcmuxrev0 I_clkmandcmuxrev0 ( .prog(progd),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]), .clk(clk),
     .clkb(clkb), .glb_netwk(glb_netwk[7:0]), .s_r(S_R),
     .glb2local(glb2local[3:0]), .cbit({cbit[2], cbit[1], cbit[0],
     cbit[27], cbit[25], cbit[26], cbit[24], cbit[23], cbit[21],
     cbit[22], cbit[20], cbit[19], cbit[17], cbit[18], cbit[16],
     cbit[15], cbit[13], cbit[14], cbit[12], cbit[31], cbit[29],
     cbit[30], cbit[28], cbit[11], cbit[9], cbit[10], cbit[8],
     cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}), .min2(min2[7:0]),
     .min1(min1[7:0]), .min0(min0[7:0]), .min3(min3[7:0]),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}));
sp12to4 I_sp12to4_7_ ( .prog(progd), .triout(sp4[7]),
     .cbitb(cbitb[62]), .drv(sp12[7]));
sp12to4 I_sp12to4_6_ ( .prog(progd), .triout(sp4[6]),
     .cbitb(cbitb[58]), .drv(sp12[6]));
sp12to4 I_sp12to4_5_ ( .prog(progd), .triout(sp4[5]),
     .cbitb(cbitb[54]), .drv(sp12[5]));
sp12to4 I_sp12to4_4_ ( .prog(progd), .triout(sp4[4]),
     .cbitb(cbitb[50]), .drv(sp12[4]));
sp12to4 I_sp12to4_3_ ( .prog(progd), .triout(sp4[3]),
     .cbitb(cbitb[46]), .drv(sp12[3]));
sp12to4 I_sp12to4_2_ ( .prog(progd), .triout(sp4[2]),
     .cbitb(cbitb[42]), .drv(sp12[2]));
sp12to4 I_sp12to4_1_ ( .prog(progd), .triout(sp4[1]), .cbitb(cbitb[5]),
     .drv(sp12[1]));
sp12to4 I_sp12to4_0_ ( .prog(progd), .triout(sp4[0]),
     .cbitb(cbitb[34]), .drv(sp12[0]));
sbox1 I_sbox1_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(progd));
sbox1 I_sbox1_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(progd));
cram16x4 I_cram16x4 ( .q(cbit[63:0]), .r_gnd(r_vdd[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));

endmodule
// Library - xpmem, Cell - cram2x2x6, View - schematic
// LAST TIME SAVED: May 11 14:44:08 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module cram2x2x6 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [23:0]  q;
output [23:0]  q_b;

inout [11:0]  bl;

input [1:0]  r_gnd;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_5_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_base, View - schematic
// LAST TIME SAVED: Nov  5 15:41:50 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_base ( lc_trk_out, sp4_out, bl, min0, min1, min2,
     min3, pgate, prog, reset_b, sp12_in, vdd_cntl, wl );


input  prog;

output [1:0]  sp4_out;
output [3:0]  lc_trk_out;

inout [11:0]  bl;

input [1:0]  vdd_cntl;
input [15:0]  min3;
input [1:0]  sp12_in;
input [15:0]  min1;
input [1:0]  reset_b;
input [15:0]  min2;
input [1:0]  pgate;
input [1:0]  wl;
input [15:0]  min0;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [23:0]  cbitb;

wire  [23:0]  cbit;



inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net60));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
g_mux I_mux2 ( .min(min2[15:0]), .prog(net60), .inmuxo(lc_trk_out[2]),
     .cbit({cbit[16], cbit[17], cbit[20], cbit[23], cbit[21]}),
     .cbitb({cbitb[16], cbitb[17], cbitb[20], cbitb[23], cbitb[21]}));
g_mux I_mux3 ( .min(min3[15:0]), .prog(net60), .inmuxo(lc_trk_out[3]),
     .cbit({cbit[18], cbit[19], cbit[22], cbit[15], cbit[13]}),
     .cbitb({cbitb[18], cbitb[19], cbitb[22], cbitb[15], cbitb[13]}));
g_mux I_mux1 ( .min(min1[15:0]), .prog(net60), .inmuxo(lc_trk_out[1]),
     .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}));
g_mux I_mux0 ( .min(min0[15:0]), .prog(net60), .inmuxo(lc_trk_out[0]),
     .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}));
cram2x2x6 I_mem2x2x6 ( .pgate(pgate[1:0]), .q(cbit[23:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[11:0]), .q_b(cbitb[23:0]));
sp12to4 I_sp12to4_1_ ( .triout(sp4_out[1]), .cbitb(cbitb[11]),
     .drv(sp12_in[1]), .prog(net60));
sp12to4 I_sp12to4_0_ ( .triout(sp4_out[0]), .cbitb(cbitb[9]),
     .drv(sp12_in[0]), .prog(net60));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0a, View - schematic
// LAST TIME SAVED: Jul 24 13:27:07 2007
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g0a ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g0;

inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;

input [7:0]  tnl_op;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[34], sp4_r_v_b[25]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[33], sp4_r_v_b[26]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[35], sp4_r_v_b[24]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[32], sp4_r_v_b[27]}),
     .sp4_out(sp4_v_b[13:12]), .sp12_in({sp12_v_b[3], sp12_v_b[1]}),
     .lc_trk_out(lc_trk_g0[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - pllcfg_sr26_40lp, View - schematic
// LAST TIME SAVED: Nov  2 13:15:11 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module pllcfg_sr26_40lp ( q, pll_sck, pll_sdi, reset );

input  pll_sck, pll_sdi, reset;

output [25:0]  q;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [25:0]  net16;



inv_hvt I472 ( .A(pll_sck), .Y(net11));
pll_ml_dff I4_25_ ( .R(reset), .D(q[24]), .CLK(net11), .QN(net16[0]),
     .Q(q[25]));
pll_ml_dff I4_24_ ( .R(reset), .D(q[23]), .CLK(net11), .QN(net16[1]),
     .Q(q[24]));
pll_ml_dff I4_23_ ( .R(reset), .D(q[22]), .CLK(net11), .QN(net16[2]),
     .Q(q[23]));
pll_ml_dff I4_22_ ( .R(reset), .D(q[21]), .CLK(net11), .QN(net16[3]),
     .Q(q[22]));
pll_ml_dff I4_21_ ( .R(reset), .D(q[20]), .CLK(net11), .QN(net16[4]),
     .Q(q[21]));
pll_ml_dff I4_20_ ( .R(reset), .D(q[19]), .CLK(net11), .QN(net16[5]),
     .Q(q[20]));
pll_ml_dff I4_19_ ( .R(reset), .D(q[18]), .CLK(net11), .QN(net16[6]),
     .Q(q[19]));
pll_ml_dff I4_18_ ( .R(reset), .D(q[17]), .CLK(net11), .QN(net16[7]),
     .Q(q[18]));
pll_ml_dff I4_17_ ( .R(reset), .D(q[16]), .CLK(net11), .QN(net16[8]),
     .Q(q[17]));
pll_ml_dff I4_16_ ( .R(reset), .D(q[15]), .CLK(net11), .QN(net16[9]),
     .Q(q[16]));
pll_ml_dff I4_15_ ( .R(reset), .D(q[14]), .CLK(net11), .QN(net16[10]),
     .Q(q[15]));
pll_ml_dff I4_14_ ( .R(reset), .D(q[13]), .CLK(net11), .QN(net16[11]),
     .Q(q[14]));
pll_ml_dff I4_13_ ( .R(reset), .D(q[12]), .CLK(net11), .QN(net16[12]),
     .Q(q[13]));
pll_ml_dff I4_12_ ( .R(reset), .D(q[11]), .CLK(net11), .QN(net16[13]),
     .Q(q[12]));
pll_ml_dff I4_11_ ( .R(reset), .D(q[10]), .CLK(net11), .QN(net16[14]),
     .Q(q[11]));
pll_ml_dff I4_10_ ( .R(reset), .D(q[9]), .CLK(net11), .QN(net16[15]),
     .Q(q[10]));
pll_ml_dff I4_9_ ( .R(reset), .D(q[8]), .CLK(net11), .QN(net16[16]),
     .Q(q[9]));
pll_ml_dff I4_8_ ( .R(reset), .D(q[7]), .CLK(net11), .QN(net16[17]),
     .Q(q[8]));
pll_ml_dff I4_7_ ( .R(reset), .D(q[6]), .CLK(net11), .QN(net16[18]),
     .Q(q[7]));
pll_ml_dff I4_6_ ( .R(reset), .D(q[5]), .CLK(net11), .QN(net16[19]),
     .Q(q[6]));
pll_ml_dff I4_5_ ( .R(reset), .D(q[4]), .CLK(net11), .QN(net16[20]),
     .Q(q[5]));
pll_ml_dff I4_4_ ( .R(reset), .D(q[3]), .CLK(net11), .QN(net16[21]),
     .Q(q[4]));
pll_ml_dff I4_3_ ( .R(reset), .D(q[2]), .CLK(net11), .QN(net16[22]),
     .Q(q[3]));
pll_ml_dff I4_2_ ( .R(reset), .D(q[1]), .CLK(net11), .QN(net16[23]),
     .Q(q[2]));
pll_ml_dff I4_1_ ( .R(reset), .D(q[0]), .CLK(net11), .QN(net16[24]),
     .Q(q[1]));
pll_ml_dff I4_0_ ( .R(reset), .D(pll_sdi), .CLK(net11), .QN(net16[25]),
     .Q(q[0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0b, View - schematic
// LAST TIME SAVED: Jul 24 13:26:14 2007
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g0b ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, glb2local, lft_op,
     pgate, prog, reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op,
     vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g0;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
input [3:0]  glb2local;
input [7:0]  bnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  top_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], glb2local[1]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], glb2local[2]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], glb2local[0]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], glb2local[3]}),
     .sp4_out(sp4_v_b[15:14]), .sp12_in({sp12_v_b[7], sp12_v_b[5]}),
     .lc_trk_out(lc_trk_g0[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1a, View - schematic
// LAST TIME SAVED: Jul 24 13:25:29 2007
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g1a ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [1:0]  wl;
input [7:0]  bnl_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[25], sp4_r_v_b[1]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[26], sp4_r_v_b[2]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[24], sp4_r_v_b[0]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[27], sp4_r_v_b[3]}),
     .sp4_out(sp4_v_b[17:16]), .sp12_in({sp12_v_b[11], sp12_v_b[9]}),
     .lc_trk_out(lc_trk_g1[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1b, View - schematic
// LAST TIME SAVED: Jul 24 13:24:39 2007
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g1b ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], sp4_r_v_b[5]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], sp4_r_v_b[6]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], sp4_r_v_b[4]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], sp4_r_v_b[7]}),
     .sp4_out(sp4_v_b[19:18]), .sp12_in({sp12_v_b[15], sp12_v_b[13]}),
     .lc_trk_out(lc_trk_g1[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2a, View - schematic
// LAST TIME SAVED: Jul 24 13:23:46 2007
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g2a ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g2;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;

input [7:0]  lft_op;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnl_op;
input [7:0]  slf_op;
input [1:0]  vdd_cntl;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  bnr_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[33], sp4_r_v_b[9]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[34], sp4_r_v_b[10]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[32], sp4_r_v_b[8]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[35], sp4_r_v_b[11]}),
     .sp4_out(sp4_v_b[21:20]), .sp12_in({sp12_v_b[19], sp12_v_b[17]}),
     .lc_trk_out(lc_trk_g2[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2b, View - schematic
// LAST TIME SAVED: Jul 24 13:22:58 2007
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g2b ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g2;

inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [7:0]  bnr_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[37], sp4_r_v_b[13]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[38], sp4_r_v_b[14]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[36], sp4_r_v_b[12]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[39], sp4_r_v_b[15]}),
     .sp4_out(sp4_v_b[23:22]), .sp12_in({sp12_v_b[23], sp12_v_b[21]}),
     .lc_trk_out(lc_trk_g2[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3a, View - schematic
// LAST TIME SAVED: May 11 14:44:38 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g3a ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g3;

inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  lft_op;
input [7:0]  bot_op;
input [7:0]  top_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
input [7:0]  tnr_op;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  bnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[41], sp4_r_v_b[17]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[42], sp4_r_v_b[18]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[40], sp4_r_v_b[16]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[43], sp4_r_v_b[19]}),
     .sp4_out(sp4_h_r[13:12]), .sp12_in({sp12_h_r[2], sp12_h_r[0]}),
     .lc_trk_out(lc_trk_g3[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3b, View - schematic
// LAST TIME SAVED: May 11 14:44:24 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4_g3b ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g3;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;

input [7:0]  top_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [7:0]  bot_op;
input [1:0]  wl;
input [7:0]  bnr_op;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [1:0]  vdd_cntl;
input [7:0]  slf_op;
input [7:0]  rgt_op;
input [7:0]  lft_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base I_gmux_12to4_g3b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[45], sp4_r_v_b[21]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[46], sp4_r_v_b[22]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[44], sp4_r_v_b[20]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[47], sp4_r_v_b[23]}),
     .sp4_out(sp4_h_r[15:14]), .sp12_in({sp12_h_r[6], sp12_h_r[4]}),
     .lc_trk_out(lc_trk_g3[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4, View - schematic
// LAST TIME SAVED: Jun  3 14:49:41 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module gmux_sp12to4 ( lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, bl,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bnl_op, bnr_op,
     bot_op, glb2local, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g3;

inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_r_v_b;

input [7:0]  rgt_op;
input [7:0]  top_op;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [7:0]  bnr_op;
input [3:0]  glb2local;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  tnr_op;
input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [7:0]  tnl_op;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_g0a I_g0_30 ( .vdd_cntl(vdd_cntl[1:0]),
     .pgate(pgate[1:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp12_v_b(sp12_v_b[23:0]), .lc_trk_g0(lc_trk_g0[3:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g0b I_g0_74 ( .vdd_cntl(vdd_cntl[3:2]),
     .pgate(pgate[3:2]), .glb2local(glb2local[3:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .lc_trk_g0(lc_trk_g0[7:4]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[3:2]), .reset_b(reset_b[3:2]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g1a I_g1_30 ( .vdd_cntl(vdd_cntl[5:4]),
     .pgate(pgate[5:4]), .bl(bl[11:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]),
     .lft_op(lft_op[7:0]), .prog(prog), .rgt_op(rgt_op[7:0]),
     .reset_b(reset_b[5:4]), .slf_op(slf_op[7:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .wl(wl[5:4]), .lc_trk_g1(lc_trk_g1[3:0]));
gmux_sp12to4_g1b I_g1_74 ( .vdd_cntl(vdd_cntl[7:6]),
     .pgate(pgate[7:6]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g1(lc_trk_g1[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g2a I_g2_30 ( .vdd_cntl(vdd_cntl[9:8]), .wl(wl[9:8]),
     .reset_b(reset_b[9:8]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[3:0]), .pgate(pgate[9:8]));
gmux_sp12to4_g2b I_g2_74 ( .vdd_cntl(vdd_cntl[11:10]),
     .pgate(pgate[11:10]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[11:10]),
     .reset_b(reset_b[11:10]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g3a I_g3_30 ( .vdd_cntl(vdd_cntl[13:12]), .wl(wl[13:12]),
     .reset_b(reset_b[13:12]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .pgate(pgate[13:12]), .lc_trk_g3(lc_trk_g3[3:0]));
gmux_sp12to4_g3b I_g3_74 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g3(lc_trk_g3[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .prog(prog),
     .bl(bl[11:0]), .reset_b(reset_b[15:14]), .wl(wl[15:14]));

endmodule
// Library - leafcell, Cell - bram_routing_tracks4_v3, View - schematic
// LAST TIME SAVED: Jan 12 15:56:31 2011
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_routing_tracks4_v3 ( bram_cbit, clk, cntl_cbit, lc_trk_g0,
     lc_trk_g1, lc_trk_g2, lc_trk_g3, s_r, bl, sp4_h_l, sp4_h_r,
     sp4_r_v_b, sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r, sp12_v_b,
     sp12_v_t, bnl_op, bnr_op, bot_op, glb_netwk, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );
output  clk, s_r;


input  prog;

output [7:0]  cntl_cbit;
output [7:0]  bram_cbit;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g3;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g1;

inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_t;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_l;
inout [23:0]  sp12_v_t;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_b;
inout [25:0]  bl;
inout [23:0]  sp12_h_r;

input [7:0]  bnr_op;
input [7:0]  bnl_op;
input [7:0]  tnl_op;
input [15:0]  pgate;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [7:0]  slf_op;
input [15:0]  vdd_cntl;
input [7:0]  glb_netwk;
input [7:0]  bot_op;
input [15:0]  wl;
input [15:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [63:0]  cbitb_c;

wire  [63:0]  cbit_c;

wire  [3:0]  net_glb2local;

wire  [1:0]  sp12_v_b_mid;

wire  [1:0]  sp12_h_r_mid;



inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(progd));
rm8w  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm8w  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm8w  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm8w  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm8w  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm8w  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm8w  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm8w  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm8w  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm8w  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm8w  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm8w  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm8w  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm8w  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm8w  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm8w  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm8w  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm8w  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm8w  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm8w  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm8w  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm8w  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm8w  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm8w  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
span4_ice8p I_sp4_sw ( .ccntrl_cbit(cntl_cbit[7:0]),
     .bram_cbit(bram_cbit[7:0]), .sp4_h_l(sp4_h_l[47:0]),
     .bl(bl[13:4]), .wl(wl[15:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_t(sp4_v_t[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .reset_b(reset_b[15:0]), .vdd_cntl(vdd_cntl[15:0]),
     .pgate(pgate[15:0]), .prog(progd));
misc_module4_v3 I_misc ( .wl(wl[15:0]), .sp12({sp12_h_r[22],
     sp12_h_r[20], sp12_h_r[18], sp12_h_r[16], sp12_h_r[14],
     sp12_h_r[12], sp12_h_r[10], sp12_h_r[8]}),
     .vdd_cntl(vdd_cntl[15:0]), .b(sp12_v_b[1:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .lc_trk_g1(lc_trk_g1[5:0]), .glb2local(net_glb2local[3:0]),
     .bl(bl[3:0]), .min3(glb_netwk[7:0]), .cbitb(cbitb_c[63:0]),
     .clk(clk), .min2(glb_netwk[7:0]), .reset_b(reset_b[15:0]),
     .prog(progd), .m(sp12_v_b_mid[1:0]), .r(sp12_h_r[1:0]), .S_R(s_r),
     .sp4(sp4_h_r[23:16]), .clkb(clkb), .cbit(cbit_c[63:0]),
     .lc_trk_g0(lc_trk_g0[5:0]), .glb_netwk(glb_netwk[7:0]),
     .min1(glb_netwk[7:0]), .min0(glb_netwk[7:0]),
     .l(sp12_h_r_mid[1:0]), .pgate(pgate[15:0]));
rm7y  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7y  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7y  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7y  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7y  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7y  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7y  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7y  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7y  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7y  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7y  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7y  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7y  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7y  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7y  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7y  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7y  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7y  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7y  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7y  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7y  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7y  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7y  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7y  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
gmux_sp12to4 I_gmux_sp12to4 ( .reset_b(reset_b[15:0]),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .lft_op(lft_op[7:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .glb2local(net_glb2local[3:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .wl(wl[15:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .bl(bl[25:14]), .lc_trk_g3(lc_trk_g3[7:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .vdd_cntl(vdd_cntl[15:0]), .prog(progd));

endmodule
// Library - leafcell, Cell - tiehis, View - schematic
// LAST TIME SAVED: May 12 18:03:23 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module tiehis ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - tiehi, View - schematic
// LAST TIME SAVED: Aug 18 15:41:32 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module tiehi ( tiehi );
output  tiehi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - odrv12_30, View - schematic
// LAST TIME SAVED: May 11 14:28:15 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module odrv12_30 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_h_r;

input  prog, slfop;

output [2:0]  sp4_h_r;
output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_r_v_b;

input [11:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



odrv12 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b[1]));
odrv12 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp12(sp12_v_b[0]));
odrv12 I70 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r));
odrv4 I69_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I71_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[2]));
odrv4 I71_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[1]));
odrv4 I71_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp4(sp4_v_b[0]));
odrv4 I73_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I73_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I73_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux3_0, View - schematic
// LAST TIME SAVED: May 12 18:06:38 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_4k_inmux3_0 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_h_r;

input  op, prog;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_h_r;

input [15:0]  min3;
input [15:0]  min0;
input [1:0]  reset_b;
input [15:0]  min2;
input [15:0]  min1;
input [15:0]  bl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [31:0]  cbitb;

wire  [31:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12_30 I_odrv74 ( .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
in_mux I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux I_in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - odrv12_74, View - schematic
// LAST TIME SAVED: May 12 12:56:34 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module odrv12_74 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_v_b;

input  prog, slfop;

output [2:0]  sp4_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_h_r;
output [2:0]  sp4_r_v_b;

input [11:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



odrv12 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp12(sp12_h_r[1]));
odrv12 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r[0]));
odrv12 I71 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b));
odrv4 I68_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I68_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I68_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I70_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp4(sp4_v_b[2]));
odrv4 I70_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[1]));
odrv4 I70_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[0]));
odrv4 I72_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux7_4, View - schematic
// LAST TIME SAVED: May 12 18:07:12 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_4k_inmux7_4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_v_b;

input  op, prog;

output [1:0]  sp12_h_r;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [2:0]  sp4_v_b;

input [15:0]  min0;
input [15:0]  min1;
input [15:0]  min3;
input [15:0]  min2;
input [15:0]  bl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [31:0]  cbitb;

wire  [31:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
odrv12_74 I_odrv74 ( .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));
in_mux I_in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux I_in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux I_in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux I_in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux_8x4, View - schematic
// LAST TIME SAVED: May 12 18:08:28 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_4k_inmux_8x4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, op, pgate, prog, reset_b, vdd_cntl, wl );

input  prog;

output [23:0]  sp4_h_r;
output [23:0]  sp4_r_v_b;
output [11:0]  sp12_v_b;
output [11:0]  sp12_h_r;
output [7:0]  in1;
output [7:0]  in2;
output [7:0]  in3;
output [7:0]  in0;
output [23:0]  sp4_v_b;

input [15:0]  bl;
input [7:0]  op;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g3;
input [7:0]  lc_trk_g2;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  reset_b;
input [15:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I81 ( .A(prog), .Y(progb));
inv I82 ( .A(progb), .Y(progd));
tiehis I10 ( .tiehi(tiehi));
bram_4k_inmux3_0 I3 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[3]), .sp12_v_b(sp12_v_b[7:6]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(progd), .pgate(pgate[7:6]),
     .op(op[3]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[11:9]), .sp4_r_v_b(sp4_r_v_b[11:9]),
     .sp4_h_r(sp4_h_r[11:9]), .in3(in3[3]), .in2(in2[3]), .in1(in1[3]),
     .in0(in0[3]));
bram_4k_inmux3_0 I2 ( .vdd_cntl(vdd_cntl[5:4]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[2]), .sp12_v_b(sp12_v_b[5:4]), .wl(wl[5:4]),
     .reset_b(reset_b[5:4]), .prog(progd), .pgate(pgate[5:4]),
     .op(op[2]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[8:6]), .sp4_r_v_b(sp4_r_v_b[8:6]),
     .sp4_h_r(sp4_h_r[8:6]), .in3(in3[2]), .in2(in2[2]), .in1(in1[2]),
     .in0(in0[2]));
bram_4k_inmux3_0 I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[1]), .sp12_v_b(sp12_v_b[3:2]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(progd), .pgate(pgate[3:2]),
     .op(op[1]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[5:3]), .sp4_r_v_b(sp4_r_v_b[5:3]),
     .sp4_h_r(sp4_h_r[5:3]), .in3(in3[1]), .in2(in2[1]), .in1(in1[1]),
     .in0(in0[1]));
bram_4k_inmux3_0 I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[0]), .sp12_v_b(sp12_v_b[1:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(progd), .pgate(pgate[1:0]),
     .op(op[0]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .in3(in3[0]), .in2(in2[0]), .in1(in1[0]),
     .in0(in0[0]));
bram_4k_inmux7_4 I6 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[15:0]),
     .wl(wl[13:12]), .reset_b(reset_b[13:12]), .prog(progd),
     .pgate(pgate[13:12]), .op(op[6]), .min3({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp12_v_b(sp12_v_b[10]), .sp12_h_r(sp12_h_r[9:8]),
     .sp4_v_b(sp4_v_b[20:18]), .sp4_r_v_b(sp4_r_v_b[20:18]),
     .sp4_h_r(sp4_h_r[20:18]), .in3(in3[6]), .in2(in2[6]),
     .in1(in1[6]), .in0(in0[6]));
bram_4k_inmux7_4 I5 ( .vdd_cntl(vdd_cntl[11:10]), .bl(bl[15:0]),
     .wl(wl[11:10]), .reset_b(reset_b[11:10]), .prog(progd),
     .pgate(pgate[11:10]), .op(op[5]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[9]), .sp12_h_r(sp12_h_r[7:6]),
     .sp4_v_b(sp4_v_b[17:15]), .sp4_r_v_b(sp4_r_v_b[17:15]),
     .sp4_h_r(sp4_h_r[17:15]), .in3(in3[5]), .in2(in2[5]),
     .in1(in1[5]), .in0(in0[5]));
bram_4k_inmux7_4 I4 ( .vdd_cntl(vdd_cntl[9:8]), .bl(bl[15:0]),
     .wl(wl[9:8]), .reset_b(reset_b[9:8]), .prog(progd),
     .pgate(pgate[9:8]), .op(op[4]), .min3({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .sp12_v_b(sp12_v_b[8]),
     .sp12_h_r(sp12_h_r[5:4]), .sp4_v_b(sp4_v_b[14:12]),
     .sp4_r_v_b(sp4_r_v_b[14:12]), .sp4_h_r(sp4_h_r[14:12]),
     .in3(in3[4]), .in2(in2[4]), .in1(in1[4]), .in0(in0[4]));
bram_4k_inmux7_4 I7 ( .vdd_cntl(vdd_cntl[15:14]), .bl(bl[15:0]),
     .wl(wl[15:14]), .reset_b(reset_b[15:14]), .prog(progd),
     .pgate(pgate[15:14]), .op(op[7]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[11]), .sp12_h_r(sp12_h_r[11:10]),
     .sp4_v_b(sp4_v_b[23:21]), .sp4_r_v_b(sp4_r_v_b[23:21]),
     .sp4_h_r(sp4_h_r[23:21]), .in3(in3[7]), .in2(in2[7]),
     .in1(in1[7]), .in0(in0[7]));

endmodule
// Library - ice1chip, Cell - bram_4kprouting_left_ice1p, View -
//schematic
// LAST TIME SAVED: Mar 31 14:01:12 2011
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_4kprouting_left_ice1p ( bm_bweb, bm_clkr2rf_n40,
     bm_clkw2rf_n40, bm_d, bm_ren2rf_n40, bm_wen2rf_n40, bram_aa,
     bram_ab, bram_cbit_bot, bram_cbit_top, cntl_cbit_bot,
     cntl_cbit_top, bl, sp4_h_l_bot, sp4_h_l_top, sp4_h_r_bot,
     sp4_h_r_top, sp4_r_v_b_bot, sp4_r_v_b_top, sp4_v_b_bot,
     sp4_v_b_top, sp4_v_t_top, sp12_h_l_bot, sp12_h_l_top,
     sp12_h_r_bot, sp12_h_r_top, sp12_v_b_bot, sp12_v_t_top,
     bnl_op_bot, bnr_op_bot, bot_op_bot, glb_netwk, lft_op_bot,
     lft_op_top, pgate_bot, pgate_top, prog, reset_b_bot, reset_b_top,
     rgt_op_bot, rgt_op_top, slf_op_bot, slf_op_top, tnl_op_top,
     tnr_op_top, top_op_top, vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top
     );
output  bm_clkr2rf_n40, bm_clkw2rf_n40, bm_ren2rf_n40, bm_wen2rf_n40;


input  prog;

output [7:0]  cntl_cbit_top;
output [10:0]  bram_aa;
output [7:0]  cntl_cbit_bot;
output [10:0]  bram_ab;
output [7:0]  bram_cbit_bot;
output [7:0]  bram_cbit_top;
output [15:0]  bm_d;
output [15:0]  bm_bweb;

inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_h_r_bot;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_top;
inout [41:0]  bl;
inout [47:0]  sp4_v_b_top;

input [7:0]  slf_op_top;
input [7:0]  rgt_op_top;
input [15:0]  pgate_top;
input [7:0]  slf_op_bot;
input [7:0]  lft_op_top;
input [7:0]  tnr_op_top;
input [15:0]  wl_bot;
input [7:0]  glb_netwk;
input [15:0]  wl_top;
input [7:0]  rgt_op_bot;
input [7:0]  tnl_op_top;
input [7:0]  bot_op_bot;
input [15:0]  vdd_cntl_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  lft_op_bot;
input [7:0]  bnr_op_bot;
input [7:0]  bnl_op_bot;
input [15:0]  reset_b_bot;
input [7:0]  top_op_top;
input [15:0]  reset_b_top;
input [15:0]  pgate_bot;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net194;

wire  [7:0]  net196;

wire  [7:0]  net229;

wire  [7:0]  net228;

wire  [7:0]  net195;

wire  [4:0]  in2_bot;

wire  [7:0]  net193;

wire  [7:0]  net226;

wire  [7:0]  net227;

wire  [4:0]  in2_top;

wire  [23:0]  sp12_v_b_top;



bram_routing_tracks4_v3 I_bram_routing_tracks4_v2_bot (
     .cntl_cbit(cntl_cbit_bot[7:0]), .bram_cbit(bram_cbit_bot[7:0]),
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .s_r(bm_wen2rf_n40), .wl({wl_bot[14],
     wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11],
     wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5],
     wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(rgt_op_top[7:0]),
     .tnl_op(lft_op_top[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3({net193[0], net193[1], net193[2], net193[3], net193[4],
     net193[5], net193[6], net193[7]}), .lc_trk_g2({net194[0],
     net194[1], net194[2], net194[3], net194[4], net194[5], net194[6],
     net194[7]}), .lc_trk_g1({net195[0], net195[1], net195[2],
     net195[3], net195[4], net195[5], net195[6], net195[7]}),
     .lc_trk_g0({net196[0], net196[1], net196[2], net196[3], net196[4],
     net196[5], net196[6], net196[7]}), .clk(bm_clkw2rf_n40),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4_v3 I_bram_routing_tracks4_v2_top (
     .cntl_cbit(cntl_cbit_top[7:0]), .bram_cbit(bram_cbit_top[7:0]),
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .s_r(bm_ren2rf_n40), .wl({wl_top[14],
     wl_top[15], wl_top[12], wl_top[13], wl_top[10], wl_top[11],
     wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5],
     wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bot_op(slf_op_bot[7:0]),
     .bnr_op(rgt_op_bot[7:0]), .bnl_op(lft_op_bot[7:0]),
     .lc_trk_g3({net226[0], net226[1], net226[2], net226[3], net226[4],
     net226[5], net226[6], net226[7]}), .lc_trk_g2({net227[0],
     net227[1], net227[2], net227[3], net227[4], net227[5], net227[6],
     net227[7]}), .lc_trk_g1({net228[0], net228[1], net228[2],
     net228[3], net228[4], net228[5], net228[6], net228[7]}),
     .lc_trk_g0({net229[0], net229[1], net229[2], net229[3], net229[4],
     net229[5], net229[6], net229[7]}), .clk(bm_clkr2rf_n40),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_bot (
     .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15], vdd_cntl_bot[12],
     vdd_cntl_bot[13], vdd_cntl_bot[10], vdd_cntl_bot[11],
     vdd_cntl_bot[8], vdd_cntl_bot[9], vdd_cntl_bot[6],
     vdd_cntl_bot[7], vdd_cntl_bot[4], vdd_cntl_bot[5],
     vdd_cntl_bot[2], vdd_cntl_bot[3], vdd_cntl_bot[0],
     vdd_cntl_bot[1]}), .bl(bl[41:26]), .wl({wl_bot[14], wl_bot[15],
     wl_bot[12], wl_bot[13], wl_bot[10], wl_bot[11], wl_bot[8],
     wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4], wl_bot[5], wl_bot[2],
     wl_bot[3], wl_bot[0], wl_bot[1]}), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .op(slf_op_bot[7:0]), .lc_trk_g3({net193[0],
     net193[1], net193[2], net193[3], net193[4], net193[5], net193[6],
     net193[7]}), .lc_trk_g2({net194[0], net194[1], net194[2],
     net194[3], net194[4], net194[5], net194[6], net194[7]}),
     .lc_trk_g1({net195[0], net195[1], net195[2], net195[3], net195[4],
     net195[5], net195[6], net195[7]}), .lc_trk_g0({net196[0],
     net196[1], net196[2], net196[3], net196[4], net196[5], net196[6],
     net196[7]}), .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6],
     sp12_h_r_bot[20], sp12_h_r_bot[4], sp12_h_r_bot[18],
     sp12_h_r_bot[2], sp12_h_r_bot[16], sp12_h_r_bot[0],
     sp12_h_r_bot[14], sp12_h_r_bot[12], sp12_h_r_bot[10],
     sp12_h_r_bot[8]}), .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30],
     sp4_v_b_bot[14], sp4_v_b_bot[44], sp4_v_b_bot[28],
     sp4_v_b_bot[12], sp4_v_b_bot[42], sp4_v_b_bot[26],
     sp4_v_b_bot[10], sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8],
     sp4_v_b_bot[38], sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36],
     sp4_v_b_bot[20], sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18],
     sp4_v_b_bot[2], sp4_v_b_bot[32], sp4_v_b_bot[16],
     sp4_v_b_bot[0]}), .sp4_r_v_b({sp4_r_v_b_bot[47],
     sp4_r_v_b_bot[31], sp4_r_v_b_bot[15], sp4_r_v_b_bot[45],
     sp4_r_v_b_bot[29], sp4_r_v_b_bot[13], sp4_r_v_b_bot[43],
     sp4_r_v_b_bot[27], sp4_r_v_b_bot[11], sp4_r_v_b_bot[41],
     sp4_r_v_b_bot[25], sp4_r_v_b_bot[9], sp4_r_v_b_bot[39],
     sp4_r_v_b_bot[23], sp4_r_v_b_bot[7], sp4_r_v_b_bot[37],
     sp4_r_v_b_bot[21], sp4_r_v_b_bot[5], sp4_r_v_b_bot[35],
     sp4_r_v_b_bot[19], sp4_r_v_b_bot[3], sp4_r_v_b_bot[33],
     sp4_r_v_b_bot[17], sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46],
     sp4_h_r_bot[30], sp4_h_r_bot[14], sp4_h_r_bot[44],
     sp4_h_r_bot[28], sp4_h_r_bot[12], sp4_h_r_bot[42],
     sp4_h_r_bot[26], sp4_h_r_bot[10], sp4_h_r_bot[40],
     sp4_h_r_bot[24], sp4_h_r_bot[8], sp4_h_r_bot[38], sp4_h_r_bot[22],
     sp4_h_r_bot[6], sp4_h_r_bot[36], sp4_h_r_bot[20], sp4_h_r_bot[4],
     sp4_h_r_bot[34], sp4_h_r_bot[18], sp4_h_r_bot[2], sp4_h_r_bot[32],
     sp4_h_r_bot[16], sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]),
     .in2({in2_bot[4:0], bram_aa[10:8]}), .in1(bm_d[7:0]),
     .in0(bram_aa[7:0]), .sp12_v_b({sp12_v_b_bot[14], sp12_v_b_bot[12],
     sp12_v_b_bot[10], sp12_v_b_bot[8], sp12_v_b_bot[22],
     sp12_v_b_bot[6], sp12_v_b_bot[20], sp12_v_b_bot[4],
     sp12_v_b_bot[18], sp12_v_b_bot[2], sp12_v_b_bot[16],
     sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I_bram_4k_inmux_8x4_top (
     .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15], vdd_cntl_top[12],
     vdd_cntl_top[13], vdd_cntl_top[10], vdd_cntl_top[11],
     vdd_cntl_top[8], vdd_cntl_top[9], vdd_cntl_top[6],
     vdd_cntl_top[7], vdd_cntl_top[4], vdd_cntl_top[5],
     vdd_cntl_top[2], vdd_cntl_top[3], vdd_cntl_top[0],
     vdd_cntl_top[1]}), .bl(bl[41:26]), .sp12_v_b({sp12_v_b_top[14],
     sp12_v_b_top[12], sp12_v_b_top[10], sp12_v_b_top[8],
     sp12_v_b_top[22], sp12_v_b_top[6], sp12_v_b_top[20],
     sp12_v_b_top[4], sp12_v_b_top[18], sp12_v_b_top[2],
     sp12_v_b_top[16], sp12_v_b_top[0]}), .wl({wl_top[14], wl_top[15],
     wl_top[12], wl_top[13], wl_top[10], wl_top[11], wl_top[8],
     wl_top[9], wl_top[6], wl_top[7], wl_top[4], wl_top[5], wl_top[2],
     wl_top[3], wl_top[0], wl_top[1]}), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .op(slf_op_top[7:0]), .lc_trk_g3({net226[0],
     net226[1], net226[2], net226[3], net226[4], net226[5], net226[6],
     net226[7]}), .lc_trk_g2({net227[0], net227[1], net227[2],
     net227[3], net227[4], net227[5], net227[6], net227[7]}),
     .lc_trk_g1({net228[0], net228[1], net228[2], net228[3], net228[4],
     net228[5], net228[6], net228[7]}), .lc_trk_g0({net229[0],
     net229[1], net229[2], net229[3], net229[4], net229[5], net229[6],
     net229[7]}), .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6],
     sp12_h_r_top[20], sp12_h_r_top[4], sp12_h_r_top[18],
     sp12_h_r_top[2], sp12_h_r_top[16], sp12_h_r_top[0],
     sp12_h_r_top[14], sp12_h_r_top[12], sp12_h_r_top[10],
     sp12_h_r_top[8]}), .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30],
     sp4_v_b_top[14], sp4_v_b_top[44], sp4_v_b_top[28],
     sp4_v_b_top[12], sp4_v_b_top[42], sp4_v_b_top[26],
     sp4_v_b_top[10], sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8],
     sp4_v_b_top[38], sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36],
     sp4_v_b_top[20], sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18],
     sp4_v_b_top[2], sp4_v_b_top[32], sp4_v_b_top[16],
     sp4_v_b_top[0]}), .sp4_r_v_b({sp4_r_v_b_top[47],
     sp4_r_v_b_top[31], sp4_r_v_b_top[15], sp4_r_v_b_top[45],
     sp4_r_v_b_top[29], sp4_r_v_b_top[13], sp4_r_v_b_top[43],
     sp4_r_v_b_top[27], sp4_r_v_b_top[11], sp4_r_v_b_top[41],
     sp4_r_v_b_top[25], sp4_r_v_b_top[9], sp4_r_v_b_top[39],
     sp4_r_v_b_top[23], sp4_r_v_b_top[7], sp4_r_v_b_top[37],
     sp4_r_v_b_top[21], sp4_r_v_b_top[5], sp4_r_v_b_top[35],
     sp4_r_v_b_top[19], sp4_r_v_b_top[3], sp4_r_v_b_top[33],
     sp4_r_v_b_top[17], sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46],
     sp4_h_r_top[30], sp4_h_r_top[14], sp4_h_r_top[44],
     sp4_h_r_top[28], sp4_h_r_top[12], sp4_h_r_top[42],
     sp4_h_r_top[26], sp4_h_r_top[10], sp4_h_r_top[40],
     sp4_h_r_top[24], sp4_h_r_top[8], sp4_h_r_top[38], sp4_h_r_top[22],
     sp4_h_r_top[6], sp4_h_r_top[36], sp4_h_r_top[20], sp4_h_r_top[4],
     sp4_h_r_top[34], sp4_h_r_top[18], sp4_h_r_top[2], sp4_h_r_top[32],
     sp4_h_r_top[16], sp4_h_r_top[0]}), .in3(bm_bweb[15:8]),
     .in2({in2_top[4:0], bram_ab[10:8]}), .in1(bm_d[15:8]),
     .in0(bram_ab[7:0]));

endmodule
// Library - leafcell, Cell - bram_2mux, View - schematic
// LAST TIME SAVED: Jan  2 17:58:11 2011
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_2mux ( out, c, in0, in1 );
output  out;

input  c, in0, in1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate I14 ( .in(in1), .out(net52), .pp(net045), .nn(c));
txgate I33 ( .in(in0), .out(net52), .pp(c), .nn(net045));
inv I15 ( .A(net52), .Y(net029));
inv I0 ( .A(net029), .Y(out));
inv_hvt I1 ( .A(c), .Y(net045));

endmodule
// Library - leafcell, Cell - bram_cascade_addr, View - schematic
// LAST TIME SAVED: Jan  2 17:57:15 2011
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_cascade_addr ( addr_2bot, addr_muxo, addr, addr_top, cbit,
     prog );

input  prog;

output [10:0]  addr_2bot;
output [10:0]  addr_muxo;

input [10:0]  addr_top;
input [10:0]  addr;
input [1:0]  cbit;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(cbit[1]), .Y(net71));
bram_bufferx4 I33 ( .in(cbit[0]), .out(net66));
nor2_hvt I65 ( .A(prog), .B(net71), .Y(net69));
spn4dbuf I_addr_2bot_10_ ( .T(net69), .A(addr_muxo[10]),
     .Y(addr_2bot[10]));
spn4dbuf I_addr_2bot_9_ ( .T(net69), .A(addr_muxo[9]),
     .Y(addr_2bot[9]));
spn4dbuf I_addr_2bot_8_ ( .T(net69), .A(addr_muxo[8]),
     .Y(addr_2bot[8]));
spn4dbuf I_addr_2bot_7_ ( .T(net69), .A(addr_muxo[7]),
     .Y(addr_2bot[7]));
spn4dbuf I_addr_2bot_6_ ( .T(net69), .A(addr_muxo[6]),
     .Y(addr_2bot[6]));
spn4dbuf I_addr_2bot_5_ ( .T(net69), .A(addr_muxo[5]),
     .Y(addr_2bot[5]));
spn4dbuf I_addr_2bot_4_ ( .T(net69), .A(addr_muxo[4]),
     .Y(addr_2bot[4]));
spn4dbuf I_addr_2bot_3_ ( .T(net69), .A(addr_muxo[3]),
     .Y(addr_2bot[3]));
spn4dbuf I_addr_2bot_2_ ( .T(net69), .A(addr_muxo[2]),
     .Y(addr_2bot[2]));
spn4dbuf I_addr_2bot_1_ ( .T(net69), .A(addr_muxo[1]),
     .Y(addr_2bot[1]));
spn4dbuf I_addr_2bot_0_ ( .T(net69), .A(addr_muxo[0]),
     .Y(addr_2bot[0]));
bram_2mux I_bram_2mux_10_ ( .c(net66), .out(addr_muxo[10]),
     .in0(addr[10]), .in1(addr_top[10]));
bram_2mux I_bram_2mux_9_ ( .c(net66), .out(addr_muxo[9]),
     .in0(addr[9]), .in1(addr_top[9]));
bram_2mux I_bram_2mux_8_ ( .c(net66), .out(addr_muxo[8]),
     .in0(addr[8]), .in1(addr_top[8]));
bram_2mux I_bram_2mux_7_ ( .c(net66), .out(addr_muxo[7]),
     .in0(addr[7]), .in1(addr_top[7]));
bram_2mux I_bram_2mux_6_ ( .c(net66), .out(addr_muxo[6]),
     .in0(addr[6]), .in1(addr_top[6]));
bram_2mux I_bram_2mux_5_ ( .c(net66), .out(addr_muxo[5]),
     .in0(addr[5]), .in1(addr_top[5]));
bram_2mux I_bram_2mux_4_ ( .c(net66), .out(addr_muxo[4]),
     .in0(addr[4]), .in1(addr_top[4]));
bram_2mux I_bram_2mux_3_ ( .c(net66), .out(addr_muxo[3]),
     .in0(addr[3]), .in1(addr_top[3]));
bram_2mux I_bram_2mux_2_ ( .c(net66), .out(addr_muxo[2]),
     .in0(addr[2]), .in1(addr_top[2]));
bram_2mux I_bram_2mux_1_ ( .c(net66), .out(addr_muxo[1]),
     .in0(addr[1]), .in1(addr_top[1]));
bram_2mux I_bram_2mux_0_ ( .c(net66), .out(addr_muxo[0]),
     .in0(addr[0]), .in1(addr_top[0]));

endmodule
// Library - leafcell, Cell - bram_2mux_lvt, View - schematic
// LAST TIME SAVED: Nov  8 18:34:36 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module bram_2mux_lvt ( out, c, in0, in1 );
output  out;

input  c, in0, in1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I14 ( .in(in1), .out(net52), .pp(net045), .nn(c));
txgate_lvt I33 ( .in(in0), .out(net52), .pp(c), .nn(net045));
inv_lvt I15 ( .A(net52), .Y(net029));
inv_lvt I0 ( .A(net029), .Y(out));
inv_hvt I1 ( .A(c), .Y(net045));

endmodule
// Library - misc, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: May 13 14:45:34 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module ml_mux2_hvt ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - tielo, View - schematic
// LAST TIME SAVED: Jul 23 17:02:44 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module tielo ( tielo );
output  tielo;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M1 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));
nch_hvt  M2 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - leafcell, Cell - rf_4k_n40, View - schematic
// LAST TIME SAVED: Aug 16 16:53:19 2010
// NETLIST TIME: May  5 11:56:41 2011
`timescale 1ns / 1ns 

module rf_4k_n40 ( Q, AA, AB, AMA, AMB, BIST, BWEB, BWEBM, CLKR, CLKW,
     D, DM, PD, REB, REBM, WEB, WEBM );

input  BIST, CLKR, CLKW, PD, REB, REBM, WEB, WEBM;

output [15:0]  Q;

input [7:0]  AMA;
input [15:0]  DM;
input [7:0]  AA;
input [15:0]  D;
input [15:0]  BWEB;
input [15:0]  BWEBM;
input [7:0]  AB;
input [7:0]  AMB;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: May 12 17:56:32 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ml_mux2_hvt_schematic ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - bram_dff_mux, View - schematic
// LAST TIME SAVED: Oct  4 14:55:56 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_dff_mux ( q, bm_q, bm_sdi, ce, clk, rcapmux_en, rst );
output  q;

input  bm_q, bm_sdi, ce, clk, rcapmux_en, rst;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_mux2_hvt I5 ( .in1(net14), .in0(q), .out(net020), .sel(ce));
ml_dff I_ml_dff ( .R(rst), .D(net020), .CLK(clk), .QN(net10), .Q(q));
ml_mux2_hvt_schematic I1 ( .in1(bm_q), .in0(bm_sdi), .out(net14),
     .sel(rcapmux_en));

endmodule
// Library - leafcell, Cell - bram_4k_sr_v1, View - schematic
// LAST TIME SAVED: Oct 29 10:24:13 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_4k_sr_v1 ( bm_dm, bm_sdo, bm_sweb, clk, rcapmux_en, rst,
     bm_q, bm_sdi, wdummymux_en );
output  bm_sdo;

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



ml_dff I_dff15 ( .R(rst), .D(bm_dm[14]), .CLK(clk), .QN(net0258),
     .Q(rdummy_reg));
ml_dff I_dff0 ( .R(rst), .D(bm_sdi), .CLK(clk), .QN(net157),
     .Q(wdummy_reg));
bram_dff_mux I_dff_mux_15_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[14]),
     .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I_dff_mux_14_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[13]),
     .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I_dff_mux_13_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[12]),
     .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I_dff_mux_12_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[11]),
     .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I_dff_mux_11_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[10]),
     .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I_dff_mux_10_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[9]),
     .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I_dff_mux_9_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[8]),
     .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I_dff_mux_8_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[7]),
     .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I_dff_mux_7_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[6]),
     .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I_dff_mux_6_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[5]),
     .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I_dff_mux_5_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[4]),
     .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I_dff_mux_4_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[3]),
     .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I_dff_mux_3_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[2]),
     .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I_dff_mux_2_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_dm[1]),
     .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I_dff_mux_1_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(net150),
     .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I_dff_mux_0_ ( .rst(rst), .ce(bm_sweb),
     .rcapmux_en(rcapmux_en), .clk(clk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[0]), .q(bm_dm[0]));
ml_mux2_hvt_schematic I_mux15 ( .in1(rdummy_reg), .in0(bm_dm[15]),
     .out(bm_sdo), .sel(rcapmux_en));
ml_mux2_hvt_schematic I_mux0 ( .in1(wdummy_reg), .in0(bm_dm[0]),
     .out(net150), .sel(wdummymux_en));

endmodule
// Library - leafcell, Cell - bram_4k_n40, View - schematic
// LAST TIME SAVED: Jan  2 17:48:30 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_4k_n40 ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_pd, bm_rcapmux_en, bm_ren, bm_sa,
     bm_sclk, bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en,
     bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_pd, bm_rcapmux_en, bm_ren,
     bm_sclk, bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en,
     bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [7:0]  bm_sa;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [7:0]  bm_aa;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  bm_dm;



bram_2mux_lvt I22 ( .c(bm_init), .out(net108), .in0(bm_clkr),
     .in1(bm_sclkrw));
bram_2mux_lvt I23 ( .c(bm_init), .out(net110), .in0(bm_clkw),
     .in1(bm_sclkrw));
inv_lvt I6 ( .A(bm_ren), .Y(reb));
inv_lvt I5 ( .A(bm_wen), .Y(web));
ml_mux2_hvt I20 ( .in1(net90), .in0(bm_pd), .out(net0118),
     .sel(bm_init));
bram_bufferx4 I19 ( .in(net0118), .out(net0111));
rf_4k_n40 I_rf_4k ( .PD(net0111), .DM(bm_dm[15:0]), .WEBM(bm_sweb),
     .WEB(web), .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]),
     .CLKW(net110), .CLKR(net108), .BWEBM({net0128, net0128, net0128,
     net0128, net0128, net0128, net0128, net0128, net0128, net0128,
     net0128, net0128, net0128, net0128, net0128, net0128}),
     .BWEB(bm_bweb[15:0]), .BIST(bm_init), .AMB(bm_sa[7:0]),
     .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]), .AA(bm_aa[7:0]),
     .Q(bm_q[15:0]));
bram_4k_sr_v1 I_bram_4k_sr ( .bm_sdo(bm_sdo), .bm_dm(bm_dm[15:0]),
     .rst(net90), .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
tielo I15 ( .tielo(net0128));
tielo I18 ( .tielo(net90));

endmodule
// Library - leafcell, Cell - o_mux_out_bram, View - schematic
// LAST TIME SAVED: Dec  3 13:44:44 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module o_mux_out_bram ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_lvt I181 ( .A(in), .Y(out));

endmodule
// Library - leafcell, Cell - bram_3muxinv, View - schematic
// LAST TIME SAVED: Nov  8 18:26:34 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_3muxinv ( out, c, .cdsNet0(in[0]), .cdsNet0(in[1]),
     .cdsNet0(in[2]) );
output  out;


input [2:0]  in;
input [1:0]  c;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  ci;

wire  [1:0]  cb;



txgate_lvt I21 ( .in(in[2]), .out(net52), .pp(cb[1]), .nn(ci[1]));
txgate_lvt I33 ( .in(in[0]), .out(net52), .pp(net048), .nn(net053));
txgate_lvt I20 ( .in(in[1]), .out(net52), .pp(net045), .nn(net051));
inv_lvt I0 ( .A(net52), .Y(out));
nand2_hvt I15 ( .A(ci[0]), .Y(net045), .B(cb[1]));
nand2_hvt I2 ( .A(cb[0]), .Y(net048), .B(cb[1]));
inv_hvt I19 ( .A(net045), .Y(net051));
inv_hvt I18 ( .A(net048), .Y(net053));
inv_hvt I14_1_ ( .A(c[1]), .Y(cb[1]));
inv_hvt I14_0_ ( .A(c[0]), .Y(cb[0]));
inv_hvt I1_1_ ( .A(cb[1]), .Y(ci[1]));
inv_hvt I1_0_ ( .A(cb[0]), .Y(ci[0]));

endmodule
// Library - leafcell, Cell - bram_2muxinv, View - schematic
// LAST TIME SAVED: Nov  8 18:25:27 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_2muxinv ( out, c, in0, in1 );
output  out;

input  c, in0, in1;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I13 ( .in(in1), .out(net52), .pp(net045), .nn(c));
txgate_lvt I33 ( .in(in0), .out(net52), .pp(c), .nn(net045));
inv_lvt I0 ( .A(net52), .Y(out));
inv_hvt I1 ( .A(c), .Y(net045));

endmodule
// Library - leafcell, Cell - bram_rd_decoder0to7, View - schematic
// LAST TIME SAVED: Jan  2 18:16:33 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_rd_decoder0to7 ( rd, c, raq, rdi );


output [7:0]  rd;

input [10:8]  raq;
input [1:0]  c;
input [7:0]  rdi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cd;

wire  [10:10]  raqb;

wire  [1:0]  cb;



nand2 I65 ( .A(mode16_b), .Y(raq8_b), .B(raq[8]));
inv I85 ( .A(raq[9]), .Y(net0245));
inv I68 ( .A(raq[10]), .Y(raqb[10]));
o_mux_out_bram I69 ( .in(net360), .out(rd[0]));
o_mux_out_bram I92 ( .out(rd[7]), .in(net378));
o_mux_out_bram I91 ( .out(rd[6]), .in(net333));
o_mux_out_bram I90 ( .out(rd[5]), .in(net372));
o_mux_out_bram I89 ( .out(rd[4]), .in(net362));
o_mux_out_bram I88 ( .out(rd[3]), .in(net390));
o_mux_out_bram I87 ( .out(rd[2]), .in(net329));
o_mux_out_bram I86 ( .out(rd[1]), .in(net384));
inv_lvt I104 ( .A(rdi[7]), .Y(net378));
nand2_hvt I106 ( .A(cd[1]), .Y(mode4_b), .B(cb[0]));
nand2_hvt I107 ( .A(cd[1]), .Y(mode2_b), .B(cd[0]));
nand2_hvt I105 ( .A(cb[1]), .Y(mode16_b), .B(cb[0]));
inv_hvt I22_1_ ( .A(cb[1]), .Y(cd[1]));
inv_hvt I22_0_ ( .A(cb[0]), .Y(cd[0]));
inv_hvt I53_1_ ( .A(c[1]), .Y(cb[1]));
inv_hvt I53_0_ ( .A(c[0]), .Y(cb[0]));
bram_3muxinv I3 ( net390, {mode2_b, raqb[10]}, net285, net357, rdi[3]);
bram_2muxinv I35 ( .in1(rdi[2]), .c(raq8_b), .out(net329),
     .in0(rdi[3]));
bram_2muxinv I36 ( .in1(rdi[4]), .c(raq8_b), .out(net362),
     .in0(rdi[5]));
bram_2muxinv I37 ( .in1(rdi[6]), .c(raq8_b), .out(net333),
     .in0(rdi[7]));
bram_2muxinv I34 ( .in1(rdi[0]), .c(raq8_b), .out(net360),
     .in0(rdi[1]));
bram_2muxinv I42 ( .in1(net360), .c(net0245), .out(net357),
     .in0(net329));
bram_2muxinv I43 ( .in1(net362), .c(net0245), .out(net285),
     .in0(net333));
bram_2muxinv I49 ( .in1(rdi[5]), .c(mode4_b), .out(net372),
     .in0(net285));
bram_2muxinv I50 ( .in1(rdi[1]), .c(mode4_b), .out(net384),
     .in0(net357));

endmodule
// Library - leafcell, Cell - bram_4muxinv, View - schematic
// LAST TIME SAVED: Jan  2 18:09:52 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_4muxinv ( out, .cdsNet0(in[0]), .cdsNet0(in[1]),
     .cdsNet0(in[2]), .cdsNet0(in[3]), sel, selb );
output  out;


input [3:0]  selb;
input [3:0]  sel;
input [3:0]  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I0 ( .A(net47), .Y(out));
txgate_lvt I19 ( .in(in[3]), .out(net47), .pp(selb[3]), .nn(sel[3]));
txgate_lvt I17 ( .in(in[2]), .out(net47), .pp(selb[2]), .nn(sel[2]));
txgate_lvt I33 ( .in(in[0]), .out(net47), .pp(selb[0]), .nn(sel[0]));
txgate_lvt I16 ( .in(in[1]), .out(net47), .pp(selb[1]), .nn(sel[1]));

endmodule
// Library - leafcell, Cell - mux4plldly, View - schematic
// LAST TIME SAVED: Jun 28 10:07:29 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module mux4plldly ( mout, cbit, min );
output  mout;


input [1:0]  cbit;
input [3:0]  min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cbit_b;



txgate_hvt I11 ( .in(net_2_0), .out(net52), .pp(cbit[1]),
     .nn(cbit_b[1]));
txgate_hvt I8 ( .in(min[1]), .out(net_2_0), .pp(cbit_b[0]),
     .nn(cbit[0]));
txgate_hvt I9 ( .in(min[2]), .out(net_2_1), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I12 ( .in(net_2_1), .out(net52), .pp(cbit_b[1]),
     .nn(cbit[1]));
txgate_hvt Itg20 ( .in(min[0]), .out(net_2_0), .pp(cbit[0]),
     .nn(cbit_b[0]));
txgate_hvt I10 ( .in(min[3]), .out(net_2_1), .pp(cbit_b[0]),
     .nn(cbit[0]));
inv_hvt I1_1_ ( .A(cbit[1]), .Y(cbit_b[1]));
inv_hvt I1_0_ ( .A(cbit[0]), .Y(cbit_b[0]));
inv_hvt I0 ( .A(net52), .Y(mout));

endmodule
// Library - leafcell, Cell - bram_wd_decoder0to7, View - schematic
// LAST TIME SAVED: Jan  2 18:06:52 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_wd_decoder0to7 ( wd, sel, wdi );


output [7:0]  wd;

input [3:0]  sel;
input [7:0]  wdi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  selb;

wire  [3:0]  net0210;

wire  [3:0]  net0202;



inv I74 ( .A(wdi[1]), .Y(net176));
inv I75 ( .A(wdi[2]), .Y(net162));
inv I76 ( .A(wdi[3]), .Y(net177));
inv I77 ( .A(wdi[3]), .Y(net159));
inv I78 ( .A(wdi[4]), .Y(net150));
inv I79 ( .A(wdi[5]), .Y(net152));
inv I80 ( .A(wdi[6]), .Y(net138));
inv I81 ( .A(wdi[7]), .Y(net132));
inv I22 ( .A(wdi[0]), .Y(net174));
bram_4muxinv I95 ( wd[5], net152, net150, net152, net159, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
bram_4muxinv I96 ( wd[6], net138, net138, net152, net159, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
bram_4muxinv I97 ( wd[7], net132, net138, net152, net159, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
bram_4muxinv I91 ( wd[1], net176, net174, net176, net177, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
bram_4muxinv I92 ( wd[2], net162, net162, net176, net177, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
bram_4muxinv I93 ( wd[3], net177, net162, net176, net159, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
bram_4muxinv I94 ( wd[4], net150, net150, net152, net159, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
bram_4muxinv I3 ( wd[0], net174, net174, net176, net177, {net0202[0],
     net0202[1], net0202[2], net0202[3]}, selb[3:0]);
inv_hvt I122_3_ ( .A(net0210[0]), .Y(net0202[0]));
inv_hvt I122_2_ ( .A(net0210[1]), .Y(net0202[1]));
inv_hvt I122_1_ ( .A(net0210[2]), .Y(net0202[2]));
inv_hvt I122_0_ ( .A(net0210[3]), .Y(net0202[3]));
inv_hvt I125_3_ ( .A(sel[3]), .Y(selb[3]));
inv_hvt I125_2_ ( .A(sel[2]), .Y(selb[2]));
inv_hvt I125_1_ ( .A(sel[1]), .Y(selb[1]));
inv_hvt I125_0_ ( .A(sel[0]), .Y(selb[0]));
inv_hvt I123_3_ ( .A(sel[3]), .Y(net0210[0]));
inv_hvt I123_2_ ( .A(sel[2]), .Y(net0210[1]));
inv_hvt I123_1_ ( .A(sel[1]), .Y(net0210[2]));
inv_hvt I123_0_ ( .A(sel[0]), .Y(net0210[3]));

endmodule
// Library - leafcell, Cell - bram_4mux, View - schematic
// LAST TIME SAVED: Jan  2 18:15:04 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_4mux ( out, .cdsNet0(in[0]), .cdsNet0(in[1]),
     .cdsNet0(in[2]), .cdsNet0(in[3]), sel, selb );
output  out;


input [3:0]  sel;
input [3:0]  in;
input [3:0]  selb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv I13 ( .A(net62), .Y(net48));
inv I14 ( .A(net48), .Y(out));
txgate_lvt I26 ( .in(in[3]), .out(net62), .pp(selb[3]), .nn(sel[3]));
txgate_lvt I33 ( .in(in[0]), .out(net62), .pp(selb[0]), .nn(sel[0]));
txgate_lvt I24 ( .in(in[1]), .out(net62), .pp(selb[1]), .nn(sel[1]));
txgate_lvt I25 ( .in(in[2]), .out(net62), .pp(selb[2]), .nn(sel[2]));

endmodule
// Library - leafcell, Cell - bram_wd_bweb, View - schematic
// LAST TIME SAVED: Jan  2 18:13:57 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_wd_bweb ( bweb, bwebi, sel, wai );


output [15:0]  bweb;

input [3:0]  sel;
input [10:8]  wai;
input [15:0]  bwebi;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  net168;

wire  [3:0]  net0282;

wire  [3:0]  selb;

wire  [10:8]  wa;

wire  [3:0]  net0226;

wire  [10:8]  wa_b;



nand2 I105 ( .A(wa[8]), .Y(nandwa89), .B(wa[9]));
nand2 I2 ( .A(wa_b[8]), .B(wa_b[9]), .Y(nandwa8b9b));
nand2 I104 ( .A(wa_b[8]), .Y(nandwa8b9), .B(wa[9]));
nand2 I103 ( .A(wa[8]), .Y(nandwa89b), .B(wa_b[9]));
nand3 I60 ( .C(wa_b[10]), .A(wa_b[8]), .Y(nandwa8b9b10b), .B(wa_b[9]));
nand3 I98 ( .Y(nandwa8910b), .B(wa[9]), .C(wa_b[10]), .A(wa[8]));
nand3 I97 ( .Y(nandwa8b910b), .B(wa[9]), .C(wa_b[10]), .A(wa_b[8]));
nand3 I96 ( .Y(nandwa89b10b), .B(wa_b[9]), .C(wa_b[10]), .A(wa[8]));
nand3 I99 ( .Y(nandwa8b9b10), .B(wa_b[9]), .C(wa[10]), .A(wa_b[8]));
nand3 I100 ( .Y(nandwa89b10), .B(wa_b[9]), .C(wa[10]), .A(wa[8]));
nand3 I101 ( .Y(nandwa8b910), .B(wa[9]), .C(wa[10]), .A(wa_b[8]));
nand3 I102 ( .Y(nandwa8910), .B(wa[9]), .C(wa[10]), .A(wa[8]));
inv I106 ( .A(wa_b[8]), .Y(wa8));
inv I71 ( .A(wa[8]), .Y(wa8b));
inv I82_2_ ( .A(wai[10]), .Y(net168[0]));
inv I82_1_ ( .A(wai[9]), .Y(net168[1]));
inv I82_0_ ( .A(wai[8]), .Y(net168[2]));
inv I95_2_ ( .A(wai[10]), .Y(wa_b[10]));
inv I95_1_ ( .A(wai[9]), .Y(wa_b[9]));
inv I95_0_ ( .A(wai[8]), .Y(wa_b[8]));
inv I83_2_ ( .A(net168[0]), .Y(wa[10]));
inv I83_1_ ( .A(net168[1]), .Y(wa[9]));
inv I83_0_ ( .A(net168[2]), .Y(wa[8]));
bram_4mux I107 ( bweb[1], bwebi[1], wa8b, nandwa89b, nandwa89b10b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I108 ( bweb[2], bwebi[2], wa8, nandwa8b9, nandwa8b910b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I109 ( bweb[3], bwebi[3], wa8b, nandwa89, nandwa8910b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I110 ( bweb[4], bwebi[4], wa8, nandwa8b9b, nandwa8b9b10,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I111 ( bweb[5], bwebi[5], wa8b, nandwa89b, nandwa89b10,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I112 ( bweb[6], bwebi[6], wa8, nandwa8b9, nandwa8b910,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I113 ( bweb[7], bwebi[7], wa8b, nandwa89, nandwa8910,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I114 ( bweb[8], bwebi[8], wa8, nandwa8b9b, nandwa8b9b10b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I115 ( bweb[9], bwebi[9], wa8b, nandwa89b, nandwa89b10b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I116 ( bweb[10], bwebi[10], wa8, nandwa8b9, nandwa8b910b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I117 ( bweb[11], bwebi[11], wa8b, nandwa89, nandwa8910b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I118 ( bweb[12], bwebi[12], wa8, nandwa8b9b, nandwa8b9b10,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I119 ( bweb[13], bwebi[13], wa8b, nandwa89b, nandwa89b10,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I120 ( bweb[14], bwebi[14], wa8, nandwa8b9, nandwa8b910,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I121 ( bweb[15], bwebi[15], wa8b, nandwa89, nandwa8910,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
bram_4mux I40 ( bweb[0], bwebi[0], wa8, nandwa8b9b, nandwa8b9b10b,
     {net0226[0], net0226[1], net0226[2], net0226[3]}, selb[3:0]);
inv_hvt I122_3_ ( .A(net0282[0]), .Y(net0226[0]));
inv_hvt I122_2_ ( .A(net0282[1]), .Y(net0226[1]));
inv_hvt I122_1_ ( .A(net0282[2]), .Y(net0226[2]));
inv_hvt I122_0_ ( .A(net0282[3]), .Y(net0226[3]));
inv_hvt I123_3_ ( .A(sel[3]), .Y(net0282[0]));
inv_hvt I123_2_ ( .A(sel[2]), .Y(net0282[1]));
inv_hvt I123_1_ ( .A(sel[1]), .Y(net0282[2]));
inv_hvt I123_0_ ( .A(sel[0]), .Y(net0282[3]));
inv_hvt I125_3_ ( .A(sel[3]), .Y(selb[3]));
inv_hvt I125_2_ ( .A(sel[2]), .Y(selb[2]));
inv_hvt I125_1_ ( .A(sel[1]), .Y(selb[1]));
inv_hvt I125_0_ ( .A(sel[0]), .Y(selb[0]));

endmodule
// Library - leafcell, Cell - bram_bufferx6, View - schematic
// LAST TIME SAVED: Jan  2 18:54:54 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_bufferx6 ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - bram_4k_buffer, View - schematic
// LAST TIME SAVED: Sep 30 18:29:20 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_4k_buffer ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;

input [7:0]  bm_sa_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I14 ( .in(bm_sdo_i), .out(bm_sdo_o));
bram_bufferx6 I6 ( .in(bm_sdi_i), .out(bm_sdi_o));
bram_bufferx6 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx6 I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx6 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx6 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx6 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx6 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx6 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx6 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx6 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx6 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx6 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx6 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx6 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx6 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx6 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbank_pbuffer_v1, View -
//schematic
// LAST TIME SAVED: Jan  2 18:54:22 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_v1 ( bm_aa_2bot, bm_ab_2bot, bm_init_o,
     bm_q, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bm_aa,
     bm_aa_top, bm_ab, bm_ab_top, bm_bweb, bm_clkr, bm_clkw, bm_d,
     bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen, cbit, prog );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen, prog;

output [10:0]  bm_aa_2bot;
output [1:0]  bm_sclkrw_o;
output [10:0]  bm_ab_2bot;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [10:0]  bm_aa_top;
input [10:0]  bm_ab_top;
input [1:0]  bm_sweb_i;
input [1:0]  bm_sdo_i;
input [10:0]  bm_aa;
input [1:0]  bm_sdi_i;
input [10:0]  bm_ab;
input [7:0]  bm_sa_i;
input [8:0]  cbit;
input [1:0]  bm_sclkrw_i;
input [15:0]  bm_d;
input [15:0]  bm_bweb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  net231;

wire  [2:0]  net200;

wire  [2:0]  net232;

wire  [15:0]  net236;

wire  [15:0]  bm_q_fromip;

wire  [8:0]  cbitb;

wire  [10:0]  bm_ab_2ip;

wire  [1:0]  cbitd;

wire  [10:0]  bm_aa_2ip;

wire  [15:0]  bm_d_2ip;

wire  [3:0]  sel;



inv_hvt I41 ( .A(net178), .Y(sel[2]));
inv_hvt I55_1_ ( .A(cbitb[1]), .Y(cbitd[1]));
inv_hvt I55_0_ ( .A(cbitb[0]), .Y(cbitd[0]));
inv_hvt I43 ( .A(cbit[8]), .Y(cbitb[8]));
inv_hvt I54_1_ ( .A(cbit[1]), .Y(cbitb[1]));
inv_hvt I54_0_ ( .A(cbit[0]), .Y(cbitb[0]));
inv_hvt I56 ( .A(net172), .Y(sel[0]));
inv_hvt I42 ( .A(net175), .Y(sel[3]));
inv_hvt I40 ( .A(net181), .Y(sel[1]));
bram_cascade_addr I_cascade_addr4ra ( .prog(prog),
     .addr_2bot(bm_ab_2bot[10:0]), .cbit(cbit[7:6]),
     .addr_top(bm_ab_top[10:0]), .addr(bm_ab[10:0]),
     .addr_muxo(bm_ab_2ip[10:0]));
bram_cascade_addr I_cascade_addr4wa ( .prog(prog),
     .addr_2bot(bm_aa_2bot[10:0]), .cbit(cbit[5:4]),
     .addr_top(bm_aa_top[10:0]), .addr(bm_aa[10:0]),
     .addr_muxo(bm_aa_2ip[10:0]));
bram_4k_n40 I_bram_4k ( .bm_pd(cbitb[8]), .bm_ab(bm_ab_2ip[7:0]),
     .bm_aa(bm_aa_2ip[7:0]), .bm_q(bm_q_fromip[15:0]),
     .bm_sclk(bm_sclk_o), .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb({net236[0], net236[1],
     net236[2], net236[3], net236[4], net236[5], net236[6], net236[7],
     net236[8], net236[9], net236[10], net236[11], net236[12],
     net236[13], net236[14], net236[15]}), .bm_ren(bm_ren),
     .bm_wen(bm_wen), .bm_clkr(bm_clkr), .bm_sweb(bm_sweb_o[0]),
     .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d_2ip[15:0]), .bm_clkw(bm_clkw),
     .bm_sdo(net246));
bram_rd_decoder0to7 I_bram_rd_decoder8to15 ( .rd(bm_q[15:8]),
     .rdi(bm_q_fromip[15:8]), .c(cbit[3:2]), .raq({net200[0],
     net200[1], net200[2]}));
bram_rd_decoder0to7 I_bram_rd_decoder0to7 ( .c(cbit[3:2]),
     .rd(bm_q[7:0]), .raq({net200[0], net200[1], net200[2]}),
     .rdi(bm_q_fromip[7:0]));
bram_wd_decoder0to7 I_bram_wd_decoder8to15 ( .wd(bm_d_2ip[15:8]),
     .wdi(bm_d[15:8]), .sel(sel[3:0]));
bram_wd_decoder0to7 I_bram_wd_decoder0to7 ( .wd(bm_d_2ip[7:0]),
     .sel(sel[3:0]), .wdi(bm_d[7:0]));
nand2_hvt I92 ( .A(cbitb[0]), .Y(net172), .B(cbitb[1]));
nand2_hvt I39 ( .A(cbitd[0]), .Y(net175), .B(cbitd[1]));
nand2_hvt I38 ( .A(cbitb[0]), .Y(net178), .B(cbitd[1]));
nand2_hvt I37 ( .A(cbitd[0]), .Y(net181), .B(cbitb[1]));
inv I46_2_ ( .A(net231[0]), .Y(net200[0]));
inv I46_1_ ( .A(net231[1]), .Y(net200[1]));
inv I46_0_ ( .A(net231[2]), .Y(net200[2]));
ml_dff I_RAQ_2_ ( .R(prog), .D(bm_ab_2ip[10]), .CLK(bm_clkr),
     .QN(net231[0]), .Q(net232[0]));
ml_dff I_RAQ_1_ ( .R(prog), .D(bm_ab_2ip[9]), .CLK(bm_clkr),
     .QN(net231[1]), .Q(net232[1]));
ml_dff I_RAQ_0_ ( .R(prog), .D(bm_ab_2ip[8]), .CLK(bm_clkr),
     .QN(net231[2]), .Q(net232[2]));
bram_wd_bweb I_bram_wd_bweb ( .sel(sel[3:0]), .wai(bm_aa_2ip[10:8]),
     .bwebi(bm_bweb[15:0]), .bweb({net236[0], net236[1], net236[2],
     net236[3], net236[4], net236[5], net236[6], net236[7], net236[8],
     net236[9], net236[10], net236[11], net236[12], net236[13],
     net236[14], net236[15]}));
bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k_buffer I_bram_4k_buffer ( .bm_sdo_o(bm_sdo_o[0]),
     .bm_sdo_i(net246), .bm_sclkrw_i(bm_sclkrw_i[0]),
     .bm_sclkrw_o(bm_sclkrw_o[0]), .bm_sdi_o(bm_sdi_o[0]),
     .bm_sdi_i(bm_sdi_i[0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - ice1chip, Cell - bram_4kprouting_ice1p, View - schematic
// LAST TIME SAVED: Apr 20 10:01:28 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram_4kprouting_ice1p ( bm_aa_2bot, bm_ab_2bot, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, cntl_cbit_bot,
     cntl_cbit_top, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_aa_top, bm_ab_top, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_bot,
     bnr_op_bot, bot_op_bot, glb_netwk, lft_op_bot, lft_op_top,
     pgate_bot, pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot,
     rgt_op_top, tnl_op_top, tnr_op_top, top_op_top, vdd_cntl_bot,
     vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sclkrw_o;
output [10:0]  bm_ab_2bot;
output [7:0]  cntl_cbit_top;
output [10:0]  bm_aa_2bot;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;
output [1:0]  bm_sweb_o;
output [7:0]  cntl_cbit_bot;

inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_h_l_top;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_h_l_top;
inout [41:0]  bl;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_h_l_bot;

input [7:0]  rgt_op_bot;
input [1:0]  bm_sweb_i;
input [15:0]  wl_bot;
input [10:0]  bm_ab_top;
input [7:0]  lft_op_bot;
input [7:0]  top_op_top;
input [15:0]  pgate_top;
input [1:0]  bm_sclkrw_i;
input [15:0]  pgate_bot;
input [7:0]  bm_sa_i;
input [1:0]  bm_sdo_i;
input [10:0]  bm_aa_top;
input [7:0]  tnl_op_top;
input [7:0]  bnr_op_bot;
input [7:0]  bnl_op_bot;
input [15:0]  wl_top;
input [15:0]  vdd_cntl_top;
input [7:0]  glb_netwk;
input [7:0]  bot_op_bot;
input [7:0]  tnr_op_top;
input [7:0]  lft_op_top;
input [15:0]  vdd_cntl_bot;
input [15:0]  reset_b_bot;
input [1:0]  bm_sdi_i;
input [7:0]  rgt_op_top;
input [15:0]  reset_b_top;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  bm_bweb;

wire  [10:0]  bram_ab;

wire  [10:0]  bram_aa;

wire  [15:0]  bm_d;

wire  [7:0]  bram_cbit_top;

wire  [7:0]  bram_cbit_bot;



bram_4kprouting_left_ice1p I22 ( .slf_op_top(slf_op_top[7:0]),
     .slf_op_bot(slf_op_bot[7:0]), .wl_bot(wl_bot[15:0]),
     .top_op_top(top_op_top[7:0]), .sp12_h_l_bot(sp12_h_l_bot[23:0]),
     .sp4_h_l_bot(sp4_h_l_bot[47:0]), .tnl_op_top(tnl_op_top[7:0]),
     .reset_b_top(reset_b_top[15:0]), .reset_b_bot(reset_b_bot[15:0]),
     .vdd_cntl_top(vdd_cntl_top[15:0]), .prog(prog),
     .pgate_top(pgate_top[15:0]), .pgate_bot(pgate_bot[15:0]),
     .lft_op_bot(lft_op_bot[7:0]), .bot_op_bot(bot_op_bot[7:0]),
     .rgt_op_bot(rgt_op_bot[7:0]), .bnl_op_bot(bnl_op_bot[7:0]),
     .sp4_h_r_top(sp4_h_r_top[47:0]),
     .sp12_v_t_top(sp12_v_t_top[23:0]),
     .sp12_v_b_bot(sp12_v_b_bot[23:0]),
     .sp4_h_r_bot(sp4_h_r_bot[47:0]),
     .sp12_h_r_bot(sp12_h_r_bot[23:0]),
     .sp4_v_t_top(sp4_v_t_top[47:0]), .sp4_v_b_bot(sp4_v_b_bot[47:0]),
     .sp12_h_r_top(sp12_h_r_top[23:0]), .bl(bl[41:0]),
     .sp4_h_l_top(sp4_h_l_top[47:0]), .lft_op_top(lft_op_top[7:0]),
     .wl_top(wl_top[15:0]), .sp12_h_l_top(sp12_h_l_top[23:0]),
     .sp4_v_b_top(sp4_v_b_top[47:0]), .rgt_op_top(rgt_op_top[7:0]),
     .vdd_cntl_bot(vdd_cntl_bot[15:0]), .bnr_op_bot(bnr_op_bot[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_bot[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_top[47:0]),
     .cntl_cbit_bot(cntl_cbit_bot[7:0]),
     .cntl_cbit_top(cntl_cbit_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bram_ab(bram_ab[10:0]), .bram_aa(bram_aa[10:0]),
     .bm_bweb(bm_bweb[15:0]), .bm_clkr2rf_n40(bm_clkr2rf_n40),
     .bm_clkw2rf_n40(bm_clkw2rf_n40), .bm_d(bm_d[15:0]),
     .bm_ren2rf_n40(bm_ren2rf_n40), .bm_wen2rf_n40(bm_wen2rf_n40),
     .bram_cbit_top(bram_cbit_top[7:0]),
     .bram_cbit_bot(bram_cbit_bot[7:0]), .tnr_op_top(tnr_op_top[7:0]));
bram_4kbank_pbuffer_v1 I_bram_4kbank_pbuffer ( .cbit({bram_cbit_bot[0],
     bram_cbit_top[7:0]}), .bm_aa(bram_aa[10:0]), .prog(prog),
     .bm_ab(bram_ab[10:0]), .bm_aa_2bot(bm_aa_2bot[10:0]),
     .bm_ab_2bot(bm_ab_2bot[10:0]), .bm_aa_top(bm_aa_top[10:0]),
     .bm_ab_top(bm_ab_top[10:0]), .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(bm_ren2rf_n40),
     .bm_wen(bm_wen2rf_n40), .bm_d(bm_d[15:0]),
     .bm_clkr(bm_clkr2rf_n40), .bm_clkw(bm_clkw2rf_n40),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));

endmodule
// Library - leafcell, Cell - clk_colbuf12k, View - schematic
// LAST TIME SAVED: Aug 20 07:53:18 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module clk_colbuf12k ( clko, cbit, clki );
output  clko;

input  cbit, clki;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_lvt I_nand2_lvt ( .A(clki), .Y(clkb), .B(cbit));
nch_lvt  M1 ( .D(clko), .B(gnd_), .G(clkb), .S(net7));
nch_lvt  M2 ( .D(net7), .B(gnd_), .G(cbit), .S(gnd_));
pch_lvt  M0 ( .D(clko), .B(vdd_), .G(clkb), .S(vdd_));

endmodule
// Library - ice8chip, Cell - clk_col_buf_x8_ice8p, View - schematic
// LAST TIME SAVED: Jan  6 15:52:04 2009
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module clk_col_buf_x8_ice8p ( col_clk, clk_in, colbuf_cntl );


output [7:0]  col_clk;

input [7:0]  colbuf_cntl;
input [7:0]  clk_in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



clk_colbuf12k I_colbuf12k_7_ ( .clki(clk_in[7]), .clko(col_clk[7]),
     .cbit(colbuf_cntl[7]));
clk_colbuf12k I_colbuf12k_6_ ( .clki(clk_in[6]), .clko(col_clk[6]),
     .cbit(colbuf_cntl[6]));
clk_colbuf12k I_colbuf12k_5_ ( .clki(clk_in[5]), .clko(col_clk[5]),
     .cbit(colbuf_cntl[5]));
clk_colbuf12k I_colbuf12k_4_ ( .clki(clk_in[4]), .clko(col_clk[4]),
     .cbit(colbuf_cntl[4]));
clk_colbuf12k I_colbuf12k_3_ ( .clki(clk_in[3]), .clko(col_clk[3]),
     .cbit(colbuf_cntl[3]));
clk_colbuf12k I_colbuf12k_2_ ( .clki(clk_in[2]), .clko(col_clk[2]),
     .cbit(colbuf_cntl[2]));
clk_colbuf12k I_colbuf12k_1_ ( .clki(clk_in[1]), .clko(col_clk[1]),
     .cbit(colbuf_cntl[1]));
clk_colbuf12k I_colbuf12k_0_ ( .clki(clk_in[0]), .clko(col_clk[0]),
     .cbit(colbuf_cntl[0]));

endmodule
// Library - ice1chip, Cell - bram1x4_ice1f, View - schematic
// LAST TIME SAVED: Apr 20 09:56:03 2011
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module bram1x4_ice1f ( bm_aa_2bot, bm_ab_2bot, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, glb_netwk_bot,
     glb_netwk_top, slf_op_01, slf_op_02, slf_op_03, slf_op_04,
     slf_op_05, slf_op_06, slf_op_07, slf_op_08, bl, pgate, reset_b,
     sp4_h_l_01, sp4_h_l_02, sp4_h_l_03, sp4_h_l_04, sp4_h_l_05,
     sp4_h_l_06, sp4_h_l_07, sp4_h_l_08, sp4_h_r_01, sp4_h_r_02,
     sp4_h_r_03, sp4_h_r_04, sp4_h_r_05, sp4_h_r_06, sp4_h_r_07,
     sp4_h_r_08, sp4_r_v_b_01, sp4_r_v_b_02, sp4_r_v_b_03,
     sp4_r_v_b_04, sp4_r_v_b_05, sp4_r_v_b_06, sp4_r_v_b_07,
     sp4_r_v_b_08, sp4_v_b_01, sp4_v_b_02, sp4_v_b_03, sp4_v_b_04,
     sp4_v_b_05, sp4_v_b_06, sp4_v_b_07, sp4_v_b_08, sp4_v_t_08,
     sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04, sp12_h_l_05,
     sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_r_01, sp12_h_r_02,
     sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06, sp12_h_r_07,
     sp12_h_r_08, sp12_v_b_01, sp12_v_t_08, vdd_cntl, wl, bm_aa_top,
     bm_ab_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_01, bnr_op_01, bot_op_01, glb_netwk_col,
     lft_op_01, lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06,
     lft_op_07, lft_op_08, prog, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, tnl_op_08,
     tnr_op_08, top_op_08 );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sweb_o;
output [10:0]  bm_aa_2bot;
output [7:0]  slf_op_08;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_05;
output [7:0]  slf_op_04;
output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [10:0]  bm_ab_2bot;
output [7:0]  slf_op_02;
output [7:0]  slf_op_07;
output [7:0]  glb_netwk_bot;
output [7:0]  slf_op_03;
output [7:0]  slf_op_01;
output [7:0]  slf_op_06;
output [7:0]  glb_netwk_top;

inout [23:0]  sp12_v_t_08;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_v_b_03;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_h_l_05;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_v_b_01;
inout [23:0]  sp12_h_l_02;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_h_l_04;
inout [47:0]  sp4_r_v_b_06;
inout [23:0]  sp12_h_l_03;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_08;
inout [23:0]  sp12_v_b_01;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_h_r_05;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_h_r_08;
inout [47:0]  sp4_h_l_08;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_h_l_03;
inout [47:0]  sp4_v_b_05;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_v_b_07;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_h_l_02;
inout [47:0]  sp4_v_t_08;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_h_l_06;
inout [23:0]  sp12_h_r_01;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_v_b_06;
inout [47:0]  sp4_r_v_b_07;
inout [23:0]  sp12_h_l_06;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_h_r_07;
inout [143:16]  pgate;
inout [47:0]  sp4_r_v_b_05;
inout [143:16]  reset_b;
inout [47:0]  sp4_h_l_01;
inout [47:0]  sp4_r_v_b_08;
inout [143:16]  vdd_cntl;
inout [47:0]  sp4_r_v_b_02;
inout [143:16]  wl;
inout [47:0]  sp4_h_r_01;

input [1:0]  bm_sclkrw_i;
input [10:0]  bm_ab_top;
input [7:0]  bnr_op_01;
input [7:0]  rgt_op_04;
input [7:0]  rgt_op_08;
input [7:0]  lft_op_08;
input [7:0]  lft_op_01;
input [7:0]  bnl_op_01;
input [7:0]  lft_op_03;
input [1:0]  bm_sdi_i;
input [7:0]  lft_op_06;
input [7:0]  lft_op_05;
input [10:0]  bm_aa_top;
input [7:0]  lft_op_02;
input [1:0]  bm_sdo_i;
input [7:0]  rgt_op_02;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_07;
input [7:0]  tnr_op_08;
input [7:0]  top_op_08;
input [7:0]  bm_sa_i;
input [7:0]  lft_op_07;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_01;
input [7:0]  glb_netwk_col;
input [7:0]  tnl_op_08;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_04;
input [7:0]  bot_op_01;
input [1:0]  bm_sweb_i;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  net1120;

wire  [1:0]  net933;

wire  [23:0]  net1023;

wire  [10:0]  net0806;

wire  [10:0]  net0875;

wire  [1:0]  net993;

wire  [1:0]  net929;

wire  [1:0]  net999;

wire  [1:0]  net994;

wire  [1:0]  net935;

wire  [7:0]  net863;

wire  [1:0]  net1121;

wire  [1:0]  net1125;

wire  [1:0]  net1127;

wire  [10:0]  net01011;

wire  [7:0]  colbuf_cntl_top;

wire  [7:0]  net1049;

wire  [1:0]  net1122;

wire  [10:0]  net0807;

wire  [7:0]  net0666;

wire  [10:0]  net01010;

wire  [1:0]  net997;

wire  [7:0]  net1177;

wire  [23:0]  net959;

wire  [7:0]  net985;

wire  [7:0]  net991;

wire  [1:0]  net930;

wire  [10:0]  net0874;

wire  [7:0]  net928;

wire  [23:0]  net1151;

wire  [7:0]  net1119;

wire  [7:0]  colbuf_cntl_bot;



bram_4kprouting_ice1p I_bram_0825_08 ( .cntl_cbit_top({net0666[0],
     net0666[1], net0666[2], net0666[3], net0666[4], net0666[5],
     net0666[6], net0666[7]}), .cntl_cbit_bot({net863[0], net863[1],
     net863[2], net863[3], net863[4], net863[5], net863[6],
     net863[7]}), .bm_aa_2bot({net0806[0], net0806[1], net0806[2],
     net0806[3], net0806[4], net0806[5], net0806[6], net0806[7],
     net0806[8], net0806[9], net0806[10]}), .bm_ab_2bot({net0807[0],
     net0807[1], net0807[2], net0807[3], net0807[4], net0807[5],
     net0807[6], net0807[7], net0807[8], net0807[9], net0807[10]}),
     .bm_aa_top(bm_aa_top[10:0]), .bm_ab_top(bm_ab_top[10:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sclkrw_i({net930[0], net930[1]}), .bm_sweb_i({net933[0],
     net933[1]}), .bm_sweb_o(bm_sweb_o[1:0]), .bm_sdi_i({net929[0],
     net929[1]}), .bm_sdo_i(bm_sdo_i[1:0]), .bm_sdo_o({net935[0],
     net935[1]}), .slf_op_top(slf_op_08[7:0]),
     .slf_op_bot(slf_op_07[7:0]), .wl_bot(wl[127:112]),
     .top_op_top(top_op_08[7:0]), .sp12_h_l_bot(sp12_h_l_07[23:0]),
     .sp4_h_l_bot(sp4_h_l_07[47:0]), .tnl_op_top(tnl_op_08[7:0]),
     .reset_b_top(reset_b[143:128]), .reset_b_bot(reset_b[127:112]),
     .vdd_cntl_top(vdd_cntl[143:128]), .prog(prog),
     .pgate_top(pgate[143:128]), .pgate_bot(pgate[127:112]),
     .lft_op_bot(lft_op_07[7:0]), .glb_netwk(glb_netwk_top[7:0]),
     .bm_wdummymux_en_i(net988), .bot_op_bot(slf_op_06[7:0]),
     .rgt_op_bot(rgt_op_07[7:0]), .bnl_op_bot(lft_op_06[7:0]),
     .sp4_h_r_top(sp4_h_r_08[47:0]), .sp12_v_t_top(sp12_v_t_08[23:0]),
     .sp12_v_b_bot({net959[0], net959[1], net959[2], net959[3],
     net959[4], net959[5], net959[6], net959[7], net959[8], net959[9],
     net959[10], net959[11], net959[12], net959[13], net959[14],
     net959[15], net959[16], net959[17], net959[18], net959[19],
     net959[20], net959[21], net959[22], net959[23]}),
     .bm_init_i(net984), .sp4_h_r_bot(sp4_h_r_07[47:0]),
     .sp12_h_r_bot(sp12_h_r_07[23:0]), .sp4_v_t_top(sp4_v_t_08[47:0]),
     .sp4_v_b_bot(sp4_v_b_07[47:0]), .sp12_h_r_top(sp12_h_r_08[23:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net983),
     .sp4_h_l_top(sp4_h_l_08[47:0]), .lft_op_top(lft_op_08[7:0]),
     .wl_top(wl[143:128]), .sp12_h_l_top(sp12_h_l_08[23:0]),
     .sp4_v_b_top(sp4_v_b_08[47:0]), .tnr_op_top(tnr_op_08[7:0]),
     .rgt_op_top(rgt_op_08[7:0]), .bm_sa_i({net985[0], net985[1],
     net985[2], net985[3], net985[4], net985[5], net985[6],
     net985[7]}), .bm_sclk_i(net986), .bm_sreb_i(net987),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .vdd_cntl_bot(vdd_cntl[127:112]), .bnr_op_bot(rgt_op_06[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_07[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_08[47:0]));
bram_4kprouting_ice1p I_bram_0825_06 ( .cntl_cbit_top({net928[0],
     net928[1], net928[2], net928[3], net928[4], net928[5], net928[6],
     net928[7]}), .cntl_cbit_bot(colbuf_cntl_top[7:0]),
     .bm_aa_2bot({net0874[0], net0874[1], net0874[2], net0874[3],
     net0874[4], net0874[5], net0874[6], net0874[7], net0874[8],
     net0874[9], net0874[10]}), .bm_ab_2bot({net0875[0], net0875[1],
     net0875[2], net0875[3], net0875[4], net0875[5], net0875[6],
     net0875[7], net0875[8], net0875[9], net0875[10]}),
     .bm_aa_top({net0806[0], net0806[1], net0806[2], net0806[3],
     net0806[4], net0806[5], net0806[6], net0806[7], net0806[8],
     net0806[9], net0806[10]}), .bm_ab_top({net0807[0], net0807[1],
     net0807[2], net0807[3], net0807[4], net0807[5], net0807[6],
     net0807[7], net0807[8], net0807[9], net0807[10]}),
     .bm_sdi_o({net929[0], net929[1]}), .bm_sclkrw_o({net930[0],
     net930[1]}), .bm_sclkrw_i({net994[0], net994[1]}),
     .bm_sweb_i({net997[0], net997[1]}), .bm_sweb_o({net933[0],
     net933[1]}), .bm_sdi_i({net993[0], net993[1]}),
     .bm_sdo_i({net935[0], net935[1]}), .bm_sdo_o({net999[0],
     net999[1]}), .slf_op_top(slf_op_06[7:0]),
     .slf_op_bot(slf_op_05[7:0]), .wl_top(wl[111:96]),
     .wl_bot(wl[95:80]), .top_op_top(slf_op_07[7:0]),
     .tnl_op_top(lft_op_07[7:0]), .reset_b_top(reset_b[111:96]),
     .reset_b_bot(reset_b[95:80]), .prog(prog),
     .pgate_top(pgate[111:96]), .pgate_bot(pgate[95:80]),
     .lft_op_top(lft_op_06[7:0]), .lft_op_bot(lft_op_05[7:0]),
     .glb_netwk(glb_netwk_top[7:0]), .bm_wdummymux_en_i(net1052),
     .bot_op_bot(slf_op_04[7:0]), .sp4_h_r_top(sp4_h_r_06[47:0]),
     .bnl_op_bot(lft_op_04[7:0]), .bnr_op_bot(rgt_op_04[7:0]),
     .sp4_h_r_bot(sp4_h_r_05[47:0]), .sp12_v_t_top({net959[0],
     net959[1], net959[2], net959[3], net959[4], net959[5], net959[6],
     net959[7], net959[8], net959[9], net959[10], net959[11],
     net959[12], net959[13], net959[14], net959[15], net959[16],
     net959[17], net959[18], net959[19], net959[20], net959[21],
     net959[22], net959[23]}), .sp12_v_b_bot({net1023[0], net1023[1],
     net1023[2], net1023[3], net1023[4], net1023[5], net1023[6],
     net1023[7], net1023[8], net1023[9], net1023[10], net1023[11],
     net1023[12], net1023[13], net1023[14], net1023[15], net1023[16],
     net1023[17], net1023[18], net1023[19], net1023[20], net1023[21],
     net1023[22], net1023[23]}), .bm_init_i(net1048),
     .sp12_h_l_top(sp12_h_l_06[23:0]),
     .sp12_h_r_bot(sp12_h_r_05[23:0]),
     .sp12_h_l_bot(sp12_h_l_05[23:0]),
     .sp12_h_r_top(sp12_h_r_06[23:0]), .sp4_v_t_top(sp4_v_b_07[47:0]),
     .sp4_v_b_top(sp4_v_b_06[47:0]), .sp4_v_b_bot(sp4_v_b_05[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_05[47:0]),
     .sp4_h_l_top(sp4_h_l_06[47:0]), .tnr_op_top(rgt_op_07[7:0]),
     .sp4_h_l_bot(sp4_h_l_05[47:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net1047), .sp4_r_v_b_top(sp4_r_v_b_06[47:0]),
     .rgt_op_bot(rgt_op_05[7:0]), .rgt_op_top(rgt_op_06[7:0]),
     .bm_sa_i({net1049[0], net1049[1], net1049[2], net1049[3],
     net1049[4], net1049[5], net1049[6], net1049[7]}),
     .bm_sclk_i(net1050), .bm_sreb_i(net1051),
     .bm_rcapmux_en_o(net983), .bm_init_o(net984), .bm_sa_o({net985[0],
     net985[1], net985[2], net985[3], net985[4], net985[5], net985[6],
     net985[7]}), .bm_sclk_o(net986), .bm_sreb_o(net987),
     .bm_wdummymux_en_o(net988), .vdd_cntl_top(vdd_cntl[111:96]),
     .vdd_cntl_bot(vdd_cntl[95:80]));
bram_4kprouting_ice1p I_bram_0825_04 (
     .cntl_cbit_top(colbuf_cntl_bot[7:0]), .cntl_cbit_bot({net991[0],
     net991[1], net991[2], net991[3], net991[4], net991[5], net991[6],
     net991[7]}), .bm_aa_2bot({net01010[0], net01010[1], net01010[2],
     net01010[3], net01010[4], net01010[5], net01010[6], net01010[7],
     net01010[8], net01010[9], net01010[10]}),
     .bm_ab_2bot({net01011[0], net01011[1], net01011[2], net01011[3],
     net01011[4], net01011[5], net01011[6], net01011[7], net01011[8],
     net01011[9], net01011[10]}), .bm_aa_top({net0874[0], net0874[1],
     net0874[2], net0874[3], net0874[4], net0874[5], net0874[6],
     net0874[7], net0874[8], net0874[9], net0874[10]}),
     .bm_ab_top({net0875[0], net0875[1], net0875[2], net0875[3],
     net0875[4], net0875[5], net0875[6], net0875[7], net0875[8],
     net0875[9], net0875[10]}), .bm_sdi_o({net993[0], net993[1]}),
     .bm_sclkrw_o({net994[0], net994[1]}), .bm_sclkrw_i({net1122[0],
     net1122[1]}), .bm_sweb_i({net1125[0], net1125[1]}),
     .bm_sweb_o({net997[0], net997[1]}), .bm_sdi_i({net1121[0],
     net1121[1]}), .bm_sdo_i({net999[0], net999[1]}),
     .bm_sdo_o({net1127[0], net1127[1]}), .slf_op_top(slf_op_04[7:0]),
     .slf_op_bot(slf_op_03[7:0]), .wl_top(wl[79:64]),
     .wl_bot(wl[63:48]), .top_op_top(slf_op_05[7:0]),
     .tnl_op_top(lft_op_05[7:0]), .reset_b_top(reset_b[79:64]),
     .reset_b_bot(reset_b[63:48]), .prog(prog),
     .pgate_top(pgate[79:64]), .pgate_bot(pgate[63:48]),
     .lft_op_top(lft_op_04[7:0]), .lft_op_bot(lft_op_03[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]), .bm_wdummymux_en_i(net1180),
     .bot_op_bot(slf_op_02[7:0]), .sp4_h_r_top(sp4_h_r_04[47:0]),
     .bnl_op_bot(lft_op_02[7:0]), .bnr_op_bot(rgt_op_02[7:0]),
     .sp4_h_r_bot(sp4_h_r_03[47:0]), .sp12_v_t_top({net1023[0],
     net1023[1], net1023[2], net1023[3], net1023[4], net1023[5],
     net1023[6], net1023[7], net1023[8], net1023[9], net1023[10],
     net1023[11], net1023[12], net1023[13], net1023[14], net1023[15],
     net1023[16], net1023[17], net1023[18], net1023[19], net1023[20],
     net1023[21], net1023[22], net1023[23]}),
     .sp12_v_b_bot({net1151[0], net1151[1], net1151[2], net1151[3],
     net1151[4], net1151[5], net1151[6], net1151[7], net1151[8],
     net1151[9], net1151[10], net1151[11], net1151[12], net1151[13],
     net1151[14], net1151[15], net1151[16], net1151[17], net1151[18],
     net1151[19], net1151[20], net1151[21], net1151[22], net1151[23]}),
     .bm_init_i(net1176), .sp12_h_l_top(sp12_h_l_04[23:0]),
     .sp12_h_r_bot(sp12_h_r_03[23:0]),
     .sp12_h_l_bot(sp12_h_l_03[23:0]),
     .sp12_h_r_top(sp12_h_r_04[23:0]), .sp4_v_t_top(sp4_v_b_05[47:0]),
     .sp4_v_b_top(sp4_v_b_04[47:0]), .sp4_v_b_bot(sp4_v_b_03[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_03[47:0]),
     .sp4_h_l_top(sp4_h_l_04[47:0]), .tnr_op_top(rgt_op_05[7:0]),
     .sp4_h_l_bot(sp4_h_l_03[47:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net1175), .sp4_r_v_b_top(sp4_r_v_b_04[47:0]),
     .rgt_op_bot(rgt_op_03[7:0]), .rgt_op_top(rgt_op_04[7:0]),
     .bm_sa_i({net1177[0], net1177[1], net1177[2], net1177[3],
     net1177[4], net1177[5], net1177[6], net1177[7]}),
     .bm_sclk_i(net1178), .bm_sreb_i(net1179),
     .bm_rcapmux_en_o(net1047), .bm_init_o(net1048),
     .bm_sa_o({net1049[0], net1049[1], net1049[2], net1049[3],
     net1049[4], net1049[5], net1049[6], net1049[7]}),
     .bm_sclk_o(net1050), .bm_sreb_o(net1051),
     .bm_wdummymux_en_o(net1052), .vdd_cntl_top(vdd_cntl[79:64]),
     .vdd_cntl_bot(vdd_cntl[63:48]));
bram_4kprouting_ice1p I_bram_0825_02 ( .cntl_cbit_top({net1120[0],
     net1120[1], net1120[2], net1120[3], net1120[4], net1120[5],
     net1120[6], net1120[7]}), .cntl_cbit_bot({net1119[0], net1119[1],
     net1119[2], net1119[3], net1119[4], net1119[5], net1119[6],
     net1119[7]}), .bm_aa_2bot(bm_aa_2bot[10:0]),
     .bm_ab_2bot(bm_ab_2bot[10:0]), .bm_aa_top({net01010[0],
     net01010[1], net01010[2], net01010[3], net01010[4], net01010[5],
     net01010[6], net01010[7], net01010[8], net01010[9],
     net01010[10]}), .bm_ab_top({net01011[0], net01011[1], net01011[2],
     net01011[3], net01011[4], net01011[5], net01011[6], net01011[7],
     net01011[8], net01011[9], net01011[10]}), .bm_sdi_o({net1121[0],
     net1121[1]}), .bm_sclkrw_o({net1122[0], net1122[1]}),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .bm_sweb_i(bm_sweb_i[1:0]),
     .bm_sweb_o({net1125[0], net1125[1]}), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sdo_i({net1127[0], net1127[1]}), .bm_sdo_o(bm_sdo_o[1:0]),
     .slf_op_top(slf_op_02[7:0]), .slf_op_bot(slf_op_01[7:0]),
     .wl_top(wl[47:32]), .wl_bot(wl[31:16]),
     .top_op_top(slf_op_03[7:0]), .tnl_op_top(lft_op_03[7:0]),
     .reset_b_top(reset_b[47:32]), .reset_b_bot(reset_b[31:16]),
     .prog(prog), .pgate_top(pgate[47:32]), .pgate_bot(pgate[31:16]),
     .lft_op_top(lft_op_02[7:0]), .lft_op_bot(lft_op_01[7:0]),
     .glb_netwk(glb_netwk_bot[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_01[7:0]), .sp4_h_r_top(sp4_h_r_02[47:0]),
     .bnl_op_bot(bnl_op_01[7:0]), .bnr_op_bot(bnr_op_01[7:0]),
     .sp4_h_r_bot(sp4_h_r_01[47:0]), .sp12_v_t_top({net1151[0],
     net1151[1], net1151[2], net1151[3], net1151[4], net1151[5],
     net1151[6], net1151[7], net1151[8], net1151[9], net1151[10],
     net1151[11], net1151[12], net1151[13], net1151[14], net1151[15],
     net1151[16], net1151[17], net1151[18], net1151[19], net1151[20],
     net1151[21], net1151[22], net1151[23]}),
     .sp12_v_b_bot(sp12_v_b_01[23:0]), .bm_init_i(bm_init_i),
     .sp12_h_l_top(sp12_h_l_02[23:0]),
     .sp12_h_r_bot(sp12_h_r_01[23:0]),
     .sp12_h_l_bot(sp12_h_l_01[23:0]),
     .sp12_h_r_top(sp12_h_r_02[23:0]), .sp4_v_t_top(sp4_v_b_03[47:0]),
     .sp4_v_b_top(sp4_v_b_02[47:0]), .sp4_v_b_bot(sp4_v_b_01[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_01[47:0]),
     .sp4_h_l_top(sp4_h_l_02[47:0]), .tnr_op_top(rgt_op_03[7:0]),
     .sp4_h_l_bot(sp4_h_l_01[47:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .sp4_r_v_b_top(sp4_r_v_b_02[47:0]), .rgt_op_bot(rgt_op_01[7:0]),
     .rgt_op_top(rgt_op_02[7:0]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(net1175), .bm_init_o(net1176),
     .bm_sa_o({net1177[0], net1177[1], net1177[2], net1177[3],
     net1177[4], net1177[5], net1177[6], net1177[7]}),
     .bm_sclk_o(net1178), .bm_sreb_o(net1179),
     .bm_wdummymux_en_o(net1180), .vdd_cntl_top(vdd_cntl[47:32]),
     .vdd_cntl_bot(vdd_cntl[31:16]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_top (
     .colbuf_cntl(colbuf_cntl_top[7:0]), .col_clk(glb_netwk_top[7:0]),
     .clk_in(glb_netwk_col[7:0]));
clk_col_buf_x8_ice8p I_clk_col_buf_x8_ice8p_bot (
     .colbuf_cntl(colbuf_cntl_bot[7:0]), .col_clk(glb_netwk_bot[7:0]),
     .clk_in(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - delay150ps, View - schematic
// LAST TIME SAVED: Dec 21 17:50:49 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module delay150ps ( out, in );
output  out;

input  in;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



inv_hvt I4 ( .A(in), .Y(net12));
inv_hvt I0 ( .A(net013), .Y(out));
inv_hvt I6 ( .A(net12), .Y(net17));
inv_hvt I2 ( .A(net17), .Y(net013));

endmodule
// Library - io, Cell - ioin_mux_v3, View - schematic
// LAST TIME SAVED: Dec  7 10:44:24 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioin_mux_v3 ( inmuxo, cbit,
     cbitb, min[7:0], prog );
output  inmuxo;

input  prog;

input [3:0]  cbitb;
input [3:0]  cbit;
input [7:0]  min;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_lvt I282 ( .A(prog), .Y(en), .B(cbitb[3]));
inv_lvt I281 ( .A(inmuxob), .Y(inmuxo));
nand2_lvt I_nand2 ( .A(st2), .Y(inmuxob), .B(en));
txgate_lvt I285 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I289 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I286 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I283 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_lvt I292 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I293 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I291 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I294 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I287 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I290 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I288 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I295 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I284 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc_v0, View - schematic
// LAST TIME SAVED: Dec  7 10:49:57 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc_v0 ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  spi;
output [1:0]  ti;

inout [5:0]  bl;

input [7:0]  min2;
input [7:0]  min1;
input [1:0]  vdd_cntl;
input [7:0]  min0;
input [1:0]  reset;
input [1:0]  padin;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



ioin_mux_v3 I_ioin_mux_bankcntl ( bankcntl, {cbit[11], cbit[8], cbit[9],
     cbit[10]}, {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0],
     prog);
ioin_mux_v3 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v3 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
inv_lvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_lvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
nor2_lvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_lvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioinmx2nand2inv_v0, View - schematic
// LAST TIME SAVED: Dec  7 10:48:43 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioinmx2nand2inv_v0 ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  reset;
input [7:0]  min0;
input [7:0]  min1;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [7:0]  ce;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;

wire  [11:0]  cbit;



ioin_mux_v3 I_ioin_mux0 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux_v3 I_ioin_mux1 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]},
     {cbitb[5], cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);
nand2_lvt I180 ( .A(update_b), .Y(updt), .B(bs_en));
inv_lvt I181 ( .A(update), .Y(update_b));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioin_mux_v2, View - schematic
// LAST TIME SAVED: Dec 23 08:37:52 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioin_mux_v2 ( inmuxo, cbit,
     cbitb, min[7:0], prog );
output  inmuxo;

input  prog;

input [3:0]  cbit;
input [7:0]  min;
input [3:0]  cbitb;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nor2_lvt I_nor2_lvt ( .A(prog), .Y(en), .B(cbitb[3]));
inv_lvt I281 ( .A(inmuxob), .Y(inmuxo));
nand2_lvt I_nand2 ( .A(st2), .Y(inmuxob), .B(en));
txgate_lvt I285 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I289 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I286 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I283 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_lvt I292 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I293 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I291 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I294 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_lvt I287 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_lvt I290 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I288 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_lvt I295 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_lvt I284 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));

endmodule
// Library - io, Cell - ioinmx1mux2_v1, View - schematic
// LAST TIME SAVED: Oct 25 17:52:38 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module ioinmx1mux2_v1 ( clk, ti, bl, ce, ceb, min, pgate, prog, reset,
     vdd_cntl, wl );
output  clk, ti;


input  ceb, prog;

inout [5:0]  bl;

input [7:0]  min;
input [1:0]  reset;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [11:0]  ce;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;

wire  [11:0]  cbit;



ioin_mux_v2 I_ioin_mux ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]},
     {cbitb[1], cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clk_mux12to1 I_clk_mux12to1 ( .prog(prog), .min(ce[11:0]), .clk(clk),
     .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7], cbitb[10],
     cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7], cbit[10],
     cbit[6], cbit[4]}), .cenb(ceb));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1mem, View - schematic
// LAST TIME SAVED: Aug  9 13:33:24 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module sbox1mem ( b, bl, l, r, t, pgate, prog, reset, vdd_cntl, wl );
inout  b, l, r, t;

input  prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  reset;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;

wire  [11:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox1m3to1 I232 ( .in2(r), .cb({cbitb[3], cbitb[6]}), .op(t), .in0(l),
     .in1(b), .c({cbit[3], cbit[6]}), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb({cbitb[1], cbitb[4]}), .op(l), .in0(b),
     .in1(t), .c({cbit[1], cbit[4]}), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb({cbitb[8], cbitb[5]}), .op(b), .in0(l),
     .in1(t), .c({cbit[8], cbit[5]}), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb({cbitb[10], cbitb[7]}), .op(r), .in0(l),
     .in1(t), .c({cbit[10], cbit[7]}), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc_v4, View - schematic
// LAST TIME SAVED: Dec  7 10:50:25 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module sbox1_colbdlc_v4 ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [5:0]  ti;

inout [5:0]  bl;
inout [3:0]  r;
inout [3:0]  l;
inout [3:0]  sp4_v_b;
inout [3:0]  t_mid;

input [1:0]  oeb;
input [7:0]  min1;
input [1:0]  padin;
input [7:0]  min3;
input [7:0]  min4;
input [7:0]  min6;
input [11:0]  clk_in;
input [1:0]  out;
input [7:0]  min0;
input [11:0]  inclk_in;
input [1:0]  spioeb;
input [1:0]  spiout;
input [7:0]  ceb_in;
input [15:0]  reset;
input [7:0]  min2;
input [15:0]  vdd_cntl;
input [7:0]  min5;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spioob;

wire  [1:0]  spioo;

wire  [1:0]  oeboo;

wire  [1:0]  oeboob;



ioinmx2nor2invx2bdlc_v0 I5 ( .vdd_cntl(vdd_cntl[5:4]),
     .min2(min6[7:0]), .bankcntl(fabric_out), .bl(bl[5:0]),
     .prog(prog), .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx2nand2inv_v0 I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
ioinmx1mux2_v1 I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .ti(ti[2]), .min(min2[7:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]));
ioinmx1mux2_v1 I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .ti(ti[5]), .min(min5[7:0]), .wl(wl[15:14]), .reset(reset[15:14]),
     .pgate(pgate[15:14]));
inv_lvt I_inv_2_1_ ( .A(spioob[1]), .Y(pado[1]));
inv_lvt I_inv_2_0_ ( .A(spioob[0]), .Y(pado[0]));
inv_lvt I9_1_ ( .A(oeboo[1]), .Y(oeboob[1]));
inv_lvt I9_0_ ( .A(oeboo[0]), .Y(oeboob[0]));
inv_lvt I8_1_ ( .A(oeboob[1]), .Y(padeb[1]));
inv_lvt I8_0_ ( .A(oeboob[0]), .Y(padeb[0]));
inv_lvt inv_1_1_ ( .A(spioo[1]), .Y(spioob[1]));
inv_lvt inv_1_0_ ( .A(spioo[0]), .Y(spioob[0]));
mux2x1_hvt I10_1_ ( .in1(oeb[1]), .in0(spioeb[1]), .out(oeboo[1]),
     .sel(cdone_in));
mux2x1_hvt I10_0_ ( .in1(oeb[0]), .in0(spioeb[0]), .out(oeboo[0]),
     .sel(cdone_in));
mux2x1_hvt I_emux_1_ ( .in1(out[1]), .in0(spiout[1]), .out(spioo[1]),
     .sel(cdone_in));
mux2x1_hvt I_emux_0_ ( .in1(out[0]), .in0(spiout[0]), .out(spioo[0]),
     .sel(cdone_in));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - io, Cell - io_gmux_x2v3, View - schematic
// LAST TIME SAVED: Aug 25 13:36:12 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_gmux_x2v3 ( .cbit_colcntl({cbit[11], cbit[9]}), gout, bl,
     min0, min1, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [11:0]  cbit;
output [1:0]  gout;

inout [5:0]  bl;

input [15:0]  min1;
input [15:0]  min0;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I_xpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 I_xpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux I_g_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux I_g_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare_v4, View - schematic
// LAST TIME SAVED: Aug 25 13:36:24 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module io_gmux_x16bare_v4 ( cbit_colcntl, lc_trk_g0, lc_trk_g1, bl,
     min0, min1, min2, min3, min4, min5, min6, min7, min8, min9, min10,
     min11, min12, min13, min14, min15, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [7:0]  cbit_colcntl;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g1;

inout [5:0]  bl;

input [15:0]  min9;
input [15:0]  min12;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min0;
input [15:0]  min7;
input [15:0]  min5;
input [15:0]  min3;
input [15:0]  min4;
input [15:0]  min10;
input [15:0]  min6;
input [15:0]  min8;
input [15:0]  min15;
input [15:0]  min14;
input [15:0]  min11;
input [15:0]  reset;
input [15:0]  min2;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [15:0]  pgate;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  net187;

wire  [1:0]  net114;

wire  [1:0]  net124;

wire  [1:0]  net188;



io_gmux_x2v3 I_io_gmux_x2_7 ( .cbit_colcntl({net114[0], net114[1]}),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[15:14]));
io_gmux_x2v3 I_io_gmux_x2_6 ( .cbit_colcntl({net124[0], net124[1]}),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[13:12]));
io_gmux_x2v3 I_io_gmux_x2_2 ( .cbit_colcntl(cbit_colcntl[5:4]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[5:4]));
io_gmux_x2v3 I_io_gmux_x2_0 ( .cbit_colcntl(cbit_colcntl[1:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[1:0]));
io_gmux_x2v3 _io_gmux_x2_1 ( .cbit_colcntl(cbit_colcntl[3:2]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[3:2]));
io_gmux_x2v3 I_io_gmux_x2_4 ( .cbit_colcntl({net187[0], net187[1]}),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[9:8]));
io_gmux_x2v3 I_io_gmux_x2_5 ( .cbit_colcntl({net188[0], net188[1]}),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[11:10]));
io_gmux_x2v3 I_io_gmux_x2_3 ( .cbit_colcntl(cbit_colcntl[7:6]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog), .bl(bl[5:0]), .vdd_cntl(vdd_cntl[7:6]));

endmodule
// Library - io, Cell - insel1_lvt_imp, View - schematic
// LAST TIME SAVED: Aug 12 13:25:22 2010
// NETLIST TIME: May  5 11:56:42 2011
`timescale 1ns / 1ns 

module insel1_lvt_imp ( out, in0, in1, in2, in3, sb, sel );
output  out;

input  in0, in1, in2, in3;

input [1:0]  sb;
input [1:0]  sel;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



txgate_lvt I39 ( .in(in3), .out(outd23), .pp(sb[0]), .nn(sel[0]));
txgate_lvt I40 ( .in(in2), .out(outd23), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I33 ( .in(outd01), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_lvt I_txgate1 ( .in(in1), .out(outd01), .pp(sb[0]),
     .nn(sel[0]));
txgate_lvt I31 ( .in(in0), .out(outd01), .pp(sel[0]), .nn(sb[0]));
txgate_lvt I34 ( .in(outd23), .out(out), .pp(sb[1]), .nn(sel[1]));

endmodule
// Library - leafcell, Cell - oa4plldly_40lp, View - schematic
// LAST TIME SAVED: Jul 23 17:36:30 2010
// NETLIST TIME: May  5 11:56:40 2011
`timescale 1ns / 1ns 

module oa4plldly_40lp ( out, cbit, fda_en, in, prog );
output  out;

input  cbit, fda_en, in, prog;
supply1 vdd_;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I7 ( .A(net9), .Y(net6), .B(cbit));
anor21_hvt I1 ( .A(net031), .B(fda_en), .Y(out), .C(net6));
inv_hvt I3 ( .A(prog), .Y(net9));
inv_hvt I23 ( .A(in), .Y(net031));

endmodule
