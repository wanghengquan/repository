module via (w, w);
inout w;
wire w;

endmodule
