// Library - leafcell, Cell - tielo, View - schematic
// LAST TIME SAVED: Jul  8 16:15:53 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module tielo ( tielo );
output  tielo;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M0 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));
nch_hvt  M1 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_gwl_drv_x57, View - schematic
// LAST TIME SAVED: Apr 30 16:01:52 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwl_drv_x57 ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25,
     gnv2_b_25, gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25,
     gnv5_b_25, gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1,
     gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25, gnv2_b_25,
     gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25, gnv5_b_25,
     gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1, gwl_misc_25,
     gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

output [56:0]  gwl_wr_25;
output [56:0]  gwl_b_25;
output [56:0]  gwp_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_gwl_drv Igwl_drv_51_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[55]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[55]), .gwl_wr_25(gwl_wr_25[55]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_50_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[54]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[54]), .gwl_wr_25(gwl_wr_25[54]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_49_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[53]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[53]), .gwl_wr_25(gwl_wr_25[53]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_48_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[52]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[52]), .gwl_wr_25(gwl_wr_25[52]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_47_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[51]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[51]), .gwl_wr_25(gwl_wr_25[51]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_46_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[50]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[50]), .gwl_wr_25(gwl_wr_25[50]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_45_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[49]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[49]), .gwl_wr_25(gwl_wr_25[49]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_44_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[48]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[48]), .gwl_wr_25(gwl_wr_25[48]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_43_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[47]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[47]), .gwl_wr_25(gwl_wr_25[47]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_42_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[46]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[46]), .gwl_wr_25(gwl_wr_25[46]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_41_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[45]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[45]), .gwl_wr_25(gwl_wr_25[45]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_40_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[44]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[44]), .gwl_wr_25(gwl_wr_25[44]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_39_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[43]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[43]), .gwl_wr_25(gwl_wr_25[43]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_38_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[42]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[42]), .gwl_wr_25(gwl_wr_25[42]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_37_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[41]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[41]), .gwl_wr_25(gwl_wr_25[41]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_36_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[40]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[40]), .gwl_wr_25(gwl_wr_25[40]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_35_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[39]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[39]), .gwl_wr_25(gwl_wr_25[39]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_34_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[38]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[38]), .gwl_wr_25(gwl_wr_25[38]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_33_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[37]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[37]), .gwl_wr_25(gwl_wr_25[37]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_32_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[36]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[36]), .gwl_wr_25(gwl_wr_25[36]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_red_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[3]),
     .radd_0_25(gred_25_0), .radd_1_25(gred_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[3]), .gwl_wr_25(gwl_wr_25[3]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_red_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[2]),
     .radd_0_25(gred_b_25_0), .radd_1_25(gred_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[2]), .gwl_wr_25(gwl_wr_25[2]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_red_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[1]),
     .radd_0_25(gred_25_0), .radd_1_25(gred_b_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[1]), .gwl_wr_25(gwl_wr_25[1]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_red_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[0]),
     .radd_0_25(gred_b_25_0), .radd_1_25(gred_b_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[0]), .gwl_wr_25(gwl_wr_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_misc_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[56]),
     .radd_0_25(vddp_tieh), .radd_1_25(vddp_tieh),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_misc_25),
     .gwp_hv(gwp_hv[56]), .gwl_wr_25(gwl_wr_25[56]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_31_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[35]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[35]), .gwl_wr_25(gwl_wr_25[35]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_30_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[34]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[34]), .gwl_wr_25(gwl_wr_25[34]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_29_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[33]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[33]), .gwl_wr_25(gwl_wr_25[33]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_28_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[32]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[32]), .gwl_wr_25(gwl_wr_25[32]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_27_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[31]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[31]), .gwl_wr_25(gwl_wr_25[31]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_26_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[30]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[30]), .gwl_wr_25(gwl_wr_25[30]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_25_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[29]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[29]), .gwl_wr_25(gwl_wr_25[29]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_24_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[28]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_25), .radd_4_25(gnv4_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[28]),
     .gwl_wr_25(gwl_wr_25[28]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_23_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[27]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[27]), .gwl_wr_25(gwl_wr_25[27]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_22_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[26]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[26]), .gwl_wr_25(gwl_wr_25[26]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_21_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[25]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[25]), .gwl_wr_25(gwl_wr_25[25]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_20_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[24]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[24]), .gwl_wr_25(gwl_wr_25[24]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_19_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[23]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[23]), .gwl_wr_25(gwl_wr_25[23]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_18_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[22]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[22]), .gwl_wr_25(gwl_wr_25[22]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_17_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[21]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[21]), .gwl_wr_25(gwl_wr_25[21]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_16_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[20]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[20]),
     .gwl_wr_25(gwl_wr_25[20]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_15_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[19]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[19]), .gwl_wr_25(gwl_wr_25[19]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_14_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[18]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[18]), .gwl_wr_25(gwl_wr_25[18]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_13_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[17]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[17]), .gwl_wr_25(gwl_wr_25[17]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_12_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[16]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[16]), .gwl_wr_25(gwl_wr_25[16]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_11_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[15]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[15]), .gwl_wr_25(gwl_wr_25[15]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_10_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[14]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[14]), .gwl_wr_25(gwl_wr_25[14]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_9_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[13]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[13]), .gwl_wr_25(gwl_wr_25[13]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_8_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[12]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[12]),
     .gwl_wr_25(gwl_wr_25[12]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_7_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[11]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[11]),
     .gwl_wr_25(gwl_wr_25[11]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_6_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[10]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[10]),
     .gwl_wr_25(gwl_wr_25[10]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_5_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[9]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[9]),
     .gwl_wr_25(gwl_wr_25[9]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_4_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[8]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[8]),
     .gwl_wr_25(gwl_wr_25[8]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[7]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[7]),
     .gwl_wr_25(gwl_wr_25[7]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[6]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[6]),
     .gwl_wr_25(gwl_wr_25[6]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[5]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[5]),
     .gwl_wr_25(gwl_wr_25[5]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[4]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25),
     .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[4]), .gwl_wr_25(gwl_wr_25[4]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM, Cell - ml_gwlwr, View - schematic
// LAST TIME SAVED: Apr 30 16:02:13 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_gwlwr ( gwl_b_25, gwp_hv, wr, gwl_b_sup_25, gwp_sup_hv,
     gnv_25, gnv_b_25, gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25,
     gwl_red_25, gwlb_dis_25, gwlb_en_25, s_25, vddp_tieh, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, wr_sup_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wr_sup_25;

output [227:0]  wr;
output [56:0]  gwp_hv;
output [56:0]  gwl_b_25;

input [3:0]  s_25;
input [1:0]  gred_25;
input [5:0]  gnv_b_25;
input [5:0]  gnv_25;
input [1:0]  gred_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [56:0]  gwl_wr_25;



ml_rock_lwldrv_wr_x228 Ilwldrv_wr_x228 ( .wr_sup_25(wr_sup_25),
     .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[56:0]), .wr(wr[227:0]));
ml_gwl_drv_x57 Igwl_drv_x57 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[56:0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25_1(gred_b_25[1]), .gred_b_25_0(gred_b_25[0]),
     .gred_25_1(gred_25[1]), .gred_25_0(gred_25[0]),
     .gnv5_b_25(gnv_b_25[5]), .gnv5_25(gnv_25[5]),
     .gnv4_b_25(gnv_b_25[4]), .gnv4_25(gnv_25[4]),
     .gnv3_b_25(gnv_b_25[3]), .gnv3_25(gnv_25[3]),
     .gnv2_b_25(gnv_b_25[2]), .gnv2_25(gnv_25[2]),
     .gnv1_b_25(gnv_b_25[1]), .gnv1_25(gnv_25[1]),
     .gnv0_b_25(gnv_b_25[0]), .gnv0_25(gnv_25[0]),
     .gwp_hv(gwp_hv[56:0]), .gwl_wr_25(gwl_wr_25[56:0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_gwlwr_top, View - schematic
// LAST TIME SAVED: May  1 11:11:13 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_gwlwr_top ( fsm_gwlbdis_b_25, gwl_b_25, gwl_b_sup_25, gwp_hv,
     pgminhi_dmmy_b_25, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wr, bgr, bl_pgm_glb, vpp_int, vpxa, fsm_coladd,
     fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_b_sup_25, pgminhi_dmmy_b_25, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25;

inout  bgr, bl_pgm_glb, vpp_int, vpxa;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [227:0]  wr;
output [4:1]  sa_ngate_25;
output [56:0]  gwp_hv;
output [4:1]  sa_pgate_vpxa;
output [56:0]  gwl_b_25;

input [3:0]  fsm_trim_ipp;
input [0:0]  fsm_coladd;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_25;

wire  [1:0]  gred_25;

wire  [1:0]  gred_b_25;

wire  [5:0]  gnv_b_25;

wire  [5:0]  gnv_25;



ml_gwlwr_ctrl Igwlwr_ctrl ( .fsm_pgmdisc(fsm_pgmdisc),
     .gwlb_en_25(gwlb_en_25), .fsm_din(fsm_din),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_allwl_l(fsm_tm_allwl_l), .fsm_tm_allwl_h(fsm_tm_allwl_h),
     .fsm_tm_allbl_l(fsm_tm_allbl_l), .fsm_tm_allbl_h(fsm_tm_allbl_h),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .s_25(s_25[3:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_red_25(gwl_red_25), .gwl_nvcm_25(gwl_nvcm_25),
     .gwl_misc_25(gwl_misc_25), .gred_b_25(gred_b_25[1:0]),
     .gred_25(gred_25[1:0]), .gnv_b_25(gnv_b_25[5:0]),
     .gnv_25(gnv_25[5:0]), .wr_sup_25(wr_sup_25), .vpxa(vpxa),
     .vpp_int(vpp_int), .vddp_tieh(vddp_tieh), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr));
ml_gwlwr Igwlwr ( .gwlb_en_25(gwlb_en_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_b_25(gwl_b_25[56:0]), .wr_sup_25(wr_sup_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]), .wr(wr[227:0]),
     .gwp_hv(gwp_hv[56:0]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_spare, View - schematic
// LAST TIME SAVED: Sep 22 17:28:46 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa_spare (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:9]  net501;



rppolywo_m  R7 ( .MINUS(net033), .PLUS(net036), .BULK(gnd_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(net033), .BULK(gnd_));
rppolywo_m  R3 ( .MINUS(net042), .PLUS(net039), .BULK(gnd_));
rppolywo_m  R4 ( .MINUS(gnd_), .PLUS(net042), .BULK(gnd_));
rppolywo_m  R5 ( .MINUS(net039), .PLUS(net045), .BULK(gnd_));
rppolywo_m  R6 ( .MINUS(net045), .PLUS(net027), .BULK(gnd_));
rppolywo_m  R9 ( .MINUS(net036), .PLUS(net030), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(net030), .PLUS(net027), .BULK(gnd_));
vdd_tielow I144_9_ ( .gnd_tiel(net501[0]));
vdd_tielow I144_8_ ( .gnd_tiel(net501[1]));
vdd_tielow I144_7_ ( .gnd_tiel(net501[2]));
vdd_tielow I144_6_ ( .gnd_tiel(net501[3]));
vdd_tielow I144_5_ ( .gnd_tiel(net501[4]));
vdd_tielow I144_4_ ( .gnd_tiel(net501[5]));
vdd_tielow I144_3_ ( .gnd_tiel(net501[6]));
vdd_tielow I144_2_ ( .gnd_tiel(net501[7]));
vdd_tielow I144_1_ ( .gnd_tiel(net501[8]));
vdd_tielow I144_0_ ( .gnd_tiel(net501[9]));

endmodule
// Library - sbtlibn65lp, Cell - oai221x2_hvt, View - schematic
// LAST TIME SAVED: May  4 14:29:05 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module oai221x2_hvt ( Y, A0, A1, B0, B1, C0 );
output  Y;

input  A0, A1, B0, B1, C0;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net040), .B(GND_), .G(A0), .S(net024));
nch_hvt  M11 ( .D(Y), .B(GND_), .G(C0), .S(net040));
nch_hvt  M8 ( .D(net040), .B(GND_), .G(A1), .S(net024));
nch_hvt  M10 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M7 ( .D(Y), .B(VDD_), .G(C0), .S(vdd_));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M4 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_ls_vdd25_nor2, View - schematic
// LAST TIME SAVED: Jan 12 15:33:21 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ls_vdd25_nor2 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_25 I79 ( .A(in), .Y(out_vddio_b), .Gb(gnd_), .G(gnd_), .Pb(sup),
     .P(sup), .B(out_vddio));
nor2_25 I151 ( .A(out_vddio_b), .Y(out_vddio), .Gb(gnd_), .G(gnd_),
     .Pb(sup), .P(sup), .B(in_b));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_logic, View - schematic
// LAST TIME SAVED: May 12 10:24:23 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_ctrl_logic ( dec_trim, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25, yp1_sel,
     yp2_sel, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, yp21_b_low_b, yp_test, fsm_blkadd,
     fsm_coladd, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, tm_tcol, ysup_25 );
output  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp21_b_low_b;

input  fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h,
     fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, tm_tcol, ysup_25;

output [7:0]  yp3_sel;
output [3:0]  sb25_high_25;
output [3:0]  sbhv_high_25;
output [3:0]  sb25_gnd_25;
output [7:0]  yp2_sel;
output [1:0]  yp_test;
output [7:5]  dec_trim;
output [5:0]  yp1_sel;
output [3:0]  sbhv_gnd_25;

input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefpgm;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net319;

wire  [7:0]  yp2_sel_b;

wire  [7:0]  yp3_sel_b;

wire  [7:5]  dec_trim_b;

wire  [2:0]  tdec_b;

wire  [2:0]  tdec;

wire  [3:0]  sb25low_b;

wire  [1:0]  yp_test_b;

wire  [0:3]  net339;

wire  [0:3]  net317;

wire  [1:0]  xadd;

wire  [3:0]  sbhvlow_b;

wire  [1:0]  xadd_b;

wire  [5:0]  yp1_sel_b;

wire  [8:0]  yadd;

wire  [8:0]  yadd_b;

wire  [0:3]  net387;

wire  [0:3]  net523;

wire  [0:3]  net407;

wire  [0:3]  net299;

wire  [0:3]  net522;

wire  [0:3]  net323;

wire  [0:3]  net393;

wire  [0:3]  net409;

wire  [0:3]  net304;

wire  [0:3]  net552;

wire  [0:3]  net546;

wire  [0:3]  net321;

wire  [0:2]  net629;

wire  [0:3]  net411;

wire  [0:3]  net391;

wire  [0:3]  net549;

wire  [0:3]  net544;



oai21x2 I36 ( .A1(fsm_pgmvfy), .A0(fsm_rd), .B0(net425),
     .Y(all_blk_sel_b));
oai221x2_hvt I86_3_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[3]),
     .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai221x2_hvt I86_2_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[2]),
     .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd_b[6]));
oai221x2_hvt I86_1_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[1]),
     .A0(yadd_b[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai221x2_hvt I86_0_ ( .C0(yadd_b[8]), .A1(net565), .Y(yp1_sel_b[0]),
     .A0(yadd_b[7]), .B0(vddp_rd_overw), .B1(yadd_b[6]));
vdd_tiehigh I198 ( .vdd_tieh(vdd_tieh));
exor2_hvt I151_3_ ( .A(net339[0]), .Y(sb25low_b[3]), .B(pgm_hvact_b));
exor2_hvt I151_2_ ( .A(net339[1]), .Y(sb25low_b[2]), .B(pgm_hvact_b));
exor2_hvt I151_1_ ( .A(net339[2]), .Y(sb25low_b[1]), .B(pgm_hvact_b));
exor2_hvt I151_0_ ( .A(net339[3]), .Y(sb25low_b[0]), .B(pgm_hvact_b));
anor21_hvt I119_1_ ( .A(fsm_rowadd[1]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I119_0_ ( .A(fsm_rowadd[0]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
anor21_hvt I109 ( .A(pgm_hvact), .B(fsm_tm_allwl_h), .Y(net394),
     .C(nvcmen_buf_b));
ml_ls_vdd2vdd25 I168_3_ ( .in(net411[0]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[3]), .out_vddio(net299[0]),
     .in_b(net552[0]));
ml_ls_vdd2vdd25 I168_2_ ( .in(net411[1]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[2]), .out_vddio(net299[1]),
     .in_b(net552[1]));
ml_ls_vdd2vdd25 I168_1_ ( .in(net411[2]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[1]), .out_vddio(net299[2]),
     .in_b(net552[2]));
ml_ls_vdd2vdd25 I168_0_ ( .in(net411[3]), .sup(vddp_),
     .out_vddio_b(sb25_high_25[0]), .out_vddio(net299[3]),
     .in_b(net552[3]));
ml_ls_vdd2vdd25 I167_3_ ( .in(net407[0]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[3]), .out_vddio(net304[0]),
     .in_b(net549[0]));
ml_ls_vdd2vdd25 I167_2_ ( .in(net407[1]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[2]), .out_vddio(net304[1]),
     .in_b(net549[1]));
ml_ls_vdd2vdd25 I167_1_ ( .in(net407[2]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[1]), .out_vddio(net304[2]),
     .in_b(net549[2]));
ml_ls_vdd2vdd25 I167_0_ ( .in(net407[3]), .sup(vddp_),
     .out_vddio_b(sb25_gnd_25[0]), .out_vddio(net304[3]),
     .in_b(net549[3]));
ml_ls_vdd2vdd25 I144_3_ ( .in(net387[0]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[3]), .out_vddio(net522[0]),
     .in_b(net544[0]));
ml_ls_vdd2vdd25 I144_2_ ( .in(net387[1]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[2]), .out_vddio(net522[1]),
     .in_b(net544[1]));
ml_ls_vdd2vdd25 I144_1_ ( .in(net387[2]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[1]), .out_vddio(net522[2]),
     .in_b(net544[2]));
ml_ls_vdd2vdd25 I144_0_ ( .in(net387[3]), .sup(vddp_),
     .out_vddio_b(sbhv_high_25[0]), .out_vddio(net522[3]),
     .in_b(net544[3]));
ml_ls_vdd2vdd25 I148_3_ ( .in(net393[0]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[3]), .out_vddio(net523[0]),
     .in_b(net546[0]));
ml_ls_vdd2vdd25 I148_2_ ( .in(net393[1]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[2]), .out_vddio(net523[1]),
     .in_b(net546[1]));
ml_ls_vdd2vdd25 I148_1_ ( .in(net393[2]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[1]), .out_vddio(net523[2]),
     .in_b(net546[2]));
ml_ls_vdd2vdd25 I148_0_ ( .in(net393[3]), .sup(vddp_),
     .out_vddio_b(sbhv_gnd_25[0]), .out_vddio(net523[3]),
     .in_b(net546[3]));
ml_pump_a_clkdly I141_3_ ( .in(net393[0]), .out(net317[0]));
ml_pump_a_clkdly I141_2_ ( .in(net393[1]), .out(net317[1]));
ml_pump_a_clkdly I141_1_ ( .in(net393[2]), .out(net317[2]));
ml_pump_a_clkdly I141_0_ ( .in(net393[3]), .out(net317[3]));
ml_pump_a_clkdly I219_3_ ( .in(net387[0]), .out(net319[0]));
ml_pump_a_clkdly I219_2_ ( .in(net387[1]), .out(net319[1]));
ml_pump_a_clkdly I219_1_ ( .in(net387[2]), .out(net319[2]));
ml_pump_a_clkdly I219_0_ ( .in(net387[3]), .out(net319[3]));
ml_pump_a_clkdly I169_3_ ( .in(net411[0]), .out(net321[0]));
ml_pump_a_clkdly I169_2_ ( .in(net411[1]), .out(net321[1]));
ml_pump_a_clkdly I169_1_ ( .in(net411[2]), .out(net321[2]));
ml_pump_a_clkdly I169_0_ ( .in(net411[3]), .out(net321[3]));
ml_pump_a_clkdly I170_3_ ( .in(net407[0]), .out(net323[0]));
ml_pump_a_clkdly I170_2_ ( .in(net407[1]), .out(net323[1]));
ml_pump_a_clkdly I170_1_ ( .in(net407[2]), .out(net323[2]));
ml_pump_a_clkdly I170_0_ ( .in(net407[3]), .out(net323[3]));
nor3_hvt I111 ( .B(fsm_tm_allbl_l), .Y(yp3_b_high_b),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_l));
nor3_hvt I112 ( .C(yp3_b_high_b), .A(nvcmen_buf_b), .B(fsm_tm_allbl_h),
     .Y(net331));
nor3_hvt I57 ( .C(fsm_tm_allbl_h), .A(fsm_tm_allbl_l),
     .B(fsm_tm_testdec), .Y(net335));
anor31_hvt I155_3_ ( .A(ensb25_dec), .D(net395), .B(xadd[1]),
     .Y(net339[0]), .C(xadd[0]));
anor31_hvt I155_2_ ( .A(ensb25_dec), .D(net395), .B(xadd[1]),
     .Y(net339[1]), .C(xadd_b[0]));
anor31_hvt I155_1_ ( .A(ensb25_dec), .D(net395), .B(xadd_b[1]),
     .Y(net339[2]), .C(xadd[0]));
anor31_hvt I155_0_ ( .A(ensb25_dec), .D(net395), .B(xadd_b[1]),
     .Y(net339[3]), .C(xadd_b[0]));
anor31_hvt I121_3_ ( .A(net397), .D(net399), .B(xadd[1]),
     .Y(sbhvlow_b[3]), .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net397), .D(net399), .B(xadd[1]),
     .Y(sbhvlow_b[2]), .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net397), .D(net399), .B(xadd_b[1]),
     .Y(sbhvlow_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net397), .D(net399), .B(xadd_b[1]),
     .Y(sbhvlow_b[0]), .C(xadd_b[0]));
anor31_hvt I107 ( .A(fsm_tm_testdec), .D(net331), .B(nvcmen_buf),
     .Y(net349), .C(yadd[0]));
anor31_hvt I108 ( .A(fsm_tm_testdec), .D(net331), .B(nvcmen_buf),
     .Y(net354), .C(yadd_b[0]));
oai22x2_hvt I93 ( .A1(net381), .Y(net357), .A0(net453),
     .B0(fsm_nv_rri_trim), .B1(fsm_nv_sisi_ui));
nand4_hvt I122 ( .D(fsm_lshven), .C(pgm_hvact), .A(tm_allwl_l_b),
     .Y(net396), .B(blk_dec));
nand4_hvt I49_7_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[7]), .B(yadd[2]));
nand4_hvt I49_6_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[6]), .B(yadd[2]));
nand4_hvt I49_5_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[5]), .B(yadd[2]));
nand4_hvt I49_4_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[4]), .B(yadd[2]));
nand4_hvt I49_3_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[3]), .B(yadd_b[2]));
nand4_hvt I49_2_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[2]), .B(yadd_b[2]));
nand4_hvt I49_1_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[1]), .B(yadd_b[2]));
nand4_hvt I49_0_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[0]), .B(yadd_b[2]));
nand4_hvt I27 ( .D(fsm_blkadd[0]), .Y(blk_dec_b), .B(fsm_blkadd[2]),
     .C(fsm_blkadd[1]), .A(fsm_blkadd[3]));
inv_hvt I207 ( .A(net0579), .Y(ref_pgm));
inv_hvt I200 ( .A(fsm_tm_testdec), .Y(net377));
inv_hvt I120_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I120_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I181 ( .A(all_blk_sel_b), .Y(net381));
inv_hvt I161 ( .A(net570), .Y(net383));
inv_hvt I158 ( .A(pgm_hvact_b), .Y(pgm_hvact));
inv_hvt I142_3_ ( .A(net544[0]), .Y(net387[0]));
inv_hvt I142_2_ ( .A(net544[1]), .Y(net387[1]));
inv_hvt I142_1_ ( .A(net544[2]), .Y(net387[2]));
inv_hvt I142_0_ ( .A(net544[3]), .Y(net387[3]));
inv_hvt I157 ( .A(fsm_pgmvfy), .Y(net389));
inv_hvt I134_3_ ( .A(sbhvlow_b[3]), .Y(net391[0]));
inv_hvt I134_2_ ( .A(sbhvlow_b[2]), .Y(net391[1]));
inv_hvt I134_1_ ( .A(sbhvlow_b[1]), .Y(net391[2]));
inv_hvt I134_0_ ( .A(sbhvlow_b[0]), .Y(net391[3]));
inv_hvt I143_3_ ( .A(net546[0]), .Y(net393[0]));
inv_hvt I143_2_ ( .A(net546[1]), .Y(net393[1]));
inv_hvt I143_1_ ( .A(net546[2]), .Y(net393[2]));
inv_hvt I143_0_ ( .A(net546[3]), .Y(net393[3]));
inv_hvt I160 ( .A(net394), .Y(net395));
inv_hvt I123 ( .A(net396), .Y(net397));
inv_hvt I125 ( .A(net490), .Y(net399));
inv_hvt I189 ( .A(fsm_nvcmen), .Y(nvcmen_buf_b));
inv_hvt I164 ( .A(net402), .Y(net403));
inv_hvt I131 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I171_3_ ( .A(net549[0]), .Y(net407[0]));
inv_hvt I171_2_ ( .A(net549[1]), .Y(net407[1]));
inv_hvt I171_1_ ( .A(net549[2]), .Y(net407[2]));
inv_hvt I171_0_ ( .A(net549[3]), .Y(net407[3]));
inv_hvt I172_3_ ( .A(sb25low_b[3]), .Y(net409[0]));
inv_hvt I172_2_ ( .A(sb25low_b[2]), .Y(net409[1]));
inv_hvt I172_1_ ( .A(sb25low_b[1]), .Y(net409[2]));
inv_hvt I172_0_ ( .A(sb25low_b[0]), .Y(net409[3]));
inv_hvt I173_3_ ( .A(net552[0]), .Y(net411[0]));
inv_hvt I173_2_ ( .A(net552[1]), .Y(net411[1]));
inv_hvt I173_1_ ( .A(net552[2]), .Y(net411[2]));
inv_hvt I173_0_ ( .A(net552[3]), .Y(net411[3]));
inv_hvt I97 ( .A(fsm_multibl_read), .Y(net413));
inv_hvt I94 ( .A(net357), .Y(vddp_rd_overw));
inv_hvt I84 ( .A(nvcmen_buf_b), .Y(nvcmen_buf));
inv_hvt I72_7_ ( .A(yp2_sel_b[7]), .Y(yp2_sel[7]));
inv_hvt I72_6_ ( .A(yp2_sel_b[6]), .Y(yp2_sel[6]));
inv_hvt I72_5_ ( .A(yp2_sel_b[5]), .Y(yp2_sel[5]));
inv_hvt I72_4_ ( .A(yp2_sel_b[4]), .Y(yp2_sel[4]));
inv_hvt I72_3_ ( .A(yp2_sel_b[3]), .Y(yp2_sel[3]));
inv_hvt I72_2_ ( .A(yp2_sel_b[2]), .Y(yp2_sel[2]));
inv_hvt I72_1_ ( .A(yp2_sel_b[1]), .Y(yp2_sel[1]));
inv_hvt I72_0_ ( .A(yp2_sel_b[0]), .Y(yp2_sel[0]));
inv_hvt I66 ( .A(net349), .Y(net622));
inv_hvt I46_8_ ( .A(fsm_coladd[8]), .Y(yadd_b[8]));
inv_hvt I46_7_ ( .A(fsm_coladd[7]), .Y(yadd_b[7]));
inv_hvt I46_6_ ( .A(fsm_coladd[6]), .Y(yadd_b[6]));
inv_hvt I46_5_ ( .A(fsm_coladd[5]), .Y(yadd_b[5]));
inv_hvt I46_4_ ( .A(fsm_coladd[4]), .Y(yadd_b[4]));
inv_hvt I46_3_ ( .A(fsm_coladd[3]), .Y(yadd_b[3]));
inv_hvt I46_2_ ( .A(fsm_coladd[2]), .Y(yadd_b[2]));
inv_hvt I46_1_ ( .A(fsm_coladd[1]), .Y(yadd_b[1]));
inv_hvt I46_0_ ( .A(fsm_coladd[0]), .Y(yadd_b[0]));
inv_hvt I201 ( .A(fsm_tm_rd_mode), .Y(net425));
inv_hvt I25_2_ ( .A(tdec_b[2]), .Y(tdec[2]));
inv_hvt I25_1_ ( .A(tdec_b[1]), .Y(tdec[1]));
inv_hvt I25_0_ ( .A(tdec_b[0]), .Y(tdec[0]));
inv_hvt I24_2_ ( .A(net629[0]), .Y(tdec_b[2]));
inv_hvt I24_1_ ( .A(net629[1]), .Y(tdec_b[1]));
inv_hvt I24_0_ ( .A(net629[2]), .Y(tdec_b[0]));
inv_hvt I38_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I38_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I38_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I40 ( .A(net591), .Y(sa_bl_to_pgm_glb));
inv_hvt I103 ( .A(net511), .Y(en_blinhi_pgm_b));
inv_hvt I47_8_ ( .A(yadd_b[8]), .Y(yadd[8]));
inv_hvt I47_7_ ( .A(yadd_b[7]), .Y(yadd[7]));
inv_hvt I47_6_ ( .A(yadd_b[6]), .Y(yadd[6]));
inv_hvt I47_5_ ( .A(yadd_b[5]), .Y(yadd[5]));
inv_hvt I47_4_ ( .A(yadd_b[4]), .Y(yadd[4]));
inv_hvt I47_3_ ( .A(yadd_b[3]), .Y(yadd[3]));
inv_hvt I47_2_ ( .A(yadd_b[2]), .Y(yadd[2]));
inv_hvt I47_1_ ( .A(yadd_b[1]), .Y(yadd[1]));
inv_hvt I47_0_ ( .A(yadd_b[0]), .Y(yadd[0]));
inv_hvt I71 ( .A(net500), .Y(yp21_b_low_b));
inv_hvt I51_7_ ( .A(yp3_sel_b[7]), .Y(yp3_sel[7]));
inv_hvt I51_6_ ( .A(yp3_sel_b[6]), .Y(yp3_sel[6]));
inv_hvt I51_5_ ( .A(yp3_sel_b[5]), .Y(yp3_sel[5]));
inv_hvt I51_4_ ( .A(yp3_sel_b[4]), .Y(yp3_sel[4]));
inv_hvt I51_3_ ( .A(yp3_sel_b[3]), .Y(yp3_sel[3]));
inv_hvt I51_2_ ( .A(yp3_sel_b[2]), .Y(yp3_sel[2]));
inv_hvt I51_1_ ( .A(yp3_sel_b[1]), .Y(yp3_sel[1]));
inv_hvt I51_0_ ( .A(yp3_sel_b[0]), .Y(yp3_sel[0]));
inv_hvt I61 ( .A(net594), .Y(net443));
inv_hvt I28 ( .A(blk_dec_b), .Y(blk_dec));
inv_hvt I69 ( .A(net354), .Y(net612));
inv_hvt I117_1_ ( .A(yp_test_b[1]), .Y(yp_test[1]));
inv_hvt I117_0_ ( .A(yp_test_b[0]), .Y(yp_test[0]));
inv_hvt I185 ( .A(tm_tcol), .Y(net451));
inv_hvt I90 ( .A(net562), .Y(net453));
inv_25 I104 ( .IN(net606), .OUT(en_blinhi_pgm_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net620), .OUT(yp3_b_high_even_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I79 ( .IN(net610), .OUT(yp3_b_high_odd_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I77 ( .IN(net615), .OUT(yp3_b_low_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
nand3_hvt I204 ( .Y(yp1_sel_b[4]), .B(yadd_b[7]), .C(yadd[8]),
     .A(yadd_b[6]));
nand3_hvt I205 ( .Y(yp1_sel_b[5]), .B(yadd_b[7]), .C(yadd[6]),
     .A(yadd[8]));
nand3_hvt I156 ( .Y(pgm_hvact_b), .B(fsm_pgm), .C(net389),
     .A(fsm_lshven));
nand3_hvt I127 ( .Y(net490), .B(pgm_hvact), .C(fsm_tm_allwl_h),
     .A(fsm_lshven));
nand3_hvt I163 ( .C(tm_allwl_l_b), .A(fsm_vpxaset), .Y(net402),
     .B(sa_bl_to_blsa));
nand3_hvt I70 ( .C(nvcmen_buf), .A(net588), .Y(net500), .B(net377));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(tdec[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(tdec[1]), .C(tdec_b[0]),
     .A(tdec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(tdec_b[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I73_7_ ( .A(yadd[5]), .C(yadd[3]), .Y(yp2_sel_b[7]),
     .B(yadd[4]));
nand3_hvt I73_6_ ( .A(yadd[5]), .C(yadd_b[3]), .Y(yp2_sel_b[6]),
     .B(yadd[4]));
nand3_hvt I73_5_ ( .A(yadd[5]), .C(yadd[3]), .Y(yp2_sel_b[5]),
     .B(yadd_b[4]));
nand3_hvt I73_4_ ( .A(yadd[5]), .C(yadd_b[3]), .Y(yp2_sel_b[4]),
     .B(yadd_b[4]));
nand3_hvt I73_3_ ( .A(yadd_b[5]), .C(yadd[3]), .Y(yp2_sel_b[3]),
     .B(yadd[4]));
nand3_hvt I73_2_ ( .A(yadd_b[5]), .C(yadd_b[3]), .Y(yp2_sel_b[2]),
     .B(yadd[4]));
nand3_hvt I73_1_ ( .A(yadd_b[5]), .C(yadd[3]), .Y(yp2_sel_b[1]),
     .B(yadd_b[4]));
nand3_hvt I73_0_ ( .A(yadd_b[5]), .C(yadd_b[3]), .Y(yp2_sel_b[0]),
     .B(yadd_b[4]));
nor4_hvt I98 ( .B(fsm_tm_allbl_l), .Y(net511), .D(nvcmen_buf_b),
     .A(net573), .C(fsm_tm_allbl_l));
nor4_hvt I52 ( .D(net580), .B(fsm_tm_allbl_h), .Y(ymux_dis_b),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_h));
nor2_hvt I202 ( .A(yp1_sel_b[4]), .B(tm_tcol), .Y(yp1_sel[4]));
nor2_hvt I203 ( .A(yp1_sel_b[5]), .B(tm_tcol), .Y(yp1_sel[5]));
nor2_hvt I195 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I128_3_ ( .B(net317[0]), .A(net391[0]), .Y(net544[0]));
nor2_hvt I128_2_ ( .B(net317[1]), .A(net391[1]), .Y(net544[1]));
nor2_hvt I128_1_ ( .B(net317[2]), .A(net391[2]), .Y(net544[2]));
nor2_hvt I128_0_ ( .B(net317[3]), .A(net391[3]), .Y(net544[3]));
nor2_hvt I140_3_ ( .A(net319[0]), .Y(net546[0]), .B(sbhvlow_b[3]));
nor2_hvt I140_2_ ( .A(net319[1]), .Y(net546[1]), .B(sbhvlow_b[2]));
nor2_hvt I140_1_ ( .A(net319[2]), .Y(net546[2]), .B(sbhvlow_b[1]));
nor2_hvt I140_0_ ( .A(net319[3]), .Y(net546[3]), .B(sbhvlow_b[0]));
nor2_hvt I176_3_ ( .A(sb25low_b[3]), .Y(net549[0]), .B(net321[0]));
nor2_hvt I176_2_ ( .A(sb25low_b[2]), .Y(net549[1]), .B(net321[1]));
nor2_hvt I176_1_ ( .A(sb25low_b[1]), .Y(net549[2]), .B(net321[2]));
nor2_hvt I176_0_ ( .A(sb25low_b[0]), .Y(net549[3]), .B(net321[3]));
nor2_hvt I177_3_ ( .A(net323[0]), .Y(net552[0]), .B(net409[0]));
nor2_hvt I177_2_ ( .A(net323[1]), .Y(net552[1]), .B(net409[1]));
nor2_hvt I177_1_ ( .A(net323[2]), .Y(net552[2]), .B(net409[2]));
nor2_hvt I177_0_ ( .A(net323[3]), .Y(net552[3]), .B(net409[3]));
nor2_hvt I114 ( .A(tm_tcol), .B(net600), .Y(ymux_en_core));
nor2_hvt I186 ( .A(net451), .B(net600), .Y(ymux_test_en));
nor2_hvt I88 ( .A(fsm_tm_rd_mode), .B(fsm_pgmvfy), .Y(net562));
nor2_hvt I96 ( .A(net357), .B(net413), .Y(net565));
nor2_hvt I75_3_ ( .A(yp1_sel_b[3]), .B(tm_tcol), .Y(yp1_sel[3]));
nor2_hvt I75_2_ ( .A(yp1_sel_b[2]), .B(tm_tcol), .Y(yp1_sel[2]));
nor2_hvt I75_1_ ( .A(yp1_sel_b[1]), .B(tm_tcol), .Y(yp1_sel[1]));
nor2_hvt I75_0_ ( .A(yp1_sel_b[0]), .B(tm_tcol), .Y(yp1_sel[0]));
nor2_hvt I206 ( .A(fsm_pgmvfy), .B(fsm_pgm), .Y(net0579));
nand2_hvt I162 ( .A(blk_dec), .Y(net570), .B(tm_allwl_l_b));
nand2_hvt I101 ( .A(pgm_hvact), .Y(net573), .B(pgm_hvact));
nand2_hvt I35 ( .B(one_blk_sel_b), .Y(sa_bl_to_blsa),
     .A(all_blk_sel_b));
nand2_hvt I53 ( .A(fsm_nvcmen), .B(fsm_lshven), .Y(net580));
nand2_hvt I116_1_ ( .A(yadd[0]), .Y(yp_test_b[1]), .B(ymux_test_en));
nand2_hvt I116_0_ ( .A(yadd_b[0]), .Y(yp_test_b[0]), .B(ymux_test_en));
nand2_hvt I59 ( .A(fsm_lshven), .Y(net588), .B(pgm_hvact));
nand2_hvt I39 ( .A(blk_dec), .Y(net591), .B(fsm_pgmien));
nand2_hvt I60 ( .A(net588), .Y(net594), .B(net335));
nand2_hvt I89 ( .A(fsm_tm_rd_mode), .Y(one_blk_sel_b), .B(blk_dec));
oai21x2_hvt I55 ( .A1(sa_bl_to_blsa), .Y(net600), .A0(blk_dec),
     .B0(ymux_dis_b));
ml_ls_vdd25_nor2 I106 ( .in(net511), .sup(ysup_25),
     .out_vddio_b(net605), .out_vddio(net606), .in_b(en_blinhi_pgm_b));
ml_ls_vdd25_nor2 I68 ( .in(net354), .sup(ysup_25),
     .out_vddio_b(net610), .out_vddio(net611), .in_b(net612));
ml_ls_vdd25_nor2 I192 ( .in(net594), .sup(ysup_25),
     .out_vddio_b(net615), .out_vddio(net616), .in_b(net443));
ml_ls_vdd25_nor2 I65 ( .in(net349), .sup(ysup_25),
     .out_vddio_b(net620), .out_vddio(net621), .in_b(net622));
mux2_hvt I152 ( .in1(net383), .in0(net403), .out(ensb25_dec),
     .sel(pgm_hvact));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net629[0]), .sel(ref_pgm));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net629[1]), .sel(ref_pgm));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net629[2]), .sel(ref_pgm));

endmodule
// Library - NVCM, Cell - ml_core_sa_resbot_m2, View - schematic
// LAST TIME SAVED: Sep  5 15:33:35 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa_resbot_m2 ( bl_in, bl_out, div_2r, div_3r, nwell,
     sa_ngate_25, sa_pgate_vpxa );
inout  bl_in, bl_out, div_2r, div_3r, nwell;


input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M4 ( .D(net115), .B(gnd_), .G(sa_ngate_25[4]), .S(bl_out));
nch_25  M3 ( .D(net090), .B(gnd_), .G(sa_ngate_25[3]), .S(net115));
nch_25  M0 ( .D(net086), .B(gnd_), .G(sa_ngate_25[2]), .S(net090));
nch_25  M32 ( .D(net111), .B(gnd_), .G(sa_ngate_25[1]), .S(net086));
pch_25  M5 ( .D(bl_out), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net115));
pch_25  M1 ( .D(net090), .B(nwell), .G(sa_pgate_vpxa[2]), .S(net086));
pch_25  M2 ( .D(net115), .B(nwell), .G(sa_pgate_vpxa[3]), .S(net090));
pch_25  M37 ( .D(net086), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net111));
rppolywo_m  R31 ( .MINUS(net099), .PLUS(div_3r), .BULK(gnd_));
rppolywo_m  R32 ( .MINUS(div_2r), .PLUS(net099), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(div_3r), .PLUS(net111), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net111), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R30 ( .MINUS(net0111), .PLUS(div_2r), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(net0111), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_gwlgnd_nor2, View - schematic
// LAST TIME SAVED: Jan 23 10:17:03 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_rock_gwlgnd_nor2 ( gwl_gnd_25, gwl_b_sup_25, gwl_b_25,
     gwl_b_gnden_25 );
output  gwl_gnd_25;

inout  gwl_b_sup_25;

input  gwl_b_25, gwl_b_gnden_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(net14), .B(GND_), .G(gwl_b_gnden_25), .S(GND_));
nch_25  M0 ( .D(gwl_gnd_25), .B(GND_), .G(gwl_b_25), .S(net14));
pch_25  M2 ( .D(gwl_gnd_25), .B(gwl_b_sup_25), .G(gwl_b_25),
     .S(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_refres, View - schematic
// LAST TIME SAVED: Sep  8 13:55:16 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa_refres ( bot, nwell, wp_ref, sa_ngate_25,
     sa_pgate_vpxa );
inout  bot, nwell, wp_ref;


input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M32 ( .D(net44), .B(gnd_), .G(sa_ngate_25[1]), .S(net40));
nch_25  M2 ( .D(net50), .B(gnd_), .G(sa_ngate_25[3]), .S(net084));
nch_25  M6 ( .D(net084), .B(gnd_), .G(sa_ngate_25[4]), .S(bot));
nch_25  M1 ( .D(net40), .B(gnd_), .G(sa_ngate_25[2]), .S(net50));
pch_25  M3 ( .D(net084), .B(nwell), .G(sa_pgate_vpxa[3]), .S(net50));
pch_25  M37 ( .D(net40), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net44));
pch_25  M5 ( .D(bot), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net084));
pch_25  M0 ( .D(net50), .B(nwell), .G(sa_pgate_vpxa[2]), .S(net40));
rppolywo_m  R2 ( .MINUS(net088), .PLUS(net090), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(bot), .PLUS(net32), .BULK(gnd_));
rppolywo_m  R6 ( .MINUS(net32), .PLUS(net088), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net090), .PLUS(net44), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net44), .PLUS(wp_ref), .BULK(gnd_));

endmodule
// Library - xpmem, Cell - ml_buf_ice5_2, View - schematic
// LAST TIME SAVED: Aug 15 18:07:29 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_buf_ice5_2 ( o, in, sel );
output  o;

input  in, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));
inv_hvt I391 ( .A(net77), .Y(o));

endmodule
// Library - NVCM, Cell - ml_core_sa_resbot, View - schematic
// LAST TIME SAVED: Apr  9 15:18:14 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa_resbot ( bl_in, bl_out, div_2r, div_3r, nwell,
     sa_ngate_25, sa_pgate_vpxa );
inout  bl_in, bl_out, div_2r, div_3r, nwell;


input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M4 ( .D(net115), .B(gnd_), .G(sa_ngate_25[4]), .S(bl_out));
nch_25  M3 ( .D(div_2r), .B(gnd_), .G(sa_ngate_25[3]), .S(net115));
nch_25  M0 ( .D(div_3r), .B(gnd_), .G(sa_ngate_25[2]), .S(div_2r));
nch_25  M32 ( .D(net111), .B(gnd_), .G(sa_ngate_25[1]), .S(div_3r));
pch_25  M5 ( .D(bl_out), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net115));
pch_25  M1 ( .D(div_2r), .B(nwell), .G(sa_pgate_vpxa[2]), .S(div_3r));
pch_25  M2 ( .D(net115), .B(nwell), .G(sa_pgate_vpxa[3]), .S(div_2r));
pch_25  M37 ( .D(div_3r), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net111));
rppolywo_m  R31 ( .MINUS(net099), .PLUS(div_3r), .BULK(gnd_));
rppolywo_m  R32 ( .MINUS(div_2r), .PLUS(net099), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(div_3r), .PLUS(net111), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net111), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R30 ( .MINUS(net115), .PLUS(div_2r), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(net115), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp, View - schematic
// LAST TIME SAVED: Jan 21 10:22:42 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp ( wp, ngate_25, gwl_b_25, gwl_gnd_25, gwp_hv,
     s_b_25, s_b_hv );
output  wp;

inout  ngate_25;

input  gwl_b_25, gwl_gnd_25, gwp_hv, s_b_25, s_b_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M6 ( .D(wp), .B(gwp_hv), .G(s_b_hv), .S(gwp_hv));
nch_25  M11 ( .D(net18), .B(GND_), .G(s_b_25), .S(gwl_gnd_25));
nch_25  M12 ( .D(wp), .B(GND_), .G(ngate_25), .S(net18));
nch_25  M10 ( .D(net18), .B(GND_), .G(gwl_b_25), .S(gwl_gnd_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp, View - schematic
// LAST TIME SAVED: Jan 21 17:21:12 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_b_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M4_1_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M0 ( .D(out_div), .B(vddp_), .G(in_div), .S(net65));
pch_25  M3 ( .D(out_ref), .B(vddp_), .G(in_ref), .S(net65));
nch_25  M1 ( .D(out_ref), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M2 ( .D(out_div), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M8 ( .D(out_ref), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M5 ( .D(out_div), .B(GND_), .G(saen_b_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_top, View - schematic
// LAST TIME SAVED: Jan 21 17:21:37 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp_top ( sa_out, in_div, in_ref, saen_25 );
output  sa_out;

input  in_div, in_ref, saen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I85 ( .IN(saen_25), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(sa_out_b_25), .OUT(net051), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net038), .OUT(sa_out), .P(vdd_), .Pb(vdd_), .G(gnd_),
     .Gb(gnd_));
nand2_25 I80 ( .G(gnd_), .Pb(vdd_), .A(net051), .Y(net038), .P(vdd_),
     .B(saen_25), .Gb(gnd_));
nand2_25 I96 ( .G(gnd_), .Pb(vddp_), .A(out_div2), .Y(sa_out_b_25),
     .P(vddp_), .B(saen_25), .Gb(gnd_));
ml_core_sa_comp Icore_sa_comp0 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp Icore_sa_comp1 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref2), .in_div(in_div2),
     .out_ref(net73), .out_div(out_div2));
nch_25  M0 ( .D(net039), .B(gnd_), .G(saen_25), .S(gnd_));
pch_25  M43 ( .D(sa_bias), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M4_4_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_3_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_2_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_1_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
rppolywo_m  R0 ( .MINUS(net039), .PLUS(net45), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net45), .PLUS(sa_bias), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa, View - schematic
// LAST TIME SAVED: Sep 11 11:12:56 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa ( nv_dataout, blsa, vpxa, dec_ok_25, dec_trim,
     fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, tm_testdec_wr );
output  nv_dataout;

inout  blsa, vpxa;

input  dec_ok_25, fsm_rst_b, fsm_sample, fsm_tm_testdec, saen_25,
     saen_b_vpxa, testdec_en_b_25, tm_testdec_wr;

input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
input [7:5]  dec_trim;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_core_sa_resbot_m2 res_bot_ref_m2 ( .div_2r(dec_ref_2r),
     .div_3r(net0155), .bl_out(net0181), .nwell(nwell),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .bl_in(blsa_ref));
nch  M1 ( .D(net0173), .B(GND_), .G(testdec_b), .S(net0269));
nch  M27 ( .D(net0103), .B(GND_), .G(vdd_tieh), .S(blsa_ref));
vdd_tielow I204 ( .gnd_tiel(gnnd_tlow));
inv_25 I38 ( .IN(testdec_en_b_25), .OUT(dec_gate_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I222 ( .IN(dec_ok_25), .OUT(net0114), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I224 ( .IN(net0114), .OUT(net098), .P(vdd_), .Pb(vdd_),
     .G(gnd_), .Gb(gnd_));
nor2_hvt I214 ( .B(high_res_b), .Y(net0132), .A(testdec));
mux2_hvt I206 ( .in1(blsa), .in0(dec_in_3r), .out(in_div),
     .sel(testdec_b));
mux2_hvt I207 ( .in1(dec_ref_2r), .in0(dec_ref_2r), .out(in_ref),
     .sel(testdec_b));
mux2_hvt I219 ( .in1(net098), .in0(sa_out), .out(net0191),
     .sel(tm_testdec_wr));
rppolywo_m  R3 ( .MINUS(net0115), .PLUS(net0112), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net0169), .PLUS(net0115), .BULK(gnd_));
ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 ( .gwl_b_gnden_25(vdd_tieh),
     .gwl_b_sup_25(vpxa), .gwl_b_25(saen_b_vpxa),
     .gwl_gnd_25(gwl_gnd_25_ref));
inv_hvt I208 ( .A(fsm_tm_testdec), .Y(testdec_b));
inv_hvt I220 ( .A(testdec_b), .Y(testdec));
inv_hvt I213 ( .A(net0132), .Y(net0120));
inv_hvt I215 ( .A(fsm_rst_b), .Y(net131));
inv_hvt I136 ( .A(rd_out_b), .Y(nv_dataout));
nor3_hvt I102 ( .B(dec_trim[6]), .Y(high_res_b), .A(dec_trim[5]),
     .C(dec_trim[7]));
vddp_tiehigh I169 ( .vddp_tieh(vddp_tieh));
vdd_tiehigh I117_2_ ( .vdd_tieh(nwell));
vdd_tiehigh I117_1_ ( .vdd_tieh(nwell));
vdd_tiehigh I117_0_ ( .vdd_tieh(nwell));
vdd_tiehigh I168 ( .vdd_tieh(vdd_tieh));
ml_core_sa_refres Irefres ( .nwell(wp_ref),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .wp_ref(wp_ref), .bot(net0173));
ml_core_sa_resbot res_bot_sen ( .div_2r(net0228), .div_3r(dec_in_3r),
     .bl_out(net0112), .nwell(nwell),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .bl_in(blsa));
ml_rock_lwldrv_wp Irock_lwldrv_wp ( .gwl_gnd_25(gwl_gnd_25_ref),
     .s_b_hv(vddp_tieh), .gwp_hv(vddp_tieh), .gwl_b_25(gnnd_tlow),
     .ngate_25(vpxa), .s_b_25(vpxa), .wp(wp_ref));
sbtlibn65lp_ml_dff_schematic I132 ( .R(net131), .D(net0191),
     .CLK(fsm_sample), .QN(rd_out_b), .Q(net135));
ml_core_sa_comp_top Icore_sa_comp_top ( .saen_25(saen_25),
     .in_ref(in_ref), .in_div(in_div), .sa_out(sa_out));
nch_hvt  M48 ( .D(net0169), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M46 ( .D(net0112), .B(GND_), .G(net0120), .S(gnd_));
nch_hvt  M45 ( .D(net0181), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M47 ( .D(net0115), .B(GND_), .G(dec_trim[5]), .S(gnd_));
nch_hvt  M14 ( .D(net184), .B(GND_), .G(vdd_tieh), .S(net0103));
nch_hvt  M16 ( .D(net208), .B(GND_), .G(vdd_tieh), .S(net184));
nch_25  M21 ( .D(blsa_ref), .B(GND_), .G(saen_b_vpxa), .S(gnd_));
nch_25  M23 ( .D(vdd_), .B(gnd_), .G(dec_gate_25), .S(net0269));
nch_25  M25 ( .D(net0269), .B(GND_), .G(vddp_tieh), .S(net208));

endmodule
// Library - NVCM, Cell - ml_core_sa_top, View - schematic
// LAST TIME SAVED: Apr 18 11:05:06 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_sa_top ( nv_dataout, bl_out, bl_pgm_glb, vpxa,
     dec_ok_25, dec_trim, fsm_rst_b, fsm_sample, fsm_tm_testdec,
     sa_bl_to_blsa, sa_bl_to_pgm_glb, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, tm_dma, tm_testdec_wr );
output  nv_dataout;

inout  bl_out, bl_pgm_glb, vpxa;

input  dec_ok_25, fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, saen_25, saen_b_vpxa, testdec_en_b_25, tm_dma,
     tm_testdec_wr;

input [7:5]  dec_trim;
input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch  M27 ( .D(bl_out), .B(GND_), .G(net81), .S(net71));
inv_hvt I108 ( .A(net063), .Y(net061));
inv_hvt I131 ( .A(tm_dma), .Y(net063));
inv_hvt I101 ( .A(net69), .Y(net77));
inv_hvt I102 ( .A(sa_bl_to_pgm_glb), .Y(net69));
inv_hvt I167 ( .A(sa_bl_to_blsa), .Y(net73));
inv_hvt I96 ( .A(net73), .Y(net81));
pch_hvt  M1 ( .D(bl_pgm_glb), .B(VDD_), .G(net69), .S(bl_out));
pch_hvt  M11 ( .D(VDD_), .B(VDD_), .G(net73), .S(VDD_));
nch_hvt  M2 ( .D(bl_out), .B(GND_), .G(net77), .S(bl_pgm_glb));
nch_hvt  M4 ( .D(net71), .B(GND_), .G(net061), .S(gnd_));
ml_core_sa Iml_core_sa ( .tm_testdec_wr(tm_testdec_wr),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_tm_testdec(fsm_tm_testdec), .dec_ok_25(dec_ok_25),
     .saen_b_vpxa(saen_b_vpxa), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .dec_trim(dec_trim[7:5]),
     .nv_dataout(nv_dataout), .vpxa(vpxa), .blsa(net71));

endmodule
// Library - NVCM, Cell - ml_s_b_hv_sw, View - schematic
// LAST TIME SAVED: May 16 11:29:12 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_s_b_hv_sw ( sbout_hv, ssup_hv, sbout_gnd_25, sbout_high_25,
     vddp_tieh );
inout  sbout_hv, ssup_hv;

input  sbout_gnd_25, sbout_high_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I114 ( .IN(sbout_high_25), .OUT(net62), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M23 ( .D(sbout_hv), .B(GND_), .G(vddp_tieh), .S(net34));
nch_25  M7 ( .D(net34), .B(GND_), .G(sbout_gnd_25), .S(gnd_));
pch_25  M5 ( .D(net46), .B(ssup_hv), .G(sbout_hv_b), .S(ssup_hv));
pch_25  M14 ( .D(sbout_hv), .B(net46), .G(sbout_gnd_25), .S(net46));
ml_hv_ls_inv Iml_hv_ls_inv_vppt ( .vddp_tieh(vddp_tieh),
     .sel_b_25(net62), .sel_25(sbout_high_25), .out_b_hv(sbout_hv_b),
     .in_hv(ssup_hv));

endmodule
// Library - NVCM, Cell - ml_wp_ctrl, View - schematic
// LAST TIME SAVED: Mar  9 16:06:25 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_wp_ctrl ( s_b_25, s_b_hv, sb25sup_25, sbhvsup_hv,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25 );
inout  sb25sup_25, sbhvsup_hv;


inout [3:0]  s_b_25;
inout [3:0]  s_b_hv;

input [3:0]  sbhv_high_25;
input [3:0]  sb25_gnd_25;
input [3:0]  sbhv_gnd_25;
input [3:0]  sb25_high_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I21_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_0_ ( .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_25_sw_3_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[3]),
     .sbout_hv(s_b_25[3]), .sbout_high_25(sb25_high_25[3]));
ml_s_b_hv_sw Iml_s_b_25_sw_2_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[2]),
     .sbout_hv(s_b_25[2]), .sbout_high_25(sb25_high_25[2]));
ml_s_b_hv_sw Iml_s_b_25_sw_1_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[1]),
     .sbout_hv(s_b_25[1]), .sbout_high_25(sb25_high_25[1]));
ml_s_b_hv_sw Iml_s_b_25_sw_0_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[0]),
     .sbout_hv(s_b_25[0]), .sbout_high_25(sb25_high_25[0]));
ml_s_b_hv_sw Iml_s_b_hv_sw_3_ ( .sbout_high_25(sbhv_high_25[3]),
     .sbout_hv(s_b_hv[3]), .sbout_gnd_25(sbhv_gnd_25[3]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_2_ ( .sbout_high_25(sbhv_high_25[2]),
     .sbout_hv(s_b_hv[2]), .sbout_gnd_25(sbhv_gnd_25[2]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_1_ ( .sbout_high_25(sbhv_high_25[1]),
     .sbout_hv(s_b_hv[1]), .sbout_gnd_25(sbhv_gnd_25[1]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_0_ ( .sbout_high_25(sbhv_high_25[0]),
     .sbout_hv(s_b_hv[0]), .sbout_gnd_25(sbhv_gnd_25[0]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_sup_25, View - schematic
// LAST TIME SAVED: Dec 18 17:40:05 2007
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module oai21x2_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
nch_25  M6 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
nch_25  M7 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));
pch_25  M4 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
pch_25  M0 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));
pch_25  M5 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yptest, View - schematic
// LAST TIME SAVED: Feb 26 14:41:48 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yptest ( yp_test_25, yp_test_b_25, yp_test,
     yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25, ysup_25 );
output  yp_test_25, yp_test_b_25;

input  yp_test, yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25,
     ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



oai21x2_sup_25 I180 ( .A1(yp_test_b_low_ysup_25), .Y(yp_test_b_25),
     .A0(net37), .B0(yp_test_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(yp_test), .sup(ysup_25),
     .out_vddio_b(net028), .out_vddio(net37), .in_b(net40));
inv_hvt I181 ( .A(yp_test), .Y(net40));
inv_25 I182 ( .IN(net028), .OUT(yp_test_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - xpmem, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jun  5 11:34:46 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yp3, View - schematic
// LAST TIME SAVED: Feb 26 14:41:31 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp3 ( yp3_25, yp3_b_25, yp3_b_high_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, ysup_25 );
output  yp3_25, yp3_b_25;

input  yp3_b_high_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I201 ( .A(yp3_sel), .Y(net075));
inv_hvt I101 ( .A(net075), .Y(net070));
oai21x2_sup_25 I202 ( .A1(yp3_b_low_ysup_25), .Y(yp3_b_25),
     .A0(net069), .B0(yp3_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(net070), .sup(ysup_25),
     .out_vddio_b(yp3_25_b), .out_vddio(net069), .in_b(net075));
inv_25 I204 ( .IN(yp3_25_b), .OUT(yp3_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yp21, View - schematic
// LAST TIME SAVED: Feb 26 14:41:20 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp21 ( yp21, yp21_b_25, yp21_b_low_b, yp21_sel,
     ysup_25 );
output  yp21, yp21_b_25;

input  yp21_b_low_b, yp21_sel, ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I206 ( .A(yp21_sel_b), .Y(net50), .B(yp21_b_low_b));
inv_hvt I207 ( .A(net50), .Y(net68));
inv_hvt I208 ( .A(yp21_sel), .Y(yp21_sel_b));
inv_hvt I209 ( .A(yp21_sel_b), .Y(yp21));
ml_ls_vdd25_nor2 I194 ( .in(net68), .sup(ysup_25),
     .out_vddio_b(yp21_b_25_b), .out_vddio(net72), .in_b(net50));
inv_25 I213 ( .IN(yp21_b_25_b), .OUT(yp21_b_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl, View - schematic
// LAST TIME SAVED: May  4 14:26:38 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl ( yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test_25, yp_test_b_25, vblinhi_pgm_25, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, yp1_b_low_b, yp1_sel, yp2_b_low_b,
     yp2_sel, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, yp_test, yp_test_b_high_b,
     yp_test_b_low_b, ysup_25 );

inout  vblinhi_pgm_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b,
     yp2_b_low_b, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp_test_b_high_b, yp_test_b_low_b, ysup_25;

output [1:0]  yp_test_b_25;
output [5:0]  yp1;
output [5:0]  yp1_b_25;
output [7:0]  yp3_b_25;
output [7:0]  yp2_b_25;
output [7:0]  yp2;
output [7:0]  yp3_25;
output [1:0]  yp_test_25;

input [5:0]  yp1_sel;
input [7:0]  yp2_sel;
input [1:0]  yp_test;
input [7:0]  yp3_sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_1_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1]), .yp_test(yp_test[1]),
     .yp_test_25(yp_test_25[1]));
ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_0_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[0]), .yp_test(yp_test[0]),
     .yp_test_25(yp_test_25[0]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_7_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[7]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[7]), .yp3_25(yp3_25[7]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_6_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[6]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[6]), .yp3_25(yp3_25[6]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_5_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[5]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[5]), .yp3_25(yp3_25[5]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_4_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[4]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[4]), .yp3_25(yp3_25[4]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_3_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[3]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[3]), .yp3_25(yp3_25[3]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_2_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[2]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[2]), .yp3_25(yp3_25[2]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_1_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[1]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[1]), .yp3_25(yp3_25[1]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_0_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[0]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[0]), .yp3_25(yp3_25[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_7_ ( .yp21_sel(yp2_sel[7]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[7]), .yp21(yp2[7]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_6_ ( .yp21_sel(yp2_sel[6]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[6]), .yp21(yp2[6]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_5_ ( .yp21_sel(yp2_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[5]), .yp21(yp2[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_4_ ( .yp21_sel(yp2_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[4]), .yp21(yp2[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_3_ ( .yp21_sel(yp2_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[3]), .yp21(yp2[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_2_ ( .yp21_sel(yp2_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[2]), .yp21(yp2[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_1_ ( .yp21_sel(yp2_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[1]), .yp21(yp2[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_0_ ( .yp21_sel(yp2_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[0]), .yp21(yp2[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_5_ ( .yp21_sel(yp1_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[5]), .yp21(yp1[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_4_ ( .yp21_sel(yp1_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[4]), .yp21(yp1[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_3_ ( .yp21_sel(yp1_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[3]), .yp21(yp1[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_2_ ( .yp21_sel(yp1_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[2]), .yp21(yp1[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_1_ ( .yp21_sel(yp1_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[1]), .yp21(yp1[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_0_ ( .yp21_sel(yp1_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[0]), .yp21(yp1[0]));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_top, View - schematic
// LAST TIME SAVED: May  4 14:26:28 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_ctrl_top ( gwl_b_gnden_25, nv_dataout, yp1, yp1_b_25,
     yp2, yp2_b_25, yp3_25, yp3_b_25, yp_test, yp_test_25,
     yp_test_b_25, bl_out, bl_pgm_glb, s_b_25, s_b_hv, sb25sup_25,
     sbhvsup_hv, vblinhi_pgm_25, vdd_tieh, vpxa, ysup_25, dec_ok_25,
     fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, tm_allbl_h, tm_allbl_l, tm_allwl_h,
     tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr );
output  gwl_b_gnden_25, nv_dataout;

inout  bl_out, bl_pgm_glb, sb25sup_25, sbhvsup_hv, vblinhi_pgm_25,
     vdd_tieh, vpxa, ysup_25;

input  dec_ok_25, fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, saen_25, saen_b_vpxa, testdec_en_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [1:0]  yp_test_b_25;
output [1:0]  yp_test;
output [1:0]  yp_test_25;
output [5:0]  yp1_b_25;
output [7:0]  yp3_25;
output [5:0]  yp1;
output [7:0]  yp2_b_25;
output [7:0]  yp3_b_25;
output [7:0]  yp2;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sb25_gnd_25;

wire  [3:0]  sbhv_gnd_25;

wire  [3:0]  sbhv_high_25;

wire  [3:0]  sb25_high_25;

wire  [7:5]  dec_trim;

wire  [7:0]  yp3_sel;

wire  [7:0]  yp2_sel;

wire  [5:0]  yp1_sel;



inv_25 I38 ( .IN(net293), .OUT(gwl_b_gnden_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I30 ( .IN(fsm_gwlbdis_b_25), .OUT(net293), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_core_ctrl_logic Icore_ctrl_logic ( .yp1_sel(yp1_sel[5:0]),
     .yp2_sel(yp2_sel[7:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_tm_allwl_l(tm_allwl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25), .tm_tcol(tm_tcol),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_allbl_l(tm_allbl_l), .fsm_pgm(fsm_pgm),
     .fsm_tm_allbl_h(tm_allbl_h), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_nvcmen(fsm_nvcmen), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd(fsm_blkadd[3:0]), .yp_test(yp_test[1:0]),
     .yp21_b_low_b(yp21_b_low_b), .yp3_sel(yp3_sel[7:0]),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .sbhv_high_25(sbhv_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sb25_gnd_25(sb25_gnd_25[3:0]),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .dec_trim(dec_trim[7:5]));
vdd_tiehigh I117_9_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_8_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_7_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_6_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_5_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_4_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_3_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_2_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_1_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_0_ ( .vdd_tieh(vdd_tieh));
ml_core_sa_top Icore_sa_top ( .tm_dma(tm_dma),
     .fsm_tm_testdec(fsm_tm_testdec), .tm_testdec_wr(tm_testdec_wr),
     .testdec_en_b_25(testdec_en_b_25), .dec_ok_25(dec_ok_25),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .dec_trim(dec_trim[7:5]),
     .nv_dataout(nv_dataout), .vpxa(vpxa), .bl_pgm_glb(bl_pgm_glb),
     .bl_out(bl_out));
ml_wp_ctrl Iml_wp_ctrl ( .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .sbhv_high_25(sbhv_high_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_gnd_25(sb25_gnd_25[3:0]), .s_b_25(s_b_25[3:0]),
     .s_b_hv(s_b_hv[3:0]));
ml_ymux_ctrl Iml_ymux_ctrl ( .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]),
     .yp1(yp1[5:0]), .yp1_b_25(yp1_b_25[5:0]), .yp2_sel(yp2_sel[7:0]),
     .yp1_sel(yp1_sel[5:0]), .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_sel(yp3_sel[7:0]), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_b_high_b(gnd_),
     .yp_test_b_low_b(gnd_), .yp_test(yp_test[1:0]),
     .yp2_b_low_b(yp21_b_low_b), .yp1_b_low_b(yp21_b_low_b),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .yp_test_25(yp_test_25[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - ROCK, Cell - nvcm_cell_1, View - schematic
// LAST TIME SAVED: May 13 16:00:35 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_1 ( bl, wp, wr );
inout  bl;

input  wp, wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nchx  NR ( .D(net1), .G(wr), .S(bl));
nchx  NP ( .D(net5), .G(wp), .S(net1));

endmodule
// Library - NVCM, Cell - nvcm_cell_2x1, View - schematic
// LAST TIME SAVED: Dec 10 15:56:30 2007
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_2x1 ( bl, wp, wr );

input  wp, wr;

inout [1:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
nvcm_cell_1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));

endmodule
// Library - NVCM, Cell - nvcm_cell_2x8, View - schematic
// LAST TIME SAVED: Feb 26 14:36:29 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_2x8 ( bl, wp, wr );


inout [1:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m7 ( .bl(bl[1:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_2x1 m6 ( .bl(bl[1:0]), .wr(wr[6]), .wp(wp[6]));
nvcm_cell_2x1 m5 ( .bl(bl[1:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_2x1 m4 ( .bl(bl[1:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_2x1 m3 ( .bl(bl[1:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_2x1 m2 ( .bl(bl[1:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM, Cell - nvcm_cell_1x8, View - schematic
// LAST TIME SAVED: Jul  5 11:06:02 2007
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_1x8 ( bl, wp, wr );

input  wp, wr;

inout [7:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
nvcm_cell_1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));
nvcm_cell_1 m2 ( .wp(wp), .wr(wr), .bl(bl[2]));
nvcm_cell_1 m3 ( .wp(wp), .wr(wr), .bl(bl[3]));
nvcm_cell_1 m4 ( .wp(wp), .wr(wr), .bl(bl[4]));
nvcm_cell_1 m5 ( .wp(wp), .wr(wr), .bl(bl[5]));
nvcm_cell_1 m6 ( .wp(wp), .wr(wr), .bl(bl[6]));
nvcm_cell_1 m7 ( .wp(wp), .wr(wr), .bl(bl[7]));

endmodule
// Library - NVCM, Cell - nvcm_cell_8x8, View - schematic
// LAST TIME SAVED: Dec 10 15:35:50 2007
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_8x8 ( bl, wp, wr );


inout [7:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 m0 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 m1 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 m2 ( .bl(bl[7:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_1x8 m3 ( .bl(bl[7:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_1x8 m7 ( .bl(bl[7:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_1x8 m4 ( .bl(bl[7:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_1x8 m5 ( .bl(bl[7:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_1x8 m6 ( .bl(bl[7:0]), .wr(wr[6]), .wp(wp[6]));

endmodule
// Library - NVCM, Cell - nvcm_cell_16x8, View - schematic
// LAST TIME SAVED: Dec 10 15:41:25 2007
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_16x8 ( bl, wp, wr );


inout [15:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_8x8 m0 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[7:0]));
nvcm_cell_8x8 m1 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[15:8]));

endmodule
// Library - xpmem, Cell - ml_rowdrv2_last, View - schematic
// LAST TIME SAVED: Sep 26 14:07:07 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_rowdrv2_last ( pgate, reset, smc_rsr_out, vddctrl, wl,
     wl_rd_sup, wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write
     );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  NM0 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
ml_dff_schematic I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));

endmodule
// Library - NVCM, Cell - nvcm_cell_336x8, View - schematic
// LAST TIME SAVED: Feb 26 14:32:20 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_336x8 ( bl, bl_dummyl, bl_dummyr, bl_test, wp, wr );


inout [1:0]  bl_test;
inout [327:0]  bl;
inout [1:0]  bl_dummyl;
inout [5:0]  bl_dummyr;

input [7:0]  wp;
input [7:0]  wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x8 Invcm_cell_2x8 ( .wp(wp[7:0]), .wr(wr[7:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_16x8 Invcm_cell_16x8_19_ ( .wp(wp[7:0]), .bl(bl[319:304]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_18_ ( .wp(wp[7:0]), .bl(bl[303:288]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_17_ ( .wp(wp[7:0]), .bl(bl[287:272]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_16_ ( .wp(wp[7:0]), .bl(bl[271:256]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_15_ ( .wp(wp[7:0]), .bl(bl[255:240]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_14_ ( .wp(wp[7:0]), .bl(bl[239:224]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_13_ ( .wp(wp[7:0]), .bl(bl[223:208]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_12_ ( .wp(wp[7:0]), .bl(bl[207:192]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_11_ ( .wp(wp[7:0]), .bl(bl[191:176]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_10_ ( .wp(wp[7:0]), .bl(bl[175:160]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_9_ ( .wp(wp[7:0]), .bl(bl[159:144]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_8_ ( .wp(wp[7:0]), .bl(bl[143:128]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_7_ ( .wp(wp[7:0]), .bl(bl[127:112]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_6_ ( .wp(wp[7:0]), .bl(bl[111:96]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_5_ ( .wp(wp[7:0]), .bl(bl[95:80]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_4_ ( .wp(wp[7:0]), .bl(bl[79:64]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_3_ ( .wp(wp[7:0]), .bl(bl[63:48]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_2_ ( .wp(wp[7:0]), .bl(bl[47:32]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_1_ ( .wp(wp[7:0]), .bl(bl[31:16]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_0_ ( .wp(wp[7:0]), .bl(bl[15:0]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_20_ ( .wp(wp[7:0]), .bl({bl_dummyr[5:0],
     bl_test[1:0], bl[327:320]}), .wr(wr[7:0]));

endmodule
// Library - NVCM, Cell - nvcm_cell_338x232, View - schematic
// LAST TIME SAVED: Feb 26 14:32:01 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module nvcm_cell_338x232 ( bl, bl_dummyl, bl_dummyr, bl_test, wp,
     wp_dummyb, wp_dummyt, wr, wr_dummyb, wr_dummyt );


inout [327:0]  bl;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;

input [1:0]  wr_dummyb;
input [227:0]  wp;
input [1:0]  wr_dummyt;
input [1:0]  wp_dummyb;
input [1:0]  wp_dummyt;
input [227:0]  wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_336x8 Invcm_cell_336x8_26_ ( .wr(wr[221:214]),
     .wp(wp[221:214]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_25_ ( .wr(wr[213:206]),
     .wp(wp[213:206]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_24_ ( .wr(wr[205:198]),
     .wp(wp[205:198]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_23_ ( .wr(wr[197:190]),
     .wp(wp[197:190]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_22_ ( .wr(wr[189:182]),
     .wp(wp[189:182]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_21_ ( .wr(wr[181:174]),
     .wp(wp[181:174]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_20_ ( .wr(wr[173:166]),
     .wp(wp[173:166]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_19_ ( .wr(wr[165:158]),
     .wp(wp[165:158]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_18_ ( .wr(wr[157:150]),
     .wp(wp[157:150]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_17_ ( .wr(wr[149:142]),
     .wp(wp[149:142]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_16_ ( .wr(wr[141:134]),
     .wp(wp[141:134]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_15_ ( .wr(wr[133:126]),
     .wp(wp[133:126]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_14_ ( .wr(wr[125:118]),
     .wp(wp[125:118]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_13_ ( .wr(wr[117:110]),
     .wp(wp[117:110]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_12_ ( .wr(wr[109:102]),
     .wp(wp[109:102]), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_11_ ( .wr(wr[101:94]),
     .wp(wp[101:94]), .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0]}), .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_10_ ( .wr(wr[93:86]), .wp(wp[93:86]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_9_ ( .wr(wr[85:78]), .wp(wp[85:78]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_8_ ( .wr(wr[77:70]), .wp(wp[77:70]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_7_ ( .wr(wr[69:62]), .wp(wp[69:62]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_6_ ( .wr(wr[61:54]), .wp(wp[61:54]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_5_ ( .wr(wr[53:46]), .wp(wp[53:46]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_4_ ( .wr(wr[45:38]), .wp(wp[45:38]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_3_ ( .wr(wr[37:30]), .wp(wp[37:30]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_2_ ( .wr(wr[29:22]), .wp(wp[29:22]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_1_ ( .wr(wr[21:14]), .wp(wp[21:14]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_0_ ( .wr(wr[13:6]), .wp(wp[13:6]),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_t ( .wr({wr[5:0], wr_dummyt[1:0]}),
     .wp({wp[5:0], wp_dummyt[1:0]}), .bl_test(bl_test[1:0]),
     .bl_dummyr({bl_dummyr[1], bl_dummyr[0], bl_dummyr[1],
     bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
nvcm_cell_336x8 Invcm_cell_336x8_b ( .wr({wr_dummyb[1:0],
     wr[227:222]}), .wp({wp_dummyb[1:0], wp[227:222]}),
     .bl_test(bl_test[1:0]), .bl_dummyr({bl_dummyr[1], bl_dummyr[0],
     bl_dummyr[1], bl_dummyr[0], bl_dummyr[1], bl_dummyr[0]}),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));

endmodule
// Library - NVCM, Cell - ml_testdec_bgen, View - schematic
// LAST TIME SAVED: Jan 21 10:19:00 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_testdec_bgen ( dec_ok_25, dec_bias_25, dec_det_25,
     testdec_en_b_25, testdec_prec_b_25 );
output  dec_ok_25;

inout  dec_bias_25, dec_det_25;

input  testdec_en_b_25, testdec_prec_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I38 ( .IN(dec_det_25), .OUT(dec_ok_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M23 ( .D(dec_det_25), .B(vddp_), .G(testdec_prec_b_25),
     .S(vddp_));
pch_25  M18_1_ ( .D(dec_bias_sup), .B(vddp_), .G(testdec_en_b_25),
     .S(vddp_));
pch_25  M18_0_ ( .D(dec_bias_sup), .B(vddp_), .G(testdec_en_b_25),
     .S(vddp_));
pch_25  M16 ( .D(net049), .B(vddp_), .G(testdec_en_b_25), .S(vddp_));
pch_25  M19 ( .D(ngate), .B(vddp_), .G(dec_bias_25), .S(net049));
pch_25  M8 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
pch_25  M9_1_ ( .D(dec_det_25), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
pch_25  M9_0_ ( .D(dec_det_25), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
nch_25  M14 ( .D(ngate), .B(GND_), .G(dec_bias_25), .S(gnd_));
nch_25  M15 ( .D(ngate), .B(GND_), .G(testdec_en_b_25), .S(gnd_));
nch_25  M10 ( .D(dec_bias_sup), .B(GND_), .G(ngate), .S(dec_bias_25));
nch_25  M13 ( .D(dec_bias_25), .B(GND_), .G(testdec_en_b_25),
     .S(gnd_));
nch_25  M4 ( .D(dec_det_25), .B(GND_), .G(testdec_en_b_25), .S(gnd_));
nch_25  M17 ( .D(dec_bias_25), .B(GND_), .G(dec_bias_25), .S(gnd_));
nch_25  M20 ( .D(dec_bias_p), .B(GND_), .G(dec_bias_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_testdec_rows, View - schematic
// LAST TIME SAVED: Feb 26 14:35:11 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_testdec_rows ( dec_bias, dec_det_25, vddp_tieh, wp, wr );
inout  dec_bias, dec_det_25;

input  vddp_tieh, wp, wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(dec_det_25), .B(GND_), .G(wr), .S(gnd_));
nch_25  M12 ( .D(net20), .B(gnd_), .G(vddp_tieh), .S(wp));
nch_25  M2 ( .D(dec_det_25), .B(GND_), .G(net20), .S(gnd_));
nch_25  M0 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(net20));
nch_25  M1 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(wr));

endmodule
// Library - NVCM, Cell - ml_testdec_rowsx228, View - schematic
// LAST TIME SAVED: Feb 26 14:34:58 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_testdec_rowsx228 ( dec_det_even_25, dec_det_odd_25,
     dec_bias_25, dec_det_25, testdec_even_b_25, testdec_odd_b_25, wp,
     wr );
output  dec_det_even_25, dec_det_odd_25;

inout  dec_bias_25, dec_det_25;

input  testdec_even_b_25, testdec_odd_b_25;

input [227:0]  wr;
input [227:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I25 ( .vddp_tieh(vddp_tiel));
nor2_25 I24 ( .A(testdec_odd_b_25), .Y(dec_det_odd_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
nor2_25 I59 ( .A(testdec_even_b_25), .Y(dec_det_even_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
ml_testdec_rows Itestdec_rows_227_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[227]), .wp(wp[227]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_226_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[226]), .wp(wp[226]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_225_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[225]), .wp(wp[225]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_224_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[224]), .wp(wp[224]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_223_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[223]), .wp(wp[223]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_222_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[222]), .wp(wp[222]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_221_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[221]), .wp(wp[221]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_220_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[220]), .wp(wp[220]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_219_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[219]), .wp(wp[219]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_218_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[218]), .wp(wp[218]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_217_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[217]), .wp(wp[217]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_216_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[216]), .wp(wp[216]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_215_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[215]), .wp(wp[215]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_214_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[214]), .wp(wp[214]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_213_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[213]), .wp(wp[213]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_212_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[212]), .wp(wp[212]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_211_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[211]), .wp(wp[211]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_210_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[210]), .wp(wp[210]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_209_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[209]), .wp(wp[209]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_208_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[208]), .wp(wp[208]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_207_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[207]), .wp(wp[207]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_206_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[206]), .wp(wp[206]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_205_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[205]), .wp(wp[205]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_204_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[204]), .wp(wp[204]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_203_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[203]), .wp(wp[203]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_202_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[202]), .wp(wp[202]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_201_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[201]), .wp(wp[201]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_200_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[200]), .wp(wp[200]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_199_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[199]), .wp(wp[199]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_198_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[198]), .wp(wp[198]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_197_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[197]), .wp(wp[197]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_196_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[196]), .wp(wp[196]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_195_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[195]), .wp(wp[195]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_194_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[194]), .wp(wp[194]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_193_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[193]), .wp(wp[193]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_192_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[192]), .wp(wp[192]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_191_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[191]), .wp(wp[191]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_190_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[190]), .wp(wp[190]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_189_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[189]), .wp(wp[189]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_188_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[188]), .wp(wp[188]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_187_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[187]), .wp(wp[187]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_186_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[186]), .wp(wp[186]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_185_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[185]), .wp(wp[185]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_184_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[184]), .wp(wp[184]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_183_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[183]), .wp(wp[183]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_182_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[182]), .wp(wp[182]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_181_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[181]), .wp(wp[181]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_180_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[180]), .wp(wp[180]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_179_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[179]), .wp(wp[179]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_178_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[178]), .wp(wp[178]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_177_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[177]), .wp(wp[177]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_176_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[176]), .wp(wp[176]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_175_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[175]), .wp(wp[175]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_174_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[174]), .wp(wp[174]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_173_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[173]), .wp(wp[173]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_172_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[172]), .wp(wp[172]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_171_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[171]), .wp(wp[171]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_170_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[170]), .wp(wp[170]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_169_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[169]), .wp(wp[169]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_168_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[168]), .wp(wp[168]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_167_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[167]), .wp(wp[167]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_166_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[166]), .wp(wp[166]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_165_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[165]), .wp(wp[165]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_164_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[164]), .wp(wp[164]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_163_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[163]), .wp(wp[163]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_162_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[162]), .wp(wp[162]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_161_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[161]), .wp(wp[161]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_160_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[160]), .wp(wp[160]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_159_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[159]), .wp(wp[159]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_158_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[158]), .wp(wp[158]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_157_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[157]), .wp(wp[157]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_156_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[156]), .wp(wp[156]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_155_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[155]), .wp(wp[155]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_154_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[154]), .wp(wp[154]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_153_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[153]), .wp(wp[153]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_152_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[152]), .wp(wp[152]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_151_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[151]), .wp(wp[151]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_150_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[150]), .wp(wp[150]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_149_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[149]), .wp(wp[149]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_148_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[148]), .wp(wp[148]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_147_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[147]), .wp(wp[147]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_146_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[146]), .wp(wp[146]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_145_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[145]), .wp(wp[145]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_144_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[144]), .wp(wp[144]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_143_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[143]), .wp(wp[143]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_142_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[142]), .wp(wp[142]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_141_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[141]), .wp(wp[141]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_140_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[140]), .wp(wp[140]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_139_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[139]), .wp(wp[139]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_138_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[138]), .wp(wp[138]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_137_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[137]), .wp(wp[137]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_136_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[136]), .wp(wp[136]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_135_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[135]), .wp(wp[135]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_134_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[134]), .wp(wp[134]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_133_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[133]), .wp(wp[133]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_132_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[132]), .wp(wp[132]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_131_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[131]), .wp(wp[131]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_130_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[130]), .wp(wp[130]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_129_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[129]), .wp(wp[129]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_128_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[128]), .wp(wp[128]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_127_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[127]), .wp(wp[127]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_126_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[126]), .wp(wp[126]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_125_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[125]), .wp(wp[125]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_124_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[124]), .wp(wp[124]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_123_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[123]), .wp(wp[123]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_122_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[122]), .wp(wp[122]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_121_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[121]), .wp(wp[121]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_120_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[120]), .wp(wp[120]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_119_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[119]), .wp(wp[119]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_118_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[118]), .wp(wp[118]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_117_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[117]), .wp(wp[117]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_116_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[116]), .wp(wp[116]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_115_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[115]), .wp(wp[115]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_114_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[114]), .wp(wp[114]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_113_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[113]), .wp(wp[113]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_112_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[112]), .wp(wp[112]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_111_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[111]), .wp(wp[111]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_110_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[110]), .wp(wp[110]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_109_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[109]), .wp(wp[109]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_108_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[108]), .wp(wp[108]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_107_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[107]), .wp(wp[107]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_106_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[106]), .wp(wp[106]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_105_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[105]), .wp(wp[105]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_104_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[104]), .wp(wp[104]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_103_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[103]), .wp(wp[103]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_102_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[102]), .wp(wp[102]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_101_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[101]), .wp(wp[101]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_100_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[100]), .wp(wp[100]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_99_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[99]), .wp(wp[99]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_98_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[98]), .wp(wp[98]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_97_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[97]), .wp(wp[97]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_96_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[96]), .wp(wp[96]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_95_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[95]), .wp(wp[95]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_94_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[94]), .wp(wp[94]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_93_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[93]), .wp(wp[93]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_92_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[92]), .wp(wp[92]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_91_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[91]), .wp(wp[91]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_90_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[90]), .wp(wp[90]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_89_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[89]), .wp(wp[89]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_88_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[88]), .wp(wp[88]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_87_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[87]), .wp(wp[87]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_86_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[86]), .wp(wp[86]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_85_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[85]), .wp(wp[85]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_84_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[84]), .wp(wp[84]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_83_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[83]), .wp(wp[83]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_82_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[82]), .wp(wp[82]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_81_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[81]), .wp(wp[81]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_80_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[80]), .wp(wp[80]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_79_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[79]), .wp(wp[79]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_78_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[78]), .wp(wp[78]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_77_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[77]), .wp(wp[77]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_76_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[76]), .wp(wp[76]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_75_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[75]), .wp(wp[75]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_74_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[74]), .wp(wp[74]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_73_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[73]), .wp(wp[73]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_72_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[72]), .wp(wp[72]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_71_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[71]), .wp(wp[71]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_70_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[70]), .wp(wp[70]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_69_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[69]), .wp(wp[69]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_68_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[68]), .wp(wp[68]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_67_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[67]), .wp(wp[67]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_66_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[66]), .wp(wp[66]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_65_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[65]), .wp(wp[65]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_64_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[64]), .wp(wp[64]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_63_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[63]), .wp(wp[63]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_62_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[62]), .wp(wp[62]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_61_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[61]), .wp(wp[61]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_60_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[60]), .wp(wp[60]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_59_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[59]), .wp(wp[59]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_58_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[58]), .wp(wp[58]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_57_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[57]), .wp(wp[57]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_56_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[56]), .wp(wp[56]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_55_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[55]), .wp(wp[55]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_54_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[54]), .wp(wp[54]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_53_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[53]), .wp(wp[53]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_52_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[52]), .wp(wp[52]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_51_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[51]), .wp(wp[51]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_50_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[50]), .wp(wp[50]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_49_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[49]), .wp(wp[49]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_48_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[48]), .wp(wp[48]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_47_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[47]), .wp(wp[47]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_46_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[46]), .wp(wp[46]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_45_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[45]), .wp(wp[45]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_44_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[44]), .wp(wp[44]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_43_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[43]), .wp(wp[43]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_42_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[42]), .wp(wp[42]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_41_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[41]), .wp(wp[41]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_40_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[40]), .wp(wp[40]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_39_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[39]), .wp(wp[39]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_38_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[38]), .wp(wp[38]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_37_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[37]), .wp(wp[37]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_36_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[36]), .wp(wp[36]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_35_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[35]), .wp(wp[35]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_34_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[34]), .wp(wp[34]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_33_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[33]), .wp(wp[33]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_32_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[32]), .wp(wp[32]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_31_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[31]), .wp(wp[31]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_30_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[30]), .wp(wp[30]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_29_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[29]), .wp(wp[29]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_28_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[28]), .wp(wp[28]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_27_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[27]), .wp(wp[27]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_26_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[26]), .wp(wp[26]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_25_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[25]), .wp(wp[25]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_24_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[24]), .wp(wp[24]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_23_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[23]), .wp(wp[23]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_22_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[22]), .wp(wp[22]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_21_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[21]), .wp(wp[21]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_20_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[20]), .wp(wp[20]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_19_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[19]), .wp(wp[19]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_18_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[18]), .wp(wp[18]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_17_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[17]), .wp(wp[17]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_16_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[16]), .wp(wp[16]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_15_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[15]), .wp(wp[15]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_14_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[14]), .wp(wp[14]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_13_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[13]), .wp(wp[13]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_12_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[12]), .wp(wp[12]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_11_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[11]), .wp(wp[11]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_10_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[10]), .wp(wp[10]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_9_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[9]), .wp(wp[9]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_8_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[8]), .wp(wp[8]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_7_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[7]), .wp(wp[7]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_6_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[6]), .wp(wp[6]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_5_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[5]), .wp(wp[5]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_4_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[4]), .wp(wp[4]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_3_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[3]), .wp(wp[3]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_2_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[2]), .wp(wp[2]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_1_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[1]), .wp(wp[1]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_0_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[0]), .wp(wp[0]),
     .dec_bias(dec_bias_25));

endmodule
// Library - NVCM, Cell - ml_testdec_columns, View - schematic
// LAST TIME SAVED: Feb 26 14:35:47 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_testdec_columns ( bl, dec_det_even_25, dec_det_odd_25 );

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(vdd_), .B(gnd_), .G(dec_det_even_25), .S(bl[0]));
nch_25  M4 ( .D(vdd_), .B(gnd_), .G(dec_det_odd_25), .S(bl[1]));

endmodule
// Library - NVCM, Cell - ml_testdec_columnsx330, View - schematic
// LAST TIME SAVED: Feb 26 14:35:34 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_testdec_columnsx330 ( bl, bl_dummyl, bl_dummyr, bl_test,
     dec_det_even_25, dec_det_odd_25 );

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl_dummyl;
inout [327:0]  bl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_testdec_columns Itestdec_columns_dml (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyl[1:0]));
ml_testdec_columns Itestdec_columns_163_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[327:326]));
ml_testdec_columns Itestdec_columns_162_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[325:324]));
ml_testdec_columns Itestdec_columns_161_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[323:322]));
ml_testdec_columns Itestdec_columns_160_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[321:320]));
ml_testdec_columns Itestdec_columns_159_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[319:318]));
ml_testdec_columns Itestdec_columns_158_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[317:316]));
ml_testdec_columns Itestdec_columns_157_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[315:314]));
ml_testdec_columns Itestdec_columns_156_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[313:312]));
ml_testdec_columns Itestdec_columns_155_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[311:310]));
ml_testdec_columns Itestdec_columns_154_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[309:308]));
ml_testdec_columns Itestdec_columns_153_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[307:306]));
ml_testdec_columns Itestdec_columns_152_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[305:304]));
ml_testdec_columns Itestdec_columns_151_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[303:302]));
ml_testdec_columns Itestdec_columns_150_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[301:300]));
ml_testdec_columns Itestdec_columns_149_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[299:298]));
ml_testdec_columns Itestdec_columns_148_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[297:296]));
ml_testdec_columns Itestdec_columns_147_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[295:294]));
ml_testdec_columns Itestdec_columns_146_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[293:292]));
ml_testdec_columns Itestdec_columns_145_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[291:290]));
ml_testdec_columns Itestdec_columns_144_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[289:288]));
ml_testdec_columns Itestdec_columns_143_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[287:286]));
ml_testdec_columns Itestdec_columns_142_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[285:284]));
ml_testdec_columns Itestdec_columns_141_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[283:282]));
ml_testdec_columns Itestdec_columns_140_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[281:280]));
ml_testdec_columns Itestdec_columns_139_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[279:278]));
ml_testdec_columns Itestdec_columns_138_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[277:276]));
ml_testdec_columns Itestdec_columns_137_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[275:274]));
ml_testdec_columns Itestdec_columns_136_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[273:272]));
ml_testdec_columns Itestdec_columns_135_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[271:270]));
ml_testdec_columns Itestdec_columns_134_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[269:268]));
ml_testdec_columns Itestdec_columns_133_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[267:266]));
ml_testdec_columns Itestdec_columns_132_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[265:264]));
ml_testdec_columns Itestdec_columns_131_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[263:262]));
ml_testdec_columns Itestdec_columns_130_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[261:260]));
ml_testdec_columns Itestdec_columns_129_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[259:258]));
ml_testdec_columns Itestdec_columns_128_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[257:256]));
ml_testdec_columns Itestdec_columns_127_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[255:254]));
ml_testdec_columns Itestdec_columns_126_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[253:252]));
ml_testdec_columns Itestdec_columns_125_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[251:250]));
ml_testdec_columns Itestdec_columns_124_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[249:248]));
ml_testdec_columns Itestdec_columns_123_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[247:246]));
ml_testdec_columns Itestdec_columns_122_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[245:244]));
ml_testdec_columns Itestdec_columns_121_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[243:242]));
ml_testdec_columns Itestdec_columns_120_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[241:240]));
ml_testdec_columns Itestdec_columns_119_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[239:238]));
ml_testdec_columns Itestdec_columns_118_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[237:236]));
ml_testdec_columns Itestdec_columns_117_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[235:234]));
ml_testdec_columns Itestdec_columns_116_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[233:232]));
ml_testdec_columns Itestdec_columns_115_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[231:230]));
ml_testdec_columns Itestdec_columns_114_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[229:228]));
ml_testdec_columns Itestdec_columns_113_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[227:226]));
ml_testdec_columns Itestdec_columns_112_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[225:224]));
ml_testdec_columns Itestdec_columns_111_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[223:222]));
ml_testdec_columns Itestdec_columns_110_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[221:220]));
ml_testdec_columns Itestdec_columns_109_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[219:218]));
ml_testdec_columns Itestdec_columns_108_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[217:216]));
ml_testdec_columns Itestdec_columns_107_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[215:214]));
ml_testdec_columns Itestdec_columns_106_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[213:212]));
ml_testdec_columns Itestdec_columns_105_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[211:210]));
ml_testdec_columns Itestdec_columns_104_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[209:208]));
ml_testdec_columns Itestdec_columns_103_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[207:206]));
ml_testdec_columns Itestdec_columns_102_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[205:204]));
ml_testdec_columns Itestdec_columns_101_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[203:202]));
ml_testdec_columns Itestdec_columns_100_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[201:200]));
ml_testdec_columns Itestdec_columns_99_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[199:198]));
ml_testdec_columns Itestdec_columns_98_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[197:196]));
ml_testdec_columns Itestdec_columns_97_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[195:194]));
ml_testdec_columns Itestdec_columns_96_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[193:192]));
ml_testdec_columns Itestdec_columns_95_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[191:190]));
ml_testdec_columns Itestdec_columns_94_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[189:188]));
ml_testdec_columns Itestdec_columns_93_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[187:186]));
ml_testdec_columns Itestdec_columns_92_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[185:184]));
ml_testdec_columns Itestdec_columns_91_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[183:182]));
ml_testdec_columns Itestdec_columns_90_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[181:180]));
ml_testdec_columns Itestdec_columns_89_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[179:178]));
ml_testdec_columns Itestdec_columns_88_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[177:176]));
ml_testdec_columns Itestdec_columns_87_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[175:174]));
ml_testdec_columns Itestdec_columns_86_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[173:172]));
ml_testdec_columns Itestdec_columns_85_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[171:170]));
ml_testdec_columns Itestdec_columns_84_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[169:168]));
ml_testdec_columns Itestdec_columns_83_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[167:166]));
ml_testdec_columns Itestdec_columns_82_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[165:164]));
ml_testdec_columns Itestdec_columns_81_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[163:162]));
ml_testdec_columns Itestdec_columns_80_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[161:160]));
ml_testdec_columns Itestdec_columns_79_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[159:158]));
ml_testdec_columns Itestdec_columns_78_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[157:156]));
ml_testdec_columns Itestdec_columns_77_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[155:154]));
ml_testdec_columns Itestdec_columns_76_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[153:152]));
ml_testdec_columns Itestdec_columns_75_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[151:150]));
ml_testdec_columns Itestdec_columns_74_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[149:148]));
ml_testdec_columns Itestdec_columns_73_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[147:146]));
ml_testdec_columns Itestdec_columns_72_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[145:144]));
ml_testdec_columns Itestdec_columns_71_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[143:142]));
ml_testdec_columns Itestdec_columns_70_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[141:140]));
ml_testdec_columns Itestdec_columns_69_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[139:138]));
ml_testdec_columns Itestdec_columns_68_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[137:136]));
ml_testdec_columns Itestdec_columns_67_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[135:134]));
ml_testdec_columns Itestdec_columns_66_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[133:132]));
ml_testdec_columns Itestdec_columns_65_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[131:130]));
ml_testdec_columns Itestdec_columns_64_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[129:128]));
ml_testdec_columns Itestdec_columns_63_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[127:126]));
ml_testdec_columns Itestdec_columns_62_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[125:124]));
ml_testdec_columns Itestdec_columns_61_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[123:122]));
ml_testdec_columns Itestdec_columns_60_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[121:120]));
ml_testdec_columns Itestdec_columns_59_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[119:118]));
ml_testdec_columns Itestdec_columns_58_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[117:116]));
ml_testdec_columns Itestdec_columns_57_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[115:114]));
ml_testdec_columns Itestdec_columns_56_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[113:112]));
ml_testdec_columns Itestdec_columns_55_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[111:110]));
ml_testdec_columns Itestdec_columns_54_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[109:108]));
ml_testdec_columns Itestdec_columns_53_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[107:106]));
ml_testdec_columns Itestdec_columns_52_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[105:104]));
ml_testdec_columns Itestdec_columns_51_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[103:102]));
ml_testdec_columns Itestdec_columns_50_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[101:100]));
ml_testdec_columns Itestdec_columns_49_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[99:98]));
ml_testdec_columns Itestdec_columns_48_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[97:96]));
ml_testdec_columns Itestdec_columns_47_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[95:94]));
ml_testdec_columns Itestdec_columns_46_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[93:92]));
ml_testdec_columns Itestdec_columns_45_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[91:90]));
ml_testdec_columns Itestdec_columns_44_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[89:88]));
ml_testdec_columns Itestdec_columns_43_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[87:86]));
ml_testdec_columns Itestdec_columns_42_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[85:84]));
ml_testdec_columns Itestdec_columns_41_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[83:82]));
ml_testdec_columns Itestdec_columns_40_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[81:80]));
ml_testdec_columns Itestdec_columns_39_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[79:78]));
ml_testdec_columns Itestdec_columns_38_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[77:76]));
ml_testdec_columns Itestdec_columns_37_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[75:74]));
ml_testdec_columns Itestdec_columns_36_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[73:72]));
ml_testdec_columns Itestdec_columns_35_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[71:70]));
ml_testdec_columns Itestdec_columns_34_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[69:68]));
ml_testdec_columns Itestdec_columns_33_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[67:66]));
ml_testdec_columns Itestdec_columns_32_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[65:64]));
ml_testdec_columns Itestdec_columns_31_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[63:62]));
ml_testdec_columns Itestdec_columns_30_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[61:60]));
ml_testdec_columns Itestdec_columns_29_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[59:58]));
ml_testdec_columns Itestdec_columns_28_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[57:56]));
ml_testdec_columns Itestdec_columns_27_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[55:54]));
ml_testdec_columns Itestdec_columns_26_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[53:52]));
ml_testdec_columns Itestdec_columns_25_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[51:50]));
ml_testdec_columns Itestdec_columns_24_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[49:48]));
ml_testdec_columns Itestdec_columns_23_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[47:46]));
ml_testdec_columns Itestdec_columns_22_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[45:44]));
ml_testdec_columns Itestdec_columns_21_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[43:42]));
ml_testdec_columns Itestdec_columns_20_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[41:40]));
ml_testdec_columns Itestdec_columns_19_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[39:38]));
ml_testdec_columns Itestdec_columns_18_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[37:36]));
ml_testdec_columns Itestdec_columns_17_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[35:34]));
ml_testdec_columns Itestdec_columns_16_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[33:32]));
ml_testdec_columns Itestdec_columns_15_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[31:30]));
ml_testdec_columns Itestdec_columns_14_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[29:28]));
ml_testdec_columns Itestdec_columns_13_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[27:26]));
ml_testdec_columns Itestdec_columns_12_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[25:24]));
ml_testdec_columns Itestdec_columns_11_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[23:22]));
ml_testdec_columns Itestdec_columns_10_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[21:20]));
ml_testdec_columns Itestdec_columns_9_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[19:18]));
ml_testdec_columns Itestdec_columns_8_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[17:16]));
ml_testdec_columns Itestdec_columns_7_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[15:14]));
ml_testdec_columns Itestdec_columns_6_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[13:12]));
ml_testdec_columns Itestdec_columns_5_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[11:10]));
ml_testdec_columns Itestdec_columns_4_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[9:8]));
ml_testdec_columns Itestdec_columns_3_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[7:6]));
ml_testdec_columns Itestdec_columns_2_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[5:4]));
ml_testdec_columns Itestdec_columns_1_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[3:2]));
ml_testdec_columns Itestdec_columns_0_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[1:0]));
ml_testdec_columns Itestdec_columns_dmr (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyr[1:0]));
ml_testdec_columns Itestdec_columns_tst (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_test[1:0]));

endmodule
// Library - NVCM, Cell - ml_ymux_yp3_x8, View - schematic
// LAST TIME SAVED: Feb 26 14:33:55 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_yp3_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M5_7_ ( .D(bl[7]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_6_ ( .D(bl[6]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_5_ ( .D(bl[5]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_4_ ( .D(bl[4]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_3_ ( .D(bl[3]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_2_ ( .D(bl[2]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_1_ ( .D(bl[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_0_ ( .D(bl[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
nch_25  M22 ( .D(bl[6]), .B(GND_), .G(yp3_25[6]), .S(bl_out));
nch_25  M1 ( .D(bl[4]), .B(GND_), .G(yp3_25[4]), .S(bl_out));
nch_25  M24 ( .D(bl[2]), .B(GND_), .G(yp3_25[2]), .S(bl_out));
nch_25  M25 ( .D(bl[0]), .B(GND_), .G(yp3_25[0]), .S(bl_out));
nch_25  M26 ( .D(bl[0]), .B(GND_), .G(yp3_b_25[0]), .S(vblinhi_rde));
nch_25  M27 ( .D(bl[1]), .B(GND_), .G(yp3_b_25[1]), .S(vblinhi_rdo));
nch_25  M28 ( .D(bl[1]), .B(GND_), .G(yp3_25[1]), .S(bl_out));
nch_25  M29 ( .D(bl[3]), .B(GND_), .G(yp3_b_25[3]), .S(vblinhi_rdo));
nch_25  M30 ( .D(bl[3]), .B(GND_), .G(yp3_25[3]), .S(bl_out));
nch_25  M31 ( .D(bl[2]), .B(GND_), .G(yp3_b_25[2]), .S(vblinhi_rde));
nch_25  M20 ( .D(bl[4]), .B(GND_), .G(yp3_b_25[4]), .S(vblinhi_rde));
nch_25  M19 ( .D(bl[5]), .B(GND_), .G(yp3_b_25[5]), .S(vblinhi_rdo));
nch_25  M21 ( .D(bl[5]), .B(GND_), .G(yp3_25[5]), .S(bl_out));
nch_25  M13 ( .D(bl[7]), .B(GND_), .G(yp3_b_25[7]), .S(vblinhi_rdo));
nch_25  M23 ( .D(bl[7]), .B(GND_), .G(yp3_25[7]), .S(bl_out));
nch_25  M18 ( .D(bl[6]), .B(GND_), .G(yp3_b_25[6]), .S(vblinhi_rde));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x8, View - schematic
// LAST TIME SAVED: May  4 13:03:21 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_dummy, View - schematic
// LAST TIME SAVED: Feb 26 14:34:35 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_dummy ( bl_dummyr, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, pgminhi_dmmy_b_25, vdd_tieh );
inout  vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo;

input  pgminhi_dmmy_b_25, vdd_tieh;

inout [1:0]  bl_dummyr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(bl_dummyr[1]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rdo));
nch_25  M18 ( .D(bl_dummyr[0]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rde));
pch_25  M8 ( .D(bl_dummyr[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M0 ( .D(bl_dummyr[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));

endmodule
// Library - xpmem, Cell - ml_rowdrvsup2, View - schematic
// LAST TIME SAVED: Aug 28 14:20:28 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_rowdrvsup2 ( wl_rd_sup, wl_rden_b );
inout  wl_rd_sup, wl_rden_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



tielo I223 ( .tielo(net059));
rppolywo_m  R10 ( .MINUS(net045), .PLUS(net0110), .BULK(gnd_));
rppolywo_m  R14 ( .MINUS(wl_rd_sup), .PLUS(net0113), .BULK(gnd_));
rppolywo_m  R12 ( .MINUS(net0104), .PLUS(wl_rd_sup), .BULK(gnd_));
rppolywo_m  R13 ( .MINUS(net0107), .PLUS(net0108), .BULK(gnd_));
rppolywo_m  R11 ( .MINUS(net0110), .PLUS(net0104), .BULK(gnd_));
rppolywo_m  R15 ( .MINUS(net0113), .PLUS(net0107), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net071), .PLUS(net077), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net0108), .PLUS(net071), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(net077), .PLUS(net083), .BULK(gnd_));
rppolywo_m  R19 ( .MINUS(net080), .PLUS(net092), .BULK(gnd_));
rppolywo_m  R20 ( .MINUS(net083), .PLUS(net086), .BULK(gnd_));
rppolywo_m  R21 ( .MINUS(net086), .PLUS(net080), .BULK(gnd_));
rppolywo_m  R22 ( .MINUS(net089), .PLUS(net095), .BULK(gnd_));
rppolywo_m  R23 ( .MINUS(net092), .PLUS(net089), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(net095), .PLUS(net0158), .BULK(gnd_));
inv_hvt I217 ( .A(wl_rden_b), .Y(net0142));
inv_hvt I220 ( .A(net0142), .Y(act_rd_b));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
nch_hvt  MN16 ( .D(wl_rd_sup), .B(gnd_), .G(act_rd_b), .S(gnd_));
nch_hvt  MN14 ( .D(net0158), .B(gnd_), .G(act_rd), .S(gnd_));
pch_hvt  MP13 ( .D(wl_rden_b), .B(vdd_), .G(net059), .S(vdd_));
pch_hvt  MP15 ( .D(net045), .B(vdd_), .G(act_rd_b), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_ymux_yp2_8, View - schematic
// LAST TIME SAVED: Jan 16 10:38:35 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_yp2_8 ( bl, bl_out, vblinhi_rde, vblinhi_rdo, yp2,
     yp2_b_25 );
inout  bl_out, vblinhi_rde, vblinhi_rdo;


inout [7:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M17 ( .D(bl[7]), .B(GND_), .G(yp2_b_25[7]), .S(vblinhi_rdo));
nch_25  M16 ( .D(bl[6]), .B(GND_), .G(yp2_b_25[6]), .S(vblinhi_rde));
nch_25  M11 ( .D(bl[1]), .B(GND_), .G(yp2_b_25[1]), .S(vblinhi_rdo));
nch_25  M20 ( .D(bl[0]), .B(GND_), .G(yp2_b_25[0]), .S(vblinhi_rde));
nch_25  M15 ( .D(bl[5]), .B(GND_), .G(yp2_b_25[5]), .S(vblinhi_rdo));
nch_25  M14 ( .D(bl[4]), .B(GND_), .G(yp2_b_25[4]), .S(vblinhi_rde));
nch_25  M13 ( .D(bl[3]), .B(GND_), .G(yp2_b_25[3]), .S(vblinhi_rdo));
nch_25  M12 ( .D(bl[2]), .B(GND_), .G(yp2_b_25[2]), .S(vblinhi_rde));
nch_hvt  M3 ( .D(bl[3]), .B(GND_), .G(yp2[3]), .S(bl_out));
nch_hvt  M1 ( .D(bl[2]), .B(GND_), .G(yp2[2]), .S(bl_out));
nch_hvt  M0 ( .D(bl[1]), .B(GND_), .G(yp2[1]), .S(bl_out));
nch_hvt  M7 ( .D(bl[7]), .B(GND_), .G(yp2[7]), .S(bl_out));
nch_hvt  M6 ( .D(bl[6]), .B(GND_), .G(yp2[6]), .S(bl_out));
nch_hvt  M5 ( .D(bl[5]), .B(GND_), .G(yp2[5]), .S(bl_out));
nch_hvt  M2 ( .D(bl[0]), .B(GND_), .G(yp2[0]), .S(bl_out));
nch_hvt  M4 ( .D(bl[4]), .B(GND_), .G(yp2[4]), .S(bl_out));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x64, View - schematic
// LAST TIME SAVED: Feb 26 14:34:16 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_x64 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp2, yp2_b_25, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [63:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
input [7:0]  yp3_25;
input [7:0]  yp3_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  bl_med;



ml_ymux_yp2_8 Iml_ymux_yp2_x8 ( .bl(bl_med[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[0]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_2 ( .vdd_tieh(vdd_tieh), .bl(bl[23:16]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[2]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_3 ( .vdd_tieh(vdd_tieh), .bl(bl[31:24]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[3]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_6 ( .vdd_tieh(vdd_tieh), .bl(bl[55:48]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[6]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_7 ( .vdd_tieh(vdd_tieh), .bl(bl[63:56]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[7]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_5 ( .vdd_tieh(vdd_tieh), .bl(bl[47:40]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[5]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_4 ( .vdd_tieh(vdd_tieh), .bl(bl[39:32]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[4]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_1 ( .vdd_tieh(vdd_tieh), .bl(bl[15:8]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[1]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x328, View - schematic
// LAST TIME SAVED: May  4 14:26:48 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_x328 ( bl, bl_dummyl, bl_dummyr, bl_out, bl_test,
     vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh,
     pgminhi_dmmy_b_25, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test, yp_test_25, yp_test_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25;

inout [1:0]  bl_dummyl;
inout [1:0]  bl_test;
inout [1:0]  bl_dummyr;
inout [327:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp2_b_25;
input [7:0]  yp2;
input [1:0]  yp_test_b_25;
input [5:0]  yp1_b_25;
input [1:0]  yp_test_25;
input [7:0]  yp3_25;
input [1:0]  yp_test;
input [5:0]  yp1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [5:5]  blx8_out;

wire  [0:4]  blx64_out;



ml_ymux_bls_x8 Iml_ymux_bls_x8 ( .bl_out(blx8_out[5]),
     .bl(bl[327:320]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_r ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyr[1:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_l ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyl[1:0]));
pch_25  M7 ( .D(bl_test[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M8 ( .D(bl_test[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
ml_ymux_bls_x64 Iml_ymux_bls_x64_0 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[0]), .bl(bl[63:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_2 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[2]), .bl(bl[191:128]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_4 ( .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]), .bl(bl[319:256]),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .bl_out(blx64_out[4]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo));
ml_ymux_bls_x64 Iml_ymux_bls_x64_1 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[1]), .bl(bl[127:64]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_3 ( .yp2(yp2[7:0]), .bl_out(blx64_out[3]),
     .bl(bl[255:192]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .yp2_b_25(yp2_b_25[7:0]), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));
nch_hvt  M21 ( .D(net224), .B(GND_), .G(yp_test[1]), .S(bl_out));
nch_hvt  M19 ( .D(net228), .B(GND_), .G(yp_test[1]), .S(net224));
nch_hvt  M23 ( .D(net232), .B(GND_), .G(yp_test[0]), .S(bl_out));
nch_hvt  M28 ( .D(net236), .B(GND_), .G(yp1[5]), .S(bl_out));
nch_hvt  M0 ( .D(blx64_out[2]), .B(GND_), .G(yp1[2]), .S(bl_out));
nch_hvt  M22 ( .D(net244), .B(GND_), .G(yp_test[0]), .S(net232));
nch_hvt  M24 ( .D(blx64_out[0]), .B(GND_), .G(yp1[0]), .S(bl_out));
nch_hvt  M30 ( .D(blx8_out[5]), .B(GND_), .G(yp1[5]), .S(net236));
nch_hvt  M3 ( .D(blx64_out[4]), .B(GND_), .G(yp1[4]), .S(bl_out));
nch_hvt  M4 ( .D(blx64_out[3]), .B(GND_), .G(yp1[3]), .S(bl_out));
nch_hvt  M2 ( .D(blx64_out[1]), .B(GND_), .G(yp1[1]), .S(bl_out));
nch_25  M27 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[0]),
     .S(blx64_out[0]));
nch_25  M26 ( .D(vblinhi_rdo), .B(GND_), .G(yp_test_b_25[1]),
     .S(bl_test[1]));
nch_25  M25 ( .D(bl_test[1]), .B(GND_), .G(yp_test_25[1]), .S(net228));
nch_25  M18 ( .D(vblinhi_rde), .B(GND_), .G(yp_test_b_25[0]),
     .S(bl_test[0]));
nch_25  M29 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[5]),
     .S(blx8_out[5]));
nch_25  M17 ( .D(bl_test[0]), .B(GND_), .G(yp_test_25[0]), .S(net244));
nch_25  M1 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[2]),
     .S(blx64_out[2]));
nch_25  M20 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[1]),
     .S(blx64_out[1]));
nch_25  M5 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[4]),
     .S(blx64_out[4]));
nch_25  M6 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[3]),
     .S(blx64_out[3]));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp_x4, View - schematic
// LAST TIME SAVED: Jan 23 10:17:05 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x4 ( wp, gwl_b_sup_25, ngate_25, gwl_b_25,
     gwl_b_gnden_25, gwp_hv, s_b_25, s_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_25, gwl_b_gnden_25, gwp_hv;

output [3:0]  wp;

input [3:0]  s_b_25;
input [3:0]  s_b_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwl_b_25(gwl_b_25), .gwl_gnd_25(gwl_gnd_25));
ml_rock_lwldrv_wp Iml_lwldrv_1 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[1]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[1]), .wp(wp[1]));
ml_rock_lwldrv_wp Iml_lwldrv_2 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[2]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[2]), .wp(wp[2]));
ml_rock_lwldrv_wp Iml_lwldrv_3 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[3]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3]), .wp(wp[3]));
ml_rock_lwldrv_wp Iml_lwldrv_0 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[0]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[0]), .wp(wp[0]));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp_x228, View - schematic
// LAST TIME SAVED: Mar 28 09:57:53 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x228 ( wp, gwl_b_sup_25, ngate_25, s_b_25,
     s_b_hv, gwl_b_25, gwl_b_gnden_25, gwp_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_gnden_25;

output [227:0]  wp;

inout [3:0]  s_b_25;
inout [3:0]  s_b_hv;

input [56:0]  gwl_b_25;
input [56:0]  gwp_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_56_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[56]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[227:224]), .gwl_b_25(gwl_b_25[56]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_55_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[55]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[223:220]), .gwl_b_25(gwl_b_25[55]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_54_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[54]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[219:216]), .gwl_b_25(gwl_b_25[54]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_53_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[53]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[215:212]), .gwl_b_25(gwl_b_25[53]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_52_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[52]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[211:208]), .gwl_b_25(gwl_b_25[52]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_51_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[51]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[207:204]), .gwl_b_25(gwl_b_25[51]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_50_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[50]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[203:200]), .gwl_b_25(gwl_b_25[50]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_49_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[49]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[199:196]), .gwl_b_25(gwl_b_25[49]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_48_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[48]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[195:192]), .gwl_b_25(gwl_b_25[48]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_47_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[47]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[191:188]), .gwl_b_25(gwl_b_25[47]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_46_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[46]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[187:184]), .gwl_b_25(gwl_b_25[46]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_45_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[45]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[183:180]), .gwl_b_25(gwl_b_25[45]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_44_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[44]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[179:176]), .gwl_b_25(gwl_b_25[44]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_43_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[43]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[175:172]), .gwl_b_25(gwl_b_25[43]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_42_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[42]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[171:168]), .gwl_b_25(gwl_b_25[42]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_41_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[41]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[167:164]), .gwl_b_25(gwl_b_25[41]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_40_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[40]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[163:160]), .gwl_b_25(gwl_b_25[40]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_39_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[39]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[159:156]), .gwl_b_25(gwl_b_25[39]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_38_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[38]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[155:152]), .gwl_b_25(gwl_b_25[38]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_37_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[37]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[151:148]), .gwl_b_25(gwl_b_25[37]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_36_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[36]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[147:144]), .gwl_b_25(gwl_b_25[36]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_35_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[35]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[143:140]), .gwl_b_25(gwl_b_25[35]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_34_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[34]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[139:136]), .gwl_b_25(gwl_b_25[34]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_33_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[33]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[135:132]), .gwl_b_25(gwl_b_25[33]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_32_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[32]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[131:128]), .gwl_b_25(gwl_b_25[32]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_31_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[31]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[127:124]), .gwl_b_25(gwl_b_25[31]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_30_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[30]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[123:120]), .gwl_b_25(gwl_b_25[30]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_29_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[29]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[119:116]), .gwl_b_25(gwl_b_25[29]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_28_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[28]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[115:112]), .gwl_b_25(gwl_b_25[28]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_27_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[27]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[111:108]), .gwl_b_25(gwl_b_25[27]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_26_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[26]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[107:104]), .gwl_b_25(gwl_b_25[26]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_25_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[25]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[103:100]), .gwl_b_25(gwl_b_25[25]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_24_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[24]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[99:96]), .gwl_b_25(gwl_b_25[24]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_23_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[23]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[95:92]), .gwl_b_25(gwl_b_25[23]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_22_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[22]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[91:88]), .gwl_b_25(gwl_b_25[22]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_21_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[21]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[87:84]), .gwl_b_25(gwl_b_25[21]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_20_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[20]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[83:80]), .gwl_b_25(gwl_b_25[20]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_19_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[19]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[79:76]), .gwl_b_25(gwl_b_25[19]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_18_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[18]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[75:72]), .gwl_b_25(gwl_b_25[18]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_17_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[17]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[71:68]), .gwl_b_25(gwl_b_25[17]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_16_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[16]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[67:64]), .gwl_b_25(gwl_b_25[16]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_15_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[15]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[63:60]), .gwl_b_25(gwl_b_25[15]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_14_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[14]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[59:56]), .gwl_b_25(gwl_b_25[14]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_13_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[13]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[55:52]), .gwl_b_25(gwl_b_25[13]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_12_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[12]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[51:48]), .gwl_b_25(gwl_b_25[12]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_11_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[11]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[47:44]), .gwl_b_25(gwl_b_25[11]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_10_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[10]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[43:40]), .gwl_b_25(gwl_b_25[10]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_9_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[9]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[39:36]), .gwl_b_25(gwl_b_25[9]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_8_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[8]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[35:32]), .gwl_b_25(gwl_b_25[8]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_7_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[7]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[31:28]), .gwl_b_25(gwl_b_25[7]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_6_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[6]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[27:24]), .gwl_b_25(gwl_b_25[6]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_5_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[5]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[23:20]), .gwl_b_25(gwl_b_25[5]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_4_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[4]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[19:16]), .gwl_b_25(gwl_b_25[4]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_3_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[3]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[15:12]), .gwl_b_25(gwl_b_25[3]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_2_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[2]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[11:8]), .gwl_b_25(gwl_b_25[2]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_1_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[1]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[7:4]), .gwl_b_25(gwl_b_25[1]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_0_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[0]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[3:0]), .gwl_b_25(gwl_b_25[0]), .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM, Cell - ml_core_338x232_top, View - schematic
// LAST TIME SAVED: Sep 22 17:27:05 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_338x232_top ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25,
     sa_ngate_25, sa_pgate_vpxa, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr, wr );
output  nv_dataout;

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     pgminhi_dmmy_b_25, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

input [56:0]  gwl_b_25;
input [56:0]  gwp_hv;
input [227:0]  wr;
input [4:1]  sa_pgate_vpxa;
input [2:0]  fsm_trim_rrefrd;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [4:1]  sa_ngate_25;
input [1:0]  fsm_rowadd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  yp_test_b_25;

wire  [1:0]  yp_test_25;

wire  [1:0]  yp_test;

wire  [7:0]  yp3_b_25;

wire  [7:0]  yp3;

wire  [7:0]  yp2;

wire  [7:0]  yp2_b_25;

wire  [5:0]  yp1_b_25;

wire  [5:0]  yp1;

wire  [327:0]  bl;

wire  [1:0]  bl_dummyr;

wire  [1:0]  bl_dummyl;

wire  [227:0]  wp;

wire  [3:0]  s_b_hv;

wire  [3:0]  s_b_25;

wire  [1:0]  bl_test;



ml_core_sa_spare Iml_core_sa_spare ( );
vdd_tielow I47 ( .gnd_tiel(net127));
inv_hvt I131 ( .A(nv_dataout_in), .Y(net129));
inv_hvt I45 ( .A(net129), .Y(nv_dataout));
ml_core_ctrl_top Icore_ctrl_top ( .yp2_b_25(yp2_b_25[7:0]),
     .yp2(yp2[7:0]), .yp1_b_25(yp1_b_25[5:0]), .yp1(yp1[5:0]),
     .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .gwl_b_gnden_25(gwl_b_gnden_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .vdd_tieh(vdd_tieh), .tm_testdec_wr(tm_testdec_wr),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .testdec_en_b_25(testdec_en_b_25),
     .saen_b_vpxa(saen_b_vpxa), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .dec_ok_25(dec_ok_25), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .nv_dataout(nv_dataout_in), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_pgm_25(vblinhi_pgm_25),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .bl_out(bl_out),
     .yp_test(yp_test[1:0]));
nvcm_cell_338x232 Invcm_cell_338x232 ( .bl_dummyr(bl_dummyr[1:0]),
     .wr_dummyt({net127, net127}), .wr_dummyb({net127, net127}),
     .wr(wr[227:0]), .wp_dummyt({net127, net127}), .wp_dummyb({net127,
     net127}), .wp(wp[227:0]), .bl_test(bl_test[1:0]),
     .bl_dummyl(bl_dummyl[1:0]), .bl(bl[327:0]));
ml_testdec_bgen Itestdec_bgen ( .dec_ok_25(dec_ok_25),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25), .dec_det_25(dec_det_25),
     .dec_bias_25(dec_bias));
ml_testdec_rowsx228 Itestdec_rowsx228 ( .dec_bias_25(dec_bias),
     .dec_det_25(dec_det_25), .wr(wr[227:0]), .wp(wp[227:0]),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25));
ml_testdec_columnsx330 Itestdec_columnsx330 (
     .bl_dummyr(bl_dummyr[1:0]), .bl_dummyl(bl_dummyl[1:0]),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[327:0]),
     .bl_test(bl_test[1:0]));
ml_ymux_bls_x328 Iml_ymux_bls_x328 ( .yp1_b_25(yp1_b_25[5:0]),
     .yp1(yp1[5:0]), .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]),
     .vdd_tieh(vdd_tieh), .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25),
     .bl_dummyl(bl_dummyl[1:0]), .bl_dummyr(bl_dummyr[1:0]),
     .bl_test(bl_test[1:0]), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp_test(yp_test[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3[7:0]),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .vblinhi_pgm_25(vblinhi_pgm_25), .bl_out(bl_out), .bl(bl[327:0]));
ml_rock_lwldrv_wp_x228 Iml_rock_lwldrv_wp_x228 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[56:0]), .gwl_b_25(gwl_b_25[56:0]), .wp(wp[227:0]),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .ngate_25(ngate_25));

endmodule
// Library - NVCM, Cell - ml_core_bank_1, View - schematic
// LAST TIME SAVED: Apr 25 16:18:29 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_bank_1 ( nv_dataout, bl_pgm_glb, gwl_b_sup_25, ngate_25,
     sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa, ysup_25,
     fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv,
     pgminhi_dmmy_b_25, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     pgminhi_dmmy_b_25, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [8:4]  nv_dataout;

input [1:0]  fsm_rowadd;
input [8:0]  fsm_coladd;
input [4:1]  sa_pgate_vpxa;
input [56:0]  gwl_b_25;
input [2:0]  fsm_trim_rrefpgm;
input [56:0]  gwp_hv;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_blkadd;
input [227:0]  wr;
input [4:1]  sa_ngate_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_core_338x232_top blk4 ( .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .nv_dataout(nv_dataout[4]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x232_top blk5 ( .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd_b[1], fsm_blkadd[0]}),
     .nv_dataout(nv_dataout[5]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x232_top blk7 ( .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd[1], fsm_blkadd[0]}),
     .nv_dataout(nv_dataout[7]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x232_top blk6 ( .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd_b[3],
     fsm_blkadd[2], fsm_blkadd[1], fsm_blkadd_b[0]}),
     .nv_dataout(nv_dataout[6]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));
ml_core_338x232_top blk8 ( .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd({fsm_blkadd[3],
     fsm_blkadd_b[2], fsm_blkadd_b[1], fsm_blkadd_b[0]}),
     .nv_dataout(nv_dataout[8]), .ysup_25(ysup_25), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb));

endmodule
// Library - NVCM, Cell - ml_core_bank_0, View - schematic
// LAST TIME SAVED: May  7 10:06:14 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core_bank_0 ( nv_dataout, bl_pgm_glb, gwl_b_sup_25, ngate_25,
     sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa, ysup_25,
     fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_gwlbdis_b_25,
     fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv,
     pgminhi_dmmy_b_25, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     pgminhi_dmmy_b_25, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr;

output [3:0]  nv_dataout;

input [4:1]  sa_ngate_25;
input [8:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefrd;
input [4:1]  sa_pgate_vpxa;
input [56:0]  gwl_b_25;
input [1:0]  fsm_rowadd;
input [56:0]  gwp_hv;
input [2:0]  fsm_trim_rrefpgm;
input [227:0]  wr;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_blkadd_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_core_338x232_top blk3 ( .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd[1],
     fsm_blkadd[0]}), .nv_dataout(nv_dataout[3]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
ml_core_338x232_top blk1 ( .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd[0]}), .nv_dataout(nv_dataout[1]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
ml_core_338x232_top blk2 ( .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd[1],
     fsm_blkadd_b[0]}), .nv_dataout(nv_dataout[2]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
ml_core_338x232_top blk0 ( .wr(wr[227:0]),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen), .tm_dma(tm_dma),
     .fsm_tm_trow(fsm_tm_trow), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_coladd(fsm_coladd[8:0]),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd_b[0]}), .nv_dataout(nv_dataout[0]), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));

endmodule
// Library - NVCM, Cell - ml_core, View - schematic
// LAST TIME SAVED: May  7 10:16:05 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_core ( nv_dataout, bgr, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpp_int, vpxa, ysup_25, fsm_blkadd,
     fsm_blkadd_b, fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven,
     fsm_multibl_read, fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_trim_ipp,
     fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo,
     vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbl_h, tm_allbl_l, tm_allwl_h,
     tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [8:0]  nv_dataout;

input [3:0]  fsm_blkadd_b;
input [8:0]  fsm_coladd;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_trim_rrefrd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [227:0]  wr;

wire  [4:1]  sa_pgate_vpxa;

wire  [4:1]  sa_ngate_25;

wire  [56:0]  gwl_b_25;

wire  [56:0]  gwp_hv;



ml_gwlwr_top Igwlwr_top ( .fsm_pgmdisc(fsm_pgmdisc), .fsm_din(fsm_din),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .fsm_wren(fsm_wren),
     .tm_testdec(fsm_tm_testdec), .fsm_tm_allbl_h(tm_allbl_h),
     .fsm_tm_allwl_l(tm_allwl_l), .fsm_tm_allwl_h(tm_allwl_h),
     .fsm_tm_allbl_l(tm_allbl_l), .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_wpen(fsm_wpen), .tm_dma(tm_dma), .gwl_b_sup_25(gwl_b_sup_25),
     .gwl_b_25(gwl_b_25[56:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .wr(wr[227:0]), .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .vpxa(vpxa), .vpp_int(vpp_int), .bl_pgm_glb(bl_pgm_glb),
     .bgr(bgr));
ml_core_bank_1 bank1 ( .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwl_b_sup_25(gwl_b_sup_25),
     .ngate_25(ngate_25), .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vpxa(vpxa), .ysup_25(ysup_25),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .fsm_nvcmen(fsm_nvcmen),
     .fsm_pgm(fsm_pgm), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_rd(fsm_rd),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rst_b(fsm_rst_b),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .fsm_vpxaset(fsm_vpxaset),
     .fsm_wpen(fsm_wpen), .fsm_ymuxdis(fsm_ymuxdis),
     .gwl_b_25(gwl_b_25[56:0]), .gwp_hv(gwp_hv[56:0]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]), .saen_25(saen_25),
     .saen_b_vpxa(saen_b_vpxa), .testdec_en_b_25(testdec_en_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_prec_b_25(testdec_prec_b_25), .tm_allbl_h(tm_allbl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allwl_l(tm_allwl_l), .tm_tcol(tm_tcol),
     .tm_testdec_wr(tm_testdec_wr), .wr(wr[227:0]),
     .fsm_blkadd(fsm_blkadd[3:0]), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .nv_dataout(nv_dataout[8:4]), .bl_pgm_glb(bl_pgm_glb));
ml_core_bank_0 bank0 ( .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .ysup_25(ysup_25),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .nv_dataout(nv_dataout[3:0]), .vpxa(vpxa),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .ngate_25(ngate_25), .gwl_b_sup_25(gwl_b_sup_25),
     .bl_pgm_glb(bl_pgm_glb), .tm_testdec_wr(tm_testdec_wr),
     .wr(wr[227:0]));

endmodule
// Library - NVCM, Cell - ml_chip_nvcm, View - schematic
// LAST TIME SAVED: Sep 19 11:56:13 2008
// NETLIST TIME: Nov 14 16:12:00 2008
`timescale 1ns / 1ns 

module ml_chip_nvcm ( nv_dataout, vpp, fsm_blkadd, fsm_blkadd_b,
     fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_trim_vbg,
     fsm_vpgmwl, fsm_vpxaset, fsm_vrdwl, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbl_h, tm_allbl_l, tm_allwl_h,
     tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl );

inout  vpp;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr, tm_wleqbl;

output [8:0]  nv_dataout;

input [3:0]  fsm_blkadd;
input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_vpgmwl;
input [2:0]  fsm_vrdwl;
input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_trim_vbg;
input [7:0]  fsm_rowadd;
input [8:0]  fsm_coladd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  fsm_trim_vbg_buf;

wire  [2:0]  fsm_vpgmwl_buf;



ml_chip_spare Iml_chip_spare ( );
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(vddp_));
ml_chip_buf_top Ichip_buf_top ( .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_pgm(fsm_pgm),
     .fsm_pgm_buf(fsm_pgm_buf), .fsm_wgnden_buf(fsm_wgnden_buf),
     .fsm_wgnden(fsm_wgnden), .fsm_vpgmwl(fsm_vpgmwl[2:0]),
     .fsm_trim_vbg(fsm_trim_vbg[3:0]), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_nvcmen(fsm_nvcmen), .fsm_lshven(fsm_lshven),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .fsm_lshven_buf(fsm_lshven_buf));
ml_vppint_top Ivppint_top ( .vpint_en(vpint_en),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .vpp_int(vpp_int), .fsm_wgnden_buf(fsm_wgnden_buf), .bgr(bgr),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf));
ml_bgr_top Ibgr_top ( .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .bgr_int(bgr_int));
ml_vpxa_top Ivpxa_top ( .fsm_pumpen(fsm_pumpen),
     .fsm_vrdwl(fsm_vrdwl[2:0]), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .bgr(bgr), .vpxa_int(vpxa));
ml_hvmux_top Ihvmux_top ( .vpint_en(vpint_en), .fsm_wpen(fsm_wpen),
     .tm_wleqbl(tm_wleqbl), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden_buf), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvpxa(fsm_tm_xvpxa), .fsm_tm_xvppint(fsm_tm_xvppint),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy_buf),
     .fsm_pgm(fsm_pgm_buf), .fsm_nvcmen(fsm_nvcmen_buf),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven_buf),
     .bgr(bgr), .bgr_int(bgr_int), .ngate_25(ngate_25),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv), .vpp(vpp),
     .vpp_int(vpp_int), .vpxa(vpxa), .vpxa_int(vpxa),
     .ysup_25(ysup_25), .vblinhi(vblinhi),
     .tm_testdec(fsm_tm_testdec));
ml_core Icore ( .fsm_pgmdisc(fsm_pgmdisc), .fsm_din(fsm_din),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol), .tm_dma(tm_dma),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[8:0]), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_blkadd(fsm_blkadd[3:0]), .bgr(bgr), .ngate_25(ngate_25),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpp_int(vpp_int),
     .vpxa(vpxa), .ysup_25(ysup_25), .nv_dataout(nv_dataout[8:0]),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));

endmodule
// Library - xpmem, Cell - ml_rowdrv2, View - schematic
// LAST TIME SAVED: Aug 23 15:16:05 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_rowdrv2 ( pgate, reset, smc_rsr_out, vddctrl, wl, wl_rd_sup,
     wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
ml_dff_schematic I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));

endmodule
// Library - misc, Cell - nvcm_top, View - schematic
// LAST TIME SAVED: Apr  7 16:06:57 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module nvcm_top ( bp0, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_redrow,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_recall,
     fsm_rowadd, fsm_sample, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_dma, fsm_tm_margin0_read,
     fsm_tm_rd_mode, fsm_tm_tcol, fsm_tm_testdec, fsm_tm_testdec_wr,
     fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvpp, fsm_tm_xvpxa, fsm_tm_xvpxa_int, fsm_trim_ipp,
     fsm_trim_multibl_read, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_trim_vbg, fsm_trim_vpgmwl, fsm_trim_vrdwl, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b, clk, icef_member_sel,
     nv_dataout, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi,
     spi_ss_b );
output  bp0, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_redrow, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_recall, fsm_sample, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_dma,
     fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_tcol, fsm_tm_testdec,
     fsm_tm_testdec_wr, fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvpp, fsm_tm_xvpxa, fsm_tm_xvpxa_int,
     fsm_trim_multibl_read, fsm_vpxaset, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy, nvcm_relextspi,
     spi_sdo, spi_sdo_oe_b;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

output [8:0]  fsm_coladd;
output [3:0]  fsm_trim_vbg;
output [8:0]  fsm_rowadd;
output [2:0]  fsm_trim_vpgmwl;
output [3:0]  fsm_blkadd;
output [2:0]  fsm_trim_vrdwl;
output [2:0]  fsm_trim_rrefrd;
output [3:0]  fsm_blkadd_b;
output [2:0]  fsm_trim_rrefpgm;
output [3:0]  fsm_trim_ipp;

input [8:0]  nv_dataout;
input [1:0]  icef_member_sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - misc, Cell - nvcm_ml_block, View - schematic
// LAST TIME SAVED: Apr 21 10:48:12 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module nvcm_ml_block ( bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b, vpp, clk,
     icef_member_sel, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi,
     spi_ss_b );
output  bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b;

inout  vpp;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

input [1:0]  icef_member_sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net212;

wire  [0:3]  net249;

wire  [0:2]  net206;

wire  [0:8]  net0144;

wire  [0:2]  net209;

wire  [0:2]  net210;

wire  [0:8]  net247;

wire  [0:2]  net207;

wire  [0:3]  net248;

wire  [8:0]  fsm_rowadd;

wire  [0:3]  net208;


/*
sg_bufx10 I217 ( .in(rst_b), .out(rst_bd));
ml_chip_nvcm Iml_chip_nvcm ( .tm_wleqbl(net217),
     .tm_testdec_wr(net219), .tm_tcol(net221), .tm_dma(net224),
     .tm_allwl_l(net225), .tm_allwl_h(net226), .tm_allbl_l(net227),
     .tm_allbl_h(net228), .fsm_ymuxdis(net200), .fsm_wren(net201),
     .fsm_wpen(net202), .fsm_wgnden(net203), .fsm_vrdwl(net206[0:2]),
     .fsm_vpxaset(net204), .fsm_vpgmwl(net207[0:2]),
     .fsm_trim_vbg(net208[0:3]), .fsm_trim_rrefrd(net209[0:2]),
     .fsm_trim_rrefpgm(net210[0:2]), .fsm_trim_ipp(net212[0:3]),
     .fsm_tm_xvpxaint(net213), .fsm_tm_xvpxa(net214),
     .fsm_tm_xvppint(net272), .fsm_tm_xvbg(net205),
     .fsm_tm_xforce(net216), .fsm_tm_trow(net218),
     .fsm_tm_testdec(net220), .fsm_tm_rd_mode(net222),
     .fsm_sample(net229), .fsm_rst_b(rst_bd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(net232),
     .fsm_pumpen(net233), .fsm_pgmvfy(net234), .fsm_pgmien(net235),
     .fsm_pgmhv(net236), .fsm_pgmdisc(net237), .fsm_pgm(net238),
     .fsm_nvcmen(net239), .fsm_nv_sisi_ui(net240),
     .fsm_nv_rrow(net242), .fsm_nv_rri_trim(net241),
     .fsm_nv_bstream(net243), .fsm_multibl_read(net211),
     .fsm_lshven(net244), .fsm_gwlbdis(net245), .fsm_din(net246),
     .fsm_coladd(net247[0:8]), .fsm_blkadd_b(net248[0:3]),
     .fsm_blkadd(net249[0:3]), .nv_dataout(net0144[0:8]), .vpp(vpp));
nvcm_top Invcm_top ( .spi_ss_b(spi_ss_b), .spi_sdi(spi_sdi),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_ce_b(nvcm_ce_b), .nv_dataout(net0144[0:8]),
     .icef_member_sel(icef_member_sel[1:0]), .clk(clk),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .nvcm_relextspi(nvcm_relextspi), .nvcm_rdy(nvcm_rdy),
     .nvcm_boot(nvcm_boot), .fsm_ymuxdis(net200), .fsm_wren(net201),
     .fsm_wpen(net202), .fsm_wgnden(net203), .fsm_vpxaset(net204),
     .fsm_tm_xvbg(net205), .fsm_trim_vrdwl(net206[0:2]),
     .fsm_trim_vpgmwl(net207[0:2]), .fsm_trim_vbg(net208[0:3]),
     .fsm_trim_rrefrd(net209[0:2]), .fsm_trim_rrefpgm(net210[0:2]),
     .fsm_trim_multibl_read(net211), .fsm_trim_ipp(net212[0:3]),
     .fsm_tm_xvpxa_int(net213), .fsm_tm_xvpxa(net214),
     .fsm_tm_xvpp(net272), .fsm_tm_xforce(net216),
     .fsm_tm_vwleqbl(net217), .fsm_tm_trow(net218),
     .fsm_tm_testdec_wr(net219), .fsm_tm_testdec(net220),
     .fsm_tm_tcol(net221), .fsm_tm_rd_mode(net222),
     .fsm_tm_margin0_read(fsm_tm_margin0_read), .fsm_tm_dma(net224),
     .fsm_tm_allwl_l(net225), .fsm_tm_allwl_h(net226),
     .fsm_tm_allbl_l(net227), .fsm_tm_allbl_h(net228),
     .fsm_sample(net229), .fsm_rowadd(fsm_rowadd[8:0]),
     .fsm_recall(fsm_recall), .fsm_rd(net232), .fsm_pumpen(net233),
     .fsm_pgmvfy(net234), .fsm_pgmien(net235), .fsm_pgmhv(net236),
     .fsm_pgmdisc(net237), .fsm_pgm(net238), .fsm_nvcmen(net239),
     .fsm_nv_sisi_ui(net240), .fsm_nv_rri_trim(net241),
     .fsm_nv_redrow(net242), .fsm_nv_bstream(net243),
     .fsm_lshven(net244), .fsm_gwlbdis(net245), .fsm_din(net246),
     .fsm_coladd(net247[0:8]), .fsm_blkadd_b(net248[0:3]),
     .fsm_blkadd(net249[0:3]), .bp0(bp0));
*/
endmodule
// Library - ice4chip, Cell - CHIP_route_left, View - schematic
// LAST TIME SAVED: Oct  7 18:00:03 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module CHIP_route_left ( cm_banksel_bltld3_1_, cm_clk_bltld3,
     cm_sdi_u1d3[1:0], cm_sdo_u1d1[1:0], core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, last_rsr[1:0],
     monitor_celld2[1:0], pgate_l[351:0], reset_l[351:0],
     smc_wdis_dclk_bltld3, vdd_cntl_l[351:0], wl_l[351:0],
     cf_lbank[300], cf_lbank[479], cm_banksel_blbld1[0],
     cm_banksel_blbld[1], cm_clk_blbld, cm_sdi_u1d[1:0],
     cm_sdo_u1[1:0], core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0 );
output  cm_banksel_bltld3_1_, cm_clk_bltld3, core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, smc_wdis_dclk_bltld3;

input  cm_clk_blbld, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;

output [351:0]  reset_l;
output [1:0]  cm_sdo_u1d1;
output [351:0]  pgate_l;
output [1:0]  last_rsr;
output [1:0]  monitor_celld2;
output [351:0]  vdd_cntl_l;
output [351:0]  wl_l;
output [1:0]  cm_sdi_u1d3;

input [1:0]  cm_sdo_u1;
input [300:479]  cf_lbank;
input [0:0]  cm_banksel_blbld1;
input [1:0]  cm_sdi_u1d;
input [1:1]  cm_banksel_blbld;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net081;

wire  [1:1]  monitor_celld1;

wire  [1:0]  cm_sdo_u1d;

wire  [1:0]  cm_sdi_u1d0;

wire  [1:1]  monitor_celld;

wire  [1:1]  cm_banksel_bltld;

wire  [1:0]  cm_sdo_u1d0;

wire  [1:0]  dff_out;



tielo I451_1_ ( .tielo(net081[0]));
tielo I451_0_ ( .tielo(net081[1]));
tielo I452 ( .tielo(net0132));
bram_bufferx16 I381 ( .in(j_rst_bl1), .out(trst_rowu0));
bram_bufferx16 I391 ( .in(j_rst_bl2), .out(trst_rowu1));
bram_bufferx16 I392 ( .in(row_testl3), .out(row_test_rowu1));
bram_bufferx16 I393 ( .in(cram_pgateoffl2), .out(cram_pgateoff_rowu1));
bram_bufferx16 I394 ( .in(cram_rstl2), .out(cram_rst_rowu1));
bram_bufferx16 I395 ( .in(cram_wl_enl2), .out(cram_wl_en_rowu1));
bram_bufferx16 I396 ( .in(smc_writel2), .out(smc_write_rowu1));
bram_bufferx16 I397 ( .in(cram_vddoffl2), .out(cram_vddoff_rowu1));
bram_bufferx16 I398 ( .in(smc_row_incl2), .out(smc_row_inc_rowu1));
bram_bufferx16 I400 ( .in(smc_rsr_rstl2), .out(smc_rsr_rst_rowu1));
bram_bufferx16 I390 ( .in(smc_rsr_rstl1), .out(smc_rsr_rst_rowu0));
bram_bufferx16 I435 ( .in(tck_padl2), .out(tck_pad_rowu1));
bram_bufferx16 I384 ( .in(cram_rstl1), .out(cram_rst_rowu0));
bram_bufferx16 I290 ( .in(cm_clk_blbld), .out(net325));
bram_bufferx16 I260 ( .in(cm_clk_blbld), .out(net347));
bram_bufferx16 I385 ( .in(cram_vddoffl1), .out(cram_vddoff_rowu0));
bram_bufferx16 I386 ( .in(cram_wl_enl1), .out(cram_wl_en_rowu0));
bram_bufferx16 I387 ( .in(smc_row_incl1), .out(smc_row_inc_rowu0));
bram_bufferx16 I388 ( .in(smc_writel1), .out(smc_write_rowu0));
bram_bufferx16 I389 ( .in(core_por_bbl1), .out(core_por_b_rowu0));
bram_bufferx16 I383 ( .in(cram_pgateoffl1), .out(cram_pgateoff_rowu0));
bram_bufferx16 I437 ( .in(tck_padl1), .out(tck_pad_rowu0));
bram_bufferx16 I382 ( .in(row_testl2), .out(row_test_rowu0));
sg_dffbuf I261_1_ ( .r(net081[0]), .dffout(dff_out[1]),
     .d(cm_sdo_u1d[1]), .clk(net347));
sg_dffbuf I261_0_ ( .r(net081[1]), .dffout(dff_out[0]),
     .d(cm_sdo_u1d[0]), .clk(net347));
sg_dffbuf I289 ( .r(net0132), .d(last_rsr[0]), .clk(net325),
     .dffout(last_rsr0));
ml_rowdrv_bank Irowul (
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu1_b),
     .smc_write(smc_write_rowu1), .smc_rsr_inc(smc_row_inc_rowu1),
     .rsr_rst(smc_rsr_rst_rowu1), .por_rst(core_por_b_rowu1),
     .cram_wl_en(cram_wl_en_rowu1), .cram_vddoff(cram_vddoff_rowu1),
     .cram_rst(cram_rst_rowu1), .cram_pgateoff(cram_pgateoff_rowu1),
     .banksel(cm_banksel_bltld3_1_), .vddctrl(vdd_cntl_l[351:176]),
     .last_rsr(last_rsr[1]), .reset(reset_l[351:176]),
     .pgate(pgate_l[351:176]), .trst_b(trst_rowu1),
     .jtag_rowtest_rst(row_test_rowu1), .jtag_clk(tck_pad_rowu1),
     .wl(wl_l[351:176]));
ml_rowdrv_bank Irowbl (
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu0_b),
     .smc_write(smc_write_rowu0), .smc_rsr_inc(smc_row_inc_rowu0),
     .rsr_rst(smc_rsr_rst_rowu0), .por_rst(core_por_b_rowu0),
     .cram_wl_en(cram_wl_en_rowu0), .cram_vddoff(cram_vddoff_rowu0),
     .cram_rst(cram_rst_rowu0), .cram_pgateoff(cram_pgateoff_rowu0),
     .banksel(cm_banksel_blbld1[0]), .vddctrl(vdd_cntl_l[175:0]),
     .last_rsr(last_rsr[0]), .reset(reset_l[175:0]),
     .pgate(pgate_l[175:0]), .trst_b(trst_rowu0),
     .jtag_rowtest_rst(row_test_rowu0), .jtag_clk(tck_pad_rowu0),
     .wl(wl_l[175:0]));
sg_bufx10 I421 ( .in(cf_lbank[479]), .out(monitor_celld[1]));
sg_bufx10 I235 ( .in(data_muxsel_bltld), .out(data_muxsel_bltld3));
sg_bufx10 I425 ( .in(monitor_celld[1]), .out(monitor_celld1[1]));
sg_bufx10 I424 ( .in(cf_lbank[300]), .out(monitor_celld2[0]));
sg_bufx10 I426 ( .in(monitor_celld1[1]), .out(monitor_celld2[1]));
sg_bufx10 I450_1_ ( .in(dff_out[1]), .out(cm_sdo_u1d1[1]));
sg_bufx10 I450_0_ ( .in(dff_out[0]), .out(cm_sdo_u1d1[0]));
sg_bufx10 I106_1_ ( .in(cm_sdo_u1[1]), .out(cm_sdo_u1d0[1]));
sg_bufx10 I106_0_ ( .in(cm_sdo_u1[0]), .out(cm_sdo_u1d0[0]));
sg_bufx10 I337 ( .in(core_por_bbl0), .out(core_por_bbl1));
sg_bufx10 I338 ( .in(smc_rsr_rstl0), .out(smc_rsr_rstl1));
sg_bufx10 I339 ( .in(row_testl1), .out(row_testl2));
sg_bufx10 I340 ( .in(j_rst_bl0), .out(j_rst_bl1));
sg_bufx10 I342 ( .in(smc_writel0), .out(smc_writel1));
sg_bufx10 I343 ( .in(smc_row_incl0), .out(smc_row_incl1));
sg_bufx10 I344 ( .in(cram_wl_enl0), .out(cram_wl_enl1));
sg_bufx10 I345 ( .in(cram_vddoffl0), .out(cram_vddoffl1));
sg_bufx10 I346 ( .in(cram_rstl0), .out(cram_rstl1));
sg_bufx10 I347 ( .in(cram_pgateoffl0), .out(cram_pgateoffl1));
sg_bufx10 I355 ( .in(cram_pgateoffl1), .out(cram_pgateoffl2));
sg_bufx10 I438 ( .in(tck_padl0), .out(tck_padl1));
sg_bufx10 I237 ( .in(data_muxsel1_bltld), .out(data_muxsel1_bltld3));
sg_bufx10 I351 ( .in(smc_row_incl1), .out(smc_row_incl2));
sg_bufx10 I368 ( .in(cram_pullup_bltld), .out(cram_pullup_bltld3));
sg_bufx10 I277 ( .in(cm_banksel_blbld[1]), .out(cm_banksel_bltld[1]));
sg_bufx10 I348 ( .in(smc_rsr_rstl1), .out(smc_rsr_rstl2));
sg_bufx10 I278_1_ ( .in(cm_sdo_u1d0[1]), .out(cm_sdo_u1d[1]));
sg_bufx10 I278_0_ ( .in(cm_sdo_u1d0[0]), .out(cm_sdo_u1d[0]));
sg_bufx10 I354 ( .in(cram_rstl1), .out(cram_rstl2));
sg_bufx10 I271 ( .in(data_muxsel1_blbld), .out(data_muxsel1_bltld));
sg_bufx10 I275 ( .in(cram_prec_blbld), .out(cram_prec_bltld));
sg_bufx10 I241 ( .in(en_8bconfig_b_bltld), .out(en_8bconfig_b_bltld3));
sg_bufx10 I353 ( .in(cram_vddoffl1), .out(cram_vddoffl2));
sg_bufx10 I357 ( .in(j_rst_bl1), .out(j_rst_bl2));
sg_bufx10 I356 ( .in(row_testl2), .out(row_testl3));
sg_bufx10 I273 ( .in(smc_wdis_dclk_blbld), .out(smc_wdis_dclk_bltld));
sg_bufx10 I279_1_ ( .in(cm_sdi_u1d[1]), .out(cm_sdi_u1d0[1]));
sg_bufx10 I279_0_ ( .in(cm_sdi_u1d[0]), .out(cm_sdi_u1d0[0]));
sg_bufx10 I272 ( .in(en_8bconfig_b_blbld), .out(en_8bconfig_b_bltld));
sg_bufx10 I274 ( .in(cram_write_blbld), .out(cram_write_bltld));
sg_bufx10 I239 ( .in(smc_wdis_dclk_bltld), .out(smc_wdis_dclk_bltld3));
sg_bufx10 I270 ( .in(data_muxsel_blbld), .out(data_muxsel_bltld));
sg_bufx10 I240 ( .in(cram_write_bltld), .out(cram_write_bltld3));
sg_bufx10 I238 ( .in(cram_prec_bltld), .out(cram_prec_bltld3));
sg_bufx10 I242 ( .in(cm_clk_bltld), .out(cm_clk_bltld3));
sg_bufx10 I236 ( .in(cm_banksel_bltld[1]), .out(cm_banksel_bltld3_1_));
sg_bufx10 I276 ( .in(cm_clk_blbld), .out(cm_clk_bltld));
sg_bufx10 I352 ( .in(cram_wl_enl1), .out(cram_wl_enl2));
sg_bufx10 I280_1_ ( .in(cm_sdi_u1d0[1]), .out(cm_sdi_u1d3[1]));
sg_bufx10 I280_0_ ( .in(cm_sdi_u1d0[0]), .out(cm_sdi_u1d3[0]));
sg_bufx10 I350 ( .in(smc_writel1), .out(smc_writel2));
sg_bufx10 I349 ( .in(core_por_bbl1), .out(core_por_b_rowu1));
sg_bufx10 I369 ( .in(cram_pullup_blbld), .out(cram_pullup_bltld));
sg_bufx10 I436 ( .in(tck_padl1), .out(tck_padl2));

endmodule
// Library - xpmem, Cell - sg_bufx10bot, View - schematic
// LAST TIME SAVED: Sep 18 11:01:27 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module sg_bufx10bot ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - bram_bufferx6, View - schematic
// LAST TIME SAVED: Jun 25 13:45:32 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module bram_bufferx6 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - creset_filter, View - schematic
// LAST TIME SAVED: Aug  4 13:06:59 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module creset_filter ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I11 ( .in(net042), .out(out));
inv_hvt I6 ( .A(net13), .Y(net042));
inv_hvt I4 ( .A(in), .Y(net9));
rppolywo_m  R0 ( .MINUS(net17), .PLUS(pbias), .BULK(gnd_));
nch_hvt  M0 ( .D(net13), .B(gnd_), .G(in), .S(gnd_));
nch_hvt  MN31 ( .D(net17), .B(gnd_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(net13), .B(vdd_), .G(net042), .S(vdd_));
pch_hvt  M2 ( .D(net13), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  M1 ( .D(vdd_), .B(vdd_), .G(net13), .S(vdd_));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - xpmem, Cell - ml_dff_bl, View - schematic
// LAST TIME SAVED: Sep  6 14:18:45 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_dff_bl ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_clk_buf, View - schematic
// LAST TIME SAVED: Sep  5 15:09:27 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_clk_buf ( o, in );
output  o;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_powersurg_buf, View - schematic
// LAST TIME SAVED: Jul 31 18:29:48 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_powersurg_buf ( o, in );
output  o;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I404 ( .A(net016), .Y(net012));
inv_hvt I405 ( .A(net012), .Y(o));
inv_hvt I391 ( .A(net77), .Y(net016));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_sch, View - schematic
// LAST TIME SAVED: Sep  6 14:30:13 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_sch ( dataout, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, datain, latch_clock, latch_reset, smc_wdic_clk );
output  dataout;

inout  bl;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, datain,
     latch_clock, latch_reset, smc_wdic_clk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_dff_bl Idff ( .R(latch_reset), .D(dff_in), .CLK(latch_clock),
     .QN(write_data_b), .Q(dff_data));
nor2_hvt I223 ( .A(net084), .B(write_data_b), .Y(n_gate));
inv_hvt I163 ( .A(write_data_b), .Y(dataout));
inv_hvt I159 ( .A(cram_prec), .Y(net0161));
inv_hvt I160 ( .A(cram_write), .Y(net084));
mux2_hvt I161 ( .in1(sa_out), .in0(datain), .out(latch_in),
     .sel(data_muxsel));
mux2_hvt I164 ( .in1(dff_data), .in0(latch_in), .out(dff_in),
     .sel(smc_wdic_clk));
nch_hvt  MN12 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN8 ( .D(sa_out), .B(gnd_), .G(cram_pullup_b), .S(gnd_));
nch_hvt  MN10 ( .D(net0166), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN13 ( .D(net0184), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN3 ( .D(sa_out), .B(gnd_), .G(bl), .S(gnd_));
nch_hvt  MN6 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
pch_hvt  MP8 ( .D(net0148), .B(vdd_), .G(dataout), .S(vdd_));
pch_hvt  MP9 ( .D(bl), .B(vdd_), .G(net084), .S(net0148));
pch_hvt  MP13 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP12 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP14 ( .D(net0208), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP4 ( .D(net0143), .B(vdd_), .G(cram_pullup_b), .S(vdd_));
pch_hvt  MP5 ( .D(sa_out), .B(vdd_), .G(bl), .S(net0143));
pch_hvt  MP15 ( .D(net0204), .B(vdd_), .G(net0161), .S(vdd_));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile_last, View - schematic
// LAST TIME SAVED: Aug  9 15:08:40 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_rowdrv_tile_last ( pgate, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  wl;
output [15:0]  reset;
output [15:0]  pgate;
output [15:0]  vddctrl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  smc_rsr_out;



nor2_hvt I211 ( .A(smc_rsr_out[15]), .Y(net049), .B(smc_rsr_inc_out));
ml_rowdrv2_last Iml_rowdrv2_last ( .smc_rsr_inc(smc_rsr_inc_last),
     .smc_rsr_in(smc_rsr_out[14]), .rsr_rst(rsr_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_rst(cram_rst_buf),
     .smc_rsr_out(smc_rsr_out[15]), .reset(reset[15]), .wl(wl[15]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]));
inv_hvt I391 ( .A(net049), .Y(smc_rsr_inc_last));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I194 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I195 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I198 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I207 ( .A(net041), .Y(por_rst_buf));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net079));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I200 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I206 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I190 ( .A(net079), .Y(smc_rsr_1st_out));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_bram, View - schematic
// LAST TIME SAVED: Sep  5 15:59:47 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tile_bram ( cram_prec_out, cram_write_out, data_out,
     para_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, para_en, para_in,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out, para_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, para_en, para_in, smc_wdic_clk;

inout [41:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  ck;

wire  [0:41]  dataout;



ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
mux2_hvt I161 ( .in1(para_in), .in0(dataout[1]), .out(data_out_mux),
     .sel(para_en));
inv_hvt I262 ( .A(data_out_mux), .Y(net59));
inv_hvt I261 ( .A(net59), .Y(dataout1_mux));
inv_hvt I175 ( .A(dataout[1]), .Y(net62));
inv_hvt I176 ( .A(net62), .Y(para_out));
inv_hvt I172 ( .A(net68), .Y(data_out));
inv_hvt I171 ( .A(dataout[41]), .Y(net68));
ml_powersurg_buf I165 ( .in(cram_prec), .o(net70));
ml_powersurg_buf I163 ( .in(net70), .o(net72));
ml_powersurg_buf I162 ( .in(net78), .o(net74));
ml_powersurg_buf I169 ( .in(net74), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(cram_write), .o(net78));
ml_powersurg_buf I168 ( .in(net72), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout1_mux), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_41_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_40_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_39_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_38_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_37_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_36_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_35_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_34_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_33_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_32_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_31_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_30_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_29_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_28_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_27_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_26_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net78), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net70));
ml_blsa_sch Iml_blsa_sch_25_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_24_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_23_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_22_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_21_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_20_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_19_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_18_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[14]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[15]),
     .dataout(dataout[15]), .cram_prec(net72));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[13]),
     .data_muxsel(data_muxsel), .cram_write(net74), .bl(bl[14]),
     .dataout(dataout[14]), .cram_prec(net72));

endmodule
// Library - xpmem, Cell - ml_blsa_tile, View - schematic
// LAST TIME SAVED: Sep  5 14:53:52 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tile ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [53:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [53:0]  dataout;

wire  [13:0]  ck;



ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
inv_hvt I172 ( .A(net48), .Y(data_out));
inv_hvt I171 ( .A(dataout[53]), .Y(net48));
ml_powersurg_buf I161 ( .in(cram_write), .o(net53));
ml_powersurg_buf I165 ( .in(net57), .o(net55));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net57));
ml_powersurg_buf I163 ( .in(net55), .o(net59));
ml_powersurg_buf I162 ( .in(net65), .o(net61));
ml_powersurg_buf I169 ( .in(net61), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net53), .o(net65));
ml_powersurg_buf I168 ( .in(net59), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_47_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[47]),
     .dataout(dataout[47]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_46_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[46]),
     .dataout(dataout[46]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_45_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[45]),
     .dataout(dataout[45]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_44_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[44]),
     .dataout(dataout[44]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_43_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[43]),
     .dataout(dataout[43]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_42_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[42]),
     .dataout(dataout[42]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_41_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_40_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_39_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_38_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_37_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_36_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_35_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_34_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_33_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_32_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net55));
ml_blsa_sch I170_53_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[52]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[53]),
     .dataout(dataout[53]), .cram_prec(net57));
ml_blsa_sch I170_52_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[51]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[52]),
     .dataout(dataout[52]), .cram_prec(net57));
ml_blsa_sch I170_51_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[50]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[51]),
     .dataout(dataout[51]), .cram_prec(net57));
ml_blsa_sch I170_50_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[49]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[50]),
     .dataout(dataout[50]), .cram_prec(net57));
ml_blsa_sch I170_49_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[48]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[49]),
     .dataout(dataout[49]), .cram_prec(net57));
ml_blsa_sch I170_48_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[47]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[48]),
     .dataout(dataout[48]), .cram_prec(net57));
ml_blsa_sch Iml_blsa_sch_31_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_30_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_29_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_28_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_27_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_26_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_25_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_24_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_23_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_22_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_21_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_20_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_19_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_18_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net59));

endmodule
// Library - xpmem, Cell - ml_blprecwrt_en, View - schematic
// LAST TIME SAVED: May 16 10:09:58 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blprecwrt_en ( data_out, action, clkin, data_in, rst );
output  data_out;

input  action, clkin, data_in, rst;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I161 ( .A(net89), .Y(net88));
inv_hvt I162 ( .A(action), .Y(net86));
inv_hvt I165 ( .A(net98), .Y(data_out));
nand3_hvt I160 ( .Y(net89), .B(data_in), .C(action), .A(clkin));
nor2_hvt I385 ( .A(net88), .B(net94), .Y(net98));
nor3_hvt I387 ( .B(net86), .Y(net94), .A(net98), .C(rst));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_bram, View - schematic
// LAST TIME SAVED: Jun 26 18:10:51 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2_bram ( data_out, latch_clock_out, para_out,
     prec_out, wrt_out, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, datain, latch_clock_in, latch_reset,
     para_en, para_in, prec_in, smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, para_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, para_en, para_in, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in;

inout [95:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile_bram Iml_blsa_tile_0 ( .para_en(para_en),
     .para_in(para_in), .para_out(para_out), .bl(bl[41:0]),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[95:42]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
inv_hvt I183 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I184 ( .A(smc_wdic_clk), .Y(net088));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_buf_ice5, View - schematic
// LAST TIME SAVED: Aug 13 13:53:01 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_buf_ice5 ( o, in, sel );
output  o;

input  in, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));
inv_hvt I391 ( .A(net77), .Y(o));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_last, View - schematic
// LAST TIME SAVED: Sep  2 16:23:45 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tile_last ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [17:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:0]  ck;

wire  [17:0]  dataout;



tiehi I185 ( .tiehi(net040));
ml_dff_bl Idff ( .R(latch_reset), .D(dataout[16]), .CLK(ck[0]),
     .QN(net50), .Q(net45));
ml_dff_bl I179 ( .R(latch_reset), .D(net58), .CLK(ck[0]), .QN(net49),
     .Q(net61));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_buf_ice5 I205 ( .in(net61), .o(data_out), .sel(net040));
mux2_hvt I174 ( .in1(net45), .in0(dataout[17]), .out(net58),
     .sel(data_muxsel));
ml_powersurg_buf I169 ( .in(cram_write), .o(cram_write_out));
ml_powersurg_buf I168 ( .in(cram_prec), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[16]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[17]), .dataout(dataout[17]));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[15]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[16]), .dataout(dataout[16]));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_last, View - schematic
// LAST TIME SAVED: Aug  9 18:13:45 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2_last ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [125:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_1 ( .latch_reset(latch_reset_buf),
     .datain(data_tile), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_1st),
     .cram_prec(prec_en_1st), .data_out(datain_io),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[107:54]), .latch_clock(latch_clock_out),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blsa_tile Iml_blsa_tile_0 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_dic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
ml_blsa_tile_last Iml_blsa_tile_last ( .bl(bl[125:108]),
     .latch_reset(latch_reset_buf), .datain(datain_io),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_1st), .cram_prec_out(prec_en_1st),
     .latch_clock(latch_clock_out), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
inv_hvt I185 ( .A(smc_wdic_clk), .Y(net091));
inv_hvt I184 ( .A(net091), .Y(smc_dic_clk_buf));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_1st, View - schematic
// LAST TIME SAVED: Sep  6 14:29:58 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tile_1st ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [55:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:4]  data_dummy_in;

wire  [1:5]  data_in;

wire  [0:55]  dataout;

wire  [0:14]  ck;



ml_dff_bl I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net132), .Q(net154));
ml_dff_bl I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net137), .Q(data_dummy_in[4]));
ml_dff_bl I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net142), .Q(data_dummy_in[2]));
ml_dff_bl I179 ( .R(latch_reset), .D(datain), .CLK(ck[14]),
     .QN(net147), .Q(data_dummy_in[1]));
ml_dff_bl I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net152), .Q(data_dummy_in[3]));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_blsa_sch Iml_blsa_sch_15_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[14]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_14_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[13]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_13_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[12]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_12_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[11]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_11_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[10]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_10_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[9]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_9_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[8]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_8_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[7]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_7_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[6]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_6_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_5_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_4_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[4]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_3_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[3]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_2_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[2]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_1_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[1]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_0_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(datain), .cram_prec(cram_prec_out),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_47_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[47]),
     .dataout(dataout[47]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_46_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[46]),
     .dataout(dataout[46]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_45_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[45]),
     .dataout(dataout[45]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_44_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[44]),
     .dataout(dataout[44]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_43_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[43]),
     .dataout(dataout[43]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_42_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[42]),
     .dataout(dataout[42]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_41_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[41]),
     .dataout(dataout[41]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_40_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[40]),
     .dataout(dataout[40]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_39_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[39]),
     .dataout(dataout[39]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_38_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[38]),
     .dataout(dataout[38]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_37_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[37]),
     .dataout(dataout[37]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_36_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[36]),
     .dataout(dataout[36]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_35_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[35]),
     .dataout(dataout[35]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_34_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[34]),
     .dataout(dataout[34]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_33_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[33]),
     .dataout(dataout[33]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_32_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[32]),
     .dataout(dataout[32]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_55_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[54]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[55]),
     .dataout(dataout[55]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_54_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[53]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[54]),
     .dataout(dataout[54]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_53_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[53]),
     .dataout(dataout[53]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_52_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[52]),
     .dataout(dataout[52]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_51_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[51]),
     .dataout(dataout[51]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_50_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[50]),
     .dataout(dataout[50]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_49_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[49]),
     .dataout(dataout[49]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_48_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[48]),
     .dataout(dataout[48]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_31_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[31]),
     .dataout(dataout[31]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_30_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[30]),
     .dataout(dataout[30]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_29_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[29]),
     .dataout(dataout[29]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_28_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[28]),
     .dataout(dataout[28]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_27_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[27]),
     .dataout(dataout[27]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_26_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[26]),
     .dataout(dataout[26]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_25_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[25]),
     .dataout(dataout[25]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_24_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[24]),
     .dataout(dataout[24]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_23_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[23]),
     .dataout(dataout[23]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_22_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[22]),
     .dataout(dataout[22]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_21_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[21]),
     .dataout(dataout[21]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_20_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[20]),
     .dataout(dataout[20]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_19_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[19]),
     .dataout(dataout[19]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_18_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[18]),
     .dataout(dataout[18]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_17_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[17]),
     .dataout(dataout[17]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_16_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[16]),
     .dataout(dataout[16]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_powersurg_buf I161 ( .in(cram_write), .o(net104));
ml_powersurg_buf I165 ( .in(net108), .o(net106));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net108));
ml_powersurg_buf I163 ( .in(net106), .o(net110));
ml_powersurg_buf I162 ( .in(net116), .o(net112));
ml_powersurg_buf I169 ( .in(net112), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net104), .o(net116));
ml_powersurg_buf I168 ( .in(net110), .o(cram_prec_out));
inv_hvt I171 ( .A(dataout[55]), .Y(net121));
inv_hvt I172 ( .A(net121), .Y(data_out));
inv_hvt I224 ( .A(net0130), .Y(ck[14]));
inv_hvt I225 ( .A(net0129), .Y(net0130));
inv_hvt I226 ( .A(net0126), .Y(net0129));
inv_hvt I229 ( .A(latch_clock), .Y(net0122));
inv_hvt I227 ( .A(net0124), .Y(net0126));
inv_hvt I228 ( .A(net0122), .Y(net0124));
mux2_hvt I197 ( .in1(net154), .in0(dataout[4]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I185 ( .in1(data_dummy_in[2]), .in0(dataout[1]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I193 ( .in1(data_dummy_in[4]), .in0(dataout[3]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I180 ( .in1(data_dummy_in[1]), .in0(dataout[0]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I188 ( .in1(data_dummy_in[3]), .in0(dataout[2]),
     .out(data_in[3]), .sel(data_muxsel1));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_1st, View - schematic
// LAST TIME SAVED: Aug 13 13:56:25 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2_1st ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [109:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I186 ( .A(data_muxsel), .Y(net55));
inv_hvt I187 ( .A(net55), .Y(data_muxsel_buf));
inv_hvt I190 ( .A(net61), .Y(cram_pullup_buf));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net61));
inv_hvt I198 ( .A(smc_wdic_clk), .Y(net63));
inv_hvt I199 ( .A(net63), .Y(smc_wdic_clk_buf));
inv_hvt I197 ( .A(latch_clock_in), .Y(net67));
inv_hvt I196 ( .A(net67), .Y(latch_clock_out));
inv_hvt I194 ( .A(latch_reset), .Y(net71));
inv_hvt I195 ( .A(net71), .Y(latch_reset_buf));
ml_blsa_tile_1st Iml_blsa_tile_1st_0 ( .bl(bl[55:0]),
     .cram_pullup_b(cram_pullup_buf), .latch_clock(latch_clock_out),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .datain(datain), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_mid),
     .cram_prec(prec_en_mid), .data_out(data_tile),
     .cram_write_out(wrt_en_last), .cram_prec_out(prec_en_last));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_wdic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[109:56]));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2, View - schematic
// LAST TIME SAVED: Jun 29 11:04:00 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2 ( data_out, latch_clock_out, prec_out, wrt_out,
     bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [107:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_0 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[107:54]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
inv_hvt I183 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I184 ( .A(smc_wdic_clk), .Y(net088));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile, View - schematic
// LAST TIME SAVED: Aug 15 11:21:19 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_rowdrv_tile ( pgate, por_rst_out, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  por_rst_out, smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  vddctrl;
output [15:0]  reset;
output [15:0]  pgate;
output [15:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



inv_hvt I207 ( .A(net041), .Y(por_rst_out));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I194 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I195 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I198 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I190 ( .A(net037), .Y(smc_rsr_1st_out));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net037));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I200 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I206 ( .A(net047), .Y(rsr_rst_buf));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_15_ ( .reset(reset[15]), .wl(wl[15]),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[14]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[15]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_bank, View - schematic
// LAST TIME SAVED: Sep  8 14:09:47 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_blsa_bank ( cm_sdo_u, bl, banksel, cm_sdi_u, cor_en_8bpcfg_b,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     latch_reset, smc_clk, smc_wdic_clk );


input  banksel, cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk;

output [1:0]  cm_sdo_u;

inout [655:0]  bl;

input [1:0]  cm_sdi_u;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



tiehi I267 ( .tiehi(net0256));
tiehi I268 ( .tiehi(net0135));
tiehi I272 ( .tiehi(net0136));
tiehi I271 ( .tiehi(net0132));
tiehi I273 ( .tiehi(net0126));
tiehi I270 ( .tiehi(net0133));
tiehi I269 ( .tiehi(net0134));
ml_dff_bl I146 ( .R(latch_reset_buf), .D(para_out), .CLK(smc_clk),
     .QN(net155), .Q(net176));
ml_blsa_tilex2_bram Itile_67 ( .para_en(cor_en_8bpcfg_buf),
     .para_in(sdi1_buf), .para_out(para_out), .bl(bl[421:326]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net315),
     .latch_clock_out(net138), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret), .wrt_in(wrt_out_89),
     .prec_in(prec_out_89), .latch_reset(latch_reset_buf),
     .datain(data_out_45), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_67),
     .prec_out(prec_out_67), .data_out(data_out_67));
nor2_hvt I254 ( .B(net163), .Y(net164), .A(cram_pullup_b));
inv_hvt I253 ( .A(cor_en_8bpcfg_b), .Y(net161));
inv_hvt I256 ( .A(banksel), .Y(net163));
inv_hvt I255 ( .A(net164), .Y(cram_pullup_logic_b));
inv_hvt I189 ( .A(smc_clk), .Y(net167));
ml_buf_ice5 I247 ( .in(cm_sdi_u[1]), .o(sdi1_buf), .sel(net0136));
ml_buf_ice5 I249 ( .in(net161), .o(cor_en_8bpcfg_buf), .sel(net0136));
ml_buf_ice5 I265 ( .in(net0136), .o(cm_sdo_u[0]), .sel(net176));
ml_buf_ice5 I257 ( .in(smc_wdic_clk), .o(smc_wdic_clk_buf),
     .sel(banksel));
ml_buf_ice5 I203 ( .in(data_muxsel1), .o(data_muxsel1_buf),
     .sel(banksel));
ml_buf_ice5 I205 ( .in(latch_reset), .o(latch_reset_buf),
     .sel(net0126));
ml_buf_ice5 I207 ( .in(cram_write), .o(cram_write_buf), .sel(banksel));
ml_buf_ice5 I208 ( .in(cram_pullup_logic_b), .o(cram_pullup_b_buf),
     .sel(cram_pullup_logic_b));
ml_buf_ice5 I201 ( .in(cram_prec), .o(cram_prec_buf), .sel(banksel));
ml_buf_ice5 I216 ( .in(net0132), .o(net196), .sel(net0132));
ml_buf_ice5 I245 ( .in(cm_sdi_u[0]), .o(sdi0_buf), .sel(net0136));
ml_buf_ice5 I187 ( .in(smc_clk), .o(smc_clk_buf), .sel(smc_clk));
ml_buf_ice5 I188 ( .in(net167), .o(smc_clk_buf_b_ret), .sel(net167));
ml_buf_ice5 I204 ( .in(data_muxsel), .o(data_muxsel_buf),
     .sel(banksel));
ml_buf_ice5 I227 ( .in(net0134), .o(net211), .sel(net0134));
nor3_hvt I217 ( .B(net0133), .Y(net214), .A(net0133), .C(net0133));
nor3_hvt I220 ( .B(net222), .Y(net218), .A(net222), .C(net222));
nor3_hvt I218 ( .B(net214), .Y(net222), .A(net214), .C(net214));
nand3_hvt I231 ( .Y(net225), .B(net229), .C(net229), .A(net229));
nand3_hvt I230 ( .Y(net229), .B(net233), .C(net233), .A(net233));
nand3_hvt I224 ( .Y(net233), .B(net0135), .C(net0135), .A(net0135));
ml_blsa_tilex2_last Itile_1011 ( .bl(bl[655:530]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(smc_clk),
     .latch_clock_out(net248), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret), .wrt_in(net0256),
     .prec_in(net0256), .latch_reset(latch_reset_buf),
     .datain(data_out_89), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_11),
     .prec_out(prec_out_10), .data_out(cm_sdo_u[1]));
ml_blsa_tilex2_1st Itile_01 ( .bl(bl[109:0]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net298),
     .latch_clock_out(net265), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf), .wrt_in(wrt_out_23),
     .prec_in(prec_out_23), .latch_reset(latch_reset_buf),
     .datain(sdi0_buf), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_01),
     .prec_out(prec_out_01), .data_out(data_out_01));
ml_blsa_tilex2 Itile_45 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(net138), .latch_clock_out(net281),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf),
     .wrt_in(wrt_out_67), .prec_in(prec_out_67),
     .latch_reset(latch_reset_buf), .datain(data_out_23),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_45), .prec_out(prec_out_45),
     .data_out(data_out_45), .bl(bl[325:218]));
ml_blsa_tilex2 Itile_23 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(net281), .latch_clock_out(net298),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf_b_ret),
     .wrt_in(wrt_out_45), .prec_in(prec_out_45),
     .latch_reset(latch_reset_buf), .datain(data_out_01),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_23), .prec_out(prec_out_23),
     .data_out(data_out_23), .bl(bl[217:110]));
ml_blsa_tilex2 Itile_89 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(net248), .latch_clock_out(net315),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf),
     .wrt_in(wrt_out_11), .prec_in(prec_out_10),
     .latch_reset(latch_reset_buf), .datain(data_out_67),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_89), .prec_out(prec_out_89),
     .data_out(data_out_89), .bl(bl[529:422]));

endmodule
// Library - ice4chip, Cell - CHIP_route_bot, View - schematic
// LAST TIME SAVED: Oct  6 12:08:35 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module CHIP_route_bot ( cm_banksel_blbld1_0_, cm_banksel_blbld_1_,
     cm_clk_blbld, cm_sdi_u1d, cm_sdo_u0d1, cm_sdo_u1d3, cm_sdo_u2d1,
     core_por_b2, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, crst_filterout, data_muxsel1_blbld,
     data_muxsel_blbld, en_8bconfig_b_blbld, j_rst_bl0, last_rsr3,
     monitor_celld4, row_testl1, smc_core_por_bottom1,
     smc_core_por_bottom2, smc_row_incl0, smc_rsr_rstl0,
     smc_wdis_dclk_blbld, smc_writel0, spi_ss_in_bbankd, tck_padl0,
     bl_bot, cm_banksel, cm_banksel_blbrd_2_, cm_clk_blbrd, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2d, cm_sdo_u1d1, core_por_b0, core_por_b_rowu2,
     core_por_bb, core_por_rowu0, cram_pgateoff, cram_prec,
     cram_prec_blbrd, cram_pullup_b, cram_pullup_b_blbrd, cram_rst,
     cram_vddoff, cram_wl_en, cram_write, cram_write_blbrd,
     creset_b_int, data_muxsel, data_muxsel1, data_muxsel1_blbrd,
     data_muxsel_blbrd, en_8bconfig_b, en_8bconfig_b_blbrd, j_rst_b,
     j_tck, last_rsr1, monitor_celld2, row_test0, smc_clk_out,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk, smc_wdis_dclk_blbrd,
     smc_write, spi_ss_in_bbank, vddio_botbank, vddio_spi );
output  cm_banksel_blbld1_0_, cm_banksel_blbld_1_, cm_clk_blbld,
     core_por_b2, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, crst_filterout, data_muxsel1_blbld,
     data_muxsel_blbld, en_8bconfig_b_blbld, j_rst_bl0, last_rsr3,
     row_testl1, smc_core_por_bottom1, smc_core_por_bottom2,
     smc_row_incl0, smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0,
     tck_padl0;


input  cm_banksel_blbrd_2_, cm_clk_blbrd, core_por_b0,
     core_por_b_rowu2, core_por_bb, core_por_rowu0, cram_pgateoff,
     cram_prec, cram_prec_blbrd, cram_pullup_b, cram_pullup_b_blbrd,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, cram_write_blbrd,
     creset_b_int, data_muxsel, data_muxsel1, data_muxsel1_blbrd,
     data_muxsel_blbrd, en_8bconfig_b, en_8bconfig_b_blbrd, j_rst_b,
     j_tck, last_rsr1, row_test0, smc_clk_out, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk, smc_wdis_dclk_blbrd, smc_write,
     vddio_botbank, vddio_spi;

output [1:0]  cm_sdo_u1d3;
output [1:0]  monitor_celld4;
output [1:0]  cm_sdi_u1d;
output [1:0]  cm_sdo_u2d1;
output [4:0]  spi_ss_in_bbankd;
output [1:0]  cm_sdo_u0d1;

inout [1311:0]  bl_bot;

input [1:0]  cm_sdi_u1;
input [1:0]  monitor_celld2;
input [1:0]  cm_sdi_u2d;
input [1:0]  cm_banksel;
input [4:0]  spi_ss_in_bbank;
input [1:0]  cm_sdi_u0;
input [1:0]  cm_sdo_u1d1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u2;

wire  [1:0]  dff_u2_d1;

wire  [1:0]  monitor_celld3;

wire  [1:0]  dff_u1_d1;

wire  [1:0]  cm_sdo_u1_buf;

wire  [1:0]  cm_sdo_u0_buf;

wire  [1:0]  dff_u0_d1;

wire  [1:0]  cm_sdo_u0;

wire  [1:0]  dff_u0_d0;

wire  [1:0]  cm_sdi_u0d1;

wire  [2:2]  cm_banksel_blbrd1;

wire  [1:0]  dff_u2_d0;

wire  [1:0]  cm_sdi_u2d_buf;

wire  [0:1]  net0200;

wire  [0:1]  net0278;

wire  [0:1]  net0376;

wire  [0:1]  net0372;

wire  [0:1]  net0260;

wire  [0:1]  net0254;

wire  [0:1]  net0388;

wire  [0:1]  net0380;

wire  [0:1]  net0384;



eh_io_pup_2_new I4 ( .core_por_b(core_por_b0), .vdd_io(vddio_botbank),
     .por_b(smc_core_por_bottom1));
eh_io_pup_2_new I5 ( .core_por_b(core_por_b0), .vdd_io(vddio_spi),
     .por_b(smc_core_por_bottom2));
tielo I559_1_ ( .tielo(net0372[0]));
tielo I559_0_ ( .tielo(net0372[1]));
tielo I562_1_ ( .tielo(net0376[0]));
tielo I562_0_ ( .tielo(net0376[1]));
tielo I564 ( .tielo(net0392));
tielo I563_1_ ( .tielo(net0384[0]));
tielo I563_0_ ( .tielo(net0384[1]));
tielo I560_1_ ( .tielo(net0380[0]));
tielo I560_0_ ( .tielo(net0380[1]));
tielo I561_1_ ( .tielo(net0388[0]));
tielo I561_0_ ( .tielo(net0388[1]));
sg_bufx10bot I531_1_ ( .in(net0200[0]), .out(net0278[0]));
sg_bufx10bot I531_0_ ( .in(net0200[1]), .out(net0278[1]));
sg_bufx10bot I175 ( .in(net272), .out(data_muxsel_blbld));
sg_bufx10bot I333 ( .in(j_rst_b), .out(j_rst_bl0));
sg_bufx10bot I486 ( .in(net270), .out(cram_prec_blbld));
sg_bufx10bot I492 ( .in(net268), .out(cram_write_blbld));
sg_bufx10bot I474 ( .in(net302), .out(net312));
sg_bufx10bot I496 ( .in(en_8bconfig_b_blbrd),
     .out(predata_en_8bconfig_b));
sg_bufx10bot I481 ( .in(net318), .out(cram_rstl0));
sg_bufx10bot I495 ( .in(net264), .out(en_8bconfig_b_blbld));
sg_bufx10bot I467 ( .in(predata_muxsel1), .out(net260));
sg_bufx10bot I466 ( .in(net260), .out(data_muxsel1_blbld));
sg_bufx10bot I429_1_ ( .in(monitor_celld3[1]),
     .out(monitor_celld4[1]));
sg_bufx10bot I429_0_ ( .in(monitor_celld3[0]),
     .out(monitor_celld4[0]));
sg_bufx10bot I523 ( .in(smc_clk_mid), .out(cm_clk_blbld));
sg_bufx10bot I489 ( .in(net256), .out(cram_pullup_blbld));
sg_bufx10bot I485 ( .in(cram_prec), .out(predata_cram_prec));
sg_bufx10bot I487 ( .in(predata_cram_prec), .out(net270));
sg_bufx10bot I533_1_ ( .in(cm_sdi_u1[1]), .out(net0200[0]));
sg_bufx10bot I533_0_ ( .in(cm_sdi_u1[0]), .out(net0200[1]));
sg_bufx10bot I527_1_ ( .in(cm_sdi_u0[1]), .out(net0260[0]));
sg_bufx10bot I527_0_ ( .in(cm_sdi_u0[0]), .out(net0260[1]));
sg_bufx10bot I520 ( .in(net282), .out(net280));
sg_bufx10bot I517 ( .in(net250), .out(net206));
sg_bufx10bot I493 ( .in(predata_cram_write), .out(net268));
sg_bufx10bot I505 ( .in(net248), .out(smc_rsr_rstl0));
sg_bufx10bot I509 ( .in(net246), .out(row_testl1));
sg_bufx10bot I519 ( .in(cm_banksel[0]), .out(net282));
sg_bufx10bot I491 ( .in(cram_write), .out(predata_cram_write));
sg_bufx10bot I504 ( .in(smc_rsr_rst), .out(net298));
sg_bufx10bot I494 ( .in(predata_en_8bconfig_b), .out(net264));
sg_bufx10bot I529_1_ ( .in(net0254[0]), .out(cm_sdi_u0d1[1]));
sg_bufx10bot I529_0_ ( .in(net0254[1]), .out(cm_sdi_u0d1[0]));
sg_bufx10bot I476 ( .in(net236), .out(cram_vddoffl0));
sg_bufx10bot I479 ( .in(cram_rst), .out(net214));
sg_bufx10bot I530_1_ ( .in(net0260[0]), .out(net0254[0]));
sg_bufx10bot I530_0_ ( .in(net0260[1]), .out(net0254[1]));
sg_bufx10bot I439 ( .in(j_tck), .out(tck_padl0));
sg_bufx10bot I510 ( .in(net276), .out(net246));
sg_bufx10bot I482 ( .in(net228), .out(cram_pgateoffl0));
sg_bufx10bot I483 ( .in(net226), .out(net228));
sg_bufx10bot I464 ( .in(predata_muxsel), .out(net272));
sg_bufx10bot I525 ( .in(cm_clk_blbrd), .out(predata_smc_clk_out));
sg_bufx10bot I503 ( .in(net298), .out(net248));
sg_bufx10bot I490 ( .in(cram_pullup_b), .out(predata_cram_pullup_b));
sg_bufx10bot I532_1_ ( .in(net0278[0]), .out(cm_sdi_u1d[1]));
sg_bufx10bot I532_0_ ( .in(net0278[1]), .out(cm_sdi_u1d[0]));
sg_bufx10bot I521 ( .in(net280), .out(cm_banksel_blbld1_0_));
sg_bufx10bot I465 ( .in(data_muxsel1_blbrd), .out(predata_muxsel1));
sg_bufx10bot I484 ( .in(cram_pgateoff), .out(net226));
sg_bufx10bot I480 ( .in(net214), .out(net318));
sg_bufx10bot I518 ( .in(cm_banksel[1]), .out(net250));
sg_bufx10bot I488 ( .in(predata_cram_pullup_b), .out(net256));
sg_bufx10bot I524 ( .in(predata_smc_clk_out), .out(smc_clk_mid));
sg_bufx10bot I516 ( .in(net206), .out(cm_banksel_blbld_1_));
sg_bufx10bot I470 ( .in(net204), .out(cram_wl_enl0));
sg_bufx10bot I293 ( .in(last_rsr1), .out(last_rsr2));
sg_bufx10bot I541_1_ ( .in(dff_u0_d1[1]), .out(cm_sdo_u0d1[1]));
sg_bufx10bot I541_0_ ( .in(dff_u0_d1[0]), .out(cm_sdo_u0d1[0]));
sg_bufx10bot I539_1_ ( .in(cm_sdo_u1d1[1]), .out(cm_sdo_u1_buf[1]));
sg_bufx10bot I539_0_ ( .in(cm_sdo_u1d1[0]), .out(cm_sdo_u1_buf[0]));
sg_bufx10bot I455 ( .in(data_muxsel_blbrd), .out(predata_muxsel));
sg_bufx10bot I475 ( .in(net312), .out(smc_writel0));
sg_bufx10bot I526_1_ ( .in(cm_sdi_u2d[1]), .out(cm_sdi_u2d_buf[1]));
sg_bufx10bot I526_0_ ( .in(cm_sdi_u2d[0]), .out(cm_sdi_u2d_buf[0]));
sg_bufx10bot I459 ( .in(smc_row_inc), .out(net316));
sg_bufx10bot I477 ( .in(net292), .out(net236));
sg_bufx10bot I543_1_ ( .in(dff_u0_d0[1]), .out(cm_sdo_u0_buf[1]));
sg_bufx10bot I543_0_ ( .in(dff_u0_d0[0]), .out(cm_sdo_u0_buf[0]));
sg_bufx10bot I469 ( .in(net274), .out(smc_row_incl0));
sg_bufx10bot I522 ( .in(cm_banksel_blbrd_2_),
     .out(cm_banksel_blbrd1[2]));
sg_bufx10bot I427_1_ ( .in(monitor_celld2[1]),
     .out(monitor_celld3[1]));
sg_bufx10bot I427_0_ ( .in(monitor_celld2[0]),
     .out(monitor_celld3[0]));
sg_bufx10bot I540_1_ ( .in(dff_u1_d1[1]), .out(cm_sdo_u1d3[1]));
sg_bufx10bot I540_0_ ( .in(dff_u1_d1[0]), .out(cm_sdo_u1d3[0]));
sg_bufx10bot I473 ( .in(smc_write), .out(net302));
sg_bufx10bot I542 ( .in(net374), .out(last_rsr3));
sg_bufx10bot I497 ( .in(smc_wdis_dclk_blbrd),
     .out(predata_smc_wdis_dclk));
sg_bufx10bot I511 ( .in(row_test0), .out(net276));
sg_bufx10bot I498 ( .in(net324), .out(smc_wdis_dclk_blbld));
sg_bufx10bot I471 ( .in(net278), .out(net204));
sg_bufx10bot I499 ( .in(predata_smc_wdis_dclk), .out(net324));
sg_bufx10bot I330 ( .in(net316), .out(net274));
sg_bufx10bot I478 ( .in(cram_vddoff), .out(net292));
sg_bufx10bot I336 ( .in(core_por_bb), .out(core_por_bbl0));
sg_bufx10bot I472 ( .in(cram_wl_en), .out(net278));
creset_filter I141 ( .in(creset_b_int), .out(crst_filterout));
ml_blsa_bank Iblbr ( .smc_wdic_clk(predata_smc_wdis_dclk),
     .smc_clk(predata_smc_clk_out), .cm_sdi_u(cm_sdi_u2d_buf[1:0]),
     .latch_reset(core_por_b_rowu2), .cm_sdo_u(cm_sdo_u2[1:0]),
     .data_muxsel1(predata_muxsel1), .data_muxsel(predata_muxsel),
     .cram_write(predata_cram_write), .cram_prec(predata_cram_prec),
     .cor_en_8bpcfg_b(predata_en_8bconfig_b),
     .cram_pullup_b(predata_cram_pullup_b),
     .banksel(cm_banksel_blbrd1[2]), .bl(bl_bot[1311:656]));
ml_blsa_bank Iblbl ( .smc_wdic_clk(smc_wdis_dclk_blbld),
     .smc_clk(cm_clk_blbld), .cm_sdi_u(cm_sdi_u0d1[1:0]),
     .latch_reset(core_por_rowu0), .cm_sdo_u(cm_sdo_u0[1:0]),
     .data_muxsel1(data_muxsel1_blbld),
     .data_muxsel(data_muxsel_blbld), .cram_write(cram_write_blbld),
     .cram_prec(cram_prec_blbld),
     .cor_en_8bpcfg_b(en_8bconfig_b_blbld),
     .cram_pullup_b(cram_pullup_blbld), .banksel(cm_banksel_blbld1_0_),
     .bl({bl_bot[0], bl_bot[1], bl_bot[2], bl_bot[3], bl_bot[4],
     bl_bot[5], bl_bot[6], bl_bot[7], bl_bot[8], bl_bot[9], bl_bot[10],
     bl_bot[11], bl_bot[12], bl_bot[13], bl_bot[14], bl_bot[15],
     bl_bot[16], bl_bot[17], bl_bot[18], bl_bot[19], bl_bot[20],
     bl_bot[21], bl_bot[22], bl_bot[23], bl_bot[24], bl_bot[25],
     bl_bot[26], bl_bot[27], bl_bot[28], bl_bot[29], bl_bot[30],
     bl_bot[31], bl_bot[32], bl_bot[33], bl_bot[34], bl_bot[35],
     bl_bot[36], bl_bot[37], bl_bot[38], bl_bot[39], bl_bot[40],
     bl_bot[41], bl_bot[42], bl_bot[43], bl_bot[44], bl_bot[45],
     bl_bot[46], bl_bot[47], bl_bot[48], bl_bot[49], bl_bot[50],
     bl_bot[51], bl_bot[52], bl_bot[53], bl_bot[54], bl_bot[55],
     bl_bot[56], bl_bot[57], bl_bot[58], bl_bot[59], bl_bot[60],
     bl_bot[61], bl_bot[62], bl_bot[63], bl_bot[64], bl_bot[65],
     bl_bot[66], bl_bot[67], bl_bot[68], bl_bot[69], bl_bot[70],
     bl_bot[71], bl_bot[72], bl_bot[73], bl_bot[74], bl_bot[75],
     bl_bot[76], bl_bot[77], bl_bot[78], bl_bot[79], bl_bot[80],
     bl_bot[81], bl_bot[82], bl_bot[83], bl_bot[84], bl_bot[85],
     bl_bot[86], bl_bot[87], bl_bot[88], bl_bot[89], bl_bot[90],
     bl_bot[91], bl_bot[92], bl_bot[93], bl_bot[94], bl_bot[95],
     bl_bot[96], bl_bot[97], bl_bot[98], bl_bot[99], bl_bot[100],
     bl_bot[101], bl_bot[102], bl_bot[103], bl_bot[104], bl_bot[105],
     bl_bot[106], bl_bot[107], bl_bot[108], bl_bot[109], bl_bot[110],
     bl_bot[111], bl_bot[112], bl_bot[113], bl_bot[114], bl_bot[115],
     bl_bot[116], bl_bot[117], bl_bot[118], bl_bot[119], bl_bot[120],
     bl_bot[121], bl_bot[122], bl_bot[123], bl_bot[124], bl_bot[125],
     bl_bot[126], bl_bot[127], bl_bot[128], bl_bot[129], bl_bot[130],
     bl_bot[131], bl_bot[132], bl_bot[133], bl_bot[134], bl_bot[135],
     bl_bot[136], bl_bot[137], bl_bot[138], bl_bot[139], bl_bot[140],
     bl_bot[141], bl_bot[142], bl_bot[143], bl_bot[144], bl_bot[145],
     bl_bot[146], bl_bot[147], bl_bot[148], bl_bot[149], bl_bot[150],
     bl_bot[151], bl_bot[152], bl_bot[153], bl_bot[154], bl_bot[155],
     bl_bot[156], bl_bot[157], bl_bot[158], bl_bot[159], bl_bot[160],
     bl_bot[161], bl_bot[162], bl_bot[163], bl_bot[164], bl_bot[165],
     bl_bot[166], bl_bot[167], bl_bot[168], bl_bot[169], bl_bot[170],
     bl_bot[171], bl_bot[172], bl_bot[173], bl_bot[174], bl_bot[175],
     bl_bot[176], bl_bot[177], bl_bot[178], bl_bot[179], bl_bot[180],
     bl_bot[181], bl_bot[182], bl_bot[183], bl_bot[184], bl_bot[185],
     bl_bot[186], bl_bot[187], bl_bot[188], bl_bot[189], bl_bot[190],
     bl_bot[191], bl_bot[192], bl_bot[193], bl_bot[194], bl_bot[195],
     bl_bot[196], bl_bot[197], bl_bot[198], bl_bot[199], bl_bot[200],
     bl_bot[201], bl_bot[202], bl_bot[203], bl_bot[204], bl_bot[205],
     bl_bot[206], bl_bot[207], bl_bot[208], bl_bot[209], bl_bot[210],
     bl_bot[211], bl_bot[212], bl_bot[213], bl_bot[214], bl_bot[215],
     bl_bot[216], bl_bot[217], bl_bot[218], bl_bot[219], bl_bot[220],
     bl_bot[221], bl_bot[222], bl_bot[223], bl_bot[224], bl_bot[225],
     bl_bot[226], bl_bot[227], bl_bot[228], bl_bot[229], bl_bot[230],
     bl_bot[231], bl_bot[232], bl_bot[233], bl_bot[234], bl_bot[235],
     bl_bot[236], bl_bot[237], bl_bot[238], bl_bot[239], bl_bot[240],
     bl_bot[241], bl_bot[242], bl_bot[243], bl_bot[244], bl_bot[245],
     bl_bot[246], bl_bot[247], bl_bot[248], bl_bot[249], bl_bot[250],
     bl_bot[251], bl_bot[252], bl_bot[253], bl_bot[254], bl_bot[255],
     bl_bot[256], bl_bot[257], bl_bot[258], bl_bot[259], bl_bot[260],
     bl_bot[261], bl_bot[262], bl_bot[263], bl_bot[264], bl_bot[265],
     bl_bot[266], bl_bot[267], bl_bot[268], bl_bot[269], bl_bot[270],
     bl_bot[271], bl_bot[272], bl_bot[273], bl_bot[274], bl_bot[275],
     bl_bot[276], bl_bot[277], bl_bot[278], bl_bot[279], bl_bot[280],
     bl_bot[281], bl_bot[282], bl_bot[283], bl_bot[284], bl_bot[285],
     bl_bot[286], bl_bot[287], bl_bot[288], bl_bot[289], bl_bot[290],
     bl_bot[291], bl_bot[292], bl_bot[293], bl_bot[294], bl_bot[295],
     bl_bot[296], bl_bot[297], bl_bot[298], bl_bot[299], bl_bot[300],
     bl_bot[301], bl_bot[302], bl_bot[303], bl_bot[304], bl_bot[305],
     bl_bot[306], bl_bot[307], bl_bot[308], bl_bot[309], bl_bot[310],
     bl_bot[311], bl_bot[312], bl_bot[313], bl_bot[314], bl_bot[315],
     bl_bot[316], bl_bot[317], bl_bot[318], bl_bot[319], bl_bot[320],
     bl_bot[321], bl_bot[322], bl_bot[323], bl_bot[324], bl_bot[325],
     bl_bot[326], bl_bot[327], bl_bot[328], bl_bot[329], bl_bot[330],
     bl_bot[331], bl_bot[332], bl_bot[333], bl_bot[334], bl_bot[335],
     bl_bot[336], bl_bot[337], bl_bot[338], bl_bot[339], bl_bot[340],
     bl_bot[341], bl_bot[342], bl_bot[343], bl_bot[344], bl_bot[345],
     bl_bot[346], bl_bot[347], bl_bot[348], bl_bot[349], bl_bot[350],
     bl_bot[351], bl_bot[352], bl_bot[353], bl_bot[354], bl_bot[355],
     bl_bot[356], bl_bot[357], bl_bot[358], bl_bot[359], bl_bot[360],
     bl_bot[361], bl_bot[362], bl_bot[363], bl_bot[364], bl_bot[365],
     bl_bot[366], bl_bot[367], bl_bot[368], bl_bot[369], bl_bot[370],
     bl_bot[371], bl_bot[372], bl_bot[373], bl_bot[374], bl_bot[375],
     bl_bot[376], bl_bot[377], bl_bot[378], bl_bot[379], bl_bot[380],
     bl_bot[381], bl_bot[382], bl_bot[383], bl_bot[384], bl_bot[385],
     bl_bot[386], bl_bot[387], bl_bot[388], bl_bot[389], bl_bot[390],
     bl_bot[391], bl_bot[392], bl_bot[393], bl_bot[394], bl_bot[395],
     bl_bot[396], bl_bot[397], bl_bot[398], bl_bot[399], bl_bot[400],
     bl_bot[401], bl_bot[402], bl_bot[403], bl_bot[404], bl_bot[405],
     bl_bot[406], bl_bot[407], bl_bot[408], bl_bot[409], bl_bot[410],
     bl_bot[411], bl_bot[412], bl_bot[413], bl_bot[414], bl_bot[415],
     bl_bot[416], bl_bot[417], bl_bot[418], bl_bot[419], bl_bot[420],
     bl_bot[421], bl_bot[422], bl_bot[423], bl_bot[424], bl_bot[425],
     bl_bot[426], bl_bot[427], bl_bot[428], bl_bot[429], bl_bot[430],
     bl_bot[431], bl_bot[432], bl_bot[433], bl_bot[434], bl_bot[435],
     bl_bot[436], bl_bot[437], bl_bot[438], bl_bot[439], bl_bot[440],
     bl_bot[441], bl_bot[442], bl_bot[443], bl_bot[444], bl_bot[445],
     bl_bot[446], bl_bot[447], bl_bot[448], bl_bot[449], bl_bot[450],
     bl_bot[451], bl_bot[452], bl_bot[453], bl_bot[454], bl_bot[455],
     bl_bot[456], bl_bot[457], bl_bot[458], bl_bot[459], bl_bot[460],
     bl_bot[461], bl_bot[462], bl_bot[463], bl_bot[464], bl_bot[465],
     bl_bot[466], bl_bot[467], bl_bot[468], bl_bot[469], bl_bot[470],
     bl_bot[471], bl_bot[472], bl_bot[473], bl_bot[474], bl_bot[475],
     bl_bot[476], bl_bot[477], bl_bot[478], bl_bot[479], bl_bot[480],
     bl_bot[481], bl_bot[482], bl_bot[483], bl_bot[484], bl_bot[485],
     bl_bot[486], bl_bot[487], bl_bot[488], bl_bot[489], bl_bot[490],
     bl_bot[491], bl_bot[492], bl_bot[493], bl_bot[494], bl_bot[495],
     bl_bot[496], bl_bot[497], bl_bot[498], bl_bot[499], bl_bot[500],
     bl_bot[501], bl_bot[502], bl_bot[503], bl_bot[504], bl_bot[505],
     bl_bot[506], bl_bot[507], bl_bot[508], bl_bot[509], bl_bot[510],
     bl_bot[511], bl_bot[512], bl_bot[513], bl_bot[514], bl_bot[515],
     bl_bot[516], bl_bot[517], bl_bot[518], bl_bot[519], bl_bot[520],
     bl_bot[521], bl_bot[522], bl_bot[523], bl_bot[524], bl_bot[525],
     bl_bot[526], bl_bot[527], bl_bot[528], bl_bot[529], bl_bot[530],
     bl_bot[531], bl_bot[532], bl_bot[533], bl_bot[534], bl_bot[535],
     bl_bot[536], bl_bot[537], bl_bot[538], bl_bot[539], bl_bot[540],
     bl_bot[541], bl_bot[542], bl_bot[543], bl_bot[544], bl_bot[545],
     bl_bot[546], bl_bot[547], bl_bot[548], bl_bot[549], bl_bot[550],
     bl_bot[551], bl_bot[552], bl_bot[553], bl_bot[554], bl_bot[555],
     bl_bot[556], bl_bot[557], bl_bot[558], bl_bot[559], bl_bot[560],
     bl_bot[561], bl_bot[562], bl_bot[563], bl_bot[564], bl_bot[565],
     bl_bot[566], bl_bot[567], bl_bot[568], bl_bot[569], bl_bot[570],
     bl_bot[571], bl_bot[572], bl_bot[573], bl_bot[574], bl_bot[575],
     bl_bot[576], bl_bot[577], bl_bot[578], bl_bot[579], bl_bot[580],
     bl_bot[581], bl_bot[582], bl_bot[583], bl_bot[584], bl_bot[585],
     bl_bot[586], bl_bot[587], bl_bot[588], bl_bot[589], bl_bot[590],
     bl_bot[591], bl_bot[592], bl_bot[593], bl_bot[594], bl_bot[595],
     bl_bot[596], bl_bot[597], bl_bot[598], bl_bot[599], bl_bot[600],
     bl_bot[601], bl_bot[602], bl_bot[603], bl_bot[604], bl_bot[605],
     bl_bot[606], bl_bot[607], bl_bot[608], bl_bot[609], bl_bot[610],
     bl_bot[611], bl_bot[612], bl_bot[613], bl_bot[614], bl_bot[615],
     bl_bot[616], bl_bot[617], bl_bot[618], bl_bot[619], bl_bot[620],
     bl_bot[621], bl_bot[622], bl_bot[623], bl_bot[624], bl_bot[625],
     bl_bot[626], bl_bot[627], bl_bot[628], bl_bot[629], bl_bot[630],
     bl_bot[631], bl_bot[632], bl_bot[633], bl_bot[634], bl_bot[635],
     bl_bot[636], bl_bot[637], bl_bot[638], bl_bot[639], bl_bot[640],
     bl_bot[641], bl_bot[642], bl_bot[643], bl_bot[644], bl_bot[645],
     bl_bot[646], bl_bot[647], bl_bot[648], bl_bot[649], bl_bot[650],
     bl_bot[651], bl_bot[652], bl_bot[653], bl_bot[654],
     bl_bot[655]}));
sg_dffbuf I535_1_ ( .r(net0372[0]), .d(cm_sdo_u0[1]), .clk(net395),
     .dffout(dff_u0_d0[1]));
sg_dffbuf I535_0_ ( .r(net0372[1]), .d(cm_sdo_u0[0]), .clk(net395),
     .dffout(dff_u0_d0[0]));
sg_dffbuf I546_1_ ( .r(net0376[0]), .d(cm_sdo_u2[1]), .clk(net400),
     .dffout(dff_u2_d0[1]));
sg_dffbuf I546_0_ ( .r(net0376[1]), .d(cm_sdo_u2[0]), .clk(net400),
     .dffout(dff_u2_d0[0]));
sg_dffbuf I537_1_ ( .r(net0380[0]), .d(cm_sdo_u1_buf[1]), .clk(net393),
     .dffout(dff_u1_d1[1]));
sg_dffbuf I537_0_ ( .r(net0380[1]), .d(cm_sdo_u1_buf[0]), .clk(net393),
     .dffout(dff_u1_d1[0]));
sg_dffbuf I545_1_ ( .r(net0384[0]), .d(dff_u2_d0[1]), .clk(net401),
     .dffout(dff_u2_d1[1]));
sg_dffbuf I545_0_ ( .r(net0384[1]), .d(dff_u2_d0[0]), .clk(net401),
     .dffout(dff_u2_d1[0]));
sg_dffbuf I462_1_ ( .r(net0388[0]), .d(cm_sdo_u0_buf[1]), .clk(net393),
     .dffout(dff_u0_d1[1]));
sg_dffbuf I462_0_ ( .r(net0388[1]), .d(cm_sdo_u0_buf[0]), .clk(net393),
     .dffout(dff_u0_d1[0]));
sg_dffbuf I512 ( .r(net0392), .d(last_rsr2), .clk(net393),
     .dffout(net374));
bram_bufferx16 I534 ( .in(smc_clk_mid), .out(net393));
bram_bufferx16 I550_1_ ( .in(dff_u2_d1[1]), .out(cm_sdo_u2d1[1]));
bram_bufferx16 I550_0_ ( .in(dff_u2_d1[0]), .out(cm_sdo_u2d1[0]));
bram_bufferx16 I549 ( .in(net400), .out(net401));
bram_bufferx16 I450_4_ ( .in(spi_ss_in_bbank[4]),
     .out(spi_ss_in_bbankd[4]));
bram_bufferx16 I450_3_ ( .in(spi_ss_in_bbank[3]),
     .out(spi_ss_in_bbankd[3]));
bram_bufferx16 I450_2_ ( .in(spi_ss_in_bbank[2]),
     .out(spi_ss_in_bbankd[2]));
bram_bufferx16 I450_1_ ( .in(spi_ss_in_bbank[1]),
     .out(spi_ss_in_bbankd[1]));
bram_bufferx16 I450_0_ ( .in(spi_ss_in_bbank[0]),
     .out(spi_ss_in_bbankd[0]));
bram_bufferx16 I548 ( .in(predata_smc_clk_out), .out(net400));
bram_bufferx16 I536 ( .in(cm_clk_blbld), .out(net395));
bram_bufferx16 I186 ( .in(core_por_b0), .out(core_por_b2));

endmodule
// Library - ice4chip, Cell - CHIP_route_top, View - schematic
// LAST TIME SAVED: Oct  7 17:57:36 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module CHIP_route_top ( cm_sdo_u1, cm_sdo_u3, bl_top,
     cm_banksel_bltld3, cm_banksel_bltrd1, cm_clk_bltld3,
     cm_clk_bltrd1, .cm_prec_bltld3(cram_prec_bltld3), cm_sdi_u1d3,
     cm_sdi_u3d2, core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3,
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1) );


input  cm_clk_bltld3, cm_clk_bltrd1, cram_prec_bltld3,
     core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1;

output [1:0]  cm_sdo_u1;
output [1:0]  cm_sdo_u3;

inout [1311:0]  bl_top;

input [3:3]  cm_banksel_bltrd1;
input [1:1]  cm_banksel_bltld3;
input [1:0]  cm_sdi_u3d2;
input [1:0]  cm_sdi_u1d3;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_bank Ibltr ( .smc_wdic_clk(smc_wdis_dclk_bltrd1),
     .smc_clk(cm_clk_bltrd1), .cm_sdi_u(cm_sdi_u3d2[1:0]),
     .latch_reset(core_por_b_rowu3), .cm_sdo_u(cm_sdo_u3[1:0]),
     .data_muxsel1(data_muxsel1_bltrd1),
     .data_muxsel(data_muxsel_bltrd1), .cram_write(cram_write_bltrd1),
     .cram_prec(cram_prec_bltrd1),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltrd1),
     .cram_pullup_b(cram_pullup_b_bltrd1),
     .banksel(cm_banksel_bltrd1[3]), .bl(bl_top[1311:656]));
ml_blsa_bank Ibltlu1 ( .smc_wdic_clk(smc_wdis_dclk_bltld3),
     .smc_clk(cm_clk_bltld3), .cm_sdi_u(cm_sdi_u1d3[1:0]),
     .latch_reset(core_por_b_rowu1), .cm_sdo_u(cm_sdo_u1[1:0]),
     .data_muxsel1(data_muxsel1_bltld3),
     .data_muxsel(data_muxsel_bltld3), .cram_write(cram_write_bltld3),
     .cram_prec(cram_prec_bltld3),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltld3),
     .cram_pullup_b(cram_pullup_bltld3),
     .banksel(cm_banksel_bltld3[1]), .bl({bl_top[0], bl_top[1],
     bl_top[2], bl_top[3], bl_top[4], bl_top[5], bl_top[6], bl_top[7],
     bl_top[8], bl_top[9], bl_top[10], bl_top[11], bl_top[12],
     bl_top[13], bl_top[14], bl_top[15], bl_top[16], bl_top[17],
     bl_top[18], bl_top[19], bl_top[20], bl_top[21], bl_top[22],
     bl_top[23], bl_top[24], bl_top[25], bl_top[26], bl_top[27],
     bl_top[28], bl_top[29], bl_top[30], bl_top[31], bl_top[32],
     bl_top[33], bl_top[34], bl_top[35], bl_top[36], bl_top[37],
     bl_top[38], bl_top[39], bl_top[40], bl_top[41], bl_top[42],
     bl_top[43], bl_top[44], bl_top[45], bl_top[46], bl_top[47],
     bl_top[48], bl_top[49], bl_top[50], bl_top[51], bl_top[52],
     bl_top[53], bl_top[54], bl_top[55], bl_top[56], bl_top[57],
     bl_top[58], bl_top[59], bl_top[60], bl_top[61], bl_top[62],
     bl_top[63], bl_top[64], bl_top[65], bl_top[66], bl_top[67],
     bl_top[68], bl_top[69], bl_top[70], bl_top[71], bl_top[72],
     bl_top[73], bl_top[74], bl_top[75], bl_top[76], bl_top[77],
     bl_top[78], bl_top[79], bl_top[80], bl_top[81], bl_top[82],
     bl_top[83], bl_top[84], bl_top[85], bl_top[86], bl_top[87],
     bl_top[88], bl_top[89], bl_top[90], bl_top[91], bl_top[92],
     bl_top[93], bl_top[94], bl_top[95], bl_top[96], bl_top[97],
     bl_top[98], bl_top[99], bl_top[100], bl_top[101], bl_top[102],
     bl_top[103], bl_top[104], bl_top[105], bl_top[106], bl_top[107],
     bl_top[108], bl_top[109], bl_top[110], bl_top[111], bl_top[112],
     bl_top[113], bl_top[114], bl_top[115], bl_top[116], bl_top[117],
     bl_top[118], bl_top[119], bl_top[120], bl_top[121], bl_top[122],
     bl_top[123], bl_top[124], bl_top[125], bl_top[126], bl_top[127],
     bl_top[128], bl_top[129], bl_top[130], bl_top[131], bl_top[132],
     bl_top[133], bl_top[134], bl_top[135], bl_top[136], bl_top[137],
     bl_top[138], bl_top[139], bl_top[140], bl_top[141], bl_top[142],
     bl_top[143], bl_top[144], bl_top[145], bl_top[146], bl_top[147],
     bl_top[148], bl_top[149], bl_top[150], bl_top[151], bl_top[152],
     bl_top[153], bl_top[154], bl_top[155], bl_top[156], bl_top[157],
     bl_top[158], bl_top[159], bl_top[160], bl_top[161], bl_top[162],
     bl_top[163], bl_top[164], bl_top[165], bl_top[166], bl_top[167],
     bl_top[168], bl_top[169], bl_top[170], bl_top[171], bl_top[172],
     bl_top[173], bl_top[174], bl_top[175], bl_top[176], bl_top[177],
     bl_top[178], bl_top[179], bl_top[180], bl_top[181], bl_top[182],
     bl_top[183], bl_top[184], bl_top[185], bl_top[186], bl_top[187],
     bl_top[188], bl_top[189], bl_top[190], bl_top[191], bl_top[192],
     bl_top[193], bl_top[194], bl_top[195], bl_top[196], bl_top[197],
     bl_top[198], bl_top[199], bl_top[200], bl_top[201], bl_top[202],
     bl_top[203], bl_top[204], bl_top[205], bl_top[206], bl_top[207],
     bl_top[208], bl_top[209], bl_top[210], bl_top[211], bl_top[212],
     bl_top[213], bl_top[214], bl_top[215], bl_top[216], bl_top[217],
     bl_top[218], bl_top[219], bl_top[220], bl_top[221], bl_top[222],
     bl_top[223], bl_top[224], bl_top[225], bl_top[226], bl_top[227],
     bl_top[228], bl_top[229], bl_top[230], bl_top[231], bl_top[232],
     bl_top[233], bl_top[234], bl_top[235], bl_top[236], bl_top[237],
     bl_top[238], bl_top[239], bl_top[240], bl_top[241], bl_top[242],
     bl_top[243], bl_top[244], bl_top[245], bl_top[246], bl_top[247],
     bl_top[248], bl_top[249], bl_top[250], bl_top[251], bl_top[252],
     bl_top[253], bl_top[254], bl_top[255], bl_top[256], bl_top[257],
     bl_top[258], bl_top[259], bl_top[260], bl_top[261], bl_top[262],
     bl_top[263], bl_top[264], bl_top[265], bl_top[266], bl_top[267],
     bl_top[268], bl_top[269], bl_top[270], bl_top[271], bl_top[272],
     bl_top[273], bl_top[274], bl_top[275], bl_top[276], bl_top[277],
     bl_top[278], bl_top[279], bl_top[280], bl_top[281], bl_top[282],
     bl_top[283], bl_top[284], bl_top[285], bl_top[286], bl_top[287],
     bl_top[288], bl_top[289], bl_top[290], bl_top[291], bl_top[292],
     bl_top[293], bl_top[294], bl_top[295], bl_top[296], bl_top[297],
     bl_top[298], bl_top[299], bl_top[300], bl_top[301], bl_top[302],
     bl_top[303], bl_top[304], bl_top[305], bl_top[306], bl_top[307],
     bl_top[308], bl_top[309], bl_top[310], bl_top[311], bl_top[312],
     bl_top[313], bl_top[314], bl_top[315], bl_top[316], bl_top[317],
     bl_top[318], bl_top[319], bl_top[320], bl_top[321], bl_top[322],
     bl_top[323], bl_top[324], bl_top[325], bl_top[326], bl_top[327],
     bl_top[328], bl_top[329], bl_top[330], bl_top[331], bl_top[332],
     bl_top[333], bl_top[334], bl_top[335], bl_top[336], bl_top[337],
     bl_top[338], bl_top[339], bl_top[340], bl_top[341], bl_top[342],
     bl_top[343], bl_top[344], bl_top[345], bl_top[346], bl_top[347],
     bl_top[348], bl_top[349], bl_top[350], bl_top[351], bl_top[352],
     bl_top[353], bl_top[354], bl_top[355], bl_top[356], bl_top[357],
     bl_top[358], bl_top[359], bl_top[360], bl_top[361], bl_top[362],
     bl_top[363], bl_top[364], bl_top[365], bl_top[366], bl_top[367],
     bl_top[368], bl_top[369], bl_top[370], bl_top[371], bl_top[372],
     bl_top[373], bl_top[374], bl_top[375], bl_top[376], bl_top[377],
     bl_top[378], bl_top[379], bl_top[380], bl_top[381], bl_top[382],
     bl_top[383], bl_top[384], bl_top[385], bl_top[386], bl_top[387],
     bl_top[388], bl_top[389], bl_top[390], bl_top[391], bl_top[392],
     bl_top[393], bl_top[394], bl_top[395], bl_top[396], bl_top[397],
     bl_top[398], bl_top[399], bl_top[400], bl_top[401], bl_top[402],
     bl_top[403], bl_top[404], bl_top[405], bl_top[406], bl_top[407],
     bl_top[408], bl_top[409], bl_top[410], bl_top[411], bl_top[412],
     bl_top[413], bl_top[414], bl_top[415], bl_top[416], bl_top[417],
     bl_top[418], bl_top[419], bl_top[420], bl_top[421], bl_top[422],
     bl_top[423], bl_top[424], bl_top[425], bl_top[426], bl_top[427],
     bl_top[428], bl_top[429], bl_top[430], bl_top[431], bl_top[432],
     bl_top[433], bl_top[434], bl_top[435], bl_top[436], bl_top[437],
     bl_top[438], bl_top[439], bl_top[440], bl_top[441], bl_top[442],
     bl_top[443], bl_top[444], bl_top[445], bl_top[446], bl_top[447],
     bl_top[448], bl_top[449], bl_top[450], bl_top[451], bl_top[452],
     bl_top[453], bl_top[454], bl_top[455], bl_top[456], bl_top[457],
     bl_top[458], bl_top[459], bl_top[460], bl_top[461], bl_top[462],
     bl_top[463], bl_top[464], bl_top[465], bl_top[466], bl_top[467],
     bl_top[468], bl_top[469], bl_top[470], bl_top[471], bl_top[472],
     bl_top[473], bl_top[474], bl_top[475], bl_top[476], bl_top[477],
     bl_top[478], bl_top[479], bl_top[480], bl_top[481], bl_top[482],
     bl_top[483], bl_top[484], bl_top[485], bl_top[486], bl_top[487],
     bl_top[488], bl_top[489], bl_top[490], bl_top[491], bl_top[492],
     bl_top[493], bl_top[494], bl_top[495], bl_top[496], bl_top[497],
     bl_top[498], bl_top[499], bl_top[500], bl_top[501], bl_top[502],
     bl_top[503], bl_top[504], bl_top[505], bl_top[506], bl_top[507],
     bl_top[508], bl_top[509], bl_top[510], bl_top[511], bl_top[512],
     bl_top[513], bl_top[514], bl_top[515], bl_top[516], bl_top[517],
     bl_top[518], bl_top[519], bl_top[520], bl_top[521], bl_top[522],
     bl_top[523], bl_top[524], bl_top[525], bl_top[526], bl_top[527],
     bl_top[528], bl_top[529], bl_top[530], bl_top[531], bl_top[532],
     bl_top[533], bl_top[534], bl_top[535], bl_top[536], bl_top[537],
     bl_top[538], bl_top[539], bl_top[540], bl_top[541], bl_top[542],
     bl_top[543], bl_top[544], bl_top[545], bl_top[546], bl_top[547],
     bl_top[548], bl_top[549], bl_top[550], bl_top[551], bl_top[552],
     bl_top[553], bl_top[554], bl_top[555], bl_top[556], bl_top[557],
     bl_top[558], bl_top[559], bl_top[560], bl_top[561], bl_top[562],
     bl_top[563], bl_top[564], bl_top[565], bl_top[566], bl_top[567],
     bl_top[568], bl_top[569], bl_top[570], bl_top[571], bl_top[572],
     bl_top[573], bl_top[574], bl_top[575], bl_top[576], bl_top[577],
     bl_top[578], bl_top[579], bl_top[580], bl_top[581], bl_top[582],
     bl_top[583], bl_top[584], bl_top[585], bl_top[586], bl_top[587],
     bl_top[588], bl_top[589], bl_top[590], bl_top[591], bl_top[592],
     bl_top[593], bl_top[594], bl_top[595], bl_top[596], bl_top[597],
     bl_top[598], bl_top[599], bl_top[600], bl_top[601], bl_top[602],
     bl_top[603], bl_top[604], bl_top[605], bl_top[606], bl_top[607],
     bl_top[608], bl_top[609], bl_top[610], bl_top[611], bl_top[612],
     bl_top[613], bl_top[614], bl_top[615], bl_top[616], bl_top[617],
     bl_top[618], bl_top[619], bl_top[620], bl_top[621], bl_top[622],
     bl_top[623], bl_top[624], bl_top[625], bl_top[626], bl_top[627],
     bl_top[628], bl_top[629], bl_top[630], bl_top[631], bl_top[632],
     bl_top[633], bl_top[634], bl_top[635], bl_top[636], bl_top[637],
     bl_top[638], bl_top[639], bl_top[640], bl_top[641], bl_top[642],
     bl_top[643], bl_top[644], bl_top[645], bl_top[646], bl_top[647],
     bl_top[648], bl_top[649], bl_top[650], bl_top[651], bl_top[652],
     bl_top[653], bl_top[654], bl_top[655]}));

endmodule
// Library - io, Cell - PRCUTSSTLSTDR, View - schematic
// LAST TIME SAVED: Oct 24 13:01:45 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module PRCUTSSTLSTDR ( VSS, VSSPST );
input  VSS, VSSPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PRCUTSSTLSTDL, View - schematic
// LAST TIME SAVED: Oct 24 13:01:45 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module PRCUTSSTLSTDL ( VSS, VSSPST );
input  VSS, VSSPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - tielo4x, View - schematic
// LAST TIME SAVED: Sep 10 09:05:31 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module tielo4x ( tielo );
output  tielo;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M0 ( .D(net4), .B(vdd_), .G(net4), .S(vdd_));
nch_hvt  M1 ( .D(tielo), .B(gnd_), .G(net4), .S(gnd_));

endmodule
// Library - leafcell, Cell - tiehi4x, View - schematic
// LAST TIME SAVED: Sep 10 09:03:54 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module tiehi4x ( tiehi );
output  tiehi;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - leafcell, Cell - bram_bufferx4x6, View - schematic
// LAST TIME SAVED: Sep 15 13:53:57 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module bram_bufferx4x6 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I4 ( .in(d1), .out(d2));
bram_bufferx4 I5 ( .in(d2), .out(d3));
bram_bufferx4 I6 ( .in(d3), .out(d4));
bram_bufferx4 I7 ( .in(d4), .out(out));
bram_bufferx4 I3 ( .in(d0), .out(d1));
bram_bufferx4 I0 ( .in(in), .out(d0));

endmodule
// Library - leafcell, Cell - lowla_modified, View - schematic
// LAST TIME SAVED: Sep 15 13:19:27 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module lowla_modified ( lao, clk, min );
output  lao;

input  clk, min;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I289 ( .A(net29), .Y(lao));
inv_hvt I290 ( .A(st2), .Y(net29));
inv_hvt I_inv ( .A(clk), .Y(cbitb));
inv_hvt I_inv3 ( .A(cbitb), .Y(clkd));
txgate_hvt I249 ( .in(lao), .out(st2), .pp(cbitb), .nn(clkd));
txgate_hvt I248 ( .in(min), .out(st2), .pp(clkd), .nn(cbitb));

endmodule
// Library - xpmem, Cell - cram2x2, View - schematic
// LAST TIME SAVED: Jul 28 08:23:43 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module cram2x2 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [3:0]  q;
output [3:0]  q_b;

inout [1:0]  bl;

input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  r_vdd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



eh_cram_cell_4 Icram_cellb831r255 ( .q_b(q_b[1]), .q(q[1]), .wl(wl[0]),
     .bl(bl[1]), .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I20 ( .q_b(q_b[2]), .q(q[2]), .wl(wl[1]), .bl(bl[0]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));
eh_cram_cell_4 I15 ( .q_b(q_b[0]), .q(q[0]), .wl(wl[0]), .bl(bl[0]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I19 ( .q_b(q_b[3]), .q(q[3]), .wl(wl[1]), .bl(bl[1]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));

endmodule
// Library - xpmem, Cell - ml_rowdrv_bank, View - schematic
// LAST TIME SAVED: Aug 28 14:16:35 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_rowdrv_bank ( jtag_rowtest_mode_b, last_rsr, pgate, reset,
     vddctrl, wl, banksel, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst,
     smc_rsr_inc, smc_write, trst_b );
output  jtag_rowtest_mode_b, last_rsr;

input  banksel, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst, smc_rsr_inc,
     smc_write, trst_b;

output [175:0]  reset;
output [175:0]  vddctrl;
output [175:0]  pgate;
output [175:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  smc_rsr_1st_out_buf;

wire  [10:0]  smc_rsr_out;

wire  [9:0]  por_rst_out;

wire  [9:0]  smc_rsr_inc_out;

wire  [0:10]  smc_rsr_1st_out;



tielo I251 ( .tielo(net0130));
tiehi I269 ( .tiehi(net0157));
tiehi I249 ( .tiehi(net0126));
tiehi I250 ( .tiehi(net0125));
ml_buf_ice5_2 I227 ( .in(net0126), .o(net185), .sel(net0126));
ml_buf_ice5_2 I216 ( .in(net0126), .o(net188), .sel(net0126));
ml_buf_ice5_2 I198 ( .sel(banksel), .in(cram_wl_en),
     .o(cram_wl_en_buf));
ml_buf_ice5_2 I196 ( .sel(banksel), .in(cram_rst), .o(cram_rst_buf));
ml_buf_ice5_2 I199 ( .sel(net0125), .in(por_rst), .o(por_rst_buf));
ml_buf_ice5_2 I197 ( .sel(banksel), .in(cram_vddoff),
     .o(cram_vddoff_buf));
ml_buf_ice5_2 I195 ( .sel(banksel), .in(cram_pgateoff),
     .o(cram_pgateoff_buf));
ml_buf_ice5_2 I201 ( .sel(banksel), .in(smc_write), .o(smc_write_buf));
ml_buf_ice5_2 I203 ( .sel(net139), .in(net139), .o(smc_rsr_inc_buf));
ml_buf_ice5_2 I213 ( .in(net0157), .o(net215), .sel(net0157));
ml_rowdrv_tile_last Iml_rowdrv_tile_last (
     .smc_rsr_inc_out(smc_rsr_inc_out_last), .pgate(pgate[175:160]),
     .wl(wl[175:160]), .vddctrl(vddctrl[175:160]),
     .reset(reset[175:160]), .smc_rsr_1st_out(smc_rsr_1st_out[10]),
     .smcc_rsr_out(smc_rsr_out[10]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_buf), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[9]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf));
nand2_hvt I233 ( .A(smc_rsr_inc), .B(banksel), .Y(net136));
mux2_hvt I161 ( .in1(jtag_clk), .in0(net250), .out(net139),
     .sel(net0246));
nand3_hvt I231 ( .Y(net141), .B(net145), .C(net145), .A(net145));
nand3_hvt I230 ( .Y(net145), .B(net150), .C(net150), .A(net150));
nand3_hvt I224 ( .B(net0126), .Y(net150), .A(net0126), .C(net0126));
nor3_hvt I238 ( .B(por_rst), .Y(net233), .A(net162), .C(trst));
nor3_hvt I232 ( .C(rsr_rst), .A(jtag_rowtest_rst), .B(net0130),
     .Y(net167));
nor3_hvt I218 ( .B(net179), .Y(net169), .A(net179), .C(net179));
nor3_hvt I220 ( .B(net169), .Y(net173), .A(net169), .C(net169));
nor3_hvt I217 ( .C(net0126), .A(net0126), .B(net0126), .Y(net179));
nor3_hvt I244 ( .B(por_rst), .Y(net181), .A(net259),
     .C(smc_rsr_1st_out_buf[0]));
ml_rowdrv_tile Iml_rowdrv_tile_9_ ( .por_rst_out(por_rst_out[9]),
     .smc_rsr_inc_out(smc_rsr_inc_out[9]),
     .smcc_rsr_out(smc_rsr_out[9]),
     .smc_rsr_1st_out(smc_rsr_1st_out[9]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out_last), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[8]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[159:144]), .vddctrl(vddctrl[159:144]),
     .reset(reset[159:144]), .pgate(pgate[159:144]));
ml_rowdrv_tile Iml_rowdrv_tile_8_ ( .por_rst_out(por_rst_out[8]),
     .smc_rsr_inc_out(smc_rsr_inc_out[8]),
     .smcc_rsr_out(smc_rsr_out[8]),
     .smc_rsr_1st_out(smc_rsr_1st_out[8]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[9]), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[7]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[143:128]), .vddctrl(vddctrl[143:128]),
     .reset(reset[143:128]), .pgate(pgate[143:128]));
ml_rowdrv_tile Iml_rowdrv_tile_7_ ( .por_rst_out(por_rst_out[7]),
     .smc_rsr_inc_out(smc_rsr_inc_out[7]),
     .smcc_rsr_out(smc_rsr_out[7]),
     .smc_rsr_1st_out(smc_rsr_1st_out[7]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[8]), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[6]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[127:112]), .vddctrl(vddctrl[127:112]),
     .reset(reset[127:112]), .pgate(pgate[127:112]));
ml_rowdrv_tile Iml_rowdrv_tile_6_ ( .por_rst_out(por_rst_out[6]),
     .smc_rsr_inc_out(smc_rsr_inc_out[6]),
     .smcc_rsr_out(smc_rsr_out[6]),
     .smc_rsr_1st_out(smc_rsr_1st_out[6]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[7]), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[5]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[111:96]), .vddctrl(vddctrl[111:96]), .reset(reset[111:96]),
     .pgate(pgate[111:96]));
ml_rowdrv_tile Iml_rowdrv_tile_5_ ( .por_rst_out(por_rst_out[5]),
     .smc_rsr_inc_out(smc_rsr_inc_out[5]),
     .smcc_rsr_out(smc_rsr_out[5]),
     .smc_rsr_1st_out(smc_rsr_1st_out[5]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[6]), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[4]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[95:80]), .vddctrl(vddctrl[95:80]), .reset(reset[95:80]),
     .pgate(pgate[95:80]));
ml_rowdrv_tile Iml_rowdrv_tile_4_ ( .por_rst_out(por_rst_out[4]),
     .smc_rsr_inc_out(smc_rsr_inc_out[4]),
     .smcc_rsr_out(smc_rsr_out[4]),
     .smc_rsr_1st_out(smc_rsr_1st_out[4]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[5]), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[3]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[79:64]), .vddctrl(vddctrl[79:64]), .reset(reset[79:64]),
     .pgate(pgate[79:64]));
ml_rowdrv_tile Iml_rowdrv_tile_3_ ( .por_rst_out(por_rst_out[3]),
     .smc_rsr_inc_out(smc_rsr_inc_out[3]),
     .smcc_rsr_out(smc_rsr_out[3]),
     .smc_rsr_1st_out(smc_rsr_1st_out[3]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[4]), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[2]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[63:48]), .vddctrl(vddctrl[63:48]), .reset(reset[63:48]),
     .pgate(pgate[63:48]));
ml_rowdrv_tile Iml_rowdrv_tile_2_ ( .por_rst_out(por_rst_out[2]),
     .smc_rsr_inc_out(smc_rsr_inc_out[2]),
     .smcc_rsr_out(smc_rsr_out[2]),
     .smc_rsr_1st_out(smc_rsr_1st_out[2]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[3]), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[1]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[47:32]), .vddctrl(vddctrl[47:32]), .reset(reset[47:32]),
     .pgate(pgate[47:32]));
ml_rowdrv_tile Iml_rowdrv_tile_1_ ( .por_rst_out(por_rst_out[1]),
     .smc_rsr_inc_out(smc_rsr_inc_out[1]),
     .smcc_rsr_out(smc_rsr_out[1]),
     .smc_rsr_1st_out(smc_rsr_1st_out[1]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[2]), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[0]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[31:16]), .vddctrl(vddctrl[31:16]), .reset(reset[31:16]),
     .pgate(pgate[31:16]));
ml_rowdrv_tile Iml_rowdrv_tile_0_ ( .por_rst_out(por_rst_out[0]),
     .smc_rsr_inc_out(smc_rsr_inc_out[0]),
     .smcc_rsr_out(smc_rsr_out[0]),
     .smc_rsr_1st_out(smc_rsr_1st_out[0]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[1]), .smc_rsr_in(smc_rsr_in_1st),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[15:0]), .vddctrl(vddctrl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]));
nor2_hvt I239 ( .A(jtag_rowtest_rst), .B(net233), .Y(net162));
nor2_hvt I193 ( .A(por_rst), .B(rsr_set_1st), .Y(net237));
nor2_hvt I245 ( .A(rsr_set_1st), .B(net181), .Y(net259));
inv_hvt I247 ( .A(net0246), .Y(jtag_rowtest_mode_b));
inv_hvt I241 ( .A(net162), .Y(net0246));
inv_hvt I192 ( .A(net167), .Y(rsr_set_1st));
inv_hvt I234 ( .A(net136), .Y(net250));
inv_hvt I35 ( .A(net241), .Y(smc_rsr_1st_out_buf[0]));
inv_hvt I240 ( .A(trst_b), .Y(trst));
inv_hvt I210 ( .A(net253), .Y(last_rsr));
inv_hvt I391 ( .A(net237), .Y(rst_row_reg));
inv_hvt I36 ( .A(smc_rsr_1st_out[0]), .Y(net241));
inv_hvt I209 ( .A(smc_rsr_out[10]), .Y(net253));
inv_hvt I205 ( .A(net259), .Y(smc_rsr_in_1st));

endmodule
// Library - io, Cell - io_odrv4x5, View - schematic
// LAST TIME SAVED: Aug 21 17:59:07 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module io_odrv4x5 ( cbit, sp4_out, bl, pgate, prog,
     reset, slfop, vdd_cntl, wl );


input  prog, slfop;

output [4:0]  sp4_out;
output [7:5]  cbit;

inout [3:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
supply0 gnd_;
supply1 vdd_;

// Buses in the design

wire  [7:0]  cbitb;

wire  [1:0]  r_vdd;

wire [7:0] cbit_int;
assign cbit[7:5] = cbit_int[7:5];


pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv4 I_odrv_4_ ( .cbitb(cbitb[4]), .sp4(sp4_out[4]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_3_ ( .cbitb(cbitb[3]), .sp4(sp4_out[3]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_2_ ( .cbitb(cbitb[2]), .sp4(sp4_out[2]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_1_ ( .cbitb(cbitb[1]), .sp4(sp4_out[1]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_0_ ( .cbitb(cbitb[0]), .sp4(sp4_out[0]), .slfop(slfop),
     .prog(prog));
cram2x2 Icram2x2_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset[1:0]), .q(cbit_int[7:4]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));
cram2x2 Icram2x2_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset[1:0]), .q(cbit_int[3:0]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - io_col_odrv4_x40bare, View - schematic
// LAST TIME SAVED: Jul 31 17:45:40 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module io_col_odrv4_x40bare ( cf, bl, sp4_h_l,
     sp4_v_b, dout0, dout1,
     pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [23:0]  cf;

inout [3:0]  bl;
inout [15:0]  sp4_v_b;
inout [47:0]  sp4_h_l;

input [0:1]  dout0;
input [0:1]  dout1;
input [15:0]  pgate;
input [15:0]  wl;
input [15:0]  reset;
input [15:0]  vdd_cntl;
supply0 gnd_;
supply1 vdd_;



io_odrv4x5 I218 ( cf[20:18], {sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6]}, bl[3:0], pgate[13:12], prog,
     reset[13:12], dout1[1], vdd_cntl[13:12], wl[13:12]);
io_odrv4x5 I217 ( cf[14:12], {sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4]}, bl[3:0], pgate[9:8], prog, reset[9:8],
     dout0[1], vdd_cntl[9:8], wl[9:8]);
io_odrv4x5 I_odrv_4x5_7 ( cf[23:21], {sp4_v_b[15], sp4_v_b[11],
     sp4_v_b[7], sp4_v_b[3], sp4_h_l[46]}, bl[3:0], pgate[15:14], prog,
     reset[15:14], dout1[1], vdd_cntl[15:14], wl[15:14]);
io_odrv4x5 I220 ( cf[11:9], {sp4_v_b[13], sp4_v_b[9], sp4_v_b[5],
     sp4_v_b[1], sp4_h_l[42]}, bl[3:0], pgate[7:6], prog, reset[7:6],
     dout1[0], vdd_cntl[7:6], wl[7:6]);
io_odrv4x5 I221 ( cf[8:6], {sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2]}, bl[3:0], pgate[5:4], prog, reset[5:4],
     dout1[0], vdd_cntl[5:4], wl[5:4]);
io_odrv4x5 I_odrv_4x5_0 ( cf[2:0], {sp4_h_l[32], sp4_h_l[24],
     sp4_h_l[16], sp4_h_l[8], sp4_h_l[0]}, bl[3:0], pgate[1:0], prog,
     reset[1:0], dout0[0], vdd_cntl[1:0], wl[1:0]);
io_odrv4x5 I223 ( cf[5:3], {sp4_v_b[12], sp4_v_b[8], sp4_v_b[4],
     sp4_v_b[0], sp4_h_l[40]}, bl[3:0], pgate[3:2], prog, reset[3:2],
     dout0[0], vdd_cntl[3:2], wl[3:2]);
io_odrv4x5 I215 ( cf[17:15], {sp4_v_b[14], sp4_v_b[10], sp4_v_b[6],
     sp4_v_b[2], sp4_h_l[44]}, bl[3:0], pgate[11:10], prog,
     reset[11:10], dout0[1], vdd_cntl[11:10], wl[11:10]);

endmodule
// Library - io, Cell - io_gmux_x2, View - schematic
// LAST TIME SAVED: Aug 21 18:00:57 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module io_gmux_x2 ( gout, bl, min0, min1, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [1:0]  gout;

inout [5:0]  bl;

input [15:0]  min1;
input [15:0]  min0;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux Ig_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux Ig_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare, View - schematic
// LAST TIME SAVED: Jul 31 17:47:21 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module io_gmux_x16bare ( lc_trk_g0, lc_trk_g1, bl, min0, min1, min2,
     min3, min4, min5, min6, min7, min8, min9, min10, min11, min12,
     min13, min14, min15, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;

inout [5:0]  bl;

input [15:0]  min3;
input [15:0]  min9;
input [15:0]  min7;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min12;
input [15:0]  min14;
input [15:0]  min6;
input [15:0]  min5;
input [15:0]  min2;
input [15:0]  min10;
input [15:0]  min15;
input [15:0]  vdd_cntl;
input [15:0]  reset;
input [15:0]  wl;
input [15:0]  min11;
input [15:0]  min0;
input [15:0]  min8;
input [15:0]  min4;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



io_gmux_x2 Iio_gmux4 ( .vdd_cntl(vdd_cntl[9:8]), .bl(bl[5:0]),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux5 ( .vdd_cntl(vdd_cntl[11:10]), .bl(bl[5:0]),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux6 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux2 ( .vdd_cntl(vdd_cntl[5:4]), .bl(bl[5:0]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux3 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux7 ( .vdd_cntl(vdd_cntl[15:14]), .bl(bl[5:0]),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog));

endmodule
// Library - io, Cell - ioin_mux, View - schematic
// LAST TIME SAVED: May 18 11:01:33 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioin_mux ( inmuxo, cbit[3], cbit[2], cbit[1], cbit[0], cbitb[3],
     cbitb[2], cbitb[1], cbitb[0], min[7:0], prog );
output  inmuxo;

input  prog;

input [0:3]  cbitb;
input [7:0]  min;
input [0:3]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I278 ( .A(net146), .Y(inmuxo));
nor2_hvt I46 ( .A(prog), .B(cbitb[3]), .Y(en));
nand2_hvt Inand2_muxo ( .A(st2), .Y(net146), .B(en));
txgate_hvt I247 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I257 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I254 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I244 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I253 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_hvt I249 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_hvt I274 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_hvt I252 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));
txgate_hvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_hvt I255 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I250 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_hvt I258 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I256 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I246 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc, View - schematic
// LAST TIME SAVED: Aug 21 18:04:33 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  ti;
output [1:0]  spi;

inout [5:0]  bl;

input [7:0]  min2;
input [1:0]  vdd_cntl;
input [7:0]  min1;
input [1:0]  reset;
input [1:0]  padin;
input [7:0]  min0;
input [1:0]  pgate;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
nor2_hvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_hvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
inv_hvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_hvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
ioin_mux I193 ( bankcntl, {cbit[11], cbit[8], cbit[9], cbit[10]},
     {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0], prog);
ioin_mux I185 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux I186 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]}, {cbitb[5],
     cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);

endmodule
// Library - io, Cell - ioinmx1mux2, View - schematic
// LAST TIME SAVED: Aug 21 18:09:41 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioinmx1mux2 ( clk, mo, ti, bl, cdone_in, ce, ceb, in, min,
     pgate, prog, reset, spi, vdd_cntl, wl );
output  clk, ti;


input  cdone_in, ceb, prog;

output [1:0]  mo;

inout [5:0]  bl;

input [7:0]  min;
input [1:0]  spi;
input [1:0]  wl;
input [1:0]  in;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [11:0]  ce;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clk_mux12to1 I298 ( .prog(prog), .min(ce[11:0]), .clk(clk),
     .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7], cbitb[10],
     cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7], cbit[10],
     cbit[6], cbit[4]}), .cenb(ceb));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
mux2x1_hvt Iemux_1_ ( .in1(in[1]), .in0(spi[1]), .out(mo[1]),
     .sel(cdone_in));
mux2x1_hvt Iemux_0_ ( .in1(in[0]), .in0(spi[0]), .out(mo[0]),
     .sel(cdone_in));
ioin_mux I185 ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);

endmodule
// Library - io, Cell - ioinmx2nand2inv, View - schematic
// LAST TIME SAVED: Sep 26 11:29:24 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioinmx2nand2inv ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  ce;
input [7:0]  min0;
input [1:0]  reset;
input [7:0]  min1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
inv_hvt I181 ( .A(update), .Y(bs_enb));
nand2_hvt I180 ( .A(bs_enb), .Y(updt), .B(bs_en));
ioin_mux I185 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux I186 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]}, {cbitb[5],
     cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);

endmodule
// Library - io, Cell - sbox1mem, View - schematic
// LAST TIME SAVED: Aug 21 18:03:06 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module sbox1mem ( b, bl, l, r, t, pgate, prog, reset, vdd_cntl, wl );
inout  b, l, r, t;

input  prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbitb;

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox1m3to1 I232 ( .in2(r), .cb({cbitb[3], cbitb[6]}), .op(t), .in0(l),
     .in1(b), .c({cbit[3], cbit[6]}), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb({cbitb[1], cbitb[4]}), .op(l), .in0(b),
     .in1(t), .c({cbit[1], cbit[4]}), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb({cbitb[8], cbitb[5]}), .op(b), .in0(l),
     .in1(t), .c({cbit[8], cbit[5]}), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb({cbitb[10], cbitb[7]}), .op(r), .in0(l),
     .in1(t), .c({cbit[10], cbit[7]}), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc, View - schematic
// LAST TIME SAVED: Aug 21 18:09:59 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module sbox1_colbdlc ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  pado;
output [1:0]  padeb;
output [5:0]  ti;
output [1:0]  spi_ss_in_b;

inout [5:0]  bl;
inout [3:0]  r;
inout [3:0]  sp4_v_b;
inout [3:0]  t_mid;
inout [3:0]  l;

input [7:0]  min1;
input [1:0]  spioeb;
input [11:0]  clk_in;
input [7:0]  ceb_in;
input [1:0]  oeb;
input [7:0]  min2;
input [7:0]  min4;
input [7:0]  min0;
input [1:0]  padin;
input [7:0]  min5;
input [7:0]  min3;
input [1:0]  spiout;
input [1:0]  out;
input [7:0]  min6;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [11:0]  inclk_in;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ioinmx2nor2invx2bdlc I5 ( .vdd_cntl(vdd_cntl[5:4]), .min2(min6[7:0]),
     .bankcntl(fabric_out), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx1mux2 I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .in(out[1:0]), .ti(ti[2]), .min(min2[7:0]), .spi(spiout[1:0]),
     .wl(wl[9:8]), .reset(reset[9:8]), .pgate(pgate[9:8]),
     .cdone_in(cdone_in), .mo(pado[1:0]));
ioinmx1mux2 I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .in(oeb[1:0]), .ti(ti[5]), .min(min5[7:0]), .spi(spioeb[1:0]),
     .wl(wl[15:14]), .reset(reset[15:14]), .pgate(pgate[15:14]),
     .cdone_in(cdone_in), .mo(padeb[1:0]));
ioinmx2nand2inv I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - leafcell, Cell - bram_bufferx4, View - schematic
// LAST TIME SAVED: Jun 25 13:46:30 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module bram_bufferx4 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - io, Cell - odrv12x3, View - schematic
// LAST TIME SAVED: Aug 23 11:52:00 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module odrv12x3 ( sp12, bl, pgate, prog, reset, slfop, vdd_cntl, wl );


input  prog;

output [2:0]  sp12;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  reset;
input [1:0]  vdd_cntl;
input [2:0]  slfop;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12_2_ ( .slfop(slfop[2]), .cbitb(cbitb[2]),
     .sp12(sp12[2]), .prog(prog));
odrv12 I_odrv12_1_ ( .slfop(slfop[1]), .cbitb(cbitb[1]),
     .sp12(sp12[1]), .prog(prog));
odrv12 I_odrv12_0_ ( .slfop(slfop[0]), .cbitb(cbitb[0]),
     .sp12(sp12[0]), .prog(prog));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - cebdffrqn, View - schematic
// LAST TIME SAVED: Jan 31 09:00:47 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module cebdffrqn ( q, qn, ceb, clk, d, r );
output  q, qn;

input  ceb, clk, d, r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I54 ( .A(net62), .B(clk), .Y(clatb), .C(ceb));
nand2_hvt I290 ( .A(clk), .Y(clkb), .B(clatb));
nand2_hvt I42 ( .A(si), .B(rstb), .Y(so));
nor2_hvt INAND2_m ( .A(r), .Y(q), .B(mi));
inv_hvt I39 ( .A(q), .Y(qn));
inv_hvt Iinv_ckfb ( .A(clatb), .Y(net62));
inv_hvt I50 ( .A(clkb), .Y(clkd));
inv_hvt I43 ( .A(so), .Y(low_s));
inv_hvt I40 ( .A(r), .Y(rstb));
txgate_hvt I44 ( .in(d), .out(si), .pp(clkd), .nn(clkb));
txgate_hvt I52 ( .in(so), .out(mi), .pp(clkb), .nn(clkd));
txgate_hvt I51 ( .in(si), .out(low_s), .pp(clkb), .nn(clkd));
txgate_hvt I53 ( .in(mi), .out(qn), .pp(clkd), .nn(clkb));

endmodule
// Library - io, Cell - outsel1_hvt, View - schematic
// LAST TIME SAVED: Jul  3 13:08:26 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module outsel1_hvt ( out, clk, in0, in1, in2, sb, sel );
output  out;

input  clk, in0, in1, in2;

input [1:0]  sel;
input [1:0]  sb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I41 ( .A(in1), .Y(net036));
inv_hvt I40 ( .A(clk), .Y(clkb));
txgate_hvt I33 ( .in(whatever), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_hvt I_txgate1 ( .in(net036), .out(whatever), .pp(sb[0]),
     .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(whatever), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(ddr), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_hvt I38 ( .in(in2), .out(ddr), .pp(clkb), .nn(clk));
txgate_hvt I39 ( .in(in1), .out(ddr), .pp(clk), .nn(clkb));

endmodule
// Library - io, Cell - dffrckb, View - schematic
// LAST TIME SAVED: May 11 14:58:52 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module dffrckb ( q, qn, clk, d, e, r );
output  q, qn;

input  clk, d, e, r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



oai21x2_hvt I57 ( .A1(clk), .Y(clat), .A0(clatb), .B0(e));
nor2_hvt I48 ( .B(clat), .A(clk), .Y(clkb));
nand2_hvt I54 ( .A(rstb), .Y(qn), .B(q));
nand2_hvt I42 ( .A(si), .B(rstb), .Y(so));
inv_hvt I55 ( .A(mi), .Y(q));
inv_hvt I50 ( .A(clkb), .Y(clkd));
inv_hvt I56 ( .A(clat), .Y(clatb));
inv_hvt I43 ( .A(so), .Y(low_s));
inv_hvt I40 ( .A(r), .Y(rstb));
txgate_hvt I59 ( .in(d), .out(si), .pp(clkb), .nn(clkd));
txgate_hvt I64 ( .in(low_s), .out(si), .pp(clkd), .nn(clkb));
txgate_hvt I62 ( .in(qn), .out(mi), .pp(clkb), .nn(clkd));
txgate_hvt I60 ( .in(so), .out(mi), .pp(clkd), .nn(clkb));

endmodule
// Library - io, Cell - out_logic_v1, View - schematic
// LAST TIME SAVED: Feb  8 11:44:57 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module out_logic_v1 ( dout, sdo, bs_en, cbit, cbitb, ceb, clk, ddr0,
     ddr1, mode, rstio, sdi, shift, tclk, ud );
output  dout, sdo;

input  bs_en, ceb, clk, ddr0, ddr1, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cebdffrqn Ireg0 ( .ceb(ceb), .clk(mux4clk), .qn(net094), .r(rstio),
     .q(sdo), .d(dd));
outsel1_hvt I169 ( .clk(ddrclk), .in2(udb), .sb(cbitb[1:0]),
     .sel(cbit[1:0]), .in1(net094), .in0(dinb), .out(muxob));
nor2_hvt I179 ( .A(mux4clk), .B(cbit[0]), .Y(ddrclk));
dffrckb Ireg1 ( .e(ud), .clk(mux4clk), .qn(udb), .r(rstio), .q(net44),
     .d(mux4d));
inv_hvt I171 ( .A(doutb), .Y(dout));
inv_hvt I172 ( .A(ddr0), .Y(dinb));
mux2x1_hvt I170 ( .sel(mode), .in1(udb), .in0(muxob), .out(doutb));
mux2x1_hvt I177 ( .in1(tclk), .in0(clk), .out(mux4clk), .sel(bs_en));
mux2x1_hvt I173 ( .in1(sdi), .in0(ddr0), .out(dd), .sel(shift));
mux2x1_hvt I176 ( .in1(sdo), .in0(ddr1), .out(mux4d), .sel(bs_en));

endmodule
// Library - io, Cell - out_logic_v3, View - schematic
// LAST TIME SAVED: Feb  8 11:47:27 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module out_logic_v3 ( dout, sdo, sp12, bl, bs_en, ceb, clk, ddr0, ddr1,
     mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk, ud,
     vdd_cntl, wl );
output  dout, sdo, sp12;


input  bs_en, ceb, clk, ddr0, ddr1, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;

wire  [3:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I181 ( .slfop(slfop), .cbitb(cbitb[1]), .sp12(sp12),
     .prog(prog));
cram2x2 I183 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
out_logic_v1 I_outlogic_v1 ( .ceb(ceb), .rstio(rstio), .ddr0(ddr0),
     .ddr1(ddr1), .shift(shift), .ud(ud), .clk(clk), .sdo(sdo),
     .sdi(sdi), .cbit({cbit[2], cbit[3]}), .cbitb({cbitb[2],
     cbitb[3]}), .dout(dout), .tclk(tclk), .bs_en(bs_en), .mode(mode));

endmodule
// Library - io, Cell - insel1_hvt, View - schematic
// LAST TIME SAVED: Jul  2 18:38:19 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module insel1_hvt ( out, in0, in1, in2, in3, sb, sel );
output  out;

input  in0, in1, in2, in3;

input [1:0]  sb;
input [1:0]  sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I39 ( .in(in3), .out(net025), .pp(sb[0]), .nn(sel[0]));
txgate_hvt I40 ( .in(in2), .out(net025), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I33 ( .in(net038), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_hvt I_txgate1 ( .in(in1), .out(net038), .pp(sb[0]),
     .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(net038), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(net025), .out(out), .pp(sb[1]), .nn(sel[1]));

endmodule
// Library - io, Cell - in_logic_v1, View - schematic
// LAST TIME SAVED: Feb  8 11:39:50 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module in_logic_v1 ( dout0, dout1, sdo, bs_en, cbit, cbitb, ceb, clk,
     cntl, din, mode, rstio, sdi, shift, tclk, ud );
output  dout0, dout1, sdo;

input  bs_en, ceb, clk, cntl, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbitb;
input [1:0]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cebdffrqn I167 ( .ceb(ceb), .clk(ck2r0), .qn(regb), .r(rstio), .q(sdo),
     .d(dd));
nand2_hvt I184 ( .A(cntl), .Y(cbit1b), .B(cbit[1]));
insel1_hvt I181 ( .in1(dinb), .in0(regb), .out(reg_), .sb({cbit1b,
     cbitb[0]}), .sel({cbit1, cbit[0]}), .in2(net037), .in3(net037));
dffrckb I168 ( .e(ud), .clk(ck2r0), .qn(udd), .r(rstio), .q(net060),
     .d(net056));
inv_hvt I171 ( .A(doutb), .Y(dout0));
inv_hvt I182 ( .A(udd), .Y(dout1));
inv_hvt I185 ( .A(cbit1b), .Y(cbit1));
inv_hvt I186 ( .A(dout0), .Y(net037));
inv_hvt I172 ( .A(din), .Y(dinb));
mux2x1_hvt I170 ( .sel(mode), .in1(udd), .in0(reg_), .out(doutb));
mux2x1_hvt I178 ( .in1(tclk), .in0(clk), .out(ck2r0), .sel(bs_en));
mux2x1_hvt I173 ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
mux2x1_hvt I179 ( .in1(sdo), .in0(din), .out(net056), .sel(bs_en));

endmodule
// Library - io, Cell - in_logic_v3, View - schematic
// LAST TIME SAVED: Feb  8 11:42:24 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module in_logic_v3 ( dout0, dout1, sdo, sp12, bl, bs_en, ceb, clk,
     cntl, din, mode, pgate, prog, reset, rstio, sdi, shift, slfop,
     tclk, ud, vdd_cntl, wl );
output  dout0, dout1, sdo, sp12;


input  bs_en, ceb, clk, cntl, din, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;

wire  [3:0]  cbit;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[3]), .sp12(sp12),
     .prog(prog));
in_logic_v1 I_in_logic ( .ceb(ceb), .rstio(rstio), .din(din),
     .cntl(cntl), .dout1(dout1), .dout0(dout0), .shift(shift), .ud(ud),
     .clk(clk), .sdo(sdo), .sdi(sdi), .cbit({cbit[0], cbit[1]}),
     .cbitb({cbitb[0], cbitb[1]}), .tclk(tclk), .bs_en(bs_en),
     .mode(mode));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioesel_hvt, View - schematic
// LAST TIME SAVED: Aug 21 18:20:13 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioesel_hvt ( out, in0, in1, sb, sel );
output  out;

input  in0, in1;

input [1:0]  sel;
input [1:0]  sb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I38 ( .A(sel[0]), .Y(net017));
txgate_hvt I33 ( .in(mid), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_hvt I_txgate1 ( .in(in1), .out(mid), .pp(sb[0]), .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(mid), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(net017), .out(out), .pp(sel[1]), .nn(sb[1]));

endmodule
// Library - xpmem, Cell - sg_dffbuf, View - schematic
// LAST TIME SAVED: Aug 28 14:33:30 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module sg_dffbuf ( dffout, clk, d, r );
output  dffout;

input  clk, d, r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I2 ( .in(net10), .out(dffout));
ml_dff I0 ( .R(r), .D(d), .CLK(clk), .QN(net9), .Q(net10));

endmodule
// Library - xpmem, Cell - sg_bufx10, View - schematic
// LAST TIME SAVED: Jul 28 19:09:08 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module sg_bufx10 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - io, Cell - ioe_logic_v1, View - schematic
// LAST TIME SAVED: Feb  8 11:28:22 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioe_logic_v1 ( outb, sdo, bs_en, cbit, cbitb, ceb, clk, din,
     mode, rstio, sdi, shift, tclk, ud );
output  outb, sdo;

input  bs_en, ceb, clk, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cebdffrqn I167 ( .ceb(ceb), .clk(net039), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I168 ( .e(ud), .clk(net039), .qn(udd), .r(rstio), .q(net44),
     .d(sdo));
inv_hvt I172 ( .A(din), .Y(dinb));
mux2x1_hvt I175 ( .in1(tclk), .in0(clk), .out(net039), .sel(bs_en));
mux2x1_hvt I170 ( .sel(mode), .in1(udd), .in0(regmuxb), .out(outb));
mux2x1_hvt I173 ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
ioesel_hvt I_ioe_mux2 ( .sb(cbitb[1:0]), .sel(cbit[1:0]), .in1(regb),
     .in0(dinb), .out(regmuxb));

endmodule
// Library - io, Cell - ioe_logic_v3, View - schematic
// LAST TIME SAVED: Feb  8 11:37:10 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioe_logic_v3 ( padeb, sdo, sp12, bl, bs_en, ceb, clk, din,
     hiz_b, mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk,
     ud, vdd_cntl, wl );
output  padeb, sdo, sp12;


input  bs_en, ceb, clk, din, hiz_b, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  reset;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbit;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[1]), .sp12(sp12),
     .prog(prog));
nand2_hvt I178 ( .A(oed), .Y(padeb), .B(hiz_b));
inv_hvt I179 ( .A(oeb), .Y(oed));
ioe_logic_v1 I_ioe_logic ( .ceb(ceb), .rstio(rstio), .cbit(cbit[3:2]),
     .cbitb(cbitb[3:2]), .outb(oeb), .bs_en(bs_en), .shift(shift),
     .ud(ud), .clk(clk), .sdo(sdo), .sdi(sdi), .din(din), .tclk(tclk),
     .mode(mode));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioe_col2, View - schematic
// LAST TIME SAVED: Feb  8 13:09:06 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ioe_col2 ( dout, padeb, pado, sdo, sp12_h_l, bl, bs_en, ceb,
     hiz_b, hold, inclk, mode, outclk, padin, pgate, prog, reset,
     rstio, sdi, shift, tclk, ti, update, vdd_cntl, wl );
output  sdo;


input  bs_en, ceb, hiz_b, hold, inclk, mode, outclk, prog, rstio, sdi,
     shift, tclk, update;

output [1:0]  pado;
output [1:0]  padeb;
output [23:0]  sp12_h_l;
output [3:0]  dout;

inout [1:0]  bl;

input [5:0]  ti;
input [1:0]  padin;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



odrv12x3 I218 ( .vdd_cntl(vdd_cntl[7:6]), .slfop({dout[1], dout[1],
     dout[1]}), .sp12({sp12_h_l[18], sp12_h_l[10], sp12_h_l[2]}),
     .bl(bl[1:0]), .wl(wl[7:6]), .reset(reset[7:6]),
     .pgate(pgate[7:6]), .prog(prog));
odrv12x3 I217 ( .vdd_cntl(vdd_cntl[9:8]), .slfop({dout[2], dout[2],
     dout[2]}), .sp12({sp12_h_l[20], sp12_h_l[12], sp12_h_l[4]}),
     .bl(bl[1:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]), .prog(prog));
out_logic_v3 I_out0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[1:0]),
     .ddr0(ti[1]), .ddr1(ti[2]), .rstio(rstio), .slfop(dout[0]),
     .sp12(sp12_h_l[0]), .dout(pado[0]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[1:0]),
     .reset(reset[1:0]), .sdo(s0), .sdi(sdi), .pgate(pgate[1:0]),
     .tclk(tclk), .bs_en(bs_en), .mode(mode));
out_logic_v3 I_out1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[11:10]),
     .ddr0(ti[4]), .ddr1(ti[5]), .rstio(rstio), .slfop(dout[3]),
     .sp12(sp12_h_l[6]), .dout(pado[1]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[11:10]),
     .reset(reset[11:10]), .sdo(s3), .sdi(s2), .pgate(pgate[11:10]),
     .tclk(tclk), .bs_en(bs_en), .mode(mode));
in_logic_v3 I_in0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[3:2]), .rstio(rstio),
     .slfop(dout[0]), .sp12(sp12_h_l[8]), .shift(shift),
     .dout1(dout[1]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[0]), .wl(wl[3:2]), .reset(reset[3:2]),
     .sdo(s1), .sdi(s0), .pgate(pgate[3:2]), .din(padin[0]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode));
in_logic_v3 I_in1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[13:12]),
     .rstio(rstio), .slfop(dout[3]), .sp12(sp12_h_l[14]),
     .shift(shift), .dout1(dout[3]), .ud(update), .bl(bl[1:0]),
     .prog(prog), .clk(inclk), .dout0(dout[2]), .wl(wl[13:12]),
     .reset(reset[13:12]), .sdo(s4), .sdi(s3), .pgate(pgate[13:12]),
     .din(padin[1]), .tclk(tclk), .bs_en(bs_en), .cntl(hold),
     .mode(mode));
ioe_logic_v3 I_ioe0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[5:4]),
     .rstio(rstio), .slfop(dout[0]), .sp12(sp12_h_l[16]),
     .hiz_b(hiz_b), .padeb(padeb[0]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[5:4]),
     .reset(reset[5:4]), .sdo(s2), .sdi(s1), .pgate(pgate[5:4]),
     .din(ti[0]), .tclk(tclk), .bs_en(bs_en), .mode(mode));
ioe_logic_v3 I_ioe1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[15:14]),
     .rstio(rstio), .slfop(dout[3]), .sp12(sp12_h_l[22]),
     .hiz_b(hiz_b), .padeb(padeb[1]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[15:14]),
     .reset(reset[15:14]), .sdo(sdo), .sdi(s4), .pgate(pgate[15:14]),
     .din(ti[3]), .tclk(tclk), .bs_en(bs_en), .mode(mode));

endmodule
// Library - io, Cell - io_col4_rowright, View - schematic
// LAST TIME SAVED: Feb  8 13:12:48 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module io_col4_rowright ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [23:0]  cf;
output [1:0]  padeb;
output [3:0]  slf_op;

inout [15:0]  sp4_v_t;
inout [17:0]  bl;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;

input [15:0]  pgate;
input [1:0]  spioeb;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [15:0]  reset;
input [1:0]  spiout;
input [1:0]  padin;
input [7:0]  glb_netwk;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  oenm;

wire  [5:0]  ti;

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



rm7  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[17:14],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, pgate[15:0], prog, reset[15:0], vdd_cntl[15:0],
     wl[15:0]);
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl(vdd_cntl[15:0]),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[13:8]), .wl(wl[15:0]),
     .reset(reset[15:0]), .pgate(pgate[15:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(prog),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl(vdd_cntl[15:0]), .outclk(outclk),
     .fabric_out(fabric_out), .min6({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .inclk_in({lc_trk_g1[3],
     lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0], glb_netwk[7:0]}),
     .ceb_in({lc_trk_g1[5], lc_trk_g1[2], lc_trk_g0[5], lc_trk_g0[2],
     glb_netwk[6], glb_netwk[4], glb_netwk[2], glb_netwk[0]}),
     .clk_in({lc_trk_g1[4], lc_trk_g1[1], lc_trk_g0[4], lc_trk_g0[1],
     glb_netwk[7:0]}), .update(update), .spiout(spiout[1:0]),
     .spioeb(spioeb[1:0]), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[7:2]), .inclk(inclk), .wl(wl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]), .prog(prog));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl(vdd_cntl[15:0]),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl(wl[15:0]), .reset(reset[15:0]), .pgate(pgate[15:0]),
     .hiz_b(hiz_b), .update(enable_update), .ti(ti[5:0]), .tclk(tclk),
     .shift(shift), .sdi(sdi), .prog(prog), .padin(padin[1:0]),
     .mode(mode), .inclk(inclk), .bs_en(bs_en),
     .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo), .pado(om[1:0]),
     .padeb(oenm[1:0]), .bl(bl[1:0]));

endmodule
// Library - io, Cell - io_col4_lb, View - schematic
// LAST TIME SAVED: Feb  8 13:17:55 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module io_col4_lb ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [23:0]  cf;
output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [1:0]  padeb;
output [3:0]  slf_op;

inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;

input [1:0]  spioeb;
input [15:0]  pgate;
input [15:0]  wl;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  tnl_op;
input [15:0]  reset;
input [1:0]  spiout;
input [15:0]  vdd_cntl;
input [1:0]  padin;
input [7:0]  glb_netwk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



rm6  R14_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R14_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R14_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R14_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R14_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R14_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R14_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R14_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R14_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R14_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R14_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R14_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R14_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R14_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R14_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R14_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[17:14],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, pgate[15:0], prog, reset[15:0], vdd_cntl[15:0],
     wl[15:0]);
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl(vdd_cntl[15:0]),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[13:8]), .wl(wl[15:0]),
     .reset(reset[15:0]), .pgate(pgate[15:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(prog),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl(vdd_cntl[15:0]), .outclk(outclk),
     .fabric_out(fabric_out), .min6({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .inclk_in({lc_trk_g1[3],
     lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0], glb_netwk[7:0]}),
     .ceb_in({lc_trk_g1[5], lc_trk_g1[2], lc_trk_g0[5], lc_trk_g0[2],
     glb_netwk[6], glb_netwk[4], glb_netwk[2], glb_netwk[0]}),
     .clk_in({lc_trk_g1[4], lc_trk_g1[1], lc_trk_g0[4], lc_trk_g0[1],
     glb_netwk[7:0]}), .update(update), .spiout(spiout[1:0]),
     .spioeb(spioeb[1:0]), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[7:2]), .inclk(inclk), .wl(wl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]), .prog(prog));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl(vdd_cntl[15:0]),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl(wl[15:0]), .reset(reset[15:0]), .pgate(pgate[15:0]),
     .hiz_b(hiz_b), .update(enable_update), .ti(ti[5:0]), .tclk(tclk),
     .shift(shift), .sdi(sdi), .prog(prog), .padin(padin[1:0]),
     .mode(mode), .inclk(inclk), .bs_en(bs_en),
     .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo), .pado(om[1:0]),
     .padeb(oenm[1:0]), .bl(bl[1:0]));

endmodule
// Library - leafcell, Cell - clk_quad_buf, View - schematic
// LAST TIME SAVED: Jul 10 09:32:37 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module clk_quad_buf ( clko, clki );
output  clko;

input  clki;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv I19 ( .A(clkb), .Y(clko));
inv I22 ( .A(clki), .Y(clkb));

endmodule
// Library - leafcell, Cell - clk_quad_bufx8, View - schematic
// LAST TIME SAVED: Jul 11 09:58:57 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module clk_quad_bufx8 ( clko, clki );


output [7:0]  clko;

input [7:0]  clki;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



clk_quad_buf iclk_colbuf_7_ ( .clki(clki[7]), .clko(clko[7]));
clk_quad_buf iclk_colbuf_6_ ( .clki(clki[6]), .clko(clko[6]));
clk_quad_buf iclk_colbuf_5_ ( .clki(clki[5]), .clko(clko[5]));
clk_quad_buf iclk_colbuf_4_ ( .clki(clki[4]), .clko(clko[4]));
clk_quad_buf iclk_colbuf_3_ ( .clki(clki[3]), .clko(clko[3]));
clk_quad_buf iclk_colbuf_2_ ( .clki(clki[2]), .clko(clko[2]));
clk_quad_buf iclk_colbuf_1_ ( .clki(clki[1]), .clko(clko[1]));
clk_quad_buf iclk_colbuf_0_ ( .clki(clki[0]), .clko(clko[0]));

endmodule
// Library - leafcell, Cell - bram_bufferx1, View - schematic
// LAST TIME SAVED: Jun 14 08:59:24 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module bram_bufferx1 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I0 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - leafcell, Cell - bram_4k_buffer, View - schematic
// LAST TIME SAVED: Aug 28 14:24:48 2008
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module bram_4k_buffer ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;

input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



tielo I21 ( .tielo(net055));
bram_bufferx1 I15 ( .in(net055), .out(net49));
bram_bufferx1 I16 ( .in(net49), .out(net52));
bram_bufferx1 I17 ( .in(net52), .out(net53));
bram_bufferx1 I18 ( .in(net53), .out(net55));
bram_bufferx6 I14 ( .in(bm_sdo_i), .out(bm_sdo_o));
bram_bufferx6 I6 ( .in(bm_sdi_i), .out(bm_sdi_o));
bram_bufferx6 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx6 I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx6 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx6 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx6 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx6 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx6 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx6 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx6 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx6 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx6 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx6 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx6 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx6 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx6 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jun  5 11:34:46 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module leafcell_ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - leafcell, Cell - bram_bufferx16, View - schematic
// LAST TIME SAVED: Jun 25 13:49:31 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module bram_bufferx16 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I0 ( .A(net07), .Y(net09));
inv_hvt I2 ( .A(in), .Y(net07));
inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(net09), .Y(net6));

endmodule
// Library - leafcell, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:59 2007
// NETLIST TIME: Nov 14 16:12:01 2008
`timescale 1ns / 1ns 

module ml_mux2_hvt_schematic ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - bram_dff_mux, View - schematic
// LAST TIME SAVED: Jul 25 16:06:22 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_dff_mux ( q, bm_q, bm_sdi, ce, clk, rcapmux_en, rst );
output  q;

input  bm_q, bm_sdi, ce, clk, rcapmux_en, rst;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



leafcell_ml_dff_schematic I2 ( .R(rst), .D(net020), .CLK(clk),
     .QN(net10), .Q(q));
ml_mux2_hvt_schematic I5 ( .in1(net14), .in0(q), .out(net020),
     .sel(ce));
ml_mux2_hvt_schematic I1 ( .in1(bm_q), .in0(bm_sdi), .out(net14),
     .sel(rcapmux_en));

endmodule
// Library - leafcell, Cell - bram_4k_sr_bankout, View - schematic
// LAST TIME SAVED: Jul 25 22:59:22 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_sr_bankout ( bm_dm, bm_sdo, bm_sweb, clk, rcapmux_en,
     rst, bm_q, bm_sdi, wdummymux_en );
output  bm_sdo;

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[0]), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));
leafcell_ml_dff_schematic I29 ( .R(rst), .D(net0151), .CLK(clk),
     .QN(net0160), .Q(bm_sdo));
leafcell_ml_dff_schematic I22 ( .R(rst), .D(bm_dm[14]), .CLK(clk),
     .QN(net165), .Q(rdummy_reg));
ml_mux2_hvt_schematic I21 ( .in1(rdummy_reg), .in0(bm_dm[15]),
     .out(net0151), .sel(rdummymux_en));
nor2_hvt I24 ( .A(bm_swe), .B(rcapmux_en), .Y(net148));
inv_hvt I19 ( .A(bm_sweb), .Y(bm_swe));
inv_hvt I23 ( .A(net148), .Y(rdummymux_en));

endmodule
// Library - leafcell, Cell - rf_4k, View - schematic
// LAST TIME SAVED: Aug 15 17:39:16 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module rf_4k ( Q, AA, AB, AMA, AMB, BIST, BWEB, BWEBM, CLKR, CLKW, D,
     DM, REB, REBM, WEB, WEBM );

input  BIST, CLKR, CLKW, REB, REBM, WEB, WEBM;

output [15:0]  Q;

input [7:0]  AMA;
input [15:0]  BWEBM;
input [15:0]  DM;
input [7:0]  AA;
input [15:0]  D;
input [15:0]  BWEB;
input [7:0]  AMB;
input [7:0]  AB;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - bram_4k_bankout, View - schematic
// LAST TIME SAVED: Aug 15 18:09:39 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_bankout ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_ab;
input [7:0]  bm_sa;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [15:0]  bm_dm;



tielo I15 ( .tielo(net092));
tielo I18 ( .tielo(net093));
bram_4k_sr_bankout I12 ( .bm_dm(bm_dm[15:0]), .rst(net093),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]), .bm_sdo(bm_sdo));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM(bm_dm[15:0]), .WEBM(bm_sweb), .WEB(web), .REBM(bm_sreb),
     .REB(reb), .D(bm_d[15:0]), .CLKW(net074), .CLKR(net072),
     .BWEBM({net092, net092, net092, net092, net092, net092, net092,
     net092, net092, net092, net092, net092, net092, net092, net092,
     net092}), .BWEB(bm_bweb[15:0]), .BIST(bm_init), .AMB(bm_sa[7:0]),
     .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]), .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net89), .out(net072));
bram_bufferx6 I8 ( .in(net85), .out(net074));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net85), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net89), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbankout_pbuffer_bot, View -
//schematic
// LAST TIME SAVED: Aug 24 17:34:26 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4kbankout_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;

input [7:0]  bm_aa;
input [15:0]  bm_bweb;
input [7:0]  bm_sa_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sclkrw_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [1:0]  bm_sweb_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankout I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - xpmem, Cell - cram2x2x6, View - schematic
// LAST TIME SAVED: Jul 28 08:29:06 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module cram2x2x6 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [23:0]  q;
output [23:0]  q_b;

inout [11:0]  bl;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  r_gnd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_5_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_base, View - schematic
// LAST TIME SAVED: Sep 13 06:51:33 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_base ( lc_trk_out, sp4_out, bl, min0, min1, min2,
     min3, pgate, prog, reset_b, sp12_in, vdd_cntl, wl );


input  prog;

output [1:0]  sp4_out;
output [3:0]  lc_trk_out;

inout [11:0]  bl;

input [1:0]  wl;
input [1:0]  sp12_in;
input [15:0]  min1;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [15:0]  min3;
input [1:0]  pgate;
input [15:0]  min0;
input [15:0]  min2;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  cbitb;

wire  [23:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
g_mux Imux2 ( .min(min2[15:0]), .prog(net60), .inmuxo(lc_trk_out[2]),
     .cbit({cbit[16], cbit[17], cbit[20], cbit[23], cbit[21]}),
     .cbitb({cbitb[16], cbitb[17], cbitb[20], cbitb[23], cbitb[21]}));
g_mux Imux3 ( .min(min3[15:0]), .prog(net60), .inmuxo(lc_trk_out[3]),
     .cbit({cbit[18], cbit[19], cbit[22], cbit[15], cbit[13]}),
     .cbitb({cbitb[18], cbitb[19], cbitb[22], cbitb[15], cbitb[13]}));
g_mux Imux1 ( .min(min1[15:0]), .prog(net60), .inmuxo(lc_trk_out[1]),
     .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}));
g_mux Imux0 ( .min(min0[15:0]), .prog(net60), .inmuxo(lc_trk_out[0]),
     .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}));
cram2x2x6 Imem2x2x6 ( .pgate(pgate[1:0]), .q(cbit[23:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[11:0]), .q_b(cbitb[23:0]));
sp12to4 Isp12to4_1_ ( .triout(sp4_out[1]), .cbitb(cbitb[11]),
     .drv(sp12_in[1]), .prog(net60));
sp12to4 Isp12to4_0_ ( .triout(sp4_out[0]), .cbitb(cbitb[9]),
     .drv(sp12_in[0]), .prog(net60));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net60));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0a, View - schematic
// LAST TIME SAVED: Jul 24 13:27:07 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g0a ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g0;

inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;

input [7:0]  tnl_op;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[34], sp4_r_v_b[25]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[33], sp4_r_v_b[26]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[35], sp4_r_v_b[24]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[32], sp4_r_v_b[27]}),
     .sp4_out(sp4_v_b[13:12]), .sp12_in({sp12_v_b[3], sp12_v_b[1]}),
     .lc_trk_out(lc_trk_g0[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0b, View - schematic
// LAST TIME SAVED: Jul 24 13:26:14 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g0b ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, glb2local, lft_op,
     pgate, prog, reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op,
     vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g0;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
input [3:0]  glb2local;
input [7:0]  bnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  top_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], glb2local[1]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], glb2local[2]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], glb2local[0]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], glb2local[3]}),
     .sp4_out(sp4_v_b[15:14]), .sp12_in({sp12_v_b[7], sp12_v_b[5]}),
     .lc_trk_out(lc_trk_g0[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - xpmem, Cell - ml_cram_logic, View - schematic
// LAST TIME SAVED: Sep 28 20:58:40 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_cram_logic ( cram_pgateoff, cram_prec, cram_pullup_b,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, smc_clk_out, por,
     smc_clk, smc_read, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rwl_en, smc_seq_rst, smc_wcram_rst, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en );
output  cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, smc_clk_out;

input  por, smc_clk, smc_read, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_write, smc_wset_prec, smc_wset_precgnd, smc_wwlwrt_dis,
     smc_wwlwrt_en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I213 ( .A(net208), .Y(net177), .B(net248));
inv_hvt I370 ( .A(net273), .Y(rst_rpull_rwl));
inv_hvt I373 ( .A(cram_rst), .Y(net257));
inv_hvt I346 ( .A(net315), .Y(net220));
inv_hvt I263 ( .A(net269), .Y(net218));
inv_hvt I266 ( .A(cram_write_int), .Y(net216));
inv_hvt I286 ( .A(net359), .Y(net299));
inv_hvt I422 ( .A(smc_rwl_en), .Y(net212));
inv_hvt I323 ( .A(net282), .Y(net210));
inv_hvt I378 ( .A(net276), .Y(net248));
inv_hvt I333 ( .A(net279), .Y(net208));
inv_hvt I324 ( .A(net210), .Y(cram_pgateoff));
inv_hvt I403 ( .A(net285), .Y(net204));
inv_hvt I292 ( .A(net200), .Y(cram_prec));
inv_hvt I267 ( .A(net303), .Y(net200));
inv_hvt I224 ( .A(net291), .Y(reset_logic));
inv_hvt I401 ( .A(net294), .Y(net196));
inv_hvt I381 ( .A(net309), .Y(net194));
inv_hvt I268 ( .A(net257), .Y(net253));
inv_hvt I293 ( .A(net236), .Y(cram_vddoff));
inv_hvt I269 ( .A(net255), .Y(net251));
inv_hvt I330 ( .A(net265), .Y(net190));
inv_hvt I374 ( .A(net253), .Y(net255));
inv_hvt I294 ( .A(cram_rst_int_b), .Y(cram_rst));
inv_hvt I375 ( .A(net252), .Y(cram_rst_dly));
inv_hvt I421 ( .A(net394), .Y(net186));
inv_hvt I249 ( .A(net262), .Y(net184));
inv_hvt I250 ( .A(net184), .Y(cram_pullup_b));
inv_hvt I359 ( .A(net179), .Y(net180));
inv_hvt I376 ( .A(net251), .Y(net252));
inv_hvt I336 ( .A(smc_clk), .Y(sm_clk_b));
inv_hvt I367 ( .A(net306), .Y(dis_pgatewrt));
inv_hvt I281 ( .A(net399), .Y(net226));
inv_hvt I399 ( .A(net300), .Y(net240));
inv_hvt I290 ( .A(net218), .Y(cram_wl_en));
inv_hvt I425 ( .A(net299), .Y(net262));
inv_hvt I337 ( .A(sm_clk_b), .Y(smc_clk_out));
inv_hvt I256 ( .A(net379), .Y(cram_write_int));
inv_hvt I291 ( .A(net216), .Y(cram_write));
inv_hvt I415 ( .A(net312), .Y(net260));
inv_hvt I312 ( .A(net177), .Y(net228));
inv_hvt I270 ( .A(net228), .Y(net236));
inv_hvt I271 ( .A(net226), .Y(cram_rst_int_b));
mux2_hvt I161 ( .in1(cram_write_int), .in0(net186), .out(net269),
     .sel(net208));
mux2_hvt I295 ( .in1(net194), .in0(net220), .out(net265),
     .sel(net208));
nor2_hvt I402 ( .A(net283), .B(smc_wset_precgnd), .Y(net285));
nor2_hvt I329 ( .A(net190), .B(smc_seq_rst), .Y(net303));
nor2_hvt I398 ( .A(smc_rpull_b), .B(net299), .Y(net300));
nor2_hvt I393 ( .A(cram_rst_dly), .B(reset_logic), .Y(net179));
nor2_hvt I364 ( .A(net389), .B(smc_seq_rst), .Y(net282));
nor2_hvt I400 ( .A(net292), .B(smc_wset_prec), .Y(net294));
nor2_hvt I366 ( .A(reset_logic), .B(net370), .Y(net306));
nor2_hvt I223 ( .A(net318), .B(por), .Y(net291));
nor2_hvt I390 ( .A(smc_write), .B(smc_seq_rst), .Y(net279));
nor2_hvt I392 ( .A(net283), .B(cram_rst), .Y(net276));
nor2_hvt I389 ( .A(net375), .B(reset_logic), .Y(net273));
nor2_hvt I385 ( .A(smc_rprec), .B(net287), .Y(net315));
nor2_hvt I414 ( .A(net310), .B(smc_wwlwrt_en), .Y(net312));
nor2_hvt I391 ( .A(net292), .B(cram_rst), .Y(net309));
nor3_hvt I220 ( .B(net322), .Y(net326), .A(net322), .C(net322));
nor3_hvt I217 ( .B(net401), .Y(net330), .A(net401), .C(net401));
nor3_hvt I386 ( .B(smc_seq_rst), .Y(net318), .A(smc_write),
     .C(smc_read));
nor3_hvt I218 ( .B(net330), .Y(net322), .A(net330), .C(net330));
nor3_hvt I387 ( .B(smc_rwl_en), .Y(net287), .A(net315),
     .C(reset_logic));
nand3_hvt I230 ( .Y(net348), .B(net344), .C(net344), .A(net344));
nand3_hvt I231 ( .Y(net352), .B(net348), .C(net348), .A(net348));
nand3_hvt I426 ( .Y(net344), .B(net401), .C(net401), .A(net401));
ml_dff_schematic I411 ( .R(reset_logic), .D(smc_wwlwrt_dis),
     .CLK(smc_clk), .QN(net369), .Q(net370));
ml_dff_schematic I408 ( .R(rst_rpull_rwl), .D(net401), .CLK(net212),
     .QN(net394), .Q(net395));
ml_dff_schematic I405 ( .R(dis_pgatewrt), .D(net401),
     .CLK(cram_rst_int_b), .QN(net389), .Q(net390));
ml_dff_schematic I412 ( .R(net180), .D(net196), .CLK(smc_clk_out),
     .QN(net337), .Q(net292));
ml_dff_schematic I410 ( .R(dis_pgatewrt), .D(net260),
     .CLK(smc_clk_out), .QN(net379), .Q(net310));
ml_dff_schematic I108 ( .R(reset_logic), .D(smc_rrst_pullwlen),
     .CLK(smc_clk_out), .QN(net343), .Q(net375));
ml_dff_schematic I413 ( .R(net180), .D(net204), .CLK(smc_clk_out),
     .QN(net333), .Q(net283));
ml_dff_schematic I407 ( .R(rst_rpull_rwl), .D(net240),
     .CLK(smc_clk_out), .QN(net359), .Q(net360));
ml_dff_schematic I406 ( .R(reset_logic), .D(smc_wcram_rst),
     .CLK(smc_clk_out), .QN(net399), .Q(net400));
tiehi I427 ( .tiehi(net401));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1a, View - schematic
// LAST TIME SAVED: Jul 24 13:25:29 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g1a ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [1:0]  wl;
input [7:0]  bnl_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[25], sp4_r_v_b[1]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[26], sp4_r_v_b[2]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[24], sp4_r_v_b[0]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[27], sp4_r_v_b[3]}),
     .sp4_out(sp4_v_b[17:16]), .sp12_in({sp12_v_b[11], sp12_v_b[9]}),
     .lc_trk_out(lc_trk_g1[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1b, View - schematic
// LAST TIME SAVED: Jul 24 13:24:39 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g1b ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], sp4_r_v_b[5]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], sp4_r_v_b[6]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], sp4_r_v_b[4]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], sp4_r_v_b[7]}),
     .sp4_out(sp4_v_b[19:18]), .sp12_in({sp12_v_b[15], sp12_v_b[13]}),
     .lc_trk_out(lc_trk_g1[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2a, View - schematic
// LAST TIME SAVED: Jul 24 13:23:46 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g2a ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g2;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;

input [7:0]  lft_op;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnl_op;
input [7:0]  slf_op;
input [1:0]  vdd_cntl;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  bnr_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[33], sp4_r_v_b[9]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[34], sp4_r_v_b[10]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[32], sp4_r_v_b[8]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[35], sp4_r_v_b[11]}),
     .sp4_out(sp4_v_b[21:20]), .sp12_in({sp12_v_b[19], sp12_v_b[17]}),
     .lc_trk_out(lc_trk_g2[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2b, View - schematic
// LAST TIME SAVED: Jul 24 13:22:58 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g2b ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g2;

inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [7:0]  bnr_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[37], sp4_r_v_b[13]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[38], sp4_r_v_b[14]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[36], sp4_r_v_b[12]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[39], sp4_r_v_b[15]}),
     .sp4_out(sp4_v_b[23:22]), .sp12_in({sp12_v_b[23], sp12_v_b[21]}),
     .lc_trk_out(lc_trk_g2[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3a, View - schematic
// LAST TIME SAVED: Jul 24 13:22:20 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g3a ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g3;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  vdd_cntl;
input [7:0]  bnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  bnl_op;
input [7:0]  tnr_op;
input [7:0]  bot_op;
input [1:0]  wl;
input [7:0]  slf_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[41], sp4_r_v_b[17]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[42], sp4_r_v_b[18]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[40], sp4_r_v_b[16]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[43], sp4_r_v_b[19]}),
     .sp4_out(sp4_h_r[13:12]), .sp12_in({sp12_h_r[2], sp12_h_r[0]}),
     .lc_trk_out(lc_trk_g3[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3b, View - schematic
// LAST TIME SAVED: Jul 24 13:21:26 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g3b ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g3;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;

input [7:0]  top_op;
input [7:0]  bnr_op;
input [1:0]  reset_b;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[45], sp4_r_v_b[21]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[46], sp4_r_v_b[22]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[44], sp4_r_v_b[20]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[47], sp4_r_v_b[23]}),
     .sp4_out(sp4_h_r[15:14]), .sp12_in({sp12_h_r[6], sp12_h_r[4]}),
     .lc_trk_out(lc_trk_g3[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4, View - schematic
// LAST TIME SAVED: Jul 25 23:13:29 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module gmux_sp12to4 ( lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, bl,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bnl_op, bnr_op,
     bot_op, glb2local, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g3;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  slf_op;
input [7:0]  top_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  bot_op;
input [7:0]  lft_op;
input [7:0]  tnl_op;
input [7:0]  bnr_op;
input [3:0]  glb2local;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  reset_b;
input [7:0]  bnl_op;
input [15:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_g0a Ig0_30 ( .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_v_b(sp12_v_b[23:0]),
     .lc_trk_g0(lc_trk_g0[3:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[1:0]), .reset_b(reset_b[1:0]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g0b Ig0_74 ( .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]),
     .glb2local(glb2local[3:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .lc_trk_g0(lc_trk_g0[7:4]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g1a Ig1_30 ( .vdd_cntl(vdd_cntl[5:4]), .pgate(pgate[5:4]),
     .bl(bl[11:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]),
     .lft_op(lft_op[7:0]), .prog(prog), .rgt_op(rgt_op[7:0]),
     .reset_b(reset_b[5:4]), .slf_op(slf_op[7:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .wl(wl[5:4]), .lc_trk_g1(lc_trk_g1[3:0]));
gmux_sp12to4_g1b Ig1_74 ( .vdd_cntl(vdd_cntl[7:6]), .pgate(pgate[7:6]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .lc_trk_g1(lc_trk_g1[7:4]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[7:6]), .reset_b(reset_b[7:6]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g2a Ig2_30 ( .vdd_cntl(vdd_cntl[9:8]), .wl(wl[9:8]),
     .reset_b(reset_b[9:8]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[3:0]), .pgate(pgate[9:8]));
gmux_sp12to4_g2b Ig2_74 ( .vdd_cntl(vdd_cntl[11:10]),
     .pgate(pgate[11:10]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[11:10]),
     .reset_b(reset_b[11:10]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g3a Ig3_30 ( .vdd_cntl(vdd_cntl[13:12]), .wl(wl[13:12]),
     .reset_b(reset_b[13:12]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .pgate(pgate[13:12]), .lc_trk_g3(lc_trk_g3[3:0]));
gmux_sp12to4_g3b Ig3_74 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g3(lc_trk_g3[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .prog(prog),
     .bl(bl[11:0]), .reset_b(reset_b[15:14]), .wl(wl[15:14]));

endmodule
// Library - xpmem, Cell - cram2x2x5, View - schematic
// LAST TIME SAVED: Jul 28 08:25:47 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module cram2x2x5 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [19:0]  q_b;
output [19:0]  q;

inout [9:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  r_gnd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - sbox11to9_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:54:03 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox11to9_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[4]), .in5(t[10]), .in4(r[2]), .in3(r[10]),
     .in2(r[7]), .in1(b[10]), .in0(b[5]), .out(l[10]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[5]), .in5(t[11]), .in4(r[3]), .in3(r[11]),
     .in2(r[8]), .in1(b[11]), .in0(b[6]), .out(l[11]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[3]), .in5(t[9]), .in4(r[1]), .in3(r[9]),
     .in2(r[6]), .in1(b[9]), .in0(b[4]), .out(l[9]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[3]), .in5(r[9]), .in4(b[1]), .in3(b[9]),
     .in2(b[6]), .in1(l[9]), .in0(l[4]), .out(t[9]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[5]), .in5(r[11]), .in4(b[3]), .in3(b[11]),
     .in2(b[8]), .in1(l[11]), .in0(l[6]), .out(t[11]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[4]), .in5(r[10]), .in4(b[2]), .in3(b[10]),
     .in2(b[7]), .in1(l[10]), .in0(l[5]), .out(t[10]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox11to9_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:53:32 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox11to9_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[4]), .in5(b[10]), .in4(l[2]), .in3(l[10]),
     .in2(l[7]), .in1(t[10]), .in0(t[5]), .out(r[10]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[5]), .in5(b[11]), .in4(l[3]), .in3(l[11]),
     .in2(l[8]), .in1(t[11]), .in0(t[6]), .out(r[11]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[3]), .in5(b[9]), .in4(l[1]), .in3(l[9]),
     .in2(l[6]), .in1(t[9]), .in0(t[4]), .out(r[9]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[4]), .in5(l[10]), .in4(t[2]), .in3(t[10]),
     .in2(t[7]), .in1(r[10]), .in0(r[5]), .out(b[10]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[5]), .in5(l[11]), .in4(t[3]), .in3(t[11]),
     .in2(t[8]), .in1(r[11]), .in0(r[6]), .out(b[11]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[3]), .in5(l[9]), .in4(t[1]), .in3(t[9]),
     .in2(t[6]), .in1(r[9]), .in0(r[4]), .out(b[9]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tiehigh, View - schematic
// LAST TIME SAVED: May  8 16:23:56 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module vdd_tiehigh ( vdd_tieh );
inout  vdd_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(vdd_tieh), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - leafcell, Cell - sbox8to6_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:52:49 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox8to6_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[1]), .in5(t[7]), .in4(r[11]), .in3(r[7]),
     .in2(r[4]), .in1(b[7]), .in0(b[2]), .out(l[7]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[2]), .in5(t[8]), .in4(r[0]), .in3(r[8]),
     .in2(r[5]), .in1(b[8]), .in0(b[3]), .out(l[8]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[0]), .in5(t[6]), .in4(r[10]), .in3(r[6]),
     .in2(r[3]), .in1(b[6]), .in0(b[1]), .out(l[6]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[0]), .in5(r[6]), .in4(b[10]), .in3(b[6]),
     .in2(b[3]), .in1(l[6]), .in0(l[1]), .out(t[6]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[2]), .in5(r[8]), .in4(b[0]), .in3(b[8]),
     .in2(b[5]), .in1(l[8]), .in0(l[3]), .out(t[8]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[1]), .in5(r[7]), .in4(b[11]), .in3(b[7]),
     .in2(b[4]), .in1(l[7]), .in0(l[2]), .out(t[7]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox8to6_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:36:51 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox8to6_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  cbit;

wire  [19:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[1]), .in5(b[7]), .in4(l[11]), .in3(l[7]),
     .in2(l[4]), .in1(t[7]), .in0(t[2]), .out(r[7]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[2]), .in5(b[8]), .in4(l[0]), .in3(l[8]),
     .in2(l[5]), .in1(t[8]), .in0(t[3]), .out(r[8]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[0]), .in5(b[6]), .in4(l[10]), .in3(l[6]),
     .in2(l[3]), .in1(t[6]), .in0(t[1]), .out(r[6]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[1]), .in5(l[7]), .in4(t[11]), .in3(t[7]),
     .in2(t[4]), .in1(r[7]), .in0(r[2]), .out(b[7]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[2]), .in5(l[8]), .in4(t[0]), .in3(t[8]),
     .in2(t[5]), .in1(r[8]), .in0(r[3]), .out(b[8]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[0]), .in5(l[6]), .in4(t[10]), .in3(t[6]),
     .in2(t[3]), .in1(r[6]), .in0(r[1]), .out(b[6]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox5to3_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:36:06 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox5to3_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  t;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[10]), .in5(t[4]), .in4(r[8]), .in3(r[4]),
     .in2(r[1]), .in1(b[4]), .in0(b[11]), .out(l[4]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[11]), .in5(t[5]), .in4(r[9]), .in3(r[5]),
     .in2(r[2]), .in1(b[5]), .in0(b[0]), .out(l[5]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[9]), .in5(t[3]), .in4(r[7]), .in3(r[3]),
     .in2(r[0]), .in1(b[3]), .in0(b[10]), .out(l[3]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[9]), .in5(r[3]), .in4(b[7]), .in3(b[3]),
     .in2(b[0]), .in1(l[3]), .in0(l[10]), .out(t[3]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[11]), .in5(r[5]), .in4(b[9]), .in3(b[5]),
     .in2(b[2]), .in1(l[5]), .in0(l[0]), .out(t[5]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[10]), .in5(r[4]), .in4(b[8]), .in3(b[4]),
     .in2(b[1]), .in1(l[4]), .in0(l[11]), .out(t[4]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 I534 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - sbox5to3_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:35:35 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox5to3_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbitb;

wire  [19:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[10]), .in5(b[4]), .in4(l[8]), .in3(l[4]),
     .in2(l[1]), .in1(t[4]), .in0(t[11]), .out(r[4]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[11]), .in5(b[5]), .in4(l[9]), .in3(l[5]),
     .in2(l[2]), .in1(t[5]), .in0(t[0]), .out(r[5]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[9]), .in5(b[3]), .in4(l[7]), .in3(l[3]),
     .in2(l[0]), .in1(t[3]), .in0(t[10]), .out(r[3]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[10]), .in5(l[4]), .in4(t[8]), .in3(t[4]),
     .in2(t[1]), .in1(r[4]), .in0(r[11]), .out(b[4]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[11]), .in5(l[5]), .in4(t[9]), .in3(t[5]),
     .in2(t[2]), .in1(r[5]), .in0(r[0]), .out(b[5]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[9]), .in5(l[3]), .in4(t[7]), .in3(t[3]),
     .in2(t[0]), .in1(r[3]), .in0(r[10]), .out(b[3]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox2to0_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:35:04 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox2to0_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  l;
inout [11:0]  b;
inout [11:0]  t;
inout [11:0]  r;

input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[7]), .in5(t[1]), .in4(r[5]), .in3(r[1]),
     .in2(r[10]), .in1(b[1]), .in0(b[8]), .out(l[1]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[8]), .in5(t[2]), .in4(r[6]), .in3(r[2]),
     .in2(r[11]), .in1(b[2]), .in0(b[9]), .out(l[2]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[6]), .in5(t[0]), .in4(r[4]), .in3(r[0]),
     .in2(r[9]), .in1(b[0]), .in0(b[7]), .out(l[0]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[6]), .in5(r[0]), .in4(b[4]), .in3(b[0]),
     .in2(b[9]), .in1(l[0]), .in0(l[7]), .out(t[0]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[8]), .in5(r[2]), .in4(b[6]), .in3(b[2]),
     .in2(b[11]), .in1(l[2]), .in0(l[9]), .out(t[2]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[7]), .in5(r[1]), .in4(b[5]), .in3(b[1]),
     .in2(b[10]), .in1(l[1]), .in0(l[8]), .out(t[1]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox2to0_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:34:25 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox2to0_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;
inout [9:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  cbit;

wire  [19:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[7]), .in5(b[1]), .in4(l[5]), .in3(l[1]),
     .in2(l[10]), .in1(t[1]), .in0(t[8]), .out(r[1]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[8]), .in5(b[2]), .in4(l[6]), .in3(l[2]),
     .in2(l[11]), .in1(t[2]), .in0(t[9]), .out(r[2]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[6]), .in5(b[0]), .in4(l[4]), .in3(l[0]),
     .in2(l[9]), .in1(t[0]), .in0(t[7]), .out(r[0]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[7]), .in5(l[1]), .in4(t[5]), .in3(t[1]),
     .in2(t[10]), .in1(r[1]), .in0(r[8]), .out(b[1]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[8]), .in5(l[2]), .in4(t[6]), .in3(t[2]),
     .in2(t[11]), .in1(r[2]), .in0(r[9]), .out(b[2]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[6]), .in5(l[0]), .in4(t[4]), .in3(t[0]),
     .in2(t[9]), .in1(r[0]), .in0(r[7]), .out(b[0]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - span4_switchandmem, View - schematic
// LAST TIME SAVED: Jul 24 12:49:53 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module span4_switchandmem ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;
inout [11:0]  r;

input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sbox11to9_220_p2 I73 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .l(l[11:0]), .r(r[11:0]), .t(t[11:0]),
     .b(b[11:0]), .prog(prog), .wl(wl[15:14]), .bl(bl[9:0]),
     .reset_b(reset_b[15:14]));
sbox11to9_220_p1 I75 ( .vdd_cntl(vdd_cntl[13:12]),
     .pgate(pgate[13:12]), .l(l[11:0]), .r(r[11:0]), .t(t[11:0]),
     .b(b[11:0]), .prog(prog), .wl(wl[13:12]), .bl(bl[9:0]),
     .reset_b(reset_b[13:12]));
sbox8to6_220_p2 I74 ( .vdd_cntl(vdd_cntl[11:10]), .pgate(pgate[11:10]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[11:10]), .bl(bl[9:0]), .reset_b(reset_b[11:10]));
sbox8to6_220_p1 I76 ( .vdd_cntl(vdd_cntl[9:8]), .pgate(pgate[9:8]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[9:8]), .bl(bl[9:0]), .reset_b(reset_b[9:8]));
sbox5to3_220_p2 I71 ( .vdd_cntl(vdd_cntl[7:6]), .pgate(pgate[7:6]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[7:6]), .bl(bl[9:0]), .reset_b(reset_b[7:6]));
sbox5to3_220_p1 I72 ( .vdd_cntl(vdd_cntl[5:4]), .pgate(pgate[5:4]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[5:4]), .bl(bl[9:0]), .reset_b(reset_b[5:4]));
sbox2to0_220_p2 I70 ( .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[3:2]), .bl(bl[9:0]), .reset_b(reset_b[3:2]));
sbox2to0_220_p1 I69 ( .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[1:0]), .bl(bl[9:0]), .reset_b(reset_b[1:0]));

endmodule
// Library - leafcell, Cell - span4, View - schematic
// LAST TIME SAVED: Sep  5 23:05:28 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module span4 ( bl, sp4_h_l, sp4_h_r, sp4_v_b, sp4_v_t, pgate, prog,
     reset_b, vdd_cntl, wl );

input  prog;

inout [47:0]  sp4_v_b;
inout [9:0]  bl;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_t;
inout [47:0]  sp4_h_r;

input [15:0]  vdd_cntl;
input [15:0]  reset_b;
input [15:0]  wl;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  sp4_h_r_mid;

wire  [11:0]  sp4_v_b_mid;



rm7  R1_27_ ( .MINUS(sp4_h_r[47]), .PLUS(sp4_h_l[34]));
rm7  R1_26_ ( .MINUS(sp4_h_r[46]), .PLUS(sp4_h_l[35]));
rm7  R1_25_ ( .MINUS(sp4_h_r[45]), .PLUS(sp4_h_l[32]));
rm7  R1_24_ ( .MINUS(sp4_h_r[44]), .PLUS(sp4_h_l[33]));
rm7  R1_23_ ( .MINUS(sp4_h_r[43]), .PLUS(sp4_h_l[30]));
rm7  R1_22_ ( .MINUS(sp4_h_r[42]), .PLUS(sp4_h_l[31]));
rm7  R1_21_ ( .MINUS(sp4_h_r[41]), .PLUS(sp4_h_l[28]));
rm7  R1_20_ ( .MINUS(sp4_h_r[40]), .PLUS(sp4_h_l[29]));
rm7  R1_19_ ( .MINUS(sp4_h_r[39]), .PLUS(sp4_h_l[26]));
rm7  R1_18_ ( .MINUS(sp4_h_r[38]), .PLUS(sp4_h_l[27]));
rm7  R1_17_ ( .MINUS(sp4_h_r[37]), .PLUS(sp4_h_l[24]));
rm7  R1_16_ ( .MINUS(sp4_h_r[36]), .PLUS(sp4_h_l[25]));
rm7  R1_15_ ( .MINUS(sp4_h_r[35]), .PLUS(sp4_h_l[22]));
rm7  R1_14_ ( .MINUS(sp4_h_r[34]), .PLUS(sp4_h_l[23]));
rm7  R1_13_ ( .MINUS(sp4_h_r[23]), .PLUS(sp4_h_l[10]));
rm7  R1_12_ ( .MINUS(sp4_h_r[22]), .PLUS(sp4_h_l[11]));
rm7  R1_11_ ( .MINUS(sp4_h_r_mid[11]), .PLUS(sp4_h_l[46]));
rm7  R1_10_ ( .MINUS(sp4_h_r_mid[10]), .PLUS(sp4_h_l[47]));
rm7  R1_9_ ( .MINUS(sp4_h_r_mid[9]), .PLUS(sp4_h_l[44]));
rm7  R1_8_ ( .MINUS(sp4_h_r_mid[8]), .PLUS(sp4_h_l[45]));
rm7  R1_7_ ( .MINUS(sp4_h_r_mid[7]), .PLUS(sp4_h_l[42]));
rm7  R1_6_ ( .MINUS(sp4_h_r_mid[6]), .PLUS(sp4_h_l[43]));
rm7  R1_5_ ( .MINUS(sp4_h_r_mid[5]), .PLUS(sp4_h_l[40]));
rm7  R1_4_ ( .MINUS(sp4_h_r_mid[4]), .PLUS(sp4_h_l[41]));
rm7  R1_3_ ( .MINUS(sp4_h_r_mid[3]), .PLUS(sp4_h_l[38]));
rm7  R1_2_ ( .MINUS(sp4_h_r_mid[2]), .PLUS(sp4_h_l[39]));
rm7  R1_1_ ( .MINUS(sp4_h_r_mid[1]), .PLUS(sp4_h_l[36]));
rm7  R1_0_ ( .MINUS(sp4_h_r_mid[0]), .PLUS(sp4_h_l[37]));
rm5  R2_19_ ( .MINUS(sp4_h_r[33]), .PLUS(sp4_h_l[20]));
rm5  R2_18_ ( .MINUS(sp4_h_r[32]), .PLUS(sp4_h_l[21]));
rm5  R2_17_ ( .MINUS(sp4_h_r[31]), .PLUS(sp4_h_l[18]));
rm5  R2_16_ ( .MINUS(sp4_h_r[30]), .PLUS(sp4_h_l[19]));
rm5  R2_15_ ( .MINUS(sp4_h_r[29]), .PLUS(sp4_h_l[16]));
rm5  R2_14_ ( .MINUS(sp4_h_r[28]), .PLUS(sp4_h_l[17]));
rm5  R2_13_ ( .MINUS(sp4_h_r[27]), .PLUS(sp4_h_l[14]));
rm5  R2_12_ ( .MINUS(sp4_h_r[26]), .PLUS(sp4_h_l[15]));
rm5  R2_11_ ( .MINUS(sp4_h_r[25]), .PLUS(sp4_h_l[12]));
rm5  R2_10_ ( .MINUS(sp4_h_r[24]), .PLUS(sp4_h_l[13]));
rm5  R2_9_ ( .MINUS(sp4_h_r[21]), .PLUS(sp4_h_l[8]));
rm5  R2_8_ ( .MINUS(sp4_h_r[20]), .PLUS(sp4_h_l[9]));
rm5  R2_7_ ( .MINUS(sp4_h_r[19]), .PLUS(sp4_h_l[6]));
rm5  R2_6_ ( .MINUS(sp4_h_r[18]), .PLUS(sp4_h_l[7]));
rm5  R2_5_ ( .MINUS(sp4_h_r[17]), .PLUS(sp4_h_l[4]));
rm5  R2_4_ ( .MINUS(sp4_h_r[16]), .PLUS(sp4_h_l[5]));
rm5  R2_3_ ( .MINUS(sp4_h_r[15]), .PLUS(sp4_h_l[2]));
rm5  R2_2_ ( .MINUS(sp4_h_r[14]), .PLUS(sp4_h_l[3]));
rm5  R2_1_ ( .MINUS(sp4_h_r[13]), .PLUS(sp4_h_l[0]));
rm5  R2_0_ ( .MINUS(sp4_h_r[12]), .PLUS(sp4_h_l[1]));
rm6  R0_47_ ( .MINUS(sp4_v_b[47]), .PLUS(sp4_v_t[34]));
rm6  R0_46_ ( .MINUS(sp4_v_b[46]), .PLUS(sp4_v_t[35]));
rm6  R0_45_ ( .MINUS(sp4_v_b[45]), .PLUS(sp4_v_t[32]));
rm6  R0_44_ ( .MINUS(sp4_v_b[44]), .PLUS(sp4_v_t[33]));
rm6  R0_43_ ( .MINUS(sp4_v_b[43]), .PLUS(sp4_v_t[30]));
rm6  R0_42_ ( .MINUS(sp4_v_b[42]), .PLUS(sp4_v_t[31]));
rm6  R0_41_ ( .MINUS(sp4_v_b[41]), .PLUS(sp4_v_t[28]));
rm6  R0_40_ ( .MINUS(sp4_v_b[40]), .PLUS(sp4_v_t[29]));
rm6  R0_39_ ( .MINUS(sp4_v_b[39]), .PLUS(sp4_v_t[26]));
rm6  R0_38_ ( .MINUS(sp4_v_b[38]), .PLUS(sp4_v_t[27]));
rm6  R0_37_ ( .MINUS(sp4_v_b[37]), .PLUS(sp4_v_t[24]));
rm6  R0_36_ ( .MINUS(sp4_v_b[36]), .PLUS(sp4_v_t[25]));
rm6  R0_35_ ( .MINUS(sp4_v_b[35]), .PLUS(sp4_v_t[22]));
rm6  R0_34_ ( .MINUS(sp4_v_b[34]), .PLUS(sp4_v_t[23]));
rm6  R0_33_ ( .MINUS(sp4_v_b[33]), .PLUS(sp4_v_t[20]));
rm6  R0_32_ ( .MINUS(sp4_v_b[32]), .PLUS(sp4_v_t[21]));
rm6  R0_31_ ( .MINUS(sp4_v_b[31]), .PLUS(sp4_v_t[18]));
rm6  R0_30_ ( .MINUS(sp4_v_b[30]), .PLUS(sp4_v_t[19]));
rm6  R0_29_ ( .MINUS(sp4_v_b[29]), .PLUS(sp4_v_t[16]));
rm6  R0_28_ ( .MINUS(sp4_v_b[28]), .PLUS(sp4_v_t[17]));
rm6  R0_27_ ( .MINUS(sp4_v_b[27]), .PLUS(sp4_v_t[14]));
rm6  R0_26_ ( .MINUS(sp4_v_b[26]), .PLUS(sp4_v_t[15]));
rm6  R0_25_ ( .MINUS(sp4_v_b[25]), .PLUS(sp4_v_t[12]));
rm6  R0_24_ ( .MINUS(sp4_v_b[24]), .PLUS(sp4_v_t[13]));
rm6  R0_23_ ( .MINUS(sp4_v_b[23]), .PLUS(sp4_v_t[10]));
rm6  R0_22_ ( .MINUS(sp4_v_b[22]), .PLUS(sp4_v_t[11]));
rm6  R0_21_ ( .MINUS(sp4_v_b[21]), .PLUS(sp4_v_t[8]));
rm6  R0_20_ ( .MINUS(sp4_v_b[20]), .PLUS(sp4_v_t[9]));
rm6  R0_19_ ( .MINUS(sp4_v_b[19]), .PLUS(sp4_v_t[6]));
rm6  R0_18_ ( .MINUS(sp4_v_b[18]), .PLUS(sp4_v_t[7]));
rm6  R0_17_ ( .MINUS(sp4_v_b[17]), .PLUS(sp4_v_t[4]));
rm6  R0_16_ ( .MINUS(sp4_v_b[16]), .PLUS(sp4_v_t[5]));
rm6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[2]));
rm6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[3]));
rm6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[0]));
rm6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[1]));
rm6  R0_11_ ( .MINUS(sp4_v_b_mid[11]), .PLUS(sp4_v_t[46]));
rm6  R0_10_ ( .MINUS(sp4_v_b_mid[10]), .PLUS(sp4_v_t[47]));
rm6  R0_9_ ( .MINUS(sp4_v_b_mid[9]), .PLUS(sp4_v_t[44]));
rm6  R0_8_ ( .MINUS(sp4_v_b_mid[8]), .PLUS(sp4_v_t[45]));
rm6  R0_7_ ( .MINUS(sp4_v_b_mid[7]), .PLUS(sp4_v_t[42]));
rm6  R0_6_ ( .MINUS(sp4_v_b_mid[6]), .PLUS(sp4_v_t[43]));
rm6  R0_5_ ( .MINUS(sp4_v_b_mid[5]), .PLUS(sp4_v_t[40]));
rm6  R0_4_ ( .MINUS(sp4_v_b_mid[4]), .PLUS(sp4_v_t[41]));
rm6  R0_3_ ( .MINUS(sp4_v_b_mid[3]), .PLUS(sp4_v_t[38]));
rm6  R0_2_ ( .MINUS(sp4_v_b_mid[2]), .PLUS(sp4_v_t[39]));
rm6  R0_1_ ( .MINUS(sp4_v_b_mid[1]), .PLUS(sp4_v_t[36]));
rm6  R0_0_ ( .MINUS(sp4_v_b_mid[0]), .PLUS(sp4_v_t[37]));
span4_switchandmem ISPAN4_SW ( .vdd_cntl(vdd_cntl[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]), .b(sp4_v_b[11:0]),
     .r(sp4_h_r[11:0]), .l(sp4_h_r_mid[11:0]), .prog(prog),
     .wl(wl[15:0]), .t(sp4_v_b_mid[11:0]), .bl(bl[9:0]));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev, View - schematic
// LAST TIME SAVED: Jul 24 09:36:22 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module clkmandcmuxrev ( cin2lcl, clk, clkb, glb2local, s_r, carry_in,
     cbit, cbitb, glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, min0, min1, min2, min3, prog );
output  cin2lcl, clk, clkb, s_r;

input  carry_in, prog;

output [3:0]  glb2local;

input [7:0]  min0;
input [7:0]  min3;
input [7:0]  glb_netwk;
input [31:0]  cbit;
input [31:0]  cbitb;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g0;
input [7:0]  min2;
input [7:0]  min1;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g3;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sr_clkm8to1 I296 ( .mout(s_r), .cbitb(cbitb[12:9]), .min({lc_trk_g3[5],
     lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4], glb_netwk[6],
     glb_netwk[4], glb_netwk[2], glb_netwk[0]}), .cbit(cbit[12:9]),
     .prog(prog));
ce_clkm8to1 I283 ( .moutb(ceb), .cbitb(cbitb[8:5]), .cbit(cbit[8:5]),
     .prog(prog), .min({lc_trk_g3[3], lc_trk_g2[2], lc_trk_g1[3],
     lc_trk_g0[2], glb_netwk[7], glb_netwk[5], glb_netwk[3],
     glb_netwk[1]}));
clk_mux12to1 I298 ( .cbitb({cbitb[31], cbitb[4], cbitb[3], cbitb[2],
     cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3], cbit[2],
     cbit[1], cbit[0]}), .prog(prog), .min({lc_trk_g3[1], lc_trk_g2[0],
     lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}), .clk(clk),
     .clkb(clkb), .cenb(ceb));
clk_mux8to1 I285 ( .min(min3[7:0]), .prog(prog), .inmuxo(glb2local[0]),
     .cbit(cbit[16:13]), .cbitb(cbitb[16:13]));
clk_mux8to1 I293 ( .prog(prog), .inmuxo(glb2local[1]), .min(min2[7:0]),
     .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I294 ( .prog(prog), .inmuxo(glb2local[2]), .min(min1[7:0]),
     .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
clk_mux8to1 I295 ( .prog(prog), .inmuxo(glb2local[3]), .min(min0[7:0]),
     .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));
mux_4carry Icarry_cnt ( .cin(carry_in), .lcl_cin(cin2lcl),
     .cbitb(cbitb[30:29]), .prog(prog), .cbit(cbit[30:29]));

endmodule
// Library - leafcell, Cell - sbox1, View - schematic
// LAST TIME SAVED: Jun  8 15:19:03 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module sbox1 ( b, l, r, t, c, cb, prog );
inout  b, l, r, t;

input  prog;

input [7:0]  cb;
input [7:0]  c;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sbox1m3to1 I232 ( .in2(r), .cb(cb[7:6]), .op(t), .in0(l), .in1(b),
     .c(c[7:6]), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb(cb[3:2]), .op(l), .in0(b), .in1(t),
     .c(c[3:2]), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb(cb[1:0]), .op(b), .in0(l), .in1(t),
     .c(c[1:0]), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb(cb[5:4]), .op(r), .in0(l), .in1(t),
     .c(c[5:4]), .prog(prog));

endmodule
// Library - EH_PUP_2, Cell - eh_io_pup_2_new, View - schematic
// LAST TIME SAVED: Oct  6 14:09:30 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module eh_io_pup_2_new ( por_b, core_por_b, vdd_io );
output  por_b;

input  core_por_b, vdd_io;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_hvt  MP8 ( .D(net104), .B(vdd_), .G(core_por_b), .S(vdd_));
pch_hvt  M4 ( .D(por_b), .B(vdd_), .G(net92), .S(vdd_));
pch_hvt  M1 ( .D(net92), .B(vdd_), .G(net84), .S(vdd_));
pch_hvt  M0 ( .D(net84), .B(vdd_), .G(net104), .S(vdd_));
nch_hvt  M5 ( .D(por_b), .B(gnd_), .G(net92), .S(gnd_));
nch_hvt  M3 ( .D(net92), .B(gnd_), .G(net84), .S(gnd_));
nch_hvt  MN1 ( .D(net80), .B(gnd_), .G(core_por_b), .S(gnd_));
nch_hvt  M2 ( .D(net84), .B(gnd_), .G(net104), .S(gnd_));
pch_25  M6 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  MP11 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
pch_25  MP13 ( .D(net124), .B(vdd_io), .G(net145), .S(net122));
pch_25  MP12 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  M7 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  MP7 ( .D(net104), .B(vdd_), .G(net124), .S(vdd_));
pch_25  MP9 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
nch_25  MN6 ( .D(net124), .B(gnd_), .G(net145), .S(gnd_));
nch_25  MN38 ( .D(net104), .B(gnd_), .G(net124), .S(net104));
nch_25  M10 ( .D(net124), .B(gnd_), .G(net147), .S(net158));
nch_25  MN39 ( .D(net104), .B(gnd_), .G(net124), .S(net80));
nch_25  M11 ( .D(net140), .B(gnd_), .G(core_por_b), .S(gnd_));
rppolywo_m  R66 ( .MINUS(gnd_), .PLUS(net145), .BULK(gnd_));
vdd_tiehigh I96 ( .vdd_tieh(net147));
nch_na25  M15 ( .D(net154), .B(gnd_), .G(net154), .S(net150));
nch_na25  M16 ( .D(net158), .B(gnd_), .G(net158), .S(net154));
nch_na25  M17 ( .D(net162), .B(gnd_), .G(net162), .S(net166));
nch_na25  M14 ( .D(net150), .B(gnd_), .G(net150), .S(net162));
nch_na25  M18 ( .D(net166), .B(gnd_), .G(net166), .S(net140));

endmodule
// Library - xpmem, Cell - cram16x4, View - schematic
// LAST TIME SAVED: Jul 28 08:31:30 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module cram16x4 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [63:0]  q_b;
output [63:0]  q;

inout [3:0]  bl;

input [15:0]  pgate;
input [15:0]  r_gnd;
input [15:0]  wl;
input [15:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 I16_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[1:0]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[15:14]));
cram2x2 I16_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[1:0]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[13:12]));
cram2x2 I16_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[1:0]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[11:10]));
cram2x2 I16_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[1:0]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[9:8]));
cram2x2 I16_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[1:0]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[7:6]));
cram2x2 I16_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[1:0]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[5:4]));
cram2x2 I16_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[1:0]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[3:2]));
cram2x2 I16_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[3:2]), .q_b(q_b[63:60]),
     .q(q[63:60]), .wl(wl[15:14]));
cram2x2 Imstake_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[3:2]), .q_b(q_b[59:56]),
     .q(q[59:56]), .wl(wl[13:12]));
cram2x2 Imstake_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[3:2]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[11:10]));
cram2x2 Imstake_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[3:2]), .q_b(q_b[51:48]), .q(q[51:48]),
     .wl(wl[9:8]));
cram2x2 Imstake_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[3:2]), .q_b(q_b[47:44]), .q(q[47:44]),
     .wl(wl[7:6]));
cram2x2 Imstake_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[3:2]), .q_b(q_b[43:40]), .q(q[43:40]),
     .wl(wl[5:4]));
cram2x2 Imstake_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[3:2]), .q_b(q_b[39:36]), .q(q[39:36]),
     .wl(wl[3:2]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[35:32]), .q(q[35:32]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - misc_module4rev, View - schematic
// LAST TIME SAVED: Aug 21 17:26:57 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module misc_module4rev ( S_R, cin2lcl, clk, clkb, glb2local, sp4, bl,
     b, carry_in, glb_netwk, l, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, m, min0, min1, min2, min3, pgate, prog, r, reset_b,
     sp12, vdd_cntl, wl );
output  S_R, cin2lcl, clk, clkb;


input  carry_in, prog;

output [7:0]  sp4;
output [3:0]  glb2local;

inout [3:0]  bl;

input [15:0]  reset_b;
input [15:0]  pgate;
input [7:0]  sp12;
input [1:0]  m;
input [7:0]  min0;
input [15:0]  vdd_cntl;
input [5:0]  lc_trk_g0;
input [1:0]  l;
input [5:0]  lc_trk_g2;
input [15:0]  wl;
input [1:0]  b;
input [7:0]  min3;
input [7:0]  glb_netwk;
input [7:0]  min1;
input [5:0]  lc_trk_g3;
input [5:0]  lc_trk_g1;
input [7:0]  min2;
input [1:0]  r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [63:0]  cbitb;

wire  [15:0]  r_vdd;

wire  [63:0]  cbit;



pch_hvt  vdd_cntrl_15_ ( .D(r_vdd[15]), .B(vdd_), .G(vdd_cntl[15]),
     .S(vdd_));
pch_hvt  vdd_cntrl_14_ ( .D(r_vdd[14]), .B(vdd_), .G(vdd_cntl[14]),
     .S(vdd_));
pch_hvt  vdd_cntrl_13_ ( .D(r_vdd[13]), .B(vdd_), .G(vdd_cntl[13]),
     .S(vdd_));
pch_hvt  vdd_cntrl_12_ ( .D(r_vdd[12]), .B(vdd_), .G(vdd_cntl[12]),
     .S(vdd_));
pch_hvt  vdd_cntrl_11_ ( .D(r_vdd[11]), .B(vdd_), .G(vdd_cntl[11]),
     .S(vdd_));
pch_hvt  vdd_cntrl_10_ ( .D(r_vdd[10]), .B(vdd_), .G(vdd_cntl[10]),
     .S(vdd_));
pch_hvt  vdd_cntrl_9_ ( .D(r_vdd[9]), .B(vdd_), .G(vdd_cntl[9]),
     .S(vdd_));
pch_hvt  vdd_cntrl_8_ ( .D(r_vdd[8]), .B(vdd_), .G(vdd_cntl[8]),
     .S(vdd_));
pch_hvt  vdd_cntrl_7_ ( .D(r_vdd[7]), .B(vdd_), .G(vdd_cntl[7]),
     .S(vdd_));
pch_hvt  vdd_cntrl_6_ ( .D(r_vdd[6]), .B(vdd_), .G(vdd_cntl[6]),
     .S(vdd_));
pch_hvt  vdd_cntrl_5_ ( .D(r_vdd[5]), .B(vdd_), .G(vdd_cntl[5]),
     .S(vdd_));
pch_hvt  vdd_cntrl_4_ ( .D(r_vdd[4]), .B(vdd_), .G(vdd_cntl[4]),
     .S(vdd_));
pch_hvt  vdd_cntrl_3_ ( .D(r_vdd[3]), .B(vdd_), .G(vdd_cntl[3]),
     .S(vdd_));
pch_hvt  vdd_cntrl_2_ ( .D(r_vdd[2]), .B(vdd_), .G(vdd_cntl[2]),
     .S(vdd_));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clkmandcmuxrev Itclkm ( .min2(min2[7:0]), .min1(min1[7:0]),
     .min0(min0[7:0]), .min3(min3[7:0]), .cbit({cbit[2], cbit[1],
     cbit[0], cbit[27], cbit[25], cbit[26], cbit[24], cbit[23],
     cbit[21], cbit[22], cbit[20], cbit[19], cbit[17], cbit[18],
     cbit[16], cbit[15], cbit[13], cbit[14], cbit[12], cbit[31],
     cbit[29], cbit[30], cbit[28], cbit[11], cbit[9], cbit[10],
     cbit[8], cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}), .glb2local(glb2local[3:0]),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .glb_netwk(glb_netwk[7:0]), .prog(prog), .cin2lcl(cin2lcl),
     .clk(clk), .clkb(clkb), .s_r(S_R), .carry_in(carry_in));
sp12to4 Isp12to4_7_ ( .triout(sp4[7]), .cbitb(cbitb[62]),
     .drv(sp12[7]), .prog(net109));
sp12to4 Isp12to4_6_ ( .triout(sp4[6]), .cbitb(cbitb[58]),
     .drv(sp12[6]), .prog(net109));
sp12to4 Isp12to4_5_ ( .triout(sp4[5]), .cbitb(cbitb[54]),
     .drv(sp12[5]), .prog(net109));
sp12to4 Isp12to4_4_ ( .triout(sp4[4]), .cbitb(cbitb[50]),
     .drv(sp12[4]), .prog(net109));
sp12to4 Isp12to4_3_ ( .triout(sp4[3]), .cbitb(cbitb[46]),
     .drv(sp12[3]), .prog(net109));
sp12to4 Isp12to4_2_ ( .triout(sp4[2]), .cbitb(cbitb[42]),
     .drv(sp12[2]), .prog(net109));
sp12to4 Isp12to4_1_ ( .triout(sp4[1]), .cbitb(cbitb[5]), .drv(sp12[1]),
     .prog(net109));
sp12to4 Isp12to4_0_ ( .triout(sp4[0]), .cbitb(cbitb[34]),
     .drv(sp12[0]), .prog(net109));
sbox1 Isp12_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(prog));
sbox1 Isp12_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(prog));
cram16x4 Ic64 ( .r_gnd(r_vdd[15:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .q(cbit[63:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net109));

endmodule
// Library - leafcell, Cell - bram_routing_tracks4rev, View - schematic
// LAST TIME SAVED: Aug 28 14:41:30 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_routing_tracks4rev ( clk, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, s_r, bl, sp4_h_l, sp4_h_r, sp4_r_v_b, sp4_v_b, sp4_v_t,
     sp12_h_l, sp12_h_r, sp12_v_b, sp12_v_t, bnl_op, bnr_op, bot_op,
     carry_in, glb_netwk, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );
output  clk, s_r;


input  carry_in, prog;

output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g3;
output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g2;

inout [23:0]  sp12_h_l;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_v_t;
inout [23:0]  sp12_v_t;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [25:0]  bl;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;

input [7:0]  rgt_op;
input [7:0]  bnl_op;
input [15:0]  reset_b;
input [7:0]  top_op;
input [15:0]  pgate;
input [7:0]  bot_op;
input [7:0]  glb_netwk;
input [7:0]  bnr_op;
input [7:0]  tnl_op;
input [7:0]  tnr_op;
input [15:0]  wl;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [15:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net_glb2local;

wire  [1:0]  sp12_h_r_mid;

wire  [1:0]  sp12_v_b_mid;



rm6  R0_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm6  R0_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm6  R0_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm6  R0_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm6  R0_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm6  R0_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm6  R0_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm6  R0_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm6  R0_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm6  R0_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm6  R0_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm6  R0_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm6  R0_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm6  R0_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm6  R0_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm6  R0_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm6  R0_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm6  R0_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm6  R0_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm6  R0_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm6  R0_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm6  R0_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm6  R0_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm6  R0_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
rm7  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
inv_hvt I89 ( .A(progb), .Y(progd));
inv_hvt I90 ( .A(prog), .Y(progb));
gmux_sp12to4 Igmux_sp12to4 ( .vdd_cntl(vdd_cntl[15:0]), .wl(wl[15:0]),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .prog(progd),
     .lft_op(lft_op[7:0]), .bnr_op(bnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .bot_op(bot_op[7:0]), .glb2local(net_glb2local[3:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]),
     .sp12_v_b(sp12_v_b[23:0]), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_r(sp4_h_r[47:0]));
span4 Isp4_sw ( .vdd_cntl(vdd_cntl[15:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_l(sp4_h_l[47:0]),
     .sp4_v_t(sp4_v_t[47:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .prog(progd), .wl(wl[15:0]), .bl(bl[21:12]));
misc_module4rev Ickmux_sp12to4_sp12sw ( .vdd_cntl(vdd_cntl[15:0]),
     .prog(progd), .carry_in(carry_in), .lc_trk_g0(lc_trk_g0[5:0]),
     .glb_netwk(glb_netwk[7:0]), .lc_trk_g2(lc_trk_g2[5:0]),
     .lc_trk_g3(lc_trk_g3[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .cin2lcl(net174), .wl(wl[15:0]), .S_R(s_r), .clkb(clkb),
     .bl(bl[25:22]), .clk(clk), .sp4(sp4_h_r[23:16]),
     .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18], sp12_h_r[16],
     sp12_h_r[14], sp12_h_r[12], sp12_h_r[10], sp12_h_r[8]}),
     .reset_b(reset_b[15:0]), .b(sp12_v_b[1:0]), .r(sp12_h_r[1:0]),
     .m(sp12_v_b_mid[1:0]), .l(sp12_h_r_mid[1:0]), .pgate(pgate[15:0]),
     .glb2local(net_glb2local[3:0]), .min2(glb_netwk[7:0]),
     .min1(glb_netwk[7:0]), .min0(glb_netwk[7:0]),
     .min3(glb_netwk[7:0]));

endmodule
// Library - leafcell, Cell - odrv12_30, View - schematic
// LAST TIME SAVED: Jun  5 15:34:53 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module odrv12_30 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_h_r;

input  prog, slfop;

output [2:0]  sp4_h_r;
output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_r_v_b;

input [11:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



odrv12 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b[1]));
odrv12 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp12(sp12_v_b[0]));
odrv12 I70 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r));
odrv4 I69_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I71_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[2]));
odrv4 I71_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[1]));
odrv4 I71_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp4(sp4_v_b[0]));
odrv4 I73_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I73_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I73_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux3_0, View - schematic
// LAST TIME SAVED: Aug 23 11:45:13 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_inmux3_0 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_h_r;

input  op, prog;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;

input [15:0]  min3;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [15:0]  min1;
input [15:0]  bl;
input [15:0]  min2;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [31:0]  cbitb;

wire  [31:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12_30 Iodrv74 ( .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
in_mux in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - odrv12_74, View - schematic
// LAST TIME SAVED: Jun  5 15:30:49 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module odrv12_74 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_v_b;

input  prog, slfop;

output [2:0]  sp4_v_b;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_h_r;

input [11:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



odrv12 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp12(sp12_h_r[1]));
odrv12 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r[0]));
odrv12 I71 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b));
odrv4 I68_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I68_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I68_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I70_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp4(sp4_v_b[2]));
odrv4 I70_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[1]));
odrv4 I70_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[0]));
odrv4 I72_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux7_4, View - schematic
// LAST TIME SAVED: Aug 23 11:44:11 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_inmux7_4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_v_b;

input  op, prog;

output [1:0]  sp12_h_r;
output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min3;
input [15:0]  min0;
input [15:0]  bl;
input [1:0]  vdd_cntl;
input [15:0]  min1;
input [1:0]  wl;
input [1:0]  pgate;
input [15:0]  min2;
input [1:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [31:0]  cbit;

wire  [31:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
odrv12_74 Iodrv74 ( .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));
in_mux in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux_8x4, View - schematic
// LAST TIME SAVED: Aug 29 16:20:56 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_inmux_8x4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, op, pgate, prog, reset_b, vdd_cntl, wl );

input  prog;

output [23:0]  sp4_r_v_b;
output [23:0]  sp4_h_r;
output [7:0]  in3;
output [7:0]  in2;
output [7:0]  in1;
output [11:0]  sp12_v_b;
output [11:0]  sp12_h_r;
output [23:0]  sp4_v_b;
output [7:0]  in0;

input [15:0]  bl;
input [7:0]  op;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g2;
input [15:0]  reset_b;
input [7:0]  lc_trk_g1;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [7:0]  lc_trk_g3;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_inmux3_0 I3 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[3]), .sp12_v_b(sp12_v_b[7:6]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(progd), .pgate(pgate[7:6]),
     .op(op[3]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[11:9]), .sp4_r_v_b(sp4_r_v_b[11:9]),
     .sp4_h_r(sp4_h_r[11:9]), .in3(in3[3]), .in2(in2[3]), .in1(in1[3]),
     .in0(in0[3]));
bram_4k_inmux3_0 I2 ( .vdd_cntl(vdd_cntl[5:4]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[2]), .sp12_v_b(sp12_v_b[5:4]), .wl(wl[5:4]),
     .reset_b(reset_b[5:4]), .prog(progd), .pgate(pgate[5:4]),
     .op(op[2]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[8:6]), .sp4_r_v_b(sp4_r_v_b[8:6]),
     .sp4_h_r(sp4_h_r[8:6]), .in3(in3[2]), .in2(in2[2]), .in1(in1[2]),
     .in0(in0[2]));
bram_4k_inmux3_0 I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[1]), .sp12_v_b(sp12_v_b[3:2]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(progd), .pgate(pgate[3:2]),
     .op(op[1]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[5:3]), .sp4_r_v_b(sp4_r_v_b[5:3]),
     .sp4_h_r(sp4_h_r[5:3]), .in3(in3[1]), .in2(in2[1]), .in1(in1[1]),
     .in0(in0[1]));
bram_4k_inmux3_0 I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[0]), .sp12_v_b(sp12_v_b[1:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(progd), .pgate(pgate[1:0]),
     .op(op[0]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .in3(in3[0]), .in2(in2[0]), .in1(in1[0]),
     .in0(in0[0]));
tiehi I10 ( .tiehi(tiehi));
bram_4k_inmux7_4 I6 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[15:0]),
     .wl(wl[13:12]), .reset_b(reset_b[13:12]), .prog(progd),
     .pgate(pgate[13:12]), .op(op[6]), .min3({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp12_v_b(sp12_v_b[10]), .sp12_h_r(sp12_h_r[9:8]),
     .sp4_v_b(sp4_v_b[20:18]), .sp4_r_v_b(sp4_r_v_b[20:18]),
     .sp4_h_r(sp4_h_r[20:18]), .in3(in3[6]), .in2(in2[6]),
     .in1(in1[6]), .in0(in0[6]));
bram_4k_inmux7_4 I5 ( .vdd_cntl(vdd_cntl[11:10]), .bl(bl[15:0]),
     .wl(wl[11:10]), .reset_b(reset_b[11:10]), .prog(progd),
     .pgate(pgate[11:10]), .op(op[5]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[9]), .sp12_h_r(sp12_h_r[7:6]),
     .sp4_v_b(sp4_v_b[17:15]), .sp4_r_v_b(sp4_r_v_b[17:15]),
     .sp4_h_r(sp4_h_r[17:15]), .in3(in3[5]), .in2(in2[5]),
     .in1(in1[5]), .in0(in0[5]));
bram_4k_inmux7_4 I4 ( .vdd_cntl(vdd_cntl[9:8]), .bl(bl[15:0]),
     .wl(wl[9:8]), .reset_b(reset_b[9:8]), .prog(progd),
     .pgate(pgate[9:8]), .op(op[4]), .min3({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .sp12_v_b(sp12_v_b[8]),
     .sp12_h_r(sp12_h_r[5:4]), .sp4_v_b(sp4_v_b[14:12]),
     .sp4_r_v_b(sp4_r_v_b[14:12]), .sp4_h_r(sp4_h_r[14:12]),
     .in3(in3[4]), .in2(in2[4]), .in1(in1[4]), .in0(in0[4]));
bram_4k_inmux7_4 I7 ( .vdd_cntl(vdd_cntl[15:14]), .bl(bl[15:0]),
     .wl(wl[15:14]), .reset_b(reset_b[15:14]), .prog(progd),
     .pgate(pgate[15:14]), .op(op[7]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[11]), .sp12_h_r(sp12_h_r[11:10]),
     .sp4_v_b(sp4_v_b[23:21]), .sp4_r_v_b(sp4_r_v_b[23:21]),
     .sp4_h_r(sp4_h_r[23:21]), .in3(in3[7]), .in2(in2[7]),
     .in1(in1[7]), .in0(in0[7]));
inv_hvt I81 ( .A(prog), .Y(progb));
inv_hvt I82 ( .A(progb), .Y(progd));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbankout, View -
//schematic
// LAST TIME SAVED: Aug 22 17:35:36 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4kprouting_bbankout ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sdi_o;

inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_h_l_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_bot;
inout [23:0]  sp12_h_l_bot;
inout [41:0]  bl;
inout [23:0]  sp12_h_l_top;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_r_top;

input [7:0]  top_op_top;
input [1:0]  bm_sweb_i;
input [7:0]  tnr_op_top;
input [7:0]  lft_op_top;
input [7:0]  tnl_op_bot;
input [7:0]  bnr_op_top;
input [15:0]  pgate_bot;
input [7:0]  glb_netwk;
input [1:0]  bm_sdi_i;
input [15:0]  pgate_top;
input [7:0]  rgt_op_bot;
input [7:0]  bot_op_bot;
input [7:0]  bnl_op_top;
input [15:0]  wl_top;
input [15:0]  vdd_cntl_bot;
input [1:0]  bm_sdo_i;
input [7:0]  bm_sa_i;
input [7:0]  bnl_op_bot;
input [15:0]  vdd_cntl_top;
input [15:0]  reset_b_bot;
input [7:0]  tnl_op_top;
input [7:0]  lft_op_bot;
input [7:0]  bnr_op_bot;
input [15:0]  reset_b_top;
input [7:0]  rgt_op_top;
input [15:0]  wl_bot;
input [7:0]  tnr_op_bot;
input [1:0]  bm_sclkrw_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net341;

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net252;

wire  [0:7]  net286;

wire  [0:7]  net320;

wire  [0:7]  net253;

wire  [0:7]  net283;

wire  [0:7]  net254;

wire  [0:7]  net285;

wire  [0:7]  net251;

wire  [0:7]  net284;



bram_4kbankout_pbuffer_bot I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net266), .bm_wen(net234),
     .bm_d(bm_d[15:0]), .bm_clkr(net287), .bm_clkw(net255),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_ab(net341[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net320[0:7]),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
tielo I14 ( .tielo(net298));
tielo I15 ( .tielo(net299));
bram_routing_tracks4rev I5 ( .vdd_cntl(vdd_cntl_bot[15:0]),
     .s_r(net234), .wl(wl_bot[15:0]), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b(reset_b_bot[15:0]), .prog(prog), .pgate(pgate_bot[15:0]),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net299), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]), .clk(net255),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[41:16]));
bram_routing_tracks4rev I3 ( .vdd_cntl(vdd_cntl_top[15:0]),
     .s_r(net266), .wl(wl_top[15:0]), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b(reset_b_top[15:0]), .prog(prog), .pgate(pgate_top[15:0]),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net298), .bot_op(slf_op_bot[7:0]),
     .bnr_op(bnr_op_top[7:0]), .bnl_op(bnl_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]), .clk(net287),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[41:16]));
bram_4k_inmux_8x4 I6 ( .vdd_cntl(vdd_cntl_bot[15:0]), .bl(bl[15:0]),
     .wl(wl_bot[15:0]), .reset_b(reset_b_bot[15:0]), .prog(prog),
     .pgate(pgate_bot[15:0]), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net320[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl(vdd_cntl_top[15:0]), .bl(bl[15:0]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl(wl_top[15:0]), .reset_b(reset_b_top[15:0]), .prog(prog),
     .pgate(pgate_top[15:0]), .op(slf_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net341[0:7]));

endmodule
// Library - leafcell, Cell - bram_4k_sr, View - schematic
// LAST TIME SAVED: Aug 15 17:41:16 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_sr ( bm_dm, bm_sweb, clk, rcapmux_en, rst, bm_q, bm_sdi,
     wdummymux_en );

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[0]), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));

endmodule
// Library - EH_PUP_2, Cell - eh_core_pup_2, View - schematic
// LAST TIME SAVED: Jul 11 11:51:16 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module eh_core_pup_2 ( por_b );
output  por_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



rppolywo  R10 ( .MINUS(net130), .PLUS(net109));
rppolywo  R12 ( .MINUS(net154), .PLUS(net157));
rppolywo  R6 ( .MINUS(out_1), .PLUS(net124));
rppolywo  R9 ( .MINUS(net118), .PLUS(net130));
rppolywo  R15 ( .MINUS(net166), .PLUS(div_1));
rppolywo  R13 ( .MINUS(net157), .PLUS(net145));
rppolywo  R1 ( .MINUS(net068), .PLUS(net048));
rppolywo  R2 ( .MINUS(net067), .PLUS(net068));
rppolywo  R4 ( .MINUS(net142), .PLUS(net148));
rppolywo  R5 ( .MINUS(div_1), .PLUS(net142));
rppolywo  R41 ( .MINUS(net039), .PLUS(net042));
rppolywo  R40 ( .MINUS(net042), .PLUS(vdd_));
rppolywo  R11 ( .MINUS(net109), .PLUS(net154));
rppolywo  R0 ( .MINUS(net048), .PLUS(net039));
rppolywo  R8 ( .MINUS(net127), .PLUS(net118));
rppolywo  R14 ( .MINUS(net145), .PLUS(net166));
rppolywo  R3 ( .MINUS(net148), .PLUS(net067));
rppolywo  R7 ( .MINUS(net124), .PLUS(net127));
nch_hvt  M0 ( .D(out_1), .B(gnd_), .G(div_1), .S(gnd_));
nch_hvt  M2 ( .D(out_1), .B(gnd_), .G(out_2), .S(gnd_));
nch_hvt  M6 ( .D(gnd_), .B(gnd_), .G(out_2), .S(gnd_));
inv_hvt I11 ( .A(out_4), .Y(net193));
inv_hvt I2 ( .A(out_3), .Y(out_4));
inv_hvt I7 ( .A(out_1), .Y(out_2));
inv_hvt I9 ( .A(out_2), .Y(out_3));
inv_hvt I6 ( .A(net193), .Y(por_b));

endmodule
// Library - leafcell, Cell - bram_4k, View - schematic
// LAST TIME SAVED: Aug 15 17:44:47 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr, bm_clkw,
     bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk, bm_sclkrw,
     bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_sa;
input [7:0]  bm_ab;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [14:0]  bm_dm;



tielo I15 ( .tielo(net101));
tielo I18 ( .tielo(net102));
bram_4k_sr I12 ( .bm_dm({bm_sdo, bm_dm[14:0]}), .rst(net102),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM({bm_sdo, bm_dm[14:0]}), .WEBM(bm_sweb), .WEB(web),
     .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]), .CLKW(net81),
     .CLKR(net79), .BWEBM({net101, net101, net101, net101, net101,
     net101, net101, net101, net101, net101, net101, net101, net101,
     net101, net101, net101}), .BWEB(bm_bweb[15:0]), .BIST(bm_init),
     .AMB(bm_sa[7:0]), .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]),
     .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net97), .out(net79));
bram_bufferx6 I8 ( .in(net93), .out(net81));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net93), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net97), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbank_pbuffer_bot, View -
//schematic
// LAST TIME SAVED: Aug 24 17:32:39 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;

input [15:0]  bm_d;
input [15:0]  bm_bweb;
input [1:0]  bm_sweb_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [1:0]  bm_sclkrw_i;
input [7:0]  bm_sa_i;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbank, View - schematic
// LAST TIME SAVED: Aug 22 17:33:36 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4kprouting_bbank ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;
output [1:0]  bm_sdo_o;

inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_l_top;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_h_r_bot;
inout [23:0]  sp12_h_l_top;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_r_top;

input [7:0]  tnr_op_top;
input [7:0]  tnr_op_bot;
input [7:0]  lft_op_top;
input [7:0]  top_op_top;
input [1:0]  bm_sweb_i;
input [7:0]  rgt_op_top;
input [7:0]  bnr_op_top;
input [15:0]  reset_b_top;
input [15:0]  wl_top;
input [15:0]  pgate_top;
input [7:0]  bot_op_bot;
input [1:0]  bm_sdo_i;
input [7:0]  bnr_op_bot;
input [7:0]  rgt_op_bot;
input [7:0]  glb_netwk;
input [7:0]  tnl_op_bot;
input [1:0]  bm_sdi_i;
input [15:0]  vdd_cntl_bot;
input [7:0]  bnl_op_top;
input [15:0]  reset_b_bot;
input [7:0]  bm_sa_i;
input [7:0]  bnl_op_bot;
input [15:0]  wl_bot;
input [7:0]  lft_op_bot;
input [15:0]  vdd_cntl_top;
input [1:0]  bm_sclkrw_i;
input [7:0]  tnl_op_top;
input [15:0]  pgate_bot;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net341;

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net286;

wire  [0:7]  net320;

wire  [0:7]  net283;

wire  [0:7]  net253;

wire  [0:7]  net254;

wire  [0:7]  net285;

wire  [0:7]  net251;

wire  [0:7]  net284;

wire  [0:7]  net252;



bram_4kbank_pbuffer_bot I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net266), .bm_wen(net234),
     .bm_d(bm_d[15:0]), .bm_clkr(net287), .bm_clkw(net255),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_ab(net341[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net320[0:7]),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
tielo I14 ( .tielo(net298));
tielo I15 ( .tielo(net299));
bram_4k_inmux_8x4 I6 ( .vdd_cntl(vdd_cntl_bot[15:0]), .bl(bl[15:0]),
     .wl(wl_bot[15:0]), .reset_b(reset_b_bot[15:0]), .prog(prog),
     .pgate(pgate_bot[15:0]), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net320[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl(vdd_cntl_top[15:0]), .bl(bl[15:0]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl(wl_top[15:0]), .reset_b(reset_b_top[15:0]), .prog(prog),
     .pgate(pgate_top[15:0]), .op(slf_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net341[0:7]));
bram_routing_tracks4rev I5 ( .vdd_cntl(vdd_cntl_bot[15:0]),
     .s_r(net234), .wl(wl_bot[15:0]), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b(reset_b_bot[15:0]), .prog(prog), .pgate(pgate_bot[15:0]),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net299), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]), .clk(net255),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[41:16]));
bram_routing_tracks4rev I3 ( .vdd_cntl(vdd_cntl_top[15:0]),
     .s_r(net266), .wl(wl_top[15:0]), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b(reset_b_top[15:0]), .prog(prog), .pgate(pgate_top[15:0]),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net298), .bot_op(slf_op_bot[7:0]),
     .bnr_op(bnr_op_top[7:0]), .bnl_op(bnl_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]), .clk(net287),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[41:16]));

endmodule
// Library - leafcell, Cell - bram_4k_sr_bankin, View - schematic
// LAST TIME SAVED: Aug 15 18:05:22 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_sr_bankin ( bm_dm, bm_sweb, clk, rcapmux_en, rst, bm_q,
     bm_sdi, wdummymux_en );

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(net150), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));
ml_mux2_hvt_schematic I20 ( .in1(wdummy_reg), .in0(bm_dm[0]),
     .out(net150), .sel(wdummymux_en));
leafcell_ml_dff_schematic I19 ( .R(rst), .D(bm_sdi), .CLK(clk),
     .QN(net157), .Q(wdummy_reg));

endmodule
// Library - leafcell, Cell - bram_4k_bankin, View - schematic
// LAST TIME SAVED: Aug 15 18:08:05 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4k_bankin ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_ab;
input [7:0]  bm_sa;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [14:0]  bm_dm;



tielo I15 ( .tielo(net102));
tielo I18 ( .tielo(net103));
bram_4k_sr_bankin I12 ( .bm_dm({bm_sdo, bm_dm[14:0]}), .rst(net103),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM({bm_sdo, bm_dm[14:0]}), .WEBM(bm_sweb), .WEB(web),
     .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]), .CLKW(net82),
     .CLKR(net80), .BWEBM({net102, net102, net102, net102, net102,
     net102, net102, net102, net102, net102, net102, net102, net102,
     net102, net102, net102}), .BWEB(bm_bweb[15:0]), .BIST(bm_init),
     .AMB(bm_sa[7:0]), .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]),
     .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net98), .out(net80));
bram_bufferx6 I8 ( .in(net94), .out(net82));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net94), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net98), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbankin_pbuffer_bot, View -
//schematic
// LAST TIME SAVED: Aug 24 17:33:35 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4kbankin_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;

input [7:0]  bm_aa;
input [15:0]  bm_bweb;
input [7:0]  bm_sa_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sclkrw_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [1:0]  bm_sweb_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankin I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbankin, View - schematic
// LAST TIME SAVED: Aug 22 17:34:31 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module bram_4kprouting_bbankin ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;
output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sweb_o;

inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_h_l_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_bot;
inout [23:0]  sp12_h_l_bot;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_v_b_top;

input [15:0]  wl_top;
input [7:0]  tnr_op_top;
input [7:0]  bot_op_bot;
input [7:0]  rgt_op_top;
input [7:0]  rgt_op_bot;
input [1:0]  bm_sdi_i;
input [15:0]  pgate_top;
input [7:0]  tnr_op_bot;
input [1:0]  bm_sdo_i;
input [7:0]  tnl_op_bot;
input [7:0]  bnr_op_top;
input [1:0]  bm_sweb_i;
input [15:0]  pgate_bot;
input [7:0]  top_op_top;
input [7:0]  lft_op_top;
input [15:0]  reset_b_top;
input [7:0]  bnl_op_top;
input [7:0]  bm_sa_i;
input [15:0]  vdd_cntl_top;
input [15:0]  reset_b_bot;
input [7:0]  lft_op_bot;
input [7:0]  bnr_op_bot;
input [7:0]  bnl_op_bot;
input [15:0]  vdd_cntl_bot;
input [15:0]  wl_bot;
input [7:0]  tnl_op_top;
input [1:0]  bm_sclkrw_i;
input [7:0]  glb_netwk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net341;

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net251;

wire  [0:7]  net283;

wire  [0:7]  net254;

wire  [0:7]  net285;

wire  [0:7]  net284;

wire  [0:7]  net320;

wire  [0:7]  net286;

wire  [0:7]  net253;

wire  [0:7]  net252;



bram_4kbankin_pbuffer_bot I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net266), .bm_wen(net234),
     .bm_d(bm_d[15:0]), .bm_clkr(net287), .bm_clkw(net255),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_ab(net341[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net320[0:7]),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl(vdd_cntl_bot[15:0]), .bl(bl[15:0]),
     .wl(wl_bot[15:0]), .reset_b(reset_b_bot[15:0]), .prog(prog),
     .pgate(pgate_bot[15:0]), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net320[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl(vdd_cntl_top[15:0]), .bl(bl[15:0]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl(wl_top[15:0]), .reset_b(reset_b_top[15:0]), .prog(prog),
     .pgate(pgate_top[15:0]), .op(slf_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net341[0:7]));
tielo I14 ( .tielo(net298));
tielo I15 ( .tielo(net299));
bram_routing_tracks4rev I5 ( .vdd_cntl(vdd_cntl_bot[15:0]),
     .s_r(net234), .wl(wl_bot[15:0]), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b(reset_b_bot[15:0]), .prog(prog), .pgate(pgate_bot[15:0]),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net299), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]), .clk(net255),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[41:16]));
bram_routing_tracks4rev I3 ( .vdd_cntl(vdd_cntl_top[15:0]),
     .s_r(net266), .wl(wl_top[15:0]), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b(reset_b_top[15:0]), .prog(prog), .pgate(pgate_top[15:0]),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net298), .bot_op(slf_op_bot[7:0]),
     .bnr_op(bnr_op_top[7:0]), .bnl_op(bnl_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]), .clk(net287),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[41:16]));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev0, View - schematic
// LAST TIME SAVED: Jun  2 13:19:45 2008
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module clkmandcmuxrev0 ( clk, clkb, glb2local, s_r, cbit, cbitb,
     glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, min0, min1,
     min2, min3, prog );
output  clk, clkb, s_r;

input  prog;

output [3:0]  glb2local;

input [7:0]  min3;
input [7:0]  min1;
input [7:0]  min0;
input [7:0]  min2;
input [31:0]  cbitb;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g0;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g3;
input [31:0]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sr_clkm8to1 I296 ( .mout(s_r), .cbitb(cbitb[12:9]), .min({lc_trk_g3[5],
     lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4], glb_netwk[6],
     glb_netwk[4], glb_netwk[2], glb_netwk[0]}), .cbit(cbit[12:9]),
     .prog(prog));
ce_clkm8to1 I283 ( .moutb(ceb), .cbitb(cbitb[8:5]), .cbit(cbit[8:5]),
     .prog(prog), .min({lc_trk_g3[3], lc_trk_g2[2], lc_trk_g1[3],
     lc_trk_g0[2], glb_netwk[7], glb_netwk[5], glb_netwk[3],
     glb_netwk[1]}));
clk_mux12to1 I298 ( .cbitb({cbitb[31], cbitb[4], cbitb[3], cbitb[2],
     cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3], cbit[2],
     cbit[1], cbit[0]}), .prog(prog), .min({lc_trk_g3[1], lc_trk_g2[0],
     lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}), .clk(clk),
     .clkb(clkb), .cenb(ceb));
clk_mux8to1 I285 ( .min(min3[7:0]), .prog(prog), .inmuxo(glb2local[0]),
     .cbit(cbit[16:13]), .cbitb(cbitb[16:13]));
clk_mux8to1 I293 ( .prog(prog), .inmuxo(glb2local[1]), .min(min2[7:0]),
     .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I294 ( .prog(prog), .inmuxo(glb2local[2]), .min(min1[7:0]),
     .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
clk_mux8to1 I295 ( .prog(prog), .inmuxo(glb2local[3]), .min(min0[7:0]),
     .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));

endmodule
// Library - leafcell, Cell - misc_module4rev2, View - schematic
// LAST TIME SAVED: Oct 10 17:39:26 2008
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module misc_module4rev2 ( S_R, cbit, cbitb, clk, clkb, glb2local, sp4,
     bl, b, glb_netwk, l, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3,
     m, min0, min1, min2, min3, pgate, prog, r, reset_b, sp12,
     vdd_cntl, wl );
output  S_R, clk, clkb;


input  prog;

output [3:0]  glb2local;
output [7:0]  sp4;
output [63:0]  cbit;
output [63:0]  cbitb;

inout [3:0]  bl;

input [7:0]  min3;
input [1:0]  b;
input [15:0]  pgate;
input [5:0]  lc_trk_g0;
input [5:0]  lc_trk_g1;
input [7:0]  glb_netwk;
input [7:0]  sp12;
input [15:0]  wl;
input [5:0]  lc_trk_g2;
input [15:0]  vdd_cntl;
input [1:0]  r;
input [7:0]  min0;
input [7:0]  min1;
input [15:0]  reset_b;
input [5:0]  lc_trk_g3;
input [7:0]  min2;
input [1:0]  l;
input [1:0]  m;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  r_vdd;



clkmandcmuxrev0 Itclkm ( .min2(min2[7:0]), .min1(min1[7:0]),
     .min0(min0[7:0]), .min3(min3[7:0]), .cbit({cbit[2], cbit[1],
     cbit[0], cbit[27], cbit[25], cbit[26], cbit[24], cbit[23],
     cbit[21], cbit[22], cbit[20], cbit[19], cbit[17], cbit[18],
     cbit[16], cbit[15], cbit[13], cbit[14], cbit[12], cbit[31],
     cbit[29], cbit[30], cbit[28], cbit[11], cbit[9], cbit[10],
     cbit[8], cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}), .glb2local(glb2local[3:0]),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .glb_netwk(glb_netwk[7:0]), .prog(prog), .clk(clk), .clkb(clkb),
     .s_r(S_R));
pch_hvt  vdd_cntrl_15_ ( .D(r_vdd[15]), .B(vdd_), .G(vdd_cntl[15]),
     .S(vdd_));
pch_hvt  vdd_cntrl_14_ ( .D(r_vdd[14]), .B(vdd_), .G(vdd_cntl[14]),
     .S(vdd_));
pch_hvt  vdd_cntrl_13_ ( .D(r_vdd[13]), .B(vdd_), .G(vdd_cntl[13]),
     .S(vdd_));
pch_hvt  vdd_cntrl_12_ ( .D(r_vdd[12]), .B(vdd_), .G(vdd_cntl[12]),
     .S(vdd_));
pch_hvt  vdd_cntrl_11_ ( .D(r_vdd[11]), .B(vdd_), .G(vdd_cntl[11]),
     .S(vdd_));
pch_hvt  vdd_cntrl_10_ ( .D(r_vdd[10]), .B(vdd_), .G(vdd_cntl[10]),
     .S(vdd_));
pch_hvt  vdd_cntrl_9_ ( .D(r_vdd[9]), .B(vdd_), .G(vdd_cntl[9]),
     .S(vdd_));
pch_hvt  vdd_cntrl_8_ ( .D(r_vdd[8]), .B(vdd_), .G(vdd_cntl[8]),
     .S(vdd_));
pch_hvt  vdd_cntrl_7_ ( .D(r_vdd[7]), .B(vdd_), .G(vdd_cntl[7]),
     .S(vdd_));
pch_hvt  vdd_cntrl_6_ ( .D(r_vdd[6]), .B(vdd_), .G(vdd_cntl[6]),
     .S(vdd_));
pch_hvt  vdd_cntrl_5_ ( .D(r_vdd[5]), .B(vdd_), .G(vdd_cntl[5]),
     .S(vdd_));
pch_hvt  vdd_cntrl_4_ ( .D(r_vdd[4]), .B(vdd_), .G(vdd_cntl[4]),
     .S(vdd_));
pch_hvt  vdd_cntrl_3_ ( .D(r_vdd[3]), .B(vdd_), .G(vdd_cntl[3]),
     .S(vdd_));
pch_hvt  vdd_cntrl_2_ ( .D(r_vdd[2]), .B(vdd_), .G(vdd_cntl[2]),
     .S(vdd_));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sp12to4 Isp12to4_7_ ( .triout(sp4[7]), .cbitb(cbitb[62]),
     .drv(sp12[7]), .prog(net109));
sp12to4 Isp12to4_6_ ( .triout(sp4[6]), .cbitb(cbitb[58]),
     .drv(sp12[6]), .prog(net109));
sp12to4 Isp12to4_5_ ( .triout(sp4[5]), .cbitb(cbitb[54]),
     .drv(sp12[5]), .prog(net109));
sp12to4 Isp12to4_4_ ( .triout(sp4[4]), .cbitb(cbitb[50]),
     .drv(sp12[4]), .prog(net109));
sp12to4 Isp12to4_3_ ( .triout(sp4[3]), .cbitb(cbitb[46]),
     .drv(sp12[3]), .prog(net109));
sp12to4 Isp12to4_2_ ( .triout(sp4[2]), .cbitb(cbitb[42]),
     .drv(sp12[2]), .prog(net109));
sp12to4 Isp12to4_1_ ( .triout(sp4[1]), .cbitb(cbitb[5]), .drv(sp12[1]),
     .prog(net109));
sp12to4 Isp12to4_0_ ( .triout(sp4[0]), .cbitb(cbitb[34]),
     .drv(sp12[0]), .prog(net109));
sbox1 Isp12_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(prog));
sbox1 Isp12_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(prog));
cram16x4 Ic64 ( .r_gnd(r_vdd[15:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .q(cbit[63:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net109));

endmodule
// Library - leafcell, Cell - logic_cell, View - schematic
// LAST TIME SAVED: Aug 28 17:23:08 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module logic_cell ( carry_out, out, carry_in, cbit, clk, clkb, in0,
     in1, in2, in3, prog, purst, s_r );
output  carry_out, out;

input  carry_in, clk, clkb, in0, in1, in2, in3, prog, purst, s_r;

input [20:0]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



coredffr REG ( .purst(purst), .d(LUT4_outd), .q(rego),
     .cbit(cbit[17:16]), .clkb(clkb), .clk(clk), .S_R(s_r));
carry_logic ICARRY_LOGIC ( .b_bar(in1b1), .carry_in(carry_in), .b(in1),
     .cout(carry_out), .a(in2), .a_bar(in2b1), .vg_en(cbit[20]));
o_mux Iomux ( .in1(rego), .out(out), .cbit(cbit[19]), .prog(prog),
     .in0(LUT4_outd));
clut4 iclut4 ( .in0b(in0b1), .in3b(in3b1), .in2b(in2b1),
     .lut4(LUT4_outd), .in1b(in1b1), .in2(in2), .in1(in1), .in0(in0),
     .in3(in3), .cbit(cbit[15:0]));
inv_hvt I163 ( .A(in3), .Y(in3b1));
inv_hvt I164 ( .A(in1), .Y(in1b1));
inv_hvt I162 ( .A(in2), .Y(in2b1));
inv_hvt I161 ( .A(in0), .Y(in0b1));

endmodule
// Library - EH_PUP_2, Cell - SMC_CORE_POR_right, View - schematic
// LAST TIME SAVED: Oct  6 14:23:47 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module SMC_CORE_POR_right ( core_por_b, smc_por_b,
     smc_core_por_bottom1, smc_core_por_bottom2, vddio_rightbank );
output  core_por_b, smc_por_b;

input  smc_core_por_bottom1, smc_core_por_bottom2, vddio_rightbank;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



eh_io_pup_2_new I0 ( .vdd_io(vddio_rightbank), .core_por_b(core_por_b),
     .por_b(net3));
nand4_hvt I2 ( .D(core_por_b), .C(smc_core_por_bottom2), .A(net3),
     .Y(net04), .B(smc_core_por_bottom1));
inv_hvt I3 ( .A(net04), .Y(smc_por_b));
eh_core_pup_2 I1 ( .por_b(core_por_b));

endmodule
// Library - xpmem, Cell - cram_2x28, View - schematic
// LAST TIME SAVED: Jul 28 08:32:33 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module cram_2x28 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [55:0]  q;
output [55:0]  q_b;

inout [27:0]  bl;

input [1:0]  wl;
input [1:0]  reset;
input [1:0]  r_vdd;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_13_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[27:26]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[1:0]));
cram2x2 Imstake_12_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[25:24]), .q_b(q_b[51:48]),
     .q(q[51:48]), .wl(wl[1:0]));
cram2x2 Imstake_11_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[23:22]), .q_b(q_b[47:44]),
     .q(q[47:44]), .wl(wl[1:0]));
cram2x2 Imstake_10_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[21:20]), .q_b(q_b[43:40]),
     .q(q[43:40]), .wl(wl[1:0]));
cram2x2 Imstake_9_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[19:18]), .q_b(q_b[39:36]),
     .q(q[39:36]), .wl(wl[1:0]));
cram2x2 Imstake_8_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[17:16]), .q_b(q_b[35:32]),
     .q(q[35:32]), .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[15:14]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[1:0]));
cram2x2 Imstake_6_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[13:12]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[1:0]));
cram2x2 Imstake_5_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - lcmuxod3_0, View - schematic
// LAST TIME SAVED: Aug 21 17:57:09 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module lcmuxod3_0 ( carry_out, op, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_h_r;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min2;
input [1:0]  wl;
input [15:0]  min3;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [27:0]  bl;
input [1:0]  pgate;
input [15:0]  min1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
odrv12_30 Iodrv30 ( .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - lcmuxod7_4, View - schematic
// LAST TIME SAVED: Aug 21 17:56:42 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module lcmuxod7_4 ( carry_out, op, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_v_b;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [1:0]  sp12_h_r;
output [2:0]  sp4_v_b;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [15:0]  min2;
input [1:0]  reset_b;
input [15:0]  min3;
input [15:0]  min0;
input [27:0]  bl;
input [15:0]  min1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
odrv12_74 Iodrv74 ( .cbitb({cbitb[53], cbitb[55], cbitb[52], cbitb[54],
     cbitb[51], cbitb[49], cbitb[44], cbitb[46], cbitb[43], cbitb[41],
     cbitb[42], cbitb[40]}), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]),
     .sp12_v_b(sp12_v_b), .sp12_h_r(sp12_h_r[1:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - lccol_rev2, View - schematic
// LAST TIME SAVED: Oct 10 17:34:46 2008
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module lccol_rev2 ( carry_out, slf_op, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, cbit_c, cbitb_c, cin2local, clk, clkb,
     lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, pgate, prog, purst,
     reset_b, s_r, vdd_cntl, wl );
output  carry_out;


input  cin2local, clk, clkb, prog, purst, s_r;

output [7:0]  slf_op;

inout [27:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;

input [15:0]  vdd_cntl;
input [1:0]  cbitb_c;
input [15:0]  reset_b;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g2;
input [7:0]  lc_trk_g3;
input [1:0]  cbit_c;
input [15:0]  pgate;
input [15:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



mux_4carry Icarry_cnt ( .cin(cin2local), .lcl_cin(cin),
     .cbitb(cbitb_c[1:0]), .prog(prog), .cbit(cbit_c[1:0]));
lcmuxod3_0 ILC_02 ( .vdd_cntl(vdd_cntl[5:4]), .purst(purst),
     .pgate(pgate[5:4]), .sp4_r_v_b({sp4_r_v_b[37], sp4_r_v_b[21],
     sp4_r_v_b[5]}), .sp12_h_r(sp12_h_r[12]), .sp12_v_b({sp12_v_b[20],
     sp12_v_b[4]}), .sp4_h_r({sp4_h_r[36], sp4_h_r[20], sp4_h_r[4]}),
     .sp4_v_b({sp4_v_b[36], sp4_v_b[20], sp4_v_b[4]}), .clk(clk),
     .carry_in(c_12), .op(slf_op[2]), .carry_out(c_23), .s_r(s_r),
     .reset_b(reset_b[5:4]), .bl(bl[27:0]), .wl(wl[5:4]),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_12}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}));
lcmuxod3_0 ILC_00 ( .vdd_cntl(vdd_cntl[1:0]), .purst(purst),
     .pgate(pgate[1:0]), .sp4_r_v_b({sp4_r_v_b[33], sp4_r_v_b[17],
     sp4_r_v_b[1]}), .sp12_h_r(sp12_h_r[8]), .sp12_v_b({sp12_v_b[16],
     sp12_v_b[0]}), .sp4_h_r({sp4_h_r[32], sp4_h_r[16], sp4_h_r[0]}),
     .sp4_v_b({sp4_v_b[32], sp4_v_b[16], sp4_v_b[0]}), .clk(clk),
     .carry_in(cin), .op(slf_op[0]), .carry_out(c_01), .s_r(s_r),
     .reset_b(reset_b[1:0]), .bl(bl[27:0]), .wl(wl[1:0]),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], cin}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}));
lcmuxod3_0 ILC_03 ( .vdd_cntl(vdd_cntl[7:6]), .purst(purst),
     .pgate(pgate[7:6]), .sp4_r_v_b({sp4_r_v_b[39], sp4_r_v_b[23],
     sp4_r_v_b[7]}), .sp12_h_r(sp12_h_r[14]), .sp12_v_b({sp12_v_b[22],
     sp12_v_b[6]}), .sp4_h_r({sp4_h_r[38], sp4_h_r[22], sp4_h_r[6]}),
     .sp4_v_b({sp4_v_b[38], sp4_v_b[22], sp4_v_b[6]}), .clk(clk),
     .carry_in(c_23), .op(slf_op[3]), .carry_out(c_34), .s_r(s_r),
     .reset_b(reset_b[7:6]), .bl(bl[27:0]), .wl(wl[7:6]),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_23}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}));
lcmuxod3_0 ILC_01 ( .vdd_cntl(vdd_cntl[3:2]), .purst(purst),
     .pgate(pgate[3:2]), .sp4_r_v_b({sp4_r_v_b[35], sp4_r_v_b[19],
     sp4_r_v_b[3]}), .sp12_h_r(sp12_h_r[10]), .sp12_v_b({sp12_v_b[18],
     sp12_v_b[2]}), .sp4_h_r({sp4_h_r[34], sp4_h_r[18], sp4_h_r[2]}),
     .sp4_v_b({sp4_v_b[34], sp4_v_b[18], sp4_v_b[2]}), .clk(clk),
     .carry_in(c_01), .op(slf_op[1]), .carry_out(c_12), .s_r(s_r),
     .reset_b(reset_b[3:2]), .bl(bl[27:0]), .wl(wl[3:2]),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_01}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}));
lcmuxod7_4 ILC_07 ( .vdd_cntl(vdd_cntl[15:14]), .purst(purst),
     .pgate(pgate[15:14]), .sp4_r_v_b({sp4_r_v_b[47], sp4_r_v_b[31],
     sp4_r_v_b[15]}), .sp12_h_r({sp12_h_r[22], sp12_h_r[6]}),
     .sp12_v_b(sp12_v_b[14]), .sp4_h_r({sp4_h_r[46], sp4_h_r[30],
     sp4_h_r[14]}), .sp4_v_b({sp4_v_b[46], sp4_v_b[30], sp4_v_b[14]}),
     .clk(clk), .carry_in(c_67), .op(slf_op[7]), .carry_out(carry_out),
     .s_r(s_r), .reset_b(reset_b[15:14]), .bl(bl[27:0]),
     .wl(wl[15:14]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_67}),
     .prog(prog), .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}));
lcmuxod7_4 ILC_06 ( .vdd_cntl(vdd_cntl[13:12]), .purst(purst),
     .pgate(pgate[13:12]), .sp4_r_v_b({sp4_r_v_b[45], sp4_r_v_b[29],
     sp4_r_v_b[13]}), .sp12_h_r({sp12_h_r[20], sp12_h_r[4]}),
     .sp12_v_b(sp12_v_b[12]), .sp4_h_r({sp4_h_r[44], sp4_h_r[28],
     sp4_h_r[12]}), .sp4_v_b({sp4_v_b[44], sp4_v_b[28], sp4_v_b[12]}),
     .clk(clk), .carry_in(c_56), .op(slf_op[6]), .carry_out(c_67),
     .s_r(s_r), .reset_b(reset_b[13:12]), .bl(bl[27:0]),
     .wl(wl[13:12]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_56}),
     .prog(prog), .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}));
lcmuxod7_4 ILC_04 ( .vdd_cntl(vdd_cntl[9:8]), .purst(purst),
     .pgate(pgate[9:8]), .sp4_r_v_b({sp4_r_v_b[41], sp4_r_v_b[25],
     sp4_r_v_b[9]}), .sp12_h_r({sp12_h_r[16], sp12_h_r[0]}),
     .sp12_v_b(sp12_v_b[8]), .sp4_h_r({sp4_h_r[40], sp4_h_r[24],
     sp4_h_r[8]}), .sp4_v_b({sp4_v_b[40], sp4_v_b[24], sp4_v_b[8]}),
     .clk(clk), .carry_in(c_34), .op(slf_op[4]), .carry_out(c_45),
     .s_r(s_r), .reset_b(reset_b[9:8]), .bl(bl[27:0]), .wl(wl[9:8]),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_34}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}));
lcmuxod7_4 ILC_05 ( .vdd_cntl(vdd_cntl[11:10]), .purst(purst),
     .pgate(pgate[11:10]), .sp4_r_v_b({sp4_r_v_b[43], sp4_r_v_b[27],
     sp4_r_v_b[11]}), .sp12_h_r({sp12_h_r[18], sp12_h_r[2]}),
     .sp12_v_b(sp12_v_b[10]), .sp4_h_r({sp4_h_r[42], sp4_h_r[26],
     sp4_h_r[10]}), .sp4_v_b({sp4_v_b[42], sp4_v_b[26], sp4_v_b[10]}),
     .clk(clk), .carry_in(c_45), .op(slf_op[5]), .carry_out(c_56),
     .s_r(s_r), .reset_b(reset_b[11:10]), .bl(bl[27:0]),
     .wl(wl[11:10]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_45}),
     .prog(prog), .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}));

endmodule
// Library - leafcell, Cell - ltile4rev, View - schematic
// LAST TIME SAVED: Oct 10 17:40:03 2008
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module ltile4rev ( carry_out, slf_op, bl, sp4_h_l, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r, sp12_v_b, sp12_v_t, bnl_op,
     bnr_op, bot_op, carry_in, glb_netwk, lft_op, pgate, prog, purst,
     reset_b, rgt_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );
output  carry_out;


input  carry_in, prog, purst;

output [7:0]  slf_op;

inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_t;
inout [23:0]  sp12_h_r;
inout [23:0]  sp12_v_t;
inout [53:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_h_l;

input [7:0]  top_op;
input [7:0]  glb_netwk;
input [7:0]  bnl_op;
input [7:0]  rgt_op;
input [7:0]  bot_op;
input [15:0]  wl;
input [7:0]  lft_op;
input [7:0]  bnr_op;
input [15:0]  reset_b;
input [15:0]  pgate;
input [7:0]  tnr_op;
input [15:0]  vdd_cntl;
input [7:0]  tnl_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  lc_trk_g0;

wire  [63:0]  cbit_c;

wire  [3:0]  net_glb2local;

wire  [7:0]  lc_trk_g1;

wire  [1:0]  sp12_h_r_mid;

wire  [63:0]  cbitb_c;

wire  [7:0]  lc_trk_g2;

wire  [7:0]  lc_trk_g3;

wire  [1:0]  sp12_v_b_mid;



misc_module4rev2 Ickmux_sp12to4_sp12sw ( .cbitb(cbitb_c[63:0]),
     .cbit(cbit_c[63:0]), .vdd_cntl(vdd_cntl[15:0]),
     .glb_netwk(glb_netwk[7:0]), .l(sp12_h_r_mid[1:0]),
     .m(sp12_v_b_mid[1:0]), .r(sp12_h_r[1:0]), .b(sp12_v_b[1:0]),
     .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18], sp12_h_r[16],
     sp12_h_r[14], sp12_h_r[12], sp12_h_r[10], sp12_h_r[8]}),
     .sp4(sp4_h_r[23:16]), .min3(glb_netwk[7:0]),
     .min0(glb_netwk[7:0]), .min1(glb_netwk[7:0]),
     .min2(glb_netwk[7:0]), .prog(progd), .lc_trk_g0(lc_trk_g0[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .lc_trk_g1(lc_trk_g1[5:0]), .wl(wl[15:0]), .S_R(net178),
     .clkb(clkb), .bl(bl[53:50]), .clk(clk), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .glb2local(net_glb2local[3:0]));
lccol_rev2 I_lcx8 ( .cbit_c(cbit_c[1:0]), .cbitb_c(cbitb_c[1:0]),
     .vdd_cntl(vdd_cntl[15:0]), .wl(wl[15:0]), .s_r(net178),
     .reset_b(reset_b[15:0]), .purst(purst), .prog(progd),
     .pgate(pgate[15:0]), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .clkb(clkb), .clk(clk),
     .cin2local(carry_in), .slf_op(slf_op[7:0]), .carry_out(carry_out),
     .sp12_v_b(sp12_v_b[23:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .bl(bl[27:0]));
rm6  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm6  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm6  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm6  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm6  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm6  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm6  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm6  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm6  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm6  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm6  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm6  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm6  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm6  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm6  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm6  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm6  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm6  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm6  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm6  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm6  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm6  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm6  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm6  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
rm7  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
span4 Isp4_sw ( .vdd_cntl(vdd_cntl[15:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_l(sp4_h_l[47:0]),
     .sp4_v_t(sp4_v_t[47:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .prog(progd), .wl(wl[15:0]), .bl(bl[49:40]));
gmux_sp12to4 Igmux_sp12to4 ( .vdd_cntl(vdd_cntl[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]),
     .glb2local(net_glb2local[3:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .lc_trk_g1(lc_trk_g1[7:0]), .lc_trk_g2(lc_trk_g2[7:0]),
     .lc_trk_g3(lc_trk_g3[7:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .bot_op(bot_op[7:0]), .wl(wl[15:0]), .top_op(top_op[7:0]),
     .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]), .slf_op(slf_op[7:0]),
     .rgt_op(rgt_op[7:0]), .prog(progd), .lft_op(lft_op[7:0]),
     .bnr_op(bnr_op[7:0]), .bnl_op(bnl_op[7:0]), .bl(bl[39:28]));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(progd));

endmodule
// Library - leafcell, Cell - clk_colbuf, View - schematic
// LAST TIME SAVED: Jul  5 14:43:37 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module clk_colbuf ( clko, clki );
output  clko;

input  clki;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv I19 ( .A(clkb), .Y(clko));
inv I22 ( .A(clki), .Y(clkb));

endmodule
// Library - leafcell, Cell - clk_colbufx8, View - schematic
// LAST TIME SAVED: Jul  5 15:04:30 2007
// NETLIST TIME: Nov 14 16:12:02 2008
`timescale 1ns / 1ns 

module clk_colbufx8 ( clko, clki );


output [7:0]  clko;

input [7:0]  clki;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



clk_colbuf iclk_colbuf_7_ ( .clki(clki[7]), .clko(clko[7]));
clk_colbuf iclk_colbuf_6_ ( .clki(clki[6]), .clko(clko[6]));
clk_colbuf iclk_colbuf_5_ ( .clki(clki[5]), .clko(clko[5]));
clk_colbuf iclk_colbuf_4_ ( .clki(clki[4]), .clko(clko[4]));
clk_colbuf iclk_colbuf_3_ ( .clki(clki[3]), .clko(clko[3]));
clk_colbuf iclk_colbuf_2_ ( .clki(clki[2]), .clko(clko[2]));
clk_colbuf iclk_colbuf_1_ ( .clki(clki[1]), .clko(clko[1]));
clk_colbuf iclk_colbuf_0_ ( .clki(clki[0]), .clko(clko[0]));

endmodule
// Library - leafcell, Cell - QUAD_BR, View - schematic
// LAST TIME SAVED: Sep 15 14:22:41 2008
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module QUAD_BR ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_13_10, carry_out_14_10,
     carry_out_15_10, carry_out_16_10, carry_out_17_10,
     carry_out_18_10, carry_out_20_10, carry_out_21_10,
     carry_out_22_10, carry_out_23_10, carry_out_24_10, ceb_o, cf_b,
     cf_r, fabric_out_94, fabric_out_98, fabric_out_122,
     fabric_out_126, fabric_out_136, fabric_out_162, hiz_b_o, mode_o,
     padeb_b, padeb_r, padin_94, padin_162, pado_b, pado_r, r_o, sdo,
     sdo_pad, shift_o, slf_op_13_00, slf_op_13_01, slf_op_13_02,
     slf_op_13_03, slf_op_13_04, slf_op_13_05, slf_op_13_06,
     slf_op_13_07, slf_op_13_08, slf_op_13_09, slf_op_13_10,
     slf_op_14_10, slf_op_15_10, slf_op_16_10, slf_op_17_10,
     slf_op_18_10, slf_op_19_10, slf_op_20_10, slf_op_21_10,
     slf_op_22_10, slf_op_23_10, slf_op_24_10, slf_op_25_10,
     spi_ss_in_b, spi_ss_in_r, tclk_o, update_o, bl, pgate, reset_b,
     sp4_h_l_13_00, sp4_h_l_13_01, sp4_h_l_13_02, sp4_h_l_13_03,
     sp4_h_l_13_04, sp4_h_l_13_05, sp4_h_l_13_06, sp4_h_l_13_07,
     sp4_h_l_13_08, sp4_h_l_13_09, sp4_h_l_13_10, sp4_v_b_13_01,
     sp4_v_b_13_02, sp4_v_b_13_03, sp4_v_b_13_04, sp4_v_b_13_05,
     sp4_v_b_13_06, sp4_v_b_13_07, sp4_v_b_13_08, sp4_v_b_13_09,
     sp4_v_b_13_10, sp4_v_t_13_10, sp4_v_t_14_10, sp4_v_t_15_10,
     sp4_v_t_16_10, sp4_v_t_17_10, sp4_v_t_18_10, sp4_v_t_19_10,
     sp4_v_t_20_10, sp4_v_t_21_10, sp4_v_t_22_10, sp4_v_t_23_10,
     sp4_v_t_24_10, sp4_v_t_25_10, sp12_h_l_13_01, sp12_h_l_13_02,
     sp12_h_l_13_03, sp12_h_l_13_04, sp12_h_l_13_05, sp12_h_l_13_06,
     sp12_h_l_13_07, sp12_h_l_13_08, sp12_h_l_13_09, sp12_h_l_13_10,
     sp12_v_t_13_10, sp12_v_t_14_10, sp12_v_t_15_10, sp12_v_t_16_10,
     sp12_v_t_17_10, sp12_v_t_18_10, sp12_v_t_19_10, sp12_v_t_20_10,
     sp12_v_t_21_10, sp12_v_t_22_10, sp12_v_t_23_10, sp12_v_t_24_10,
     vdd_cntl, wl, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_13_01, bs_en_i, bs_en_mi,
     cdone_in_bot_r, cdone_in_rgt_b, ceb_i, ceb_mi, glb_in, hiz_b_i,
     hiz_b_mi, hold_b_r, hold_r_b, lft_op_13_01, lft_op_13_02,
     lft_op_13_03, lft_op_13_04, lft_op_13_05, lft_op_13_06,
     lft_op_13_07, lft_op_13_08, lft_op_13_09, lft_op_13_10, mode_i,
     mode_mi, padin_b, padin_r, prog, purst, r_i, r_mi, sdi, sdi_pad,
     shift_i, shift_mi, spioeb_b, spioeb_r, spiout_b, spiout_r, tclk_i,
     tclk_mi, tiegnd, tnl_op_13_10, tnl_op_14_10, tnl_op_15_10,
     tnl_op_16_10, tnl_op_17_10, tnl_op_18_10, tnl_op_19_10,
     tnl_op_20_10, tnl_op_21_10, tnl_op_22_10, tnl_op_23_10,
     tnl_op_24_10, tnl_op_25_10, tnr_op_13_10, tnr_op_14_10,
     tnr_op_15_10, tnr_op_16_10, tnr_op_17_10, tnr_op_18_10,
     tnr_op_19_10, tnr_op_20_10, tnr_op_21_10, tnr_op_22_10,
     tnr_op_23_10, tnr_op_24_10, top_op_13_10, top_op_14_10,
     top_op_15_10, top_op_16_10, top_op_17_10, top_op_18_10,
     top_op_19_10, top_op_20_10, top_op_21_10, top_op_22_10,
     top_op_23_10, top_op_24_10, update_i, update_mi );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_13_10, carry_out_14_10,
     carry_out_15_10, carry_out_16_10, carry_out_17_10,
     carry_out_18_10, carry_out_20_10, carry_out_21_10,
     carry_out_22_10, carry_out_23_10, carry_out_24_10, ceb_o,
     fabric_out_94, fabric_out_98, fabric_out_122, fabric_out_126,
     fabric_out_136, fabric_out_162, hiz_b_o, mode_o, padin_94,
     padin_162, r_o, sdo, sdo_pad, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, bs_en_mi, ceb_i, ceb_mi, hiz_b_i,
     hiz_b_mi, hold_b_r, hold_r_b, mode_i, mode_mi, prog, purst, r_i,
     r_mi, sdi, sdi_pad, shift_i, shift_mi, tclk_i, tclk_mi, tiegnd,
     update_i, update_mi;

output [1:0]  bm_sdo_o;
output [7:0]  slf_op_13_06;
output [7:0]  slf_op_23_10;
output [7:0]  slf_op_21_10;
output [7:0]  slf_op_14_10;
output [7:0]  slf_op_13_07;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_17_10;
output [3:0]  slf_op_25_10;
output [7:0]  slf_op_24_10;
output [7:0]  slf_op_16_10;
output [19:0]  padeb_r;
output [7:0]  slf_op_19_10;
output [7:0]  slf_op_13_10;
output [1:0]  bm_sweb_o;
output [575:288]  cf_b;
output [47:24]  padeb_b;
output [47:24]  spi_ss_in_b;
output [7:0]  slf_op_13_01;
output [7:0]  slf_op_20_10;
output [1:0]  bm_sdi_o;
output [19:0]  spi_ss_in_r;
output [7:0]  slf_op_15_10;
output [7:0]  slf_op_13_04;
output [239:0]  cf_r;
output [7:0]  slf_op_13_05;
output [3:0]  slf_op_13_00;
output [7:0]  slf_op_13_09;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_13_03;
output [7:0]  slf_op_22_10;
output [19:0]  pado_r;
output [47:24]  pado_b;
output [7:0]  slf_op_13_08;
output [7:0]  slf_op_18_10;
output [7:0]  slf_op_13_02;

inout [47:0]  sp4_v_t_18_10;
inout [23:0]  sp12_h_l_13_07;
inout [23:0]  sp12_h_l_13_04;
inout [23:0]  sp12_v_t_13_10;
inout [23:0]  sp12_h_l_13_01;
inout [47:0]  sp4_v_t_24_10;
inout [47:0]  sp4_h_l_13_02;
inout [23:0]  sp12_v_t_15_10;
inout [47:0]  sp4_v_b_13_03;
inout [47:0]  sp4_v_t_15_10;
inout [47:0]  sp4_v_t_19_10;
inout [47:0]  sp4_v_b_13_09;
inout [47:0]  sp4_v_t_16_10;
inout [47:0]  sp4_h_l_13_03;
inout [23:0]  sp12_v_t_14_10;
inout [23:0]  sp12_v_t_21_10;
inout [47:0]  sp4_h_l_13_05;
inout [23:0]  sp12_h_l_13_08;
inout [47:0]  sp4_v_b_13_10;
inout [47:0]  sp4_h_l_13_09;
inout [47:0]  sp4_v_t_23_10;
inout [47:0]  sp4_h_l_13_04;
inout [175:0]  pgate;
inout [47:0]  sp4_v_t_20_10;
inout [1311:658]  bl;
inout [15:0]  sp4_h_l_13_00;
inout [47:0]  sp4_v_t_21_10;
inout [23:0]  sp12_h_l_13_02;
inout [23:0]  sp12_v_t_18_10;
inout [23:0]  sp12_h_l_13_03;
inout [47:0]  sp4_v_t_14_10;
inout [47:0]  sp4_v_b_13_01;
inout [23:0]  sp12_h_l_13_05;
inout [47:0]  sp4_v_b_13_06;
inout [23:0]  sp12_h_l_13_06;
inout [47:0]  sp4_v_t_13_10;
inout [23:0]  sp12_v_t_16_10;
inout [23:0]  sp12_v_t_17_10;
inout [23:0]  sp12_v_t_22_10;
inout [23:0]  sp12_v_t_23_10;
inout [47:0]  sp4_v_b_13_08;
inout [47:0]  sp4_h_l_13_06;
inout [23:0]  sp12_v_t_19_10;
inout [47:0]  sp4_h_l_13_10;
inout [47:0]  sp4_v_b_13_02;
inout [23:0]  sp12_h_l_13_10;
inout [47:0]  sp4_v_b_13_05;
inout [175:0]  wl;
inout [23:0]  sp12_h_l_13_09;
inout [47:0]  sp4_h_l_13_08;
inout [47:0]  sp4_v_b_13_04;
inout [47:0]  sp4_h_l_13_01;
inout [47:0]  sp4_h_l_13_07;
inout [47:0]  sp4_v_t_17_10;
inout [47:0]  sp4_v_b_13_07;
inout [15:0]  sp4_v_t_25_10;
inout [175:0]  vdd_cntl;
inout [23:0]  sp12_v_t_20_10;
inout [47:0]  sp4_v_t_22_10;
inout [175:0]  reset_b;
inout [23:0]  sp12_v_t_24_10;

input [7:0]  tnl_op_24_10;
input [7:0]  lft_op_13_01;
input [7:0]  lft_op_13_03;
input [7:0]  top_op_18_10;
input [7:0]  lft_op_13_04;
input [7:0]  tnr_op_14_10;
input [7:0]  tnl_op_23_10;
input [7:0]  top_op_17_10;
input [7:0]  tnr_op_23_10;
input [7:0]  top_op_20_10;
input [7:0]  tnr_op_13_10;
input [7:0]  glb_in;
input [1:0]  bm_sdo_i;
input [7:0]  lft_op_13_05;
input [19:0]  padin_r;
input [7:0]  tnl_op_21_10;
input [7:0]  lft_op_13_07;
input [7:0]  tnr_op_17_10;
input [47:24]  spiout_b;
input [7:0]  bm_sa_i;
input [47:24]  spioeb_b;
input [7:0]  lft_op_13_02;
input [7:0]  tnr_op_21_10;
input [7:0]  top_op_16_10;
input [7:0]  tnl_op_19_10;
input [3:0]  bnl_op_13_01;
input [7:0]  top_op_15_10;
input [9:0]  cdone_in_rgt_b;
input [7:0]  tnl_op_18_10;
input [7:0]  tnl_op_15_10;
input [7:0]  tnl_op_20_10;
input [7:0]  tnr_op_19_10;
input [7:0]  lft_op_13_08;
input [7:0]  tnl_op_25_10;
input [47:24]  padin_b;
input [7:0]  lft_op_13_09;
input [7:0]  tnr_op_20_10;
input [7:0]  tnl_op_22_10;
input [7:0]  top_op_23_10;
input [1:0]  bm_sclkrw_i;
input [7:0]  top_op_21_10;
input [7:0]  tnl_op_17_10;
input [7:0]  top_op_24_10;
input [7:0]  lft_op_13_10;
input [7:0]  top_op_22_10;
input [7:0]  tnl_op_16_10;
input [7:0]  tnl_op_13_10;
input [1:0]  bm_sdi_i;
input [3:0]  tnr_op_24_10;
input [19:0]  spioeb_r;
input [7:0]  top_op_13_10;
input [7:0]  tnr_op_18_10;
input [7:0]  lft_op_13_06;
input [7:0]  tnr_op_15_10;
input [7:0]  tnr_op_16_10;
input [7:0]  tnl_op_14_10;
input [7:0]  top_op_14_10;
input [1:0]  bm_sweb_i;
input [11:0]  cdone_in_bot_r;
input [7:0]  top_op_19_10;
input [7:0]  tnr_op_22_10;
input [19:0]  spiout_r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:47]  net_7493;

wire  [0:7]  net_6024;

wire  [0:7]  net_5022;

wire  [0:47]  net_6292;

wire  [0:47]  net_4984;

wire  [0:47]  net_8196;

wire  [0:23]  net_8082;

wire  [0:7]  net_6808;

wire  [3:0]  io_r_07;

wire  [0:23]  net_5758;

wire  [0:7]  net_7732;

wire  [0:7]  net_7872;

wire  [0:23]  net_7130;

wire  [0:1]  net_4929;

wire  [3:0]  io_r_05;

wire  [0:47]  net_7997;

wire  [3:0]  io_r_06;

wire  [0:47]  net_6289;

wire  [3:0]  io_r_04;

wire  [3:0]  io_r_03;

wire  [0:47]  net_5956;

wire  [3:0]  io_r_02;

wire  [3:0]  io_r_01;

wire  [0:23]  net_6540;

wire  [0:23]  net_4849;

wire  [0:7]  net_7648;

wire  [3:0]  io_r_08;

wire  [3:0]  io_r_00;

wire  [3:0]  io_b_46;

wire  [3:0]  io_b_44;

wire  [3:0]  io_b_42;

wire  [3:0]  io_b_40;

wire  [0:23]  net_7268;

wire  [3:0]  io_b_38;

wire  [7:0]  glb_netwk_io_r;

wire  [3:0]  io_b_28;

wire  [3:0]  io_b_30;

wire  [3:0]  io_b_32;

wire  [3:0]  io_b_26;

wire  [7:0]  net2col_drivers;

wire  [0:7]  net_5744;

wire  [0:15]  net_4513;

wire  [7:0]  glb_netwk_13;

wire  [7:0]  glb_netwk_14;

wire  [7:0]  glb_netwk_15;

wire  [7:0]  glb_netwk_16;

wire  [7:0]  glb_netwk_17;

wire  [7:0]  glb_netwk_18;

wire  [7:0]  glb_netwk_19;

wire  [7:0]  glb_netwk_20;

wire  [7:0]  glb_netwk_21;

wire  [7:0]  glb_netwk_22;

wire  [7:0]  glb_netwk_23;

wire  [7:0]  glb_netwk_24;

wire  [3:0]  io_b_36;

wire  [3:0]  io_b_34;

wire  [0:7]  net_5240;

wire  [0:7]  net_4926;

wire  [0:23]  net_5170;

wire  [0:23]  net_6346;

wire  [0:7]  net_7032;

wire  [0:23]  net_4437;

wire  [0:47]  net_7748;

wire  [0:47]  net_6628;

wire  [0:23]  net_6288;

wire  [0:47]  net_6096;

wire  [0:47]  net_6009;

wire  [0:23]  net_8080;

wire  [0:23]  net_5786;

wire  [0:7]  net_4510;

wire  [0:47]  net_5844;

wire  [0:47]  net_7664;

wire  [0:15]  net_4231;

wire  [0:23]  net_5840;

wire  [0:47]  net_6961;

wire  [0:1]  net_4915;

wire  [0:23]  net_5280;

wire  [0:47]  net_6681;

wire  [0:47]  net_5337;

wire  [0:7]  net_5856;

wire  [0:23]  net_5224;

wire  [0:47]  net_8168;

wire  [0:47]  net_7328;

wire  [0:7]  net_5912;

wire  [0:47]  net_7552;

wire  [0:47]  net_7801;

wire  [0:23]  net_7688;

wire  [0:23]  net_5842;

wire  [0:47]  net_7241;

wire  [0:23]  net_5016;

wire  [0:23]  net_6568;

wire  [0:47]  net_5645;

wire  [0:23]  net_5618;

wire  [0:7]  net_5380;

wire  [0:23]  net_8138;

wire  [0:47]  net_7213;

wire  [0:47]  net_6852;

wire  [0:47]  net_6320;

wire  [0:23]  net_6066;

wire  [0:47]  net_8165;

wire  [0:23]  net_7744;

wire  [0:15]  net_4717;

wire  [0:7]  net_7788;

wire  [0:47]  net_6572;

wire  [0:47]  net_5704;

wire  [0:47]  net_7829;

wire  [0:23]  net_7464;

wire  [0:47]  net_7045;

wire  [0:47]  net_5396;

wire  [0:47]  net_6877;

wire  [0:47]  net_5760;

wire  [0:23]  net_7436;

wire  [0:7]  net_7984;

wire  [0:7]  net_8152;

wire  [0:23]  net_5308;

wire  [0:7]  net_7144;

wire  [0:47]  net_6765;

wire  [0:23]  net_5702;

wire  [0:23]  net_7716;

wire  [0:23]  net_4977;

wire  [0:47]  net_6989;

wire  [0:47]  net_5312;

wire  [0:47]  net_7549;

wire  [0:23]  net_5366;

wire  [0:47]  net_5508;

wire  [0:23]  net_7632;

wire  [0:23]  net_7324;

wire  [0:47]  net_6740;

wire  [0:47]  net_6180;

wire  [0:23]  net_7380;

wire  [0:23]  net_5392;

wire  [0:47]  net_6936;

wire  [0:23]  net_6484;

wire  [0:7]  net_6108;

wire  [0:47]  net_7524;

wire  [0:23]  net_5101;

wire  [0:7]  net_5268;

wire  [0:1]  net_5052;

wire  [0:23]  net_7354;

wire  [0:23]  net_6456;

wire  [0:7]  net_7228;

wire  [0:1]  net_4882;

wire  [0:47]  net_6737;

wire  [0:23]  net_6514;

wire  [0:47]  net_7916;

wire  [0:47]  net_5225;

wire  [0:47]  net_6541;

wire  [0:23]  net_5140;

wire  [0:47]  net_6205;

wire  [0:47]  net_5020;

wire  [0:23]  net_4905;

wire  [0:23]  net_5336;

wire  [0:47]  net_6152;

wire  [0:47]  net_5200;

wire  [0:47]  net_5841;

wire  [0:47]  net_5676;

wire  [0:23]  net_5812;

wire  [0:23]  net_7128;

wire  [0:1]  net_4865;

wire  [0:47]  net_5393;

wire  [0:1]  net_4932;

wire  [0:23]  net_7942;

wire  [0:7]  net_5062;

wire  [0:47]  net_7661;

wire  [0:47]  net_7353;

wire  [0:23]  net_5616;

wire  [0:23]  net_7270;

wire  [0:47]  net_7300;

wire  [0:47]  net_4983;

wire  [0:15]  net_4581;

wire  [0:23]  net_5506;

wire  [0:47]  net_5309;

wire  [0:7]  net_5013;

wire  [0:23]  net_5926;

wire  [0:47]  net_5107;

wire  [0:23]  net_6344;

wire  [0:47]  net_7885;

wire  [0:7]  net_6276;

wire  [0:47]  net_6992;

wire  [0:23]  net_4369;

wire  [0:47]  net_7521;

wire  [0:23]  net_4539;

wire  [0:23]  net_6150;

wire  [0:47]  net_7185;

wire  [0:7]  net_6584;

wire  [0:23]  net_7828;

wire  [0:7]  net_7368;

wire  [0:47]  net_5813;

wire  [0:23]  net_7102;

wire  [0:47]  net_5477;

wire  [0:47]  net_5928;

wire  [0:47]  net_7717;

wire  [0:7]  net_6360;

wire  [0:23]  net_7158;

wire  [0:23]  net_7970;

wire  [0:23]  net_6038;

wire  [0:47]  net_5365;

wire  [0:7]  net_7118;

wire  [0:23]  net_4743;

wire  [0:23]  net_5728;

wire  [0:47]  net_8109;

wire  [0:7]  net_5604;

wire  [0:23]  net_6120;

wire  [0:47]  net_6404;

wire  [0:47]  net_5816;

wire  [0:47]  net_8112;

wire  [0:47]  net_7636;

wire  [0:47]  net_4986;

wire  [0:23]  net_7576;

wire  [0:23]  net_5338;

wire  [0:47]  net_6460;

wire  [0:7]  net_7200;

wire  [0:7]  net_6332;

wire  [0:23]  net_8136;

wire  [0:7]  net_7536;

wire  [0:47]  net_6516;

wire  [0:15]  net_4129;

wire  [0:47]  net_4860;

wire  [0:23]  net_6400;

wire  [0:23]  net_7550;

wire  [0:7]  net_6192;

wire  [0:23]  net_5730;

wire  [0:23]  net_6904;

wire  [0:23]  net_5784;

wire  [0:23]  net_5814;

wire  [0:23]  net_7604;

wire  [0:7]  net_6752;

wire  [0:23]  net_6990;

wire  [0:23]  net_5560;

wire  [0:47]  net_5869;

wire  [0:1]  net_4879;

wire  [0:7]  net_6976;

wire  [0:23]  net_7408;

wire  [0:23]  net_4641;

wire  [0:23]  net_6428;

wire  [0:23]  net_6064;

wire  [0:7]  net_5958;

wire  [0:23]  net_5478;

wire  [0:47]  net_6345;

wire  [0:47]  net_7860;

wire  [0:15]  net_4683;

wire  [0:23]  net_6822;

wire  [0:7]  net_6864;

wire  [0:23]  net_5868;

wire  [0:47]  net_5533;

wire  [0:47]  net_5017;

wire  [0:47]  net_5197;

wire  [0:15]  net_4615;

wire  [0:47]  net_6012;

wire  [0:23]  net_7884;

wire  [0:47]  net_5109;

wire  [0:23]  net_7156;

wire  [0:47]  net_6488;

wire  [0:23]  net_6652;

wire  [0:23]  net_7772;

wire  [0:23]  net_7184;

wire  [0:23]  net_7242;

wire  [0:15]  net_4547;

wire  [0:23]  net_8110;

wire  [0:7]  net_5940;

wire  [0:23]  net_7634;

wire  [0:23]  net_6092;

wire  [0:47]  net_4943;

wire  [0:23]  net_6176;

wire  [0:47]  net_6824;

wire  [0:15]  net_4445;

wire  [0:47]  net_4944;

wire  [0:23]  net_5100;

wire  [0:47]  net_5144;

wire  [0:47]  net_8140;

wire  [0:47]  net_5284;

wire  [0:47]  net_8025;

wire  [0:7]  net_4936;

wire  [0:23]  net_6094;

wire  [0:7]  net_5800;

wire  [0:23]  net_5041;

wire  [0:15]  net_4751;

wire  [0:23]  net_5870;

wire  [0:7]  net_5828;

wire  [0:47]  net_6065;

wire  [0:23]  net_5644;

wire  [0:47]  net_6768;

wire  [0:47]  net_6908;

wire  [0:7]  net_6668;

wire  [0:15]  net_4479;

wire  [0:47]  net_6121;

wire  [0:23]  net_5196;

wire  [0:23]  net_5674;

wire  [0:47]  net_8081;

wire  [0:47]  net_7773;

wire  [0:23]  net_8054;

wire  [0:23]  net_7072;

wire  [0:47]  net_6880;

wire  [0:47]  net_8028;

wire  [0:23]  net_7044;

wire  [0:47]  net_4859;

wire  [0:47]  net_6684;

wire  [0:47]  net_5021;

wire  [0:23]  net_6626;

wire  [0:23]  net_5756;

wire  [0:23]  net_5646;

wire  [0:47]  net_8193;

wire  [0:23]  net_7018;

wire  [0:23]  net_5142;

wire  [0:23]  net_4573;

wire  [0:23]  net_5924;

wire  [0:23]  net_8052;

wire  [0:7]  net_5632;

wire  [0:7]  net_8040;

wire  [0:7]  net_7256;

wire  [0:15]  net_4027;

wire  [0:47]  net_7381;

wire  [0:47]  net_7269;

wire  [0:23]  net_5198;

wire  [0:7]  net_5466;

wire  [0:15]  net_4411;

wire  [0:47]  net_8053;

wire  [0:23]  net_7466;

wire  [0:47]  net_7496;

wire  [0:47]  net_7944;

wire  [0:23]  net_6542;

wire  [0:47]  net_4940;

wire  [0:23]  net_6204;

wire  [0:23]  net_5168;

wire  [0:47]  net_6656;

wire  [0:47]  net_5561;

wire  [0:7]  net_7088;

wire  [0:7]  net_7592;

wire  [0:47]  net_7244;

wire  [0:7]  net_5184;

wire  [0:23]  net_6624;

wire  [0:23]  net_5450;

wire  [0:23]  net_6932;

wire  [0:47]  net_7073;

wire  [0:47]  net_6600;

wire  [0:23]  net_6960;

wire  [0:23]  net_4505;

wire  [0:47]  net_7132;

wire  [0:7]  net_5688;

wire  [0:23]  net_6512;

wire  [0:47]  net_5536;

wire  [0:47]  net_6429;

wire  [0:23]  net_6402;

wire  [0:23]  net_6710;

wire  [0:23]  net_6680;

wire  [0:7]  net_7284;

wire  [0:23]  net_7718;

wire  [0:23]  net_5982;

wire  [0:7]  net_5548;

wire  [0:47]  net_5984;

wire  [0:47]  net_7129;

wire  [0:23]  net_4675;

wire  [0:23]  net_4471;

wire  [0:7]  net_6612;

wire  [0:23]  net_7886;

wire  [0:47]  net_7272;

wire  [0:47]  net_5729;

wire  [0:23]  net_5590;

wire  [0:7]  net_6724;

wire  [0:47]  net_7776;

wire  [0:23]  net_7998;

wire  [0:7]  net_6528;

wire  [0:23]  net_6596;

wire  [0:15]  net_4095;

wire  [0:47]  net_7689;

wire  [0:47]  net_6432;

wire  [0:7]  net_7902;

wire  [0:7]  net_6472;

wire  [0:7]  net_6556;

wire  [0:47]  net_5897;

wire  [0:7]  net_4748;

wire  [0:7]  net_8068;

wire  [0:47]  net_7913;

wire  [0:47]  net_7692;

wire  [0:47]  net_6264;

wire  [0:23]  net_6010;

wire  [0:23]  net_7326;

wire  [0:47]  net_7101;

wire  [0:23]  net_7856;

wire  [0:23]  net_6820;

wire  [0:23]  net_5588;

wire  [0:23]  net_8166;

wire  [0:7]  net_7676;

wire  [0:47]  net_5981;

wire  [0:47]  net_7468;

wire  [0:1]  net_5051;

wire  [0:23]  net_5310;

wire  [0:7]  net_7844;

wire  [0:23]  net_6736;

wire  [0:7]  net_5408;

wire  [0:47]  net_7076;

wire  [0:23]  net_7382;

wire  [0:7]  net_6416;

wire  [0:47]  net_6821;

wire  [0:47]  net_6317;

wire  [0:7]  net_7816;

wire  [0:1]  net_4990;

wire  [0:15]  net_4061;

wire  [0:7]  net_6892;

wire  [0:7]  net_5716;

wire  [0:23]  net_7522;

wire  [0:47]  net_5424;

wire  [0:23]  net_5015;

wire  [0:47]  net_5788;

wire  [0:47]  net_6124;

wire  [0:23]  net_5562;

wire  [0:7]  net_6500;

wire  [0:47]  net_6037;

wire  [0:23]  net_7016;

wire  [0:7]  net_5660;

wire  [0:23]  net_7438;

wire  [0:23]  net_5952;

wire  [0:7]  net_8012;

wire  [0:15]  net_4377;

wire  [0:7]  net_5884;

wire  [0:23]  net_7352;

wire  [0:47]  net_5925;

wire  [0:7]  net_5094;

wire  [0:47]  net_6373;

wire  [0:47]  net_7409;

wire  [0:47]  net_7972;

wire  [0:7]  net_6248;

wire  [0:47]  net_6625;

wire  [0:23]  net_7046;

wire  [0:47]  net_7941;

wire  [0:7]  net_4876;

wire  [0:47]  net_5732;

wire  [0:7]  net_4945;

wire  [0:23]  net_8024;

wire  [0:23]  net_6878;

wire  [0:7]  net_7172;

wire  [0:7]  net_6444;

wire  [0:15]  net_4333;

wire  [0:15]  net_4299;

wire  [0:47]  net_5340;

wire  [0:23]  net_6486;

wire  [0:47]  net_5449;

wire  [0:47]  net_5018;

wire  [0:23]  net_5394;

wire  [0:47]  net_5281;

wire  [0:47]  net_5757;

wire  [0:23]  net_7212;

wire  [0:47]  net_5592;

wire  [0:47]  net_7104;

wire  [0:23]  net_7746;

wire  [0:23]  net_8164;

wire  [0:47]  net_5480;

wire  [0:15]  net_4163;

wire  [0:47]  net_5172;

wire  [0:23]  net_5476;

wire  [0:47]  net_4985;

wire  [0:23]  net_8192;

wire  [0:47]  net_6796;

wire  [0:7]  net_6220;

wire  [0:47]  net_7577;

wire  [0:47]  net_7216;

wire  [0:7]  net_7004;

wire  [0:47]  net_7048;

wire  [0:7]  net_7340;

wire  [0:23]  net_7074;

wire  [0:47]  net_5169;

wire  [0:47]  net_7440;

wire  [0:47]  net_5617;

wire  [0:47]  net_7832;

wire  [0:23]  net_7690;

wire  [0:23]  net_6876;

wire  [0:23]  net_5422;

wire  [0:47]  net_7720;

wire  [0:47]  net_7888;

wire  [0:47]  net_7608;

wire  [0:47]  net_6597;

wire  [0:23]  net_6962;

wire  [0:23]  net_5448;

wire  [0:23]  net_5226;

wire  [0:23]  net_4607;

wire  [0:23]  net_6316;

wire  [0:47]  net_6093;

wire  [0:23]  net_6792;

wire  [0:23]  net_7606;

wire  [0:23]  net_4403;

wire  [0:7]  net_7704;

wire  [0:47]  net_6236;

wire  [0:23]  net_7774;

wire  [0:23]  net_6850;

wire  [0:7]  net_5968;

wire  [0:23]  net_5532;

wire  [0:23]  net_6848;

wire  [0:23]  net_7940;

wire  [0:23]  net_6934;

wire  [0:23]  net_7410;

wire  [0:23]  net_5898;

wire  [0:47]  net_6485;

wire  [0:7]  net_8124;

wire  [0:23]  net_4852;

wire  [0:47]  net_6457;

wire  [0:23]  net_5252;

wire  [0:23]  net_4938;

wire  [0:47]  net_6376;

wire  [0:23]  net_7660;

wire  [0:47]  net_7297;

wire  [0:7]  net_6052;

wire  [0:23]  net_7912;

wire  [0:47]  net_7633;

wire  [0:23]  net_7548;

wire  [0:47]  net_7605;

wire  [0:23]  net_7996;

wire  [0:47]  net_6513;

wire  [0:23]  net_6148;

wire  [0:47]  net_5900;

wire  [0:23]  net_7578;

wire  [0:47]  net_6544;

wire  [0:23]  net_5896;

wire  [0:7]  net_7760;

wire  [0:7]  net_6640;

wire  [0:23]  net_6260;

wire  [0:23]  net_4939;

wire  [0:23]  net_7298;

wire  [0:23]  net_7968;

wire  [0:23]  net_5420;

wire  [0:47]  net_6149;

wire  [0:47]  net_5953;

wire  [0:23]  net_6654;

wire  [0:23]  net_7214;

wire  [0:47]  net_6040;

wire  [0:47]  net_7857;

wire  [0:47]  net_5108;

wire  [0:47]  net_6964;

wire  [0:23]  net_7186;

wire  [0:47]  net_5701;

wire  [0:47]  net_5648;

wire  [0:47]  net_8000;

wire  [0:47]  net_5368;

wire  [0:23]  net_4973;

wire  [0:47]  net_7969;

wire  [0:47]  net_7745;

wire  [0:47]  net_8056;

wire  [0:47]  net_4862;

wire  [0:23]  net_6008;

wire  [0:23]  net_7800;

wire  [0:47]  net_8084;

wire  [0:47]  net_4861;

wire  [0:23]  net_6708;

wire  [0:1]  net_4989;

wire  [0:7]  net_5510;

wire  [0:7]  net_5000;

wire  [0:23]  net_6764;

wire  [0:47]  net_5110;

wire  [0:47]  net_5872;

wire  [0:1]  net_5003;

wire  [0:23]  net_4976;

wire  [0:7]  net_6304;

wire  [0:15]  net_4649;

wire  [0:1]  net_5065;

wire  [0:23]  net_7520;

wire  [0:47]  net_6933;

wire  [0:23]  net_7100;

wire  [0:23]  net_5980;

wire  [0:47]  net_7160;

wire  [0:47]  net_7412;

wire  [0:47]  net_7580;

wire  [0:47]  net_7437;

wire  [0:23]  net_7914;

wire  [0:47]  net_5589;

wire  [0:7]  net_6136;

wire  [0:47]  net_5421;

wire  [0:23]  net_6906;

wire  [0:23]  net_5954;

wire  [0:7]  net_7424;

wire  [0:23]  net_5504;

wire  [0:1]  net_4866;

wire  [0:7]  net_6836;

wire  [0:7]  net_7620;

wire  [0:1]  net_5068;

wire  [0:47]  net_7465;

wire  [0:23]  net_5282;

wire  [0:23]  net_8108;

wire  [0:47]  net_6793;

wire  [0:47]  net_7017;

wire  [0:47]  net_5253;

wire  [0:7]  net_7956;

wire  [0:47]  net_6208;

wire  [0:47]  net_7384;

wire  [0:23]  net_7858;

wire  [0:23]  net_6262;

wire  [0:47]  net_6905;

wire  [0:47]  net_7157;

wire  [0:23]  net_7662;

wire  [0:47]  net_6177;

wire  [0:47]  net_6401;

wire  [0:23]  net_6766;

wire  [0:7]  net_5520;

wire  [0:23]  net_5672;

wire  [0:47]  net_6569;

wire  [0:1]  net_5006;

wire  [0:47]  net_5505;

wire  [0:23]  net_6206;

wire  [0:7]  net_4970;

wire  [0:47]  net_5452;

wire  [0:7]  net_6948;

wire  [0:47]  net_7356;

wire  [0:7]  net_5996;

wire  [0:23]  net_4853;

wire  [0:47]  net_6709;

wire  [0:47]  net_7804;

wire  [0:23]  net_5364;

wire  [0:23]  net_7492;

wire  [0:23]  net_6178;

wire  [0:47]  net_7020;

wire  [0:47]  net_5785;

wire  [0:23]  net_7802;

wire  [0:7]  net_7060;

wire  [0:23]  net_8026;

wire  [0:47]  net_6068;

wire  [0:47]  net_5564;

wire  [0:47]  net_6348;

wire  [0:47]  net_7325;

wire  [0:23]  net_6372;

wire  [0:7]  net_4829;

wire  [0:23]  net_5534;

wire  [0:47]  net_6233;

wire  [0:23]  net_7494;

wire  [0:47]  net_5141;

wire  [0:23]  net_6232;

wire  [0:47]  net_5228;

wire  [0:47]  net_6261;

wire  [0:47]  net_8137;

wire  [0:7]  net_6920;

wire  [0:23]  net_6988;

wire  [0:1]  net_4916;

wire  [0:7]  net_4953;

wire  [0:47]  net_6849;

wire  [0:23]  net_6122;

wire  [0:7]  net_8208;

wire  [0:23]  net_5700;

wire  [0:47]  net_5620;

wire  [0:47]  net_7188;

wire  [0:23]  net_6036;

wire  [0:23]  net_8194;

wire  [0:23]  net_7296;

wire  [0:47]  net_5256;

wire  [0:47]  net_4941;

wire  [0:47]  net_6653;

wire  [0:15]  net_4265;

wire  [0:47]  net_5673;

wire  [0:23]  net_5254;

wire  [0:23]  net_7240;

wire  [0:47]  net_6712;

wire  [0:23]  net_4709;

wire  [0:23]  net_7830;



bram_bufferx4x6 I904 ( .in(sdpp), .out(sdpd));
bram_bufferx4x6 I905 ( .in(sdi), .out(net_04047));
bram_bufferx4x6 I906 ( .in(sdi_pad), .out(net_04056));
lowla_modified I903 ( .clk(net_4785), .min(sdpd), .lao(sdo_pad));
lowla_modified I886 ( .clk(tclk_mi), .min(net_04056), .lao(net_4013));
lowla_modified I895 ( .clk(tclk_i), .min(net_04047), .lao(net_4759));
io_col4_rowright I_25_01_ior01 ( .ceb(ceb_o), .cf(cf_r[23:0]),
     .vdd_cntl(vdd_cntl[31:16]), .hold(hold_r_b),
     .fabric_out(net_4011), .sdo(net_4012), .sdi(net_4013),
     .spiout(spiout_r[1:0]), .cdone_in(cdone_in_rgt_b[0]),
     .spioeb(spioeb_r[1:0]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[1:0]), .pado(pado_r[1:0]),
     .padeb(padeb_r[1:0]), .sp4_v_t(net_4027[0:15]),
     .sp4_h_l(net_7549[0:47]), .sp12_h_l(net_7548[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[1:0]), .tnl_op(net_8068[0:7]),
     .lft_op(net_7592[0:7]), .bnl_op({io_b_46[3], io_b_46[2],
     io_b_46[1], io_b_46[0], io_b_46[3], io_b_46[2], io_b_46[1],
     io_b_46[0]}), .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(net_4717[0:15]), .wl(wl[31:16]), .bl(bl[1311:1294]),
     .slf_op(io_r_00[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_02_ior02 ( .ceb(ceb_o), .cf(cf_r[47:24]),
     .vdd_cntl(vdd_cntl[47:32]), .hold(hold_r_b),
     .fabric_out(net_8276), .sdo(net_4285), .sdi(net_4012),
     .spiout(spiout_r[3:2]), .cdone_in(cdone_in_rgt_b[1]),
     .spioeb(spioeb_r[3:2]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[3:2]), .pado(pado_r[3:2]),
     .padeb(padeb_r[3:2]), .sp4_v_t(net_4061[0:15]),
     .sp4_h_l(net_7465[0:47]), .sp12_h_l(net_7464[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[3:2]), .tnl_op(net_8208[0:7]),
     .lft_op(net_8068[0:7]), .bnl_op(net_7592[0:7]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net_4027[0:15]), .wl(wl[47:32]), .bl(bl[1311:1294]),
     .slf_op(io_r_01[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_05_ior09 ( .ceb(ceb_o), .cf(cf_r[119:96]),
     .vdd_cntl(vdd_cntl[95:80]), .hold(hold_r_b),
     .fabric_out(net_8269), .sdo(net_4080), .sdi(net_4318),
     .spiout(spiout_r[9:8]), .cdone_in(cdone_in_rgt_b[4]),
     .spioeb(spioeb_r[9:8]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[9:8]), .pado(pado_r[9:8]),
     .padeb(padeb_r[9:8]), .sp4_v_t(net_4095[0:15]),
     .sp4_h_l(net_6149[0:47]), .sp12_h_l(net_6148[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[9:8]), .tnl_op(net_7284[0:7]),
     .lft_op(net_6192[0:7]), .bnl_op(net_6052[0:7]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net_4333[0:15]), .wl(wl[95:80]), .bl(bl[1311:1294]),
     .slf_op(io_r_04[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_06_ior11 ( .ceb(ceb_o), .cf(cf_r[143:120]),
     .vdd_cntl(vdd_cntl[111:96]), .hold(hold_r_b),
     .fabric_out(net_8263), .sdo(net_4217), .sdi(net_4080),
     .spiout(spiout_r[11:10]), .cdone_in(cdone_in_rgt_b[5]),
     .spioeb(spioeb_r[11:10]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[11:10]), .pado(pado_r[11:10]),
     .padeb(padeb_r[11:10]), .sp4_v_t(net_4129[0:15]),
     .sp4_h_l(net_6065[0:47]), .sp12_h_l(net_6064[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[11:10]), .tnl_op(net_7424[0:7]),
     .lft_op(net_7284[0:7]), .bnl_op(net_6192[0:7]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net_4095[0:15]), .wl(wl[111:96]), .bl(bl[1311:1294]),
     .slf_op(io_r_05[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_09_ior17 ( .ceb(ceb_o), .cf(cf_r[215:192]),
     .vdd_cntl(vdd_cntl[159:144]), .hold(hold_r_b),
     .fabric_out(net_4147), .sdo(net_4148), .sdi(net_4250),
     .spiout(spiout_r[17:16]), .cdone_in(cdone_in_rgt_b[8]),
     .spioeb(spioeb_r[17:16]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[17:16]), .pado(pado_r[17:16]),
     .padeb(padeb_r[17:16]), .sp4_v_t(net_4163[0:15]),
     .sp4_h_l(net_6765[0:47]), .sp12_h_l(net_6764[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[17:16]), .tnl_op(slf_op_24_10[7:0]),
     .lft_op(net_6808[0:7]), .bnl_op(net_6668[0:7]),
     .pgate(pgate[159:144]), .reset(reset_b[159:144]),
     .sp4_v_b(net_4265[0:15]), .wl(wl[159:144]), .bl(bl[1311:1294]),
     .slf_op(io_r_08[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_10_ior19 ( .ceb(ceb_o), .cf(cf_r[239:216]),
     .vdd_cntl(vdd_cntl[175:160]), .hold(hold_r_b),
     .fabric_out(net_4181), .sdo(sdo), .sdi(net_4148),
     .spiout(spiout_r[19:18]), .cdone_in(cdone_in_rgt_b[9]),
     .spioeb(spioeb_r[19:18]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[19:18]), .pado(pado_r[19:18]),
     .padeb(padeb_r[19:18]), .sp4_v_t(sp4_v_t_25_10[15:0]),
     .sp4_h_l(net_6681[0:47]), .sp12_h_l(net_6680[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[19:18]), .tnl_op(tnl_op_25_10[7:0]),
     .lft_op(slf_op_24_10[7:0]), .bnl_op(net_6808[0:7]),
     .pgate(pgate[175:160]), .reset(reset_b[175:160]),
     .sp4_v_b(net_4163[0:15]), .wl(wl[175:160]), .bl(bl[1311:1294]),
     .slf_op(slf_op_25_10[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_07_ior13 ( .ceb(ceb_o), .cf(cf_r[167:144]),
     .vdd_cntl(vdd_cntl[127:112]), .hold(hold_r_b),
     .fabric_out(net_8266), .sdo(net_4216), .sdi(net_4217),
     .spiout(spiout_r[13:12]), .cdone_in(cdone_in_rgt_b[6]),
     .spioeb(spioeb_r[13:12]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[13:12]), .pado(pado_r[13:12]),
     .padeb(padeb_r[13:12]), .sp4_v_t(net_4231[0:15]),
     .sp4_h_l(net_7381[0:47]), .sp12_h_l(net_7380[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[13:12]), .tnl_op(net_6668[0:7]),
     .lft_op(net_7424[0:7]), .bnl_op(net_7284[0:7]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net_4129[0:15]), .wl(wl[127:112]), .bl(bl[1311:1294]),
     .slf_op(io_r_06[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_08_ior15 ( .ceb(ceb_o), .cf(cf_r[191:168]),
     .vdd_cntl(vdd_cntl[143:128]), .hold(hold_r_b),
     .fabric_out(net_4249), .sdo(net_4250), .sdi(net_4216),
     .spiout(spiout_r[15:14]), .cdone_in(cdone_in_rgt_b[7]),
     .spioeb(spioeb_r[15:14]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[15:14]), .pado(pado_r[15:14]),
     .padeb(padeb_r[15:14]), .sp4_v_t(net_4265[0:15]),
     .sp4_h_l(net_7297[0:47]), .sp12_h_l(net_7296[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[15:14]), .tnl_op(net_6808[0:7]),
     .lft_op(net_6668[0:7]), .bnl_op(net_7424[0:7]),
     .pgate(pgate[143:128]), .reset(reset_b[143:128]),
     .sp4_v_b(net_4231[0:15]), .wl(wl[143:128]), .bl(bl[1311:1294]),
     .slf_op(io_r_07[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_03_ior05 ( .ceb(ceb_o), .cf(cf_r[71:48]),
     .vdd_cntl(vdd_cntl[63:48]), .hold(hold_r_b),
     .fabric_out(net_4283), .sdo(net_4284), .sdi(net_4285),
     .spiout(spiout_r[5:4]), .cdone_in(cdone_in_rgt_b[2]),
     .spioeb(spioeb_r[5:4]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[5:4]), .pado(pado_r[5:4]),
     .padeb(padeb_r[5:4]), .sp4_v_t(net_4299[0:15]),
     .sp4_h_l(net_8165[0:47]), .sp12_h_l(net_8164[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[5:4]), .tnl_op(net_6052[0:7]),
     .lft_op(net_8208[0:7]), .bnl_op(net_8068[0:7]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net_4061[0:15]), .wl(wl[63:48]), .bl(bl[1311:1294]),
     .slf_op(io_r_02[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_04_ior07 ( .ceb(ceb_o), .cf(cf_r[95:72]),
     .vdd_cntl(vdd_cntl[79:64]), .hold(hold_r_b),
     .fabric_out(net_4317), .sdo(net_4318), .sdi(net_4284),
     .spiout(spiout_r[7:6]), .cdone_in(cdone_in_rgt_b[3]),
     .spioeb(spioeb_r[7:6]), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_r[7:6]), .pado(pado_r[7:6]),
     .padeb(padeb_r[7:6]), .sp4_v_t(net_4333[0:15]),
     .sp4_h_l(net_8081[0:47]), .sp12_h_l(net_8080[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[7:6]), .tnl_op(net_6192[0:7]),
     .lft_op(net_6052[0:7]), .bnl_op(net_8208[0:7]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net_4299[0:15]), .wl(wl[79:64]), .bl(bl[1311:1294]),
     .slf_op(io_r_03[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_lb I_23_00_iob45 ( .ceb(net_04788), .cf(cf_b[551:528]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_4351),
     .sdo(net_4352), .sdi(net_4386), .spiout(spiout_b[45:44]),
     .cdone_in(cdone_in_bot_r[10]), .spioeb(spioeb_b[45:44]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[45:44]), .pado(pado_b[45:44]),
     .padeb(padeb_b[45:44]), .sp4_v_t(net_4411[0:15]),
     .sp4_h_l(net_7496[0:47]), .sp12_h_l(net_4369[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[45:44]), .tnl_op(net_5548[0:7]),
     .lft_op(net_7536[0:7]), .bnl_op(net_7592[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4377[0:15]), .wl(wl[15:0]), .bl({bl[1187], bl[1186],
     bl[1225], bl[1223], bl[1214], bl[1220], bl[1219], bl[1218],
     bl[1217], bl[1216], bl[1197], bl[1196], bl[1195], bl[1194],
     bl[1193], bl[1192], bl[1227], bl[1226]}), .slf_op(io_b_44[3:0]),
     .glb_netwk(glb_netwk_23[7:0]));
io_col4_lb I_22_00_iob43 ( .ceb(net_04788), .cf(cf_b[527:504]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8278),
     .sdo(net_4386), .sdi(net_4420), .spiout(spiout_b[43:42]),
     .cdone_in(cdone_in_bot_r[9]), .spioeb(spioeb_b[43:42]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[43:42]), .pado(pado_b[43:42]),
     .padeb(padeb_b[43:42]), .sp4_v_t(net_4445[0:15]),
     .sp4_h_l(net_5564[0:47]), .sp12_h_l(net_4403[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[43:42]), .tnl_op(net_5520[0:7]),
     .lft_op(net_5548[0:7]), .bnl_op(net_7536[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4411[0:15]), .wl(wl[15:0]), .bl({bl[1133], bl[1132],
     bl[1171], bl[1169], bl[1160], bl[1166], bl[1165], bl[1164],
     bl[1163], bl[1162], bl[1143], bl[1142], bl[1141], bl[1140],
     bl[1139], bl[1138], bl[1173], bl[1172]}), .slf_op(io_b_42[3:0]),
     .glb_netwk(glb_netwk_22[7:0]));
io_col4_lb I_21_00_iob41 ( .ceb(net_04788), .cf(cf_b[503:480]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8270),
     .sdo(net_4420), .sdi(net_4454), .spiout(spiout_b[41:40]),
     .cdone_in(cdone_in_bot_r[8]), .spioeb(spioeb_b[41:40]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[41:40]), .pado(pado_b[41:40]),
     .padeb(padeb_b[41:40]), .sp4_v_t(net_4479[0:15]),
     .sp4_h_l(net_5480[0:47]), .sp12_h_l(net_4437[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[41:40]), .tnl_op(net_4748[0:7]),
     .lft_op(net_5520[0:7]), .bnl_op(net_5548[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4445[0:15]), .wl(wl[15:0]), .bl({bl[1079], bl[1078],
     bl[1117], bl[1115], bl[1106], bl[1112], bl[1111], bl[1110],
     bl[1109], bl[1108], bl[1089], bl[1088], bl[1087], bl[1086],
     bl[1085], bl[1084], bl[1119], bl[1118]}), .slf_op(io_b_40[3:0]),
     .glb_netwk(glb_netwk_21[7:0]));
io_col4_lb I_20_00_iob39 ( .ceb(net_04788), .cf(cf_b[479:456]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8250),
     .sdo(net_4454), .sdi(net_4726), .spiout(spiout_b[39:38]),
     .cdone_in(cdone_in_bot_r[7]), .spioeb(spioeb_b[39:38]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[39:38]), .pado(pado_b[39:38]),
     .padeb(padeb_b[39:38]), .sp4_v_t(net_4751[0:15]),
     .sp4_h_l(net_4860[0:47]), .sp12_h_l(net_4471[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[39:38]), .tnl_op(net_4510[0:7]),
     .lft_op(net_4748[0:7]), .bnl_op(net_5520[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4479[0:15]), .wl(wl[15:0]), .bl({bl[1025], bl[1024],
     bl[1063], bl[1061], bl[1052], bl[1058], bl[1057], bl[1056],
     bl[1055], bl[1054], bl[1035], bl[1034], bl[1033], bl[1032],
     bl[1031], bl[1030], bl[1065], bl[1064]}), .slf_op(io_b_38[3:0]),
     .glb_netwk(glb_netwk_20[7:0]));
io_col4_lb I_18_00_iob35 ( .ceb(net_04788), .cf(cf_b[431:408]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8272),
     .sdo(net_4488), .sdi(net_4522), .spiout(spiout_b[35:34]),
     .cdone_in(cdone_in_bot_r[5]), .spioeb(spioeb_b[35:34]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[35:34]), .pado(pado_b[35:34]),
     .padeb(padeb_b[35:34]), .sp4_v_t(net_4547[0:15]),
     .sp4_h_l(net_5144[0:47]), .sp12_h_l(net_4505[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[35:34]), .tnl_op(net_5268[0:7]),
     .lft_op(net_5184[0:7]), .bnl_op(net_4510[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4513[0:15]), .wl(wl[15:0]), .bl({bl[929], bl[928],
     bl[967], bl[965], bl[956], bl[962], bl[961], bl[960], bl[959],
     bl[958], bl[939], bl[938], bl[937], bl[936], bl[935], bl[934],
     bl[969], bl[968]}), .slf_op(io_b_34[3:0]),
     .glb_netwk(glb_netwk_18[7:0]));
io_col4_lb I_17_00_iob33 ( .ceb(net_04788), .cf(cf_b[407:384]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8280),
     .sdo(net_4522), .sdi(net_4556), .spiout(spiout_b[33:32]),
     .cdone_in(cdone_in_bot_r[4]), .spioeb(spioeb_b[33:32]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[33:32]), .pado(pado_b[33:32]),
     .padeb(padeb_b[33:32]), .sp4_v_t(net_4581[0:15]),
     .sp4_h_l(net_5284[0:47]), .sp12_h_l(net_4539[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[33:32]), .tnl_op(net_5240[0:7]),
     .lft_op(net_5268[0:7]), .bnl_op(net_5184[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4547[0:15]), .wl(wl[15:0]), .bl({bl[875], bl[874],
     bl[913], bl[911], bl[902], bl[908], bl[907], bl[906], bl[905],
     bl[904], bl[885], bl[884], bl[883], bl[882], bl[881], bl[880],
     bl[915], bl[914]}), .slf_op(io_b_32[3:0]),
     .glb_netwk(glb_netwk_17[7:0]));
io_col4_lb I_16_00_iob31 ( .ceb(net_04788), .cf(cf_b[383:360]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8260),
     .sdo(net_4556), .sdi(net_4590), .spiout(spiout_b[31:30]),
     .cdone_in(cdone_in_bot_r[3]), .spioeb(spioeb_b[31:30]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[31:30]), .pado(pado_b[31:30]),
     .padeb(padeb_b[31:30]), .sp4_v_t(net_4615[0:15]),
     .sp4_h_l(net_5200[0:47]), .sp12_h_l(net_4573[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[31:30]), .tnl_op(net_5380[0:7]),
     .lft_op(net_5240[0:7]), .bnl_op(net_5268[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4581[0:15]), .wl(wl[15:0]), .bl({bl[821], bl[820],
     bl[859], bl[857], bl[848], bl[854], bl[853], bl[852], bl[851],
     bl[850], bl[831], bl[830], bl[829], bl[828], bl[827], bl[826],
     bl[861], bl[860]}), .slf_op(io_b_30[3:0]),
     .glb_netwk(glb_netwk_16[7:0]));
io_col4_lb I_15_00_iob29 ( .ceb(net_04788), .cf(cf_b[359:336]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8255),
     .sdo(net_4590), .sdi(net_4624), .spiout(spiout_b[29:28]),
     .cdone_in(cdone_in_bot_r[2]), .spioeb(spioeb_b[29:28]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[29:28]), .pado(pado_b[29:28]),
     .padeb(padeb_b[29:28]), .sp4_v_t(net_4649[0:15]),
     .sp4_h_l(net_5340[0:47]), .sp12_h_l(net_4607[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[29:28]), .tnl_op(net_5408[0:7]),
     .lft_op(net_5380[0:7]), .bnl_op(net_5240[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4615[0:15]), .wl(wl[15:0]), .bl({bl[767], bl[766],
     bl[805], bl[803], bl[794], bl[800], bl[799], bl[798], bl[797],
     bl[796], bl[777], bl[776], bl[775], bl[774], bl[773], bl[772],
     bl[807], bl[806]}), .slf_op(io_b_28[3:0]),
     .glb_netwk(glb_netwk_15[7:0]));
io_col4_lb I_14_00_iob27 ( .ceb(net_04788), .cf(cf_b[335:312]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_4806),
     .sdo(net_4624), .sdi(net_4658), .spiout(spiout_b[27:26]),
     .cdone_in(cdone_in_bot_r[1]), .spioeb(spioeb_b[27:26]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[27:26]), .pado(pado_b[27:26]),
     .padeb(padeb_b[27:26]), .sp4_v_t(net_4683[0:15]),
     .sp4_h_l(net_5424[0:47]), .sp12_h_l(net_4641[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[27:26]), .tnl_op(slf_op_13_01[7:0]),
     .lft_op(net_5408[0:7]), .bnl_op(net_5380[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4649[0:15]), .wl(wl[15:0]), .bl({bl[713], bl[712],
     bl[751], bl[749], bl[740], bl[746], bl[745], bl[744], bl[743],
     bl[742], bl[723], bl[722], bl[721], bl[720], bl[719], bl[718],
     bl[753], bl[752]}), .slf_op(io_b_26[3:0]),
     .glb_netwk(glb_netwk_14[7:0]));
io_col4_lb I_13_00_iob25 ( .ceb(net_04788), .cf(cf_b[311:288]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_4657),
     .sdo(net_4658), .sdi(net_4759), .spiout(spiout_b[25:24]),
     .cdone_in(cdone_in_bot_r[0]), .spioeb(spioeb_b[25:24]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[25:24]), .pado(pado_b[25:24]),
     .padeb(padeb_b[25:24]), .sp4_v_t(sp4_h_l_13_00[15:0]),
     .sp4_h_l(sp4_v_b_13_01[47:0]), .sp12_h_l(net_4675[0:23]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[25:24]),
     .tnl_op(lft_op_13_01[7:0]), .lft_op(slf_op_13_01[7:0]),
     .bnl_op(net_5408[0:7]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(net_4683[0:15]), .wl(wl[15:0]),
     .bl({bl[659], bl[658], bl[697], bl[695], bl[686], bl[692],
     bl[691], bl[690], bl[689], bl[688], bl[669], bl[668], bl[667],
     bl[666], bl[665], bl[664], bl[699], bl[698]}),
     .slf_op(slf_op_13_00[3:0]), .glb_netwk(glb_netwk_13[7:0]));
io_col4_lb I_24_00_iob47 ( .ceb(net_04788), .cf(cf_b[575:552]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_4792),
     .sdo(sdpp), .sdi(net_4352), .spiout(spiout_b[47:46]),
     .cdone_in(cdone_in_bot_r[11]), .spioeb(spioeb_b[47:46]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[47:46]), .pado(pado_b[47:46]),
     .padeb(padeb_b[47:46]), .sp4_v_t(net_4377[0:15]),
     .sp4_h_l(net_7440[0:47]), .sp12_h_l(net_4709[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[47:46]), .tnl_op(net_7536[0:7]),
     .lft_op(net_7592[0:7]), .bnl_op({io_r_00[3], io_r_00[2],
     io_r_00[1], io_r_00[0], io_r_00[3], io_r_00[2], io_r_00[1],
     io_r_00[0]}), .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4717[0:15]), .wl(wl[15:0]), .bl({bl[1241], bl[1240],
     bl[1279], bl[1277], bl[1268], bl[1274], bl[1273], bl[1272],
     bl[1271], bl[1270], bl[1251], bl[1250], bl[1249], bl[1248],
     bl[1247], bl[1246], bl[1281], bl[1280]}), .slf_op(io_b_46[3:0]),
     .glb_netwk(glb_netwk_24[7:0]));
io_col4_lb I_19_00_iob37 ( .ceb(net_04788), .cf(cf_b[455:432]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_r), .fabric_out(net_8258),
     .sdo(net_4726), .sdi(net_4488), .spiout(spiout_b[37:36]),
     .cdone_in(cdone_in_bot_r[6]), .spioeb(spioeb_b[37:36]),
     .mode(net_4775), .shift(net_4783), .hiz_b(net_4779), .r(net_4777),
     .bs_en(net_4787), .tclk(net_4785), .update(net_4781),
     .padin(padin_b[37:36]), .pado(pado_b[37:36]),
     .padeb(padeb_b[37:36]), .sp4_v_t(net_4513[0:15]),
     .sp4_h_l(net_5452[0:47]), .sp12_h_l(net_4743[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[37:36]), .tnl_op(net_5184[0:7]),
     .lft_op(net_4510[0:7]), .bnl_op(net_4748[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net_4751[0:15]), .wl(wl[15:0]), .bl({bl[983], bl[982],
     bl[1009], bl[1007], bl[998], bl[1004], bl[1003], bl[1002],
     bl[1001], bl[1000], bl[993], bl[992], bl[991], bl[990], bl[989],
     bl[988], bl[1011], bl[1010]}), .slf_op(io_b_36[3:0]),
     .glb_netwk(glb_netwk_19[7:0]));
bram_bufferx4 I879 ( .in(shift_mi), .out(shift_o));
bram_bufferx4 I878 ( .in(mode_mi), .out(mode_o));
bram_bufferx4 I880 ( .in(hiz_b_mi), .out(hiz_b_o));
bram_bufferx4 I881 ( .in(update_mi), .out(update_o));
bram_bufferx4 I882 ( .in(r_mi), .out(r_o));
bram_bufferx4 I883 ( .in(bs_en_mi), .out(bs_en_o));
bram_bufferx4 I885 ( .in(tclk_mi), .out(tclk_o));
bram_bufferx4 I900 ( .in(ceb_mi), .out(ceb_o));
bram_bufferx4 I901 ( .in(ceb_i), .out(net_04788));
bram_bufferx4 I887 ( .in(mode_i), .out(net_4775));
bram_bufferx4 I892 ( .in(r_i), .out(net_4777));
bram_bufferx4 I891 ( .in(hiz_b_i), .out(net_4779));
bram_bufferx4 I889 ( .in(update_i), .out(net_4781));
bram_bufferx4 I890 ( .in(shift_i), .out(net_4783));
bram_bufferx4 I888 ( .in(tclk_i), .out(net_4785));
bram_bufferx4 I893 ( .in(bs_en_i), .out(net_4787));
inv_hvt I1014 ( .A(net_4793), .Y(fabric_out_126));
inv_hvt I856 ( .A(net_4790), .Y(padin_94));
inv_hvt I1013 ( .A(net_4792), .Y(net_4793));
inv_hvt I857 ( .A(padin_b[24]), .Y(net_4790));
inv_hvt I848 ( .A(net_4351), .Y(net_4797));
inv_hvt I849 ( .A(net_4797), .Y(fabric_out_122));
inv_hvt I850 ( .A(net_4803), .Y(fabric_out_136));
inv_hvt I851 ( .A(net_4011), .Y(net_4803));
inv_hvt I860 ( .A(net_4807), .Y(fabric_out_98));
inv_hvt I861 ( .A(net_4806), .Y(net_4807));
inv_hvt I858 ( .A(padin_r[19]), .Y(net_4809));
inv_hvt I859 ( .A(net_4809), .Y(padin_162));
inv_hvt I855 ( .A(net_4819), .Y(fabric_out_94));
inv_hvt I853 ( .A(net_4817), .Y(fabric_out_162));
inv_hvt I852 ( .A(net_4181), .Y(net_4817));
inv_hvt I854 ( .A(net_4657), .Y(net_4819));
clk_quad_bufx8 I_quad_driver ( .clko(net2col_drivers[7:0]),
     .clki(glb_in[7:0]));
bram_4kprouting_bbankout I_bram1901 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_bot(vdd_cntl[31:16]), .vdd_cntl_top(vdd_cntl[47:32]),
     .slf_op_top(net_5466[0:7]), .slf_op_bot(net_4510[0:7]),
     .wl_top(wl[47:32]), .wl_bot(wl[31:16]),
     .top_op_top(net_4829[0:7]), .tnr_op_top(net_5510[0:7]),
     .tnr_op_bot(net_5022[0:7]), .tnl_op_top(net_7760[0:7]),
     .tnl_op_bot(net_7732[0:7]), .rgt_op_top(net_5022[0:7]),
     .rgt_op_bot(net_4748[0:7]), .reset_b_top(reset_b[47:32]),
     .reset_b_bot(reset_b[31:16]), .prog(prog),
     .pgate_top(pgate[47:32]), .pgate_bot(pgate[31:16]),
     .lft_op_top(net_7732[0:7]), .lft_op_bot(net_5184[0:7]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bot_op_bot({io_b_36[3],
     io_b_36[2], io_b_36[1], io_b_36[0], io_b_36[3], io_b_36[2],
     io_b_36[1], io_b_36[0]}), .bnr_op_top(net_4748[0:7]),
     .bnr_op_bot({io_b_38[3], io_b_38[2], io_b_38[1], io_b_38[0],
     io_b_38[3], io_b_38[2], io_b_38[1], io_b_38[0]}),
     .bnl_op_top(net_5184[0:7]), .bnl_op_bot({io_b_34[3], io_b_34[2],
     io_b_34[1], io_b_34[0], io_b_34[3], io_b_34[2], io_b_34[1],
     io_b_34[0]}), .sp12_v_t_top(net_4849[0:23]),
     .sp12_v_b_bot(net_4743[0:23]), .bm_init_i(bm_init_i),
     .sp12_h_r_top(net_4852[0:23]), .sp12_h_r_bot(net_4853[0:23]),
     .sp12_h_l_top(net_5308[0:23]), .sp12_h_l_bot(net_5448[0:23]),
     .sp4_v_t_top(net_7916[0:47]), .sp4_v_b_top(net_5312[0:47]),
     .sp4_v_b_bot(net_5452[0:47]), .sp4_r_v_b_top(net_4859[0:47]),
     .sp4_r_v_b_bot(net_4860[0:47]), .sp4_h_r_top(net_4861[0:47]),
     .sp4_h_r_bot(net_4862[0:47]), .sp4_h_l_top(net_5309[0:47]),
     .sp4_h_l_bot(net_5449[0:47]), .bm_sdi_o(net_4865[0:1]),
     .bm_sclkrw_o(net_4866[0:1]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i[1:0]),
     .bm_rcapmux_en_o(net_4874), .bm_init_o(net_4875),
     .bm_sa_o(net_4876[0:7]), .bm_sclk_o(net_4877),
     .bm_sreb_o(net_4878), .bm_sweb_o(net_4879[0:1]),
     .bm_wdummymux_en_o(net_4880), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sdo_i(net_4882[0:1]), .bm_sdo_o(bm_sdo_o[1:0]));
bram_4kprouting_bbank I_bram1907 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_top(vdd_cntl[143:128]),
     .vdd_cntl_bot(vdd_cntl[127:112]), .slf_op_top(net_6528[0:7]),
     .slf_op_bot(net_4953[0:7]), .wl_top(wl[143:128]),
     .wl_bot(wl[127:112]), .top_op_top(net_7118[0:7]),
     .tnl_op_top(net_6248[0:7]), .tnl_op_bot(net_6220[0:7]),
     .reset_b_top(reset_b[143:128]), .reset_b_bot(reset_b[127:112]),
     .prog(prog), .pgate_top(pgate[143:128]),
     .pgate_bot(pgate[127:112]), .lft_op_top(net_6220[0:7]),
     .lft_op_bot(net_6976[0:7]), .bm_wdummymux_en_i(net_5004),
     .bot_op_bot(net_7144[0:7]), .bnl_op_top(net_6976[0:7]),
     .bnl_op_bot(net_6948[0:7]), .sp12_v_t_top(net_4905[0:23]),
     .sp12_v_b_bot(net_4973[0:23]), .bm_init_i(net_4999),
     .sp12_h_l_top(net_7100[0:23]), .sp12_h_l_bot(net_7128[0:23]),
     .sp4_v_t_top(net_6516[0:47]), .sp4_v_b_top(net_7104[0:47]),
     .sp4_v_b_bot(net_7132[0:47]), .sp4_h_l_top(net_7101[0:47]),
     .sp4_h_l_bot(net_7129[0:47]), .bm_sdi_o(net_4915[0:1]),
     .bm_sclkrw_o(net_4916[0:1]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(net_4998), .bm_sa_i(net_5000[0:7]),
     .bm_sclk_i(net_5001), .bm_sclkrw_i(net_4990[0:1]),
     .bm_sreb_i(net_5002), .bm_sweb_i(net_5003[0:1]),
     .bm_rcapmux_en_o(net_4924), .bm_init_o(net_4925),
     .bm_sa_o(net_4926[0:7]), .bm_sclk_o(net_4927),
     .bm_sreb_o(net_4928), .bm_sweb_o(net_4929[0:1]),
     .bm_wdummymux_en_o(net_4930), .bm_sdi_i(net_4989[0:1]),
     .bm_sdo_i(net_4932[0:1]), .bm_sdo_o(net_5006[0:1]),
     .bnr_op_top(net_5958[0:7]), .rgt_op_top(net_5094[0:7]),
     .tnr_op_top(net_4936[0:7]), .tnr_op_bot(net_5094[0:7]),
     .sp12_h_r_top(net_4938[0:23]), .sp12_h_r_bot(net_4939[0:23]),
     .sp4_h_r_bot(net_4940[0:47]), .sp4_h_r_top(net_4941[0:47]),
     .rgt_op_bot(net_5958[0:7]), .sp4_r_v_b_top(net_4943[0:47]),
     .sp4_r_v_b_bot(net_4944[0:47]), .bnr_op_bot(net_4945[0:7]));
bram_4kprouting_bbank I_bram1905 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_bot(vdd_cntl[95:80]), .vdd_cntl_top(vdd_cntl[111:96]),
     .slf_op_top(net_7144[0:7]), .slf_op_bot(net_7902[0:7]),
     .wl_top(wl[111:96]), .wl_bot(wl[95:80]),
     .top_op_top(net_4953[0:7]), .tnr_op_top(net_5958[0:7]),
     .tnr_op_bot(net_4945[0:7]), .tnl_op_top(net_6976[0:7]),
     .tnl_op_bot(net_6948[0:7]), .rgt_op_top(net_4945[0:7]),
     .rgt_op_bot(net_5013[0:7]), .reset_b_top(reset_b[111:96]),
     .reset_b_bot(reset_b[95:80]), .prog(prog),
     .pgate_top(pgate[111:96]), .pgate_bot(pgate[95:80]),
     .lft_op_top(net_6948[0:7]), .lft_op_bot(net_5632[0:7]),
     .bm_wdummymux_en_i(net_5066), .bot_op_bot(net_5912[0:7]),
     .bnr_op_top(net_5013[0:7]), .bnr_op_bot(net_4970[0:7]),
     .bnl_op_top(net_5632[0:7]), .bnl_op_bot(net_5604[0:7]),
     .sp12_v_t_top(net_4973[0:23]), .sp12_v_b_bot(net_5041[0:23]),
     .bm_init_i(net_5061), .sp12_h_r_top(net_4976[0:23]),
     .sp12_h_r_bot(net_4977[0:23]), .sp12_h_l_top(net_5756[0:23]),
     .sp12_h_l_bot(net_5896[0:23]), .sp4_v_t_top(net_7132[0:47]),
     .sp4_v_b_top(net_5760[0:47]), .sp4_v_b_bot(net_5900[0:47]),
     .sp4_r_v_b_top(net_4983[0:47]), .sp4_r_v_b_bot(net_4984[0:47]),
     .sp4_h_r_top(net_4985[0:47]), .sp4_h_r_bot(net_4986[0:47]),
     .sp4_h_l_top(net_5757[0:47]), .sp4_h_l_bot(net_5897[0:47]),
     .bm_sdi_o(net_4989[0:1]), .bm_sclkrw_o(net_4990[0:1]),
     .bl(bl[1023:982]), .bm_rcapmux_en_i(net_5060),
     .bm_sa_i(net_5062[0:7]), .bm_sclk_i(net_5063),
     .bm_sclkrw_i(net_5052[0:1]), .bm_sreb_i(net_5064),
     .bm_sweb_i(net_5065[0:1]), .bm_rcapmux_en_o(net_4998),
     .bm_init_o(net_4999), .bm_sa_o(net_5000[0:7]),
     .bm_sclk_o(net_5001), .bm_sreb_o(net_5002),
     .bm_sweb_o(net_5003[0:1]), .bm_wdummymux_en_o(net_5004),
     .bm_sdi_i(net_5051[0:1]), .bm_sdo_i(net_5006[0:1]),
     .bm_sdo_o(net_5068[0:1]));
bram_4kprouting_bbank I_bram1903 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_top(vdd_cntl[79:64]), .vdd_cntl_bot(vdd_cntl[63:48]),
     .bnr_op_top(net_5510[0:7]), .rgt_op_top(net_4970[0:7]),
     .tnr_op_top(net_5013[0:7]), .tnr_op_bot(net_4970[0:7]),
     .sp12_h_r_top(net_5015[0:23]), .sp12_h_r_bot(net_5016[0:23]),
     .sp4_h_r_bot(net_5017[0:47]), .sp4_h_r_top(net_5018[0:47]),
     .rgt_op_bot(net_5510[0:7]), .sp4_r_v_b_top(net_5020[0:47]),
     .sp4_r_v_b_bot(net_5021[0:47]), .bnr_op_bot(net_5022[0:7]),
     .slf_op_top(net_5912[0:7]), .slf_op_bot(net_4829[0:7]),
     .wl_top(wl[79:64]), .wl_bot(wl[63:48]),
     .top_op_top(net_7902[0:7]), .tnl_op_top(net_5632[0:7]),
     .tnl_op_bot(net_5604[0:7]), .reset_b_top(reset_b[79:64]),
     .reset_b_bot(reset_b[63:48]), .prog(prog),
     .pgate_top(pgate[79:64]), .pgate_bot(pgate[63:48]),
     .lft_op_top(net_5604[0:7]), .lft_op_bot(net_7760[0:7]),
     .bm_wdummymux_en_i(net_4880), .bot_op_bot(net_5466[0:7]),
     .bnl_op_top(net_7760[0:7]), .bnl_op_bot(net_7732[0:7]),
     .sp12_v_t_top(net_5041[0:23]), .sp12_v_b_bot(net_4849[0:23]),
     .bm_init_i(net_4875), .sp12_h_l_top(net_7884[0:23]),
     .sp12_h_l_bot(net_7912[0:23]), .sp4_v_t_top(net_5900[0:47]),
     .sp4_v_b_top(net_7888[0:47]), .sp4_v_b_bot(net_7916[0:47]),
     .sp4_h_l_top(net_7885[0:47]), .sp4_h_l_bot(net_7913[0:47]),
     .bm_sdi_o(net_5051[0:1]), .bm_sclkrw_o(net_5052[0:1]),
     .bl(bl[1023:982]), .bm_rcapmux_en_i(net_4874),
     .bm_sa_i(net_4876[0:7]), .bm_sclk_i(net_4877),
     .bm_sclkrw_i(net_4866[0:1]), .bm_sreb_i(net_4878),
     .bm_sweb_i(net_4879[0:1]), .bm_rcapmux_en_o(net_5060),
     .bm_init_o(net_5061), .bm_sa_o(net_5062[0:7]),
     .bm_sclk_o(net_5063), .bm_sreb_o(net_5064),
     .bm_sweb_o(net_5065[0:1]), .bm_wdummymux_en_o(net_5066),
     .bm_sdi_i(net_4865[0:1]), .bm_sdo_i(net_5068[0:1]),
     .bm_sdo_o(net_4882[0:1]));
bram_4kprouting_bbankin I_bram1909 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_top(vdd_cntl[175:160]),
     .vdd_cntl_bot(vdd_cntl[159:144]), .slf_op_top(slf_op_19_10[7:0]),
     .slf_op_bot(net_7118[0:7]), .wl_top(wl[175:160]),
     .wl_bot(wl[159:144]), .top_op_top(top_op_19_10[7:0]),
     .tnr_op_top(tnr_op_19_10[7:0]), .tnr_op_bot(slf_op_20_10[7:0]),
     .tnl_op_top(tnl_op_19_10[7:0]), .tnl_op_bot(slf_op_18_10[7:0]),
     .rgt_op_top(slf_op_20_10[7:0]), .rgt_op_bot(net_4936[0:7]),
     .reset_b_top(reset_b[175:160]), .reset_b_bot(reset_b[159:144]),
     .prog(prog), .pgate_top(pgate[175:160]),
     .pgate_bot(pgate[159:144]), .lft_op_top(slf_op_18_10[7:0]),
     .lft_op_bot(net_6248[0:7]), .bm_wdummymux_en_i(net_4930),
     .bot_op_bot(net_6528[0:7]), .bnr_op_top(net_4936[0:7]),
     .bnr_op_bot(net_5094[0:7]), .bnl_op_top(net_6248[0:7]),
     .bnl_op_bot(net_6220[0:7]), .sp12_v_t_top(sp12_v_t_19_10[23:0]),
     .sp12_v_b_bot(net_4905[0:23]), .bm_init_i(net_4925),
     .sp12_h_r_top(net_5100[0:23]), .sp12_h_r_bot(net_5101[0:23]),
     .sp12_h_l_top(net_6372[0:23]), .sp12_h_l_bot(net_6512[0:23]),
     .sp4_v_t_top(sp4_v_t_19_10[47:0]), .sp4_v_b_top(net_6376[0:47]),
     .sp4_v_b_bot(net_6516[0:47]), .sp4_r_v_b_top(net_5107[0:47]),
     .sp4_r_v_b_bot(net_5108[0:47]), .sp4_h_r_top(net_5109[0:47]),
     .sp4_h_r_bot(net_5110[0:47]), .sp4_h_l_top(net_6373[0:47]),
     .sp4_h_l_bot(net_6513[0:47]), .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(net_4924), .bm_sa_i(net_4926[0:7]),
     .bm_sclk_i(net_4927), .bm_sclkrw_i(net_4916[0:1]),
     .bm_sreb_i(net_4928), .bm_sweb_i(net_4929[0:1]),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sdi_i(net_4915[0:1]),
     .bm_sdo_i(bm_sdo_i[1:0]), .bm_sdo_o(net_4932[0:1]));
ltile4rev I_17_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5134), .lft_op(net_5240[0:7]),
     .sp12_h_l(net_5280[0:23]), .sp4_h_l(net_5281[0:47]),
     .sp4_v_b(net_5284[0:47]), .sp12_v_b(net_4539[0:23]),
     .sp12_h_r(net_5140[0:23]), .sp4_h_r(net_5141[0:47]),
     .sp12_v_t(net_5142[0:23]), .sp4_v_t(net_5256[0:47]),
     .sp4_r_v_b(net_5144[0:47]), .wl(wl[31:16]),
     .top_op(net_7872[0:7]), .rgt_op(net_5184[0:7]),
     .bot_op({io_b_32[3], io_b_32[2], io_b_32[1], io_b_32[0],
     io_b_32[3], io_b_32[2], io_b_32[1], io_b_32[0]}),
     .bl(bl[927:874]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_17[7:0]), .carry_in(net_5152), .purst(purst),
     .slf_op(net_5268[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_34[3],
     io_b_34[2], io_b_34[1], io_b_34[0], io_b_34[3], io_b_34[2],
     io_b_34[1], io_b_34[0]}), .bnl_op({io_b_30[3], io_b_30[2],
     io_b_30[1], io_b_30[0], io_b_30[3], io_b_30[2], io_b_30[1],
     io_b_30[0]}), .tnr_op(net_7732[0:7]), .tnl_op(net_7788[0:7]));
ltile4rev I_17_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5162), .lft_op(net_7788[0:7]),
     .sp12_h_l(net_5252[0:23]), .sp4_h_l(net_5253[0:47]),
     .sp4_v_b(net_5256[0:47]), .sp12_v_b(net_5142[0:23]),
     .sp12_h_r(net_5168[0:23]), .sp4_h_r(net_5169[0:47]),
     .sp12_v_t(net_5170[0:23]), .sp4_v_t(net_7860[0:47]),
     .sp4_r_v_b(net_5172[0:47]), .wl(wl[47:32]),
     .top_op(net_7844[0:7]), .rgt_op(net_7732[0:7]),
     .bot_op(net_5268[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_5134), .purst(purst), .slf_op(net_7872[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_5184[0:7]),
     .bnl_op(net_5240[0:7]), .tnr_op(net_7760[0:7]),
     .tnl_op(net_7816[0:7]));
ltile4rev I_15_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5190), .lft_op(net_5408[0:7]),
     .sp12_h_l(net_5336[0:23]), .sp4_h_l(net_5337[0:47]),
     .sp4_v_b(net_5340[0:47]), .sp12_v_b(net_4607[0:23]),
     .sp12_h_r(net_5196[0:23]), .sp4_h_r(net_5197[0:47]),
     .sp12_v_t(net_5198[0:23]), .sp4_v_t(net_5368[0:47]),
     .sp4_r_v_b(net_5200[0:47]), .wl(wl[31:16]),
     .top_op(net_7704[0:7]), .rgt_op(net_5240[0:7]),
     .bot_op({io_b_28[3], io_b_28[2], io_b_28[1], io_b_28[0],
     io_b_28[3], io_b_28[2], io_b_28[1], io_b_28[0]}),
     .bl(bl[819:766]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_15[7:0]), .carry_in(net_5208), .purst(purst),
     .slf_op(net_5380[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_30[3],
     io_b_30[2], io_b_30[1], io_b_30[0], io_b_30[3], io_b_30[2],
     io_b_30[1], io_b_30[0]}), .bnl_op({io_b_26[3], io_b_26[2],
     io_b_26[1], io_b_26[0], io_b_26[3], io_b_26[2], io_b_26[1],
     io_b_26[0]}), .tnr_op(net_7788[0:7]), .tnl_op(net_7620[0:7]));
ltile4rev I_15_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5218), .lft_op(net_7620[0:7]),
     .sp12_h_l(net_5364[0:23]), .sp4_h_l(net_5365[0:47]),
     .sp4_v_b(net_5368[0:47]), .sp12_v_b(net_5198[0:23]),
     .sp12_h_r(net_5224[0:23]), .sp4_h_r(net_5225[0:47]),
     .sp12_v_t(net_5226[0:23]), .sp4_v_t(net_7692[0:47]),
     .sp4_r_v_b(net_5228[0:47]), .wl(wl[47:32]),
     .top_op(net_7676[0:7]), .rgt_op(net_7788[0:7]),
     .bot_op(net_5380[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_5190), .purst(purst), .slf_op(net_7704[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_5240[0:7]),
     .bnl_op(net_5408[0:7]), .tnr_op(net_7816[0:7]),
     .tnl_op(net_7648[0:7]));
ltile4rev I_16_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5246), .lft_op(net_7704[0:7]),
     .sp12_h_l(net_5224[0:23]), .sp4_h_l(net_5225[0:47]),
     .sp4_v_b(net_5228[0:47]), .sp12_v_b(net_5282[0:23]),
     .sp12_h_r(net_5252[0:23]), .sp4_h_r(net_5253[0:47]),
     .sp12_v_t(net_5254[0:23]), .sp4_v_t(net_7776[0:47]),
     .sp4_r_v_b(net_5256[0:47]), .wl(wl[47:32]),
     .top_op(net_7816[0:7]), .rgt_op(net_7872[0:7]),
     .bot_op(net_5240[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_5274), .purst(purst), .slf_op(net_7788[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_5268[0:7]),
     .bnl_op(net_5380[0:7]), .tnr_op(net_7844[0:7]),
     .tnl_op(net_7676[0:7]));
ltile4rev I_16_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5274), .lft_op(net_5380[0:7]),
     .sp12_h_l(net_5196[0:23]), .sp4_h_l(net_5197[0:47]),
     .sp4_v_b(net_5200[0:47]), .sp12_v_b(net_4573[0:23]),
     .sp12_h_r(net_5280[0:23]), .sp4_h_r(net_5281[0:47]),
     .sp12_v_t(net_5282[0:23]), .sp4_v_t(net_5228[0:47]),
     .sp4_r_v_b(net_5284[0:47]), .wl(wl[31:16]),
     .top_op(net_7788[0:7]), .rgt_op(net_5268[0:7]),
     .bot_op({io_b_30[3], io_b_30[2], io_b_30[1], io_b_30[0],
     io_b_30[3], io_b_30[2], io_b_30[1], io_b_30[0]}),
     .bl(bl[873:820]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_16[7:0]), .carry_in(net_5292), .purst(purst),
     .slf_op(net_5240[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_32[3],
     io_b_32[2], io_b_32[1], io_b_32[0], io_b_32[3], io_b_32[2],
     io_b_32[1], io_b_32[0]}), .bnl_op({io_b_28[3], io_b_28[2],
     io_b_28[1], io_b_28[0], io_b_28[3], io_b_28[2], io_b_28[1],
     io_b_28[0]}), .tnr_op(net_7872[0:7]), .tnl_op(net_7704[0:7]));
ltile4rev I_18_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5302), .lft_op(net_7872[0:7]),
     .sp12_h_l(net_5168[0:23]), .sp4_h_l(net_5169[0:47]),
     .sp4_v_b(net_5172[0:47]), .sp12_v_b(net_5450[0:23]),
     .sp12_h_r(net_5308[0:23]), .sp4_h_r(net_5309[0:47]),
     .sp12_v_t(net_5310[0:23]), .sp4_v_t(net_7720[0:47]),
     .sp4_r_v_b(net_5312[0:47]), .wl(wl[47:32]),
     .top_op(net_7760[0:7]), .rgt_op(net_5466[0:7]),
     .bot_op(net_5184[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_5442), .purst(purst), .slf_op(net_7732[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_4510[0:7]),
     .bnl_op(net_5268[0:7]), .tnr_op(net_4829[0:7]),
     .tnl_op(net_7844[0:7]));
ltile4rev I_14_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5330), .lft_op(slf_op_13_01[7:0]),
     .sp12_h_l(net_5420[0:23]), .sp4_h_l(net_5421[0:47]),
     .sp4_v_b(net_5424[0:47]), .sp12_v_b(net_4641[0:23]),
     .sp12_h_r(net_5336[0:23]), .sp4_h_r(net_5337[0:47]),
     .sp12_v_t(net_5338[0:23]), .sp4_v_t(net_5396[0:47]),
     .sp4_r_v_b(net_5340[0:47]), .wl(wl[31:16]),
     .top_op(net_7620[0:7]), .rgt_op(net_5380[0:7]),
     .bot_op({io_b_26[3], io_b_26[2], io_b_26[1], io_b_26[0],
     io_b_26[3], io_b_26[2], io_b_26[1], io_b_26[0]}),
     .bl(bl[765:712]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_14[7:0]), .carry_in(net_5348), .purst(purst),
     .slf_op(net_5408[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_28[3],
     io_b_28[2], io_b_28[1], io_b_28[0], io_b_28[3], io_b_28[2],
     io_b_28[1], io_b_28[0]}), .bnl_op({slf_op_13_00[3],
     slf_op_13_00[2], slf_op_13_00[1], slf_op_13_00[0],
     slf_op_13_00[3], slf_op_13_00[2], slf_op_13_00[1],
     slf_op_13_00[0]}), .tnr_op(net_7704[0:7]),
     .tnl_op(slf_op_13_02[7:0]));
ltile4rev I_14_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5358), .lft_op(slf_op_13_02[7:0]),
     .sp12_h_l(net_5392[0:23]), .sp4_h_l(net_5393[0:47]),
     .sp4_v_b(net_5396[0:47]), .sp12_v_b(net_5338[0:23]),
     .sp12_h_r(net_5364[0:23]), .sp4_h_r(net_5365[0:47]),
     .sp12_v_t(net_5366[0:23]), .sp4_v_t(net_7608[0:47]),
     .sp4_r_v_b(net_5368[0:47]), .wl(wl[47:32]),
     .top_op(net_7648[0:7]), .rgt_op(net_7704[0:7]),
     .bot_op(net_5408[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_5330), .purst(purst), .slf_op(net_7620[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_5380[0:7]),
     .bnl_op(slf_op_13_01[7:0]), .tnr_op(net_7676[0:7]),
     .tnl_op(slf_op_13_03[7:0]));
ltile4rev I_13_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5386), .lft_op(lft_op_13_02[7:0]),
     .sp12_h_l(sp12_h_l_13_02[23:0]), .sp4_h_l(sp4_h_l_13_02[47:0]),
     .sp4_v_b(sp4_v_b_13_02[47:0]), .sp12_v_b(net_5422[0:23]),
     .sp12_h_r(net_5392[0:23]), .sp4_h_r(net_5393[0:47]),
     .sp12_v_t(net_5394[0:23]), .sp4_v_t(sp4_v_b_13_03[47:0]),
     .sp4_r_v_b(net_5396[0:47]), .wl(wl[47:32]),
     .top_op(slf_op_13_03[7:0]), .rgt_op(net_7620[0:7]),
     .bot_op(slf_op_13_01[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5414), .purst(purst), .slf_op(slf_op_13_02[7:0]),
     .pgate(pgate[47:32]), .bnr_op(net_5408[0:7]),
     .bnl_op(lft_op_13_01[7:0]), .tnr_op(net_7648[0:7]),
     .tnl_op(lft_op_13_03[7:0]));
ltile4rev I_13_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5414), .lft_op(lft_op_13_01[7:0]),
     .sp12_h_l(sp12_h_l_13_01[23:0]), .sp4_h_l(sp4_h_l_13_01[47:0]),
     .sp4_v_b(sp4_v_b_13_01[47:0]), .sp12_v_b(net_4675[0:23]),
     .sp12_h_r(net_5420[0:23]), .sp4_h_r(net_5421[0:47]),
     .sp12_v_t(net_5422[0:23]), .sp4_v_t(sp4_v_b_13_02[47:0]),
     .sp4_r_v_b(net_5424[0:47]), .wl(wl[31:16]),
     .top_op(slf_op_13_02[7:0]), .rgt_op(net_5408[0:7]),
     .bot_op({slf_op_13_00[3], slf_op_13_00[2], slf_op_13_00[1],
     slf_op_13_00[0], slf_op_13_00[3], slf_op_13_00[2],
     slf_op_13_00[1], slf_op_13_00[0]}), .bl(bl[711:658]),
     .reset_b(reset_b[31:16]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5432), .purst(purst), .slf_op(slf_op_13_01[7:0]),
     .pgate(pgate[31:16]), .bnr_op({io_b_26[3], io_b_26[2], io_b_26[1],
     io_b_26[0], io_b_26[3], io_b_26[2], io_b_26[1], io_b_26[0]}),
     .bnl_op({bnl_op_13_01[3], bnl_op_13_01[2], bnl_op_13_01[1],
     bnl_op_13_01[0], bnl_op_13_01[3], bnl_op_13_01[2],
     bnl_op_13_01[1], bnl_op_13_01[0]}), .tnr_op(net_7620[0:7]),
     .tnl_op(lft_op_13_02[7:0]));
ltile4rev I_18_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5442), .lft_op(net_5268[0:7]),
     .sp12_h_l(net_5140[0:23]), .sp4_h_l(net_5141[0:47]),
     .sp4_v_b(net_5144[0:47]), .sp12_v_b(net_4505[0:23]),
     .sp12_h_r(net_5448[0:23]), .sp4_h_r(net_5449[0:47]),
     .sp12_v_t(net_5450[0:23]), .sp4_v_t(net_5172[0:47]),
     .sp4_r_v_b(net_5452[0:47]), .wl(wl[31:16]),
     .top_op(net_7732[0:7]), .rgt_op(net_4510[0:7]),
     .bot_op({io_b_34[3], io_b_34[2], io_b_34[1], io_b_34[0],
     io_b_34[3], io_b_34[2], io_b_34[1], io_b_34[0]}),
     .bl(bl[981:928]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_18[7:0]), .carry_in(net_5460), .purst(purst),
     .slf_op(net_5184[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_36[3],
     io_b_36[2], io_b_36[1], io_b_36[0], io_b_36[3], io_b_36[2],
     io_b_36[1], io_b_36[0]}), .bnl_op({io_b_32[3], io_b_32[2],
     io_b_32[1], io_b_32[0], io_b_32[3], io_b_32[2], io_b_32[1],
     io_b_32[0]}), .tnr_op(net_5466[0:7]), .tnl_op(net_7872[0:7]));
ltile4rev I_20_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5470), .lft_op(net_4510[0:7]),
     .sp12_h_l(net_4853[0:23]), .sp4_h_l(net_4862[0:47]),
     .sp4_v_b(net_4860[0:47]), .sp12_v_b(net_4471[0:23]),
     .sp12_h_r(net_5476[0:23]), .sp4_h_r(net_5477[0:47]),
     .sp12_v_t(net_5478[0:23]), .sp4_v_t(net_4859[0:47]),
     .sp4_r_v_b(net_5480[0:47]), .wl(wl[31:16]),
     .top_op(net_5022[0:7]), .rgt_op(net_5520[0:7]),
     .bot_op({io_b_38[3], io_b_38[2], io_b_38[1], io_b_38[0],
     io_b_38[3], io_b_38[2], io_b_38[1], io_b_38[0]}),
     .bl(bl[1077:1024]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_20[7:0]), .carry_in(net_5488), .purst(purst),
     .slf_op(net_4748[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_40[3],
     io_b_40[2], io_b_40[1], io_b_40[0], io_b_40[3], io_b_40[2],
     io_b_40[1], io_b_40[0]}), .bnl_op({io_b_36[3], io_b_36[2],
     io_b_36[1], io_b_36[0], io_b_36[3], io_b_36[2], io_b_36[1],
     io_b_36[0]}), .tnr_op(net_7956[0:7]), .tnl_op(net_5466[0:7]));
ltile4rev I_20_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5498), .lft_op(net_5466[0:7]),
     .sp12_h_l(net_4852[0:23]), .sp4_h_l(net_4861[0:47]),
     .sp4_v_b(net_4859[0:47]), .sp12_v_b(net_5478[0:23]),
     .sp12_h_r(net_5504[0:23]), .sp4_h_r(net_5505[0:47]),
     .sp12_v_t(net_5506[0:23]), .sp4_v_t(net_5021[0:47]),
     .sp4_r_v_b(net_5508[0:47]), .wl(wl[47:32]),
     .top_op(net_5510[0:7]), .rgt_op(net_7956[0:7]),
     .bot_op(net_4748[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_5470), .purst(purst), .slf_op(net_5022[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_5520[0:7]),
     .bnl_op(net_4510[0:7]), .tnr_op(net_7984[0:7]),
     .tnl_op(net_4829[0:7]));
ltile4rev I_21_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_5526), .lft_op(net_5022[0:7]),
     .sp12_h_l(net_5504[0:23]), .sp4_h_l(net_5505[0:47]),
     .sp4_v_b(net_5508[0:47]), .sp12_v_b(net_5562[0:23]),
     .sp12_h_r(net_5532[0:23]), .sp4_h_r(net_5533[0:47]),
     .sp12_v_t(net_5534[0:23]), .sp4_v_t(net_7944[0:47]),
     .sp4_r_v_b(net_5536[0:47]), .wl(wl[47:32]),
     .top_op(net_7984[0:7]), .rgt_op(net_8040[0:7]),
     .bot_op(net_5520[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_5554), .purst(purst), .slf_op(net_7956[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_5548[0:7]),
     .bnl_op(net_4748[0:7]), .tnr_op(net_8012[0:7]),
     .tnl_op(net_5510[0:7]));
ltile4rev I_21_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_5554), .lft_op(net_4748[0:7]),
     .sp12_h_l(net_5476[0:23]), .sp4_h_l(net_5477[0:47]),
     .sp4_v_b(net_5480[0:47]), .sp12_v_b(net_4437[0:23]),
     .sp12_h_r(net_5560[0:23]), .sp4_h_r(net_5561[0:47]),
     .sp12_v_t(net_5562[0:23]), .sp4_v_t(net_5508[0:47]),
     .sp4_r_v_b(net_5564[0:47]), .wl(wl[31:16]),
     .top_op(net_7956[0:7]), .rgt_op(net_5548[0:7]),
     .bot_op({io_b_40[3], io_b_40[2], io_b_40[1], io_b_40[0],
     io_b_40[3], io_b_40[2], io_b_40[1], io_b_40[0]}),
     .bl(bl[1131:1078]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_21[7:0]), .carry_in(net_5572), .purst(purst),
     .slf_op(net_5520[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_42[3],
     io_b_42[2], io_b_42[1], io_b_42[0], io_b_42[3], io_b_42[2],
     io_b_42[1], io_b_42[0]}), .bnl_op({io_b_38[3], io_b_38[2],
     io_b_38[1], io_b_38[0], io_b_38[3], io_b_38[2], io_b_38[1],
     io_b_38[0]}), .tnr_op(net_8040[0:7]), .tnl_op(net_5022[0:7]));
ltile4rev I_17_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_5582), .lft_op(net_5688[0:7]),
     .sp12_h_l(net_5728[0:23]), .sp4_h_l(net_5729[0:47]),
     .sp4_v_b(net_5732[0:47]), .sp12_v_b(net_7746[0:23]),
     .sp12_h_r(net_5588[0:23]), .sp4_h_r(net_5589[0:47]),
     .sp12_v_t(net_5590[0:23]), .sp4_v_t(net_5704[0:47]),
     .sp4_r_v_b(net_5592[0:47]), .wl(wl[95:80]),
     .top_op(net_7088[0:7]), .rgt_op(net_5632[0:7]),
     .bot_op(net_5744[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_7738), .purst(purst), .slf_op(net_5716[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_5604[0:7]),
     .bnl_op(net_5660[0:7]), .tnr_op(net_6948[0:7]),
     .tnl_op(net_7004[0:7]));
ltile4rev I_17_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5610), .lft_op(net_7004[0:7]),
     .sp12_h_l(net_5700[0:23]), .sp4_h_l(net_5701[0:47]),
     .sp4_v_b(net_5704[0:47]), .sp12_v_b(net_5590[0:23]),
     .sp12_h_r(net_5616[0:23]), .sp4_h_r(net_5617[0:47]),
     .sp12_v_t(net_5618[0:23]), .sp4_v_t(net_7076[0:47]),
     .sp4_r_v_b(net_5620[0:47]), .wl(wl[111:96]),
     .top_op(net_7060[0:7]), .rgt_op(net_6948[0:7]),
     .bot_op(net_5716[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_5582), .purst(purst), .slf_op(net_7088[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_5632[0:7]),
     .bnl_op(net_5688[0:7]), .tnr_op(net_6976[0:7]),
     .tnl_op(net_7032[0:7]));
ltile4rev I_15_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_5638), .lft_op(net_5856[0:7]),
     .sp12_h_l(net_5784[0:23]), .sp4_h_l(net_5785[0:47]),
     .sp4_v_b(net_5788[0:47]), .sp12_v_b(net_7802[0:23]),
     .sp12_h_r(net_5644[0:23]), .sp4_h_r(net_5645[0:47]),
     .sp12_v_t(net_5646[0:23]), .sp4_v_t(net_5816[0:47]),
     .sp4_r_v_b(net_5648[0:47]), .wl(wl[95:80]),
     .top_op(net_6920[0:7]), .rgt_op(net_5688[0:7]),
     .bot_op(net_5800[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_7794), .purst(purst), .slf_op(net_5828[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_5660[0:7]),
     .bnl_op(net_5884[0:7]), .tnr_op(net_7004[0:7]),
     .tnl_op(net_6836[0:7]));
ltile4rev I_15_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5666), .lft_op(net_6836[0:7]),
     .sp12_h_l(net_5812[0:23]), .sp4_h_l(net_5813[0:47]),
     .sp4_v_b(net_5816[0:47]), .sp12_v_b(net_5646[0:23]),
     .sp12_h_r(net_5672[0:23]), .sp4_h_r(net_5673[0:47]),
     .sp12_v_t(net_5674[0:23]), .sp4_v_t(net_6908[0:47]),
     .sp4_r_v_b(net_5676[0:47]), .wl(wl[111:96]),
     .top_op(net_6892[0:7]), .rgt_op(net_7004[0:7]),
     .bot_op(net_5828[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_5638), .purst(purst), .slf_op(net_6920[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_5688[0:7]),
     .bnl_op(net_5856[0:7]), .tnr_op(net_7032[0:7]),
     .tnl_op(net_6864[0:7]));
ltile4rev I_16_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5694), .lft_op(net_6920[0:7]),
     .sp12_h_l(net_5672[0:23]), .sp4_h_l(net_5673[0:47]),
     .sp4_v_b(net_5676[0:47]), .sp12_v_b(net_5730[0:23]),
     .sp12_h_r(net_5700[0:23]), .sp4_h_r(net_5701[0:47]),
     .sp12_v_t(net_5702[0:23]), .sp4_v_t(net_6992[0:47]),
     .sp4_r_v_b(net_5704[0:47]), .wl(wl[111:96]),
     .top_op(net_7032[0:7]), .rgt_op(net_7088[0:7]),
     .bot_op(net_5688[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_5722), .purst(purst), .slf_op(net_7004[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_5716[0:7]),
     .bnl_op(net_5828[0:7]), .tnr_op(net_7060[0:7]),
     .tnl_op(net_6892[0:7]));
ltile4rev I_16_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_5722), .lft_op(net_5828[0:7]),
     .sp12_h_l(net_5644[0:23]), .sp4_h_l(net_5645[0:47]),
     .sp4_v_b(net_5648[0:47]), .sp12_v_b(net_7830[0:23]),
     .sp12_h_r(net_5728[0:23]), .sp4_h_r(net_5729[0:47]),
     .sp12_v_t(net_5730[0:23]), .sp4_v_t(net_5676[0:47]),
     .sp4_r_v_b(net_5732[0:47]), .wl(wl[95:80]),
     .top_op(net_7004[0:7]), .rgt_op(net_5716[0:7]),
     .bot_op(net_5660[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_7822), .purst(purst), .slf_op(net_5688[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_5744[0:7]),
     .bnl_op(net_5800[0:7]), .tnr_op(net_7088[0:7]),
     .tnl_op(net_6920[0:7]));
ltile4rev I_18_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5750), .lft_op(net_7088[0:7]),
     .sp12_h_l(net_5616[0:23]), .sp4_h_l(net_5617[0:47]),
     .sp4_v_b(net_5620[0:47]), .sp12_v_b(net_5898[0:23]),
     .sp12_h_r(net_5756[0:23]), .sp4_h_r(net_5757[0:47]),
     .sp12_v_t(net_5758[0:23]), .sp4_v_t(net_6936[0:47]),
     .sp4_r_v_b(net_5760[0:47]), .wl(wl[111:96]),
     .top_op(net_6976[0:7]), .rgt_op(net_7144[0:7]),
     .bot_op(net_5632[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_5890), .purst(purst), .slf_op(net_6948[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_7902[0:7]),
     .bnl_op(net_5716[0:7]), .tnr_op(net_4953[0:7]),
     .tnl_op(net_7060[0:7]));
ltile4rev I_14_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_5778), .lft_op(slf_op_13_05[7:0]),
     .sp12_h_l(net_5868[0:23]), .sp4_h_l(net_5869[0:47]),
     .sp4_v_b(net_5872[0:47]), .sp12_v_b(net_7662[0:23]),
     .sp12_h_r(net_5784[0:23]), .sp4_h_r(net_5785[0:47]),
     .sp12_v_t(net_5786[0:23]), .sp4_v_t(net_5844[0:47]),
     .sp4_r_v_b(net_5788[0:47]), .wl(wl[95:80]),
     .top_op(net_6836[0:7]), .rgt_op(net_5828[0:7]),
     .bot_op(net_5884[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_7654), .purst(purst), .slf_op(net_5856[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_5800[0:7]),
     .bnl_op(slf_op_13_04[7:0]), .tnr_op(net_6920[0:7]),
     .tnl_op(slf_op_13_06[7:0]));
ltile4rev I_14_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5806), .lft_op(slf_op_13_06[7:0]),
     .sp12_h_l(net_5840[0:23]), .sp4_h_l(net_5841[0:47]),
     .sp4_v_b(net_5844[0:47]), .sp12_v_b(net_5786[0:23]),
     .sp12_h_r(net_5812[0:23]), .sp4_h_r(net_5813[0:47]),
     .sp12_v_t(net_5814[0:23]), .sp4_v_t(net_6824[0:47]),
     .sp4_r_v_b(net_5816[0:47]), .wl(wl[111:96]),
     .top_op(net_6864[0:7]), .rgt_op(net_6920[0:7]),
     .bot_op(net_5856[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_5778), .purst(purst), .slf_op(net_6836[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_5828[0:7]),
     .bnl_op(slf_op_13_05[7:0]), .tnr_op(net_6892[0:7]),
     .tnl_op(slf_op_13_07[7:0]));
ltile4rev I_13_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5834), .lft_op(lft_op_13_06[7:0]),
     .sp12_h_l(sp12_h_l_13_06[23:0]), .sp4_h_l(sp4_h_l_13_06[47:0]),
     .sp4_v_b(sp4_v_b_13_06[47:0]), .sp12_v_b(net_5870[0:23]),
     .sp12_h_r(net_5840[0:23]), .sp4_h_r(net_5841[0:47]),
     .sp12_v_t(net_5842[0:23]), .sp4_v_t(sp4_v_b_13_07[47:0]),
     .sp4_r_v_b(net_5844[0:47]), .wl(wl[111:96]),
     .top_op(slf_op_13_07[7:0]), .rgt_op(net_6836[0:7]),
     .bot_op(slf_op_13_05[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5862), .purst(purst), .slf_op(slf_op_13_06[7:0]),
     .pgate(pgate[111:96]), .bnr_op(net_5856[0:7]),
     .bnl_op(lft_op_13_05[7:0]), .tnr_op(net_6864[0:7]),
     .tnl_op(lft_op_13_07[7:0]));
ltile4rev I_13_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_5862), .lft_op(lft_op_13_05[7:0]),
     .sp12_h_l(sp12_h_l_13_05[23:0]), .sp4_h_l(sp4_h_l_13_05[47:0]),
     .sp4_v_b(sp4_v_b_13_05[47:0]), .sp12_v_b(net_7634[0:23]),
     .sp12_h_r(net_5868[0:23]), .sp4_h_r(net_5869[0:47]),
     .sp12_v_t(net_5870[0:23]), .sp4_v_t(sp4_v_b_13_06[47:0]),
     .sp4_r_v_b(net_5872[0:47]), .wl(wl[95:80]),
     .top_op(slf_op_13_06[7:0]), .rgt_op(net_5856[0:7]),
     .bot_op(slf_op_13_04[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_7626), .purst(purst), .slf_op(slf_op_13_05[7:0]),
     .pgate(pgate[95:80]), .bnr_op(net_5884[0:7]),
     .bnl_op(lft_op_13_04[7:0]), .tnr_op(net_6836[0:7]),
     .tnl_op(lft_op_13_06[7:0]));
ltile4rev I_18_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_5890), .lft_op(net_5716[0:7]),
     .sp12_h_l(net_5588[0:23]), .sp4_h_l(net_5589[0:47]),
     .sp4_v_b(net_5592[0:47]), .sp12_v_b(net_7886[0:23]),
     .sp12_h_r(net_5896[0:23]), .sp4_h_r(net_5897[0:47]),
     .sp12_v_t(net_5898[0:23]), .sp4_v_t(net_5620[0:47]),
     .sp4_r_v_b(net_5900[0:47]), .wl(wl[95:80]),
     .top_op(net_6948[0:7]), .rgt_op(net_7902[0:7]),
     .bot_op(net_5604[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_7878), .purst(purst), .slf_op(net_5632[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_5912[0:7]),
     .bnl_op(net_5744[0:7]), .tnr_op(net_7144[0:7]),
     .tnl_op(net_7088[0:7]));
ltile4rev I_20_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_5918), .lft_op(net_7902[0:7]),
     .sp12_h_l(net_4977[0:23]), .sp4_h_l(net_4986[0:47]),
     .sp4_v_b(net_4984[0:47]), .sp12_v_b(net_7970[0:23]),
     .sp12_h_r(net_5924[0:23]), .sp4_h_r(net_5925[0:47]),
     .sp12_v_t(net_5926[0:23]), .sp4_v_t(net_4983[0:47]),
     .sp4_r_v_b(net_5928[0:47]), .wl(wl[95:80]),
     .top_op(net_4945[0:7]), .rgt_op(net_5968[0:7]),
     .bot_op(net_4970[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_7962), .purst(purst), .slf_op(net_5013[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_5940[0:7]),
     .bnl_op(net_5912[0:7]), .tnr_op(net_7172[0:7]),
     .tnl_op(net_7144[0:7]));
ltile4rev I_20_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5946), .lft_op(net_7144[0:7]),
     .sp12_h_l(net_4976[0:23]), .sp4_h_l(net_4985[0:47]),
     .sp4_v_b(net_4983[0:47]), .sp12_v_b(net_5926[0:23]),
     .sp12_h_r(net_5952[0:23]), .sp4_h_r(net_5953[0:47]),
     .sp12_v_t(net_5954[0:23]), .sp4_v_t(net_4944[0:47]),
     .sp4_r_v_b(net_5956[0:47]), .wl(wl[111:96]),
     .top_op(net_5958[0:7]), .rgt_op(net_7172[0:7]),
     .bot_op(net_5013[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_5918), .purst(purst), .slf_op(net_4945[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_5968[0:7]),
     .bnl_op(net_7902[0:7]), .tnr_op(net_7200[0:7]),
     .tnl_op(net_4953[0:7]));
ltile4rev I_21_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_5974), .lft_op(net_4945[0:7]),
     .sp12_h_l(net_5952[0:23]), .sp4_h_l(net_5953[0:47]),
     .sp4_v_b(net_5956[0:47]), .sp12_v_b(net_6010[0:23]),
     .sp12_h_r(net_5980[0:23]), .sp4_h_r(net_5981[0:47]),
     .sp12_v_t(net_5982[0:23]), .sp4_v_t(net_7160[0:47]),
     .sp4_r_v_b(net_5984[0:47]), .wl(wl[111:96]),
     .top_op(net_7200[0:7]), .rgt_op(net_7256[0:7]),
     .bot_op(net_5968[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_6002), .purst(purst), .slf_op(net_7172[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_5996[0:7]),
     .bnl_op(net_5013[0:7]), .tnr_op(net_7228[0:7]),
     .tnl_op(net_5958[0:7]));
ltile4rev I_21_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_6002), .lft_op(net_5013[0:7]),
     .sp12_h_l(net_5924[0:23]), .sp4_h_l(net_5925[0:47]),
     .sp4_v_b(net_5928[0:47]), .sp12_v_b(net_7998[0:23]),
     .sp12_h_r(net_6008[0:23]), .sp4_h_r(net_6009[0:47]),
     .sp12_v_t(net_6010[0:23]), .sp4_v_t(net_5956[0:47]),
     .sp4_r_v_b(net_6012[0:47]), .wl(wl[95:80]),
     .top_op(net_7172[0:7]), .rgt_op(net_5996[0:7]),
     .bot_op(net_5940[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_7990), .purst(purst), .slf_op(net_5968[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_6024[0:7]),
     .bnl_op(net_4970[0:7]), .tnr_op(net_7256[0:7]),
     .tnl_op(net_4945[0:7]));
ltile4rev I_23_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_6030), .lft_op(net_5996[0:7]),
     .sp12_h_l(net_6092[0:23]), .sp4_h_l(net_6093[0:47]),
     .sp4_v_b(net_6096[0:47]), .sp12_v_b(net_8194[0:23]),
     .sp12_h_r(net_6036[0:23]), .sp4_h_r(net_6037[0:47]),
     .sp12_v_t(net_6038[0:23]), .sp4_v_t(net_6124[0:47]),
     .sp4_r_v_b(net_6040[0:47]), .wl(wl[95:80]),
     .top_op(net_7340[0:7]), .rgt_op(net_6192[0:7]),
     .bot_op(net_6108[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_8186), .purst(purst), .slf_op(net_6136[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_6052[0:7]),
     .bnl_op(net_6024[0:7]), .tnr_op(net_7284[0:7]),
     .tnl_op(net_7256[0:7]));
ltile4rev I_24_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_6058), .lft_op(net_7340[0:7]),
     .sp12_h_l(net_6176[0:23]), .sp4_h_l(net_6177[0:47]),
     .sp4_v_b(net_6180[0:47]), .sp12_v_b(net_6150[0:23]),
     .sp12_h_r(net_6064[0:23]), .sp4_h_r(net_6065[0:47]),
     .sp12_v_t(net_6066[0:23]), .sp4_v_t(net_7272[0:47]),
     .sp4_r_v_b(net_6068[0:47]), .wl(wl[111:96]),
     .top_op(net_7424[0:7]), .rgt_op({io_r_05[3], io_r_05[2],
     io_r_05[1], io_r_05[0], io_r_05[3], io_r_05[2], io_r_05[1],
     io_r_05[0]}), .bot_op(net_6192[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_6142), .purst(purst), .slf_op(net_7284[0:7]),
     .pgate(pgate[111:96]), .bnr_op({io_r_04[3], io_r_04[2],
     io_r_04[1], io_r_04[0], io_r_04[3], io_r_04[2], io_r_04[1],
     io_r_04[0]}), .bnl_op(net_6136[0:7]), .tnr_op({io_r_06[3],
     io_r_06[2], io_r_06[1], io_r_06[0], io_r_06[3], io_r_06[2],
     io_r_06[1], io_r_06[0]}), .tnl_op(net_7368[0:7]));
ltile4rev I_22_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_6086), .lft_op(net_5968[0:7]),
     .sp12_h_l(net_6008[0:23]), .sp4_h_l(net_6009[0:47]),
     .sp4_v_b(net_6012[0:47]), .sp12_v_b(net_8138[0:23]),
     .sp12_h_r(net_6092[0:23]), .sp4_h_r(net_6093[0:47]),
     .sp12_v_t(net_6094[0:23]), .sp4_v_t(net_5984[0:47]),
     .sp4_r_v_b(net_6096[0:47]), .wl(wl[95:80]),
     .top_op(net_7256[0:7]), .rgt_op(net_6136[0:7]),
     .bot_op(net_6024[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_8130), .purst(purst), .slf_op(net_5996[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net_6108[0:7]),
     .bnl_op(net_5940[0:7]), .tnr_op(net_7340[0:7]),
     .tnl_op(net_7172[0:7]));
ltile4rev I_22_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_6114), .lft_op(net_7172[0:7]),
     .sp12_h_l(net_5980[0:23]), .sp4_h_l(net_5981[0:47]),
     .sp4_v_b(net_5984[0:47]), .sp12_v_b(net_6094[0:23]),
     .sp12_h_r(net_6120[0:23]), .sp4_h_r(net_6121[0:47]),
     .sp12_v_t(net_6122[0:23]), .sp4_v_t(net_7244[0:47]),
     .sp4_r_v_b(net_6124[0:47]), .wl(wl[111:96]),
     .top_op(net_7228[0:7]), .rgt_op(net_7340[0:7]),
     .bot_op(net_5996[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_6086), .purst(purst), .slf_op(net_7256[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_6136[0:7]),
     .bnl_op(net_5968[0:7]), .tnr_op(net_7368[0:7]),
     .tnl_op(net_7200[0:7]));
ltile4rev I_24_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net_6142), .lft_op(net_6136[0:7]),
     .sp12_h_l(net_6036[0:23]), .sp4_h_l(net_6037[0:47]),
     .sp4_v_b(net_6040[0:47]), .sp12_v_b(net_8082[0:23]),
     .sp12_h_r(net_6148[0:23]), .sp4_h_r(net_6149[0:47]),
     .sp12_v_t(net_6150[0:23]), .sp4_v_t(net_6180[0:47]),
     .sp4_r_v_b(net_6152[0:47]), .wl(wl[95:80]),
     .top_op(net_7284[0:7]), .rgt_op({io_r_04[3], io_r_04[2],
     io_r_04[1], io_r_04[0], io_r_04[3], io_r_04[2], io_r_04[1],
     io_r_04[0]}), .bot_op(net_6052[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_8074), .purst(purst), .slf_op(net_6192[0:7]),
     .pgate(pgate[95:80]), .bnr_op({io_r_03[3], io_r_03[2], io_r_03[1],
     io_r_03[0], io_r_03[3], io_r_03[2], io_r_03[1], io_r_03[0]}),
     .bnl_op(net_6108[0:7]), .tnr_op({io_r_05[3], io_r_05[2],
     io_r_05[1], io_r_05[0], io_r_05[3], io_r_05[2], io_r_05[1],
     io_r_05[0]}), .tnl_op(net_7340[0:7]));
ltile4rev I_23_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net_6170), .lft_op(net_7256[0:7]),
     .sp12_h_l(net_6120[0:23]), .sp4_h_l(net_6121[0:47]),
     .sp4_v_b(net_6124[0:47]), .sp12_v_b(net_6038[0:23]),
     .sp12_h_r(net_6176[0:23]), .sp4_h_r(net_6177[0:47]),
     .sp12_v_t(net_6178[0:23]), .sp4_v_t(net_7328[0:47]),
     .sp4_r_v_b(net_6180[0:47]), .wl(wl[111:96]),
     .top_op(net_7368[0:7]), .rgt_op(net_7284[0:7]),
     .bot_op(net_6136[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_6030), .purst(purst), .slf_op(net_7340[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net_6192[0:7]),
     .bnl_op(net_5996[0:7]), .tnr_op(net_7424[0:7]),
     .tnl_op(net_7228[0:7]));
ltile4rev I_17_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6198), .lft_op(net_6304[0:7]),
     .sp12_h_l(net_6344[0:23]), .sp4_h_l(net_6345[0:47]),
     .sp4_v_b(net_6348[0:47]), .sp12_v_b(net_6962[0:23]),
     .sp12_h_r(net_6204[0:23]), .sp4_h_r(net_6205[0:47]),
     .sp12_v_t(net_6206[0:23]), .sp4_v_t(net_6320[0:47]),
     .sp4_r_v_b(net_6208[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_17_10[7:0]), .rgt_op(net_6248[0:7]),
     .bot_op(net_6360[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_6954), .purst(purst), .slf_op(net_6332[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6220[0:7]),
     .bnl_op(net_6276[0:7]), .tnr_op(slf_op_18_10[7:0]),
     .tnl_op(slf_op_16_10[7:0]));
ltile4rev I_17_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_17_10), .lft_op(slf_op_16_10[7:0]),
     .sp12_h_l(net_6316[0:23]), .sp4_h_l(net_6317[0:47]),
     .sp4_v_b(net_6320[0:47]), .sp12_v_b(net_6206[0:23]),
     .sp12_h_r(net_6232[0:23]), .sp4_h_r(net_6233[0:47]),
     .sp12_v_t(sp12_v_t_17_10[23:0]), .sp4_v_t(sp4_v_t_17_10[47:0]),
     .sp4_r_v_b(net_6236[0:47]), .wl(wl[175:160]),
     .top_op(top_op_17_10[7:0]), .rgt_op(slf_op_18_10[7:0]),
     .bot_op(net_6332[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_6198), .purst(purst), .slf_op(slf_op_17_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6248[0:7]),
     .bnl_op(net_6304[0:7]), .tnr_op(tnr_op_17_10[7:0]),
     .tnl_op(tnl_op_17_10[7:0]));
ltile4rev I_15_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6254), .lft_op(net_6472[0:7]),
     .sp12_h_l(net_6400[0:23]), .sp4_h_l(net_6401[0:47]),
     .sp4_v_b(net_6404[0:47]), .sp12_v_b(net_7018[0:23]),
     .sp12_h_r(net_6260[0:23]), .sp4_h_r(net_6261[0:47]),
     .sp12_v_t(net_6262[0:23]), .sp4_v_t(net_6432[0:47]),
     .sp4_r_v_b(net_6264[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_15_10[7:0]), .rgt_op(net_6304[0:7]),
     .bot_op(net_6416[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_7010), .purst(purst), .slf_op(net_6444[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6276[0:7]),
     .bnl_op(net_6500[0:7]), .tnr_op(slf_op_16_10[7:0]),
     .tnl_op(slf_op_14_10[7:0]));
ltile4rev I_15_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_15_10), .lft_op(slf_op_14_10[7:0]),
     .sp12_h_l(net_6428[0:23]), .sp4_h_l(net_6429[0:47]),
     .sp4_v_b(net_6432[0:47]), .sp12_v_b(net_6262[0:23]),
     .sp12_h_r(net_6288[0:23]), .sp4_h_r(net_6289[0:47]),
     .sp12_v_t(sp12_v_t_15_10[23:0]), .sp4_v_t(sp4_v_t_15_10[47:0]),
     .sp4_r_v_b(net_6292[0:47]), .wl(wl[175:160]),
     .top_op(top_op_15_10[7:0]), .rgt_op(slf_op_16_10[7:0]),
     .bot_op(net_6444[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_6254), .purst(purst), .slf_op(slf_op_15_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6304[0:7]),
     .bnl_op(net_6472[0:7]), .tnr_op(tnr_op_15_10[7:0]),
     .tnl_op(tnl_op_15_10[7:0]));
ltile4rev I_16_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_16_10), .lft_op(slf_op_15_10[7:0]),
     .sp12_h_l(net_6288[0:23]), .sp4_h_l(net_6289[0:47]),
     .sp4_v_b(net_6292[0:47]), .sp12_v_b(net_6346[0:23]),
     .sp12_h_r(net_6316[0:23]), .sp4_h_r(net_6317[0:47]),
     .sp12_v_t(sp12_v_t_16_10[23:0]), .sp4_v_t(sp4_v_t_16_10[47:0]),
     .sp4_r_v_b(net_6320[0:47]), .wl(wl[175:160]),
     .top_op(top_op_16_10[7:0]), .rgt_op(slf_op_17_10[7:0]),
     .bot_op(net_6304[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_6338), .purst(purst), .slf_op(slf_op_16_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6332[0:7]),
     .bnl_op(net_6444[0:7]), .tnr_op(tnr_op_16_10[7:0]),
     .tnl_op(tnl_op_16_10[7:0]));
ltile4rev I_16_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6338), .lft_op(net_6444[0:7]),
     .sp12_h_l(net_6260[0:23]), .sp4_h_l(net_6261[0:47]),
     .sp4_v_b(net_6264[0:47]), .sp12_v_b(net_7046[0:23]),
     .sp12_h_r(net_6344[0:23]), .sp4_h_r(net_6345[0:47]),
     .sp12_v_t(net_6346[0:23]), .sp4_v_t(net_6292[0:47]),
     .sp4_r_v_b(net_6348[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_16_10[7:0]), .rgt_op(net_6332[0:7]),
     .bot_op(net_6276[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_7038), .purst(purst), .slf_op(net_6304[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6360[0:7]),
     .bnl_op(net_6416[0:7]), .tnr_op(slf_op_17_10[7:0]),
     .tnl_op(slf_op_15_10[7:0]));
ltile4rev I_18_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_18_10), .lft_op(slf_op_17_10[7:0]),
     .sp12_h_l(net_6232[0:23]), .sp4_h_l(net_6233[0:47]),
     .sp4_v_b(net_6236[0:47]), .sp12_v_b(net_6514[0:23]),
     .sp12_h_r(net_6372[0:23]), .sp4_h_r(net_6373[0:47]),
     .sp12_v_t(sp12_v_t_18_10[23:0]), .sp4_v_t(sp4_v_t_18_10[47:0]),
     .sp4_r_v_b(net_6376[0:47]), .wl(wl[175:160]),
     .top_op(top_op_18_10[7:0]), .rgt_op(slf_op_19_10[7:0]),
     .bot_op(net_6248[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_6506), .purst(purst), .slf_op(slf_op_18_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_7118[0:7]),
     .bnl_op(net_6332[0:7]), .tnr_op(tnr_op_18_10[7:0]),
     .tnl_op(tnl_op_18_10[7:0]));
ltile4rev I_14_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6394), .lft_op(slf_op_13_09[7:0]),
     .sp12_h_l(net_6484[0:23]), .sp4_h_l(net_6485[0:47]),
     .sp4_v_b(net_6488[0:47]), .sp12_v_b(net_6878[0:23]),
     .sp12_h_r(net_6400[0:23]), .sp4_h_r(net_6401[0:47]),
     .sp12_v_t(net_6402[0:23]), .sp4_v_t(net_6460[0:47]),
     .sp4_r_v_b(net_6404[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_14_10[7:0]), .rgt_op(net_6444[0:7]),
     .bot_op(net_6500[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_6870), .purst(purst), .slf_op(net_6472[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6416[0:7]),
     .bnl_op(slf_op_13_08[7:0]), .tnr_op(slf_op_15_10[7:0]),
     .tnl_op(slf_op_13_10[7:0]));
ltile4rev I_14_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_14_10), .lft_op(slf_op_13_10[7:0]),
     .sp12_h_l(net_6456[0:23]), .sp4_h_l(net_6457[0:47]),
     .sp4_v_b(net_6460[0:47]), .sp12_v_b(net_6402[0:23]),
     .sp12_h_r(net_6428[0:23]), .sp4_h_r(net_6429[0:47]),
     .sp12_v_t(sp12_v_t_14_10[23:0]), .sp4_v_t(sp4_v_t_14_10[47:0]),
     .sp4_r_v_b(net_6432[0:47]), .wl(wl[175:160]),
     .top_op(top_op_14_10[7:0]), .rgt_op(slf_op_15_10[7:0]),
     .bot_op(net_6472[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_6394), .purst(purst), .slf_op(slf_op_14_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6444[0:7]),
     .bnl_op(slf_op_13_09[7:0]), .tnr_op(tnr_op_14_10[7:0]),
     .tnl_op(tnl_op_14_10[7:0]));
ltile4rev I_13_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_13_10), .lft_op(lft_op_13_10[7:0]),
     .sp12_h_l(sp12_h_l_13_10[23:0]), .sp4_h_l(sp4_h_l_13_10[47:0]),
     .sp4_v_b(sp4_v_b_13_10[47:0]), .sp12_v_b(net_6486[0:23]),
     .sp12_h_r(net_6456[0:23]), .sp4_h_r(net_6457[0:47]),
     .sp12_v_t(sp12_v_t_13_10[23:0]), .sp4_v_t(sp4_v_t_13_10[47:0]),
     .sp4_r_v_b(net_6460[0:47]), .wl(wl[175:160]),
     .top_op(top_op_13_10[7:0]), .rgt_op(slf_op_14_10[7:0]),
     .bot_op(slf_op_13_09[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_6478), .purst(purst), .slf_op(slf_op_13_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6472[0:7]),
     .bnl_op(lft_op_13_09[7:0]), .tnr_op(tnr_op_13_10[7:0]),
     .tnl_op(tnl_op_13_10[7:0]));
ltile4rev I_13_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6478), .lft_op(lft_op_13_09[7:0]),
     .sp12_h_l(sp12_h_l_13_09[23:0]), .sp4_h_l(sp4_h_l_13_09[47:0]),
     .sp4_v_b(sp4_v_b_13_09[47:0]), .sp12_v_b(net_6850[0:23]),
     .sp12_h_r(net_6484[0:23]), .sp4_h_r(net_6485[0:47]),
     .sp12_v_t(net_6486[0:23]), .sp4_v_t(sp4_v_b_13_10[47:0]),
     .sp4_r_v_b(net_6488[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_13_10[7:0]), .rgt_op(net_6472[0:7]),
     .bot_op(slf_op_13_08[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_6842), .purst(purst), .slf_op(slf_op_13_09[7:0]),
     .pgate(pgate[159:144]), .bnr_op(net_6500[0:7]),
     .bnl_op(lft_op_13_08[7:0]), .tnr_op(slf_op_14_10[7:0]),
     .tnl_op(lft_op_13_10[7:0]));
ltile4rev I_18_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6506), .lft_op(net_6332[0:7]),
     .sp12_h_l(net_6204[0:23]), .sp4_h_l(net_6205[0:47]),
     .sp4_v_b(net_6208[0:47]), .sp12_v_b(net_7102[0:23]),
     .sp12_h_r(net_6512[0:23]), .sp4_h_r(net_6513[0:47]),
     .sp12_v_t(net_6514[0:23]), .sp4_v_t(net_6236[0:47]),
     .sp4_r_v_b(net_6516[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_18_10[7:0]), .rgt_op(net_7118[0:7]),
     .bot_op(net_6220[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_7094), .purst(purst), .slf_op(net_6248[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6528[0:7]),
     .bnl_op(net_6360[0:7]), .tnr_op(slf_op_19_10[7:0]),
     .tnl_op(slf_op_17_10[7:0]));
ltile4rev I_20_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6534), .lft_op(net_7118[0:7]),
     .sp12_h_l(net_5101[0:23]), .sp4_h_l(net_5110[0:47]),
     .sp4_v_b(net_5108[0:47]), .sp12_v_b(net_7186[0:23]),
     .sp12_h_r(net_6540[0:23]), .sp4_h_r(net_6541[0:47]),
     .sp12_v_t(net_6542[0:23]), .sp4_v_t(net_5107[0:47]),
     .sp4_r_v_b(net_6544[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_20_10[7:0]), .rgt_op(net_6584[0:7]),
     .bot_op(net_5094[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_7178), .purst(purst), .slf_op(net_4936[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6556[0:7]),
     .bnl_op(net_6528[0:7]), .tnr_op(slf_op_21_10[7:0]),
     .tnl_op(slf_op_19_10[7:0]));
ltile4rev I_20_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_20_10), .lft_op(slf_op_19_10[7:0]),
     .sp12_h_l(net_5100[0:23]), .sp4_h_l(net_5109[0:47]),
     .sp4_v_b(net_5107[0:47]), .sp12_v_b(net_6542[0:23]),
     .sp12_h_r(net_6568[0:23]), .sp4_h_r(net_6569[0:47]),
     .sp12_v_t(sp12_v_t_20_10[23:0]), .sp4_v_t(sp4_v_t_20_10[47:0]),
     .sp4_r_v_b(net_6572[0:47]), .wl(wl[175:160]),
     .top_op(top_op_20_10[7:0]), .rgt_op(slf_op_21_10[7:0]),
     .bot_op(net_4936[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_6534), .purst(purst), .slf_op(slf_op_20_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6584[0:7]),
     .bnl_op(net_7118[0:7]), .tnr_op(tnr_op_20_10[7:0]),
     .tnl_op(tnl_op_20_10[7:0]));
ltile4rev I_21_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_21_10), .lft_op(slf_op_20_10[7:0]),
     .sp12_h_l(net_6568[0:23]), .sp4_h_l(net_6569[0:47]),
     .sp4_v_b(net_6572[0:47]), .sp12_v_b(net_6626[0:23]),
     .sp12_h_r(net_6596[0:23]), .sp4_h_r(net_6597[0:47]),
     .sp12_v_t(sp12_v_t_21_10[23:0]), .sp4_v_t(sp4_v_t_21_10[47:0]),
     .sp4_r_v_b(net_6600[0:47]), .wl(wl[175:160]),
     .top_op(top_op_21_10[7:0]), .rgt_op(slf_op_22_10[7:0]),
     .bot_op(net_6584[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_6618), .purst(purst), .slf_op(slf_op_21_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6612[0:7]),
     .bnl_op(net_4936[0:7]), .tnr_op(tnr_op_21_10[7:0]),
     .tnl_op(tnl_op_21_10[7:0]));
ltile4rev I_21_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6618), .lft_op(net_4936[0:7]),
     .sp12_h_l(net_6540[0:23]), .sp4_h_l(net_6541[0:47]),
     .sp4_v_b(net_6544[0:47]), .sp12_v_b(net_7214[0:23]),
     .sp12_h_r(net_6624[0:23]), .sp4_h_r(net_6625[0:47]),
     .sp12_v_t(net_6626[0:23]), .sp4_v_t(net_6572[0:47]),
     .sp4_r_v_b(net_6628[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_21_10[7:0]), .rgt_op(net_6612[0:7]),
     .bot_op(net_6556[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_7206), .purst(purst), .slf_op(net_6584[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6640[0:7]),
     .bnl_op(net_5094[0:7]), .tnr_op(slf_op_22_10[7:0]),
     .tnl_op(slf_op_20_10[7:0]));
ltile4rev I_23_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6646), .lft_op(net_6612[0:7]),
     .sp12_h_l(net_6708[0:23]), .sp4_h_l(net_6709[0:47]),
     .sp4_v_b(net_6712[0:47]), .sp12_v_b(net_7410[0:23]),
     .sp12_h_r(net_6652[0:23]), .sp4_h_r(net_6653[0:47]),
     .sp12_v_t(net_6654[0:23]), .sp4_v_t(net_6740[0:47]),
     .sp4_r_v_b(net_6656[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_23_10[7:0]), .rgt_op(net_6808[0:7]),
     .bot_op(net_6724[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_7402), .purst(purst), .slf_op(net_6752[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6668[0:7]),
     .bnl_op(net_6640[0:7]), .tnr_op(slf_op_24_10[7:0]),
     .tnl_op(slf_op_22_10[7:0]));
ltile4rev I_24_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_24_10), .lft_op(slf_op_23_10[7:0]),
     .sp12_h_l(net_6792[0:23]), .sp4_h_l(net_6793[0:47]),
     .sp4_v_b(net_6796[0:47]), .sp12_v_b(net_6766[0:23]),
     .sp12_h_r(net_6680[0:23]), .sp4_h_r(net_6681[0:47]),
     .sp12_v_t(sp12_v_t_24_10[23:0]), .sp4_v_t(sp4_v_t_24_10[47:0]),
     .sp4_r_v_b(net_6684[0:47]), .wl(wl[175:160]),
     .top_op(top_op_24_10[7:0]), .rgt_op({slf_op_25_10[3],
     slf_op_25_10[2], slf_op_25_10[1], slf_op_25_10[0],
     slf_op_25_10[3], slf_op_25_10[2], slf_op_25_10[1],
     slf_op_25_10[0]}), .bot_op(net_6808[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_6758), .purst(purst), .slf_op(slf_op_24_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op({io_r_08[3], io_r_08[2],
     io_r_08[1], io_r_08[0], io_r_08[3], io_r_08[2], io_r_08[1],
     io_r_08[0]}), .bnl_op(net_6752[0:7]), .tnr_op({tnr_op_24_10[3:0],
     tnr_op_24_10[3:0]}), .tnl_op(tnl_op_24_10[7:0]));
ltile4rev I_22_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6702), .lft_op(net_6584[0:7]),
     .sp12_h_l(net_6624[0:23]), .sp4_h_l(net_6625[0:47]),
     .sp4_v_b(net_6628[0:47]), .sp12_v_b(net_7354[0:23]),
     .sp12_h_r(net_6708[0:23]), .sp4_h_r(net_6709[0:47]),
     .sp12_v_t(net_6710[0:23]), .sp4_v_t(net_6600[0:47]),
     .sp4_r_v_b(net_6712[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_22_10[7:0]), .rgt_op(net_6752[0:7]),
     .bot_op(net_6640[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_7346), .purst(purst), .slf_op(net_6612[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net_6724[0:7]),
     .bnl_op(net_6556[0:7]), .tnr_op(slf_op_23_10[7:0]),
     .tnl_op(slf_op_21_10[7:0]));
ltile4rev I_22_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_22_10), .lft_op(slf_op_21_10[7:0]),
     .sp12_h_l(net_6596[0:23]), .sp4_h_l(net_6597[0:47]),
     .sp4_v_b(net_6600[0:47]), .sp12_v_b(net_6710[0:23]),
     .sp12_h_r(net_6736[0:23]), .sp4_h_r(net_6737[0:47]),
     .sp12_v_t(sp12_v_t_22_10[23:0]), .sp4_v_t(sp4_v_t_22_10[47:0]),
     .sp4_r_v_b(net_6740[0:47]), .wl(wl[175:160]),
     .top_op(top_op_22_10[7:0]), .rgt_op(slf_op_23_10[7:0]),
     .bot_op(net_6612[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_6702), .purst(purst), .slf_op(slf_op_22_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6752[0:7]),
     .bnl_op(net_6584[0:7]), .tnr_op(tnr_op_22_10[7:0]),
     .tnl_op(tnl_op_22_10[7:0]));
ltile4rev I_24_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net_6758), .lft_op(net_6752[0:7]),
     .sp12_h_l(net_6652[0:23]), .sp4_h_l(net_6653[0:47]),
     .sp4_v_b(net_6656[0:47]), .sp12_v_b(net_7298[0:23]),
     .sp12_h_r(net_6764[0:23]), .sp4_h_r(net_6765[0:47]),
     .sp12_v_t(net_6766[0:23]), .sp4_v_t(net_6796[0:47]),
     .sp4_r_v_b(net_6768[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_24_10[7:0]), .rgt_op({io_r_08[3], io_r_08[2],
     io_r_08[1], io_r_08[0], io_r_08[3], io_r_08[2], io_r_08[1],
     io_r_08[0]}), .bot_op(net_6668[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_7290), .purst(purst), .slf_op(net_6808[0:7]),
     .pgate(pgate[159:144]), .bnr_op({io_r_07[3], io_r_07[2],
     io_r_07[1], io_r_07[0], io_r_07[3], io_r_07[2], io_r_07[1],
     io_r_07[0]}), .bnl_op(net_6724[0:7]), .tnr_op({slf_op_25_10[3],
     slf_op_25_10[2], slf_op_25_10[1], slf_op_25_10[0],
     slf_op_25_10[3], slf_op_25_10[2], slf_op_25_10[1],
     slf_op_25_10[0]}), .tnl_op(slf_op_23_10[7:0]));
ltile4rev I_23_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_23_10), .lft_op(slf_op_22_10[7:0]),
     .sp12_h_l(net_6736[0:23]), .sp4_h_l(net_6737[0:47]),
     .sp4_v_b(net_6740[0:47]), .sp12_v_b(net_6654[0:23]),
     .sp12_h_r(net_6792[0:23]), .sp4_h_r(net_6793[0:47]),
     .sp12_v_t(sp12_v_t_23_10[23:0]), .sp4_v_t(sp4_v_t_23_10[47:0]),
     .sp4_r_v_b(net_6796[0:47]), .wl(wl[175:160]),
     .top_op(top_op_23_10[7:0]), .rgt_op(slf_op_24_10[7:0]),
     .bot_op(net_6752[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_6646), .purst(purst), .slf_op(slf_op_23_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net_6808[0:7]),
     .bnl_op(net_6612[0:7]), .tnr_op(tnr_op_23_10[7:0]),
     .tnl_op(tnl_op_23_10[7:0]));
ltile4rev I_13_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_6814), .lft_op(lft_op_13_07[7:0]),
     .sp12_h_l(sp12_h_l_13_07[23:0]), .sp4_h_l(sp4_h_l_13_07[47:0]),
     .sp4_v_b(sp4_v_b_13_07[47:0]), .sp12_v_b(net_5842[0:23]),
     .sp12_h_r(net_6820[0:23]), .sp4_h_r(net_6821[0:47]),
     .sp12_v_t(net_6822[0:23]), .sp4_v_t(sp4_v_b_13_08[47:0]),
     .sp4_r_v_b(net_6824[0:47]), .wl(wl[127:112]),
     .top_op(slf_op_13_08[7:0]), .rgt_op(net_6864[0:7]),
     .bot_op(slf_op_13_06[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5834), .purst(purst), .slf_op(slf_op_13_07[7:0]),
     .pgate(pgate[127:112]), .bnr_op(net_6836[0:7]),
     .bnl_op(lft_op_13_06[7:0]), .tnr_op(net_6500[0:7]),
     .tnl_op(lft_op_13_08[7:0]));
ltile4rev I_13_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_6842), .lft_op(lft_op_13_08[7:0]),
     .sp12_h_l(sp12_h_l_13_08[23:0]), .sp4_h_l(sp4_h_l_13_08[47:0]),
     .sp4_v_b(sp4_v_b_13_08[47:0]), .sp12_v_b(net_6822[0:23]),
     .sp12_h_r(net_6848[0:23]), .sp4_h_r(net_6849[0:47]),
     .sp12_v_t(net_6850[0:23]), .sp4_v_t(sp4_v_b_13_09[47:0]),
     .sp4_r_v_b(net_6852[0:47]), .wl(wl[143:128]),
     .top_op(slf_op_13_09[7:0]), .rgt_op(net_6500[0:7]),
     .bot_op(slf_op_13_07[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_6814), .purst(purst), .slf_op(slf_op_13_08[7:0]),
     .pgate(pgate[143:128]), .bnr_op(net_6864[0:7]),
     .bnl_op(lft_op_13_07[7:0]), .tnr_op(net_6472[0:7]),
     .tnl_op(lft_op_13_09[7:0]));
ltile4rev I_14_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_6870), .lft_op(slf_op_13_08[7:0]),
     .sp12_h_l(net_6848[0:23]), .sp4_h_l(net_6849[0:47]),
     .sp4_v_b(net_6852[0:47]), .sp12_v_b(net_6906[0:23]),
     .sp12_h_r(net_6876[0:23]), .sp4_h_r(net_6877[0:47]),
     .sp12_v_t(net_6878[0:23]), .sp4_v_t(net_6488[0:47]),
     .sp4_r_v_b(net_6880[0:47]), .wl(wl[143:128]),
     .top_op(net_6472[0:7]), .rgt_op(net_6416[0:7]),
     .bot_op(net_6864[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_6898), .purst(purst), .slf_op(net_6500[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_6892[0:7]),
     .bnl_op(slf_op_13_07[7:0]), .tnr_op(net_6444[0:7]),
     .tnl_op(slf_op_13_09[7:0]));
ltile4rev I_14_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_6898), .lft_op(slf_op_13_07[7:0]),
     .sp12_h_l(net_6820[0:23]), .sp4_h_l(net_6821[0:47]),
     .sp4_v_b(net_6824[0:47]), .sp12_v_b(net_5814[0:23]),
     .sp12_h_r(net_6904[0:23]), .sp4_h_r(net_6905[0:47]),
     .sp12_v_t(net_6906[0:23]), .sp4_v_t(net_6852[0:47]),
     .sp4_r_v_b(net_6908[0:47]), .wl(wl[127:112]),
     .top_op(net_6500[0:7]), .rgt_op(net_6892[0:7]),
     .bot_op(net_6836[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_5806), .purst(purst), .slf_op(net_6864[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_6920[0:7]),
     .bnl_op(slf_op_13_06[7:0]), .tnr_op(net_6416[0:7]),
     .tnl_op(slf_op_13_08[7:0]));
ltile4rev I_17_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_6926), .lft_op(net_7032[0:7]),
     .sp12_h_l(net_7072[0:23]), .sp4_h_l(net_7073[0:47]),
     .sp4_v_b(net_7076[0:47]), .sp12_v_b(net_5618[0:23]),
     .sp12_h_r(net_6932[0:23]), .sp4_h_r(net_6933[0:47]),
     .sp12_v_t(net_6934[0:23]), .sp4_v_t(net_7048[0:47]),
     .sp4_r_v_b(net_6936[0:47]), .wl(wl[127:112]),
     .top_op(net_6360[0:7]), .rgt_op(net_6976[0:7]),
     .bot_op(net_7088[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_5610), .purst(purst), .slf_op(net_7060[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_6948[0:7]),
     .bnl_op(net_7004[0:7]), .tnr_op(net_6220[0:7]),
     .tnl_op(net_6276[0:7]));
ltile4rev I_17_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_6954), .lft_op(net_6276[0:7]),
     .sp12_h_l(net_7044[0:23]), .sp4_h_l(net_7045[0:47]),
     .sp4_v_b(net_7048[0:47]), .sp12_v_b(net_6934[0:23]),
     .sp12_h_r(net_6960[0:23]), .sp4_h_r(net_6961[0:47]),
     .sp12_v_t(net_6962[0:23]), .sp4_v_t(net_6348[0:47]),
     .sp4_r_v_b(net_6964[0:47]), .wl(wl[143:128]),
     .top_op(net_6332[0:7]), .rgt_op(net_6220[0:7]),
     .bot_op(net_7060[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_6926), .purst(purst), .slf_op(net_6360[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_6976[0:7]),
     .bnl_op(net_7032[0:7]), .tnr_op(net_6248[0:7]),
     .tnl_op(net_6304[0:7]));
ltile4rev I_15_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_6982), .lft_op(net_6864[0:7]),
     .sp12_h_l(net_6904[0:23]), .sp4_h_l(net_6905[0:47]),
     .sp4_v_b(net_6908[0:47]), .sp12_v_b(net_5674[0:23]),
     .sp12_h_r(net_6988[0:23]), .sp4_h_r(net_6989[0:47]),
     .sp12_v_t(net_6990[0:23]), .sp4_v_t(net_6880[0:47]),
     .sp4_r_v_b(net_6992[0:47]), .wl(wl[127:112]),
     .top_op(net_6416[0:7]), .rgt_op(net_7032[0:7]),
     .bot_op(net_6920[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_5666), .purst(purst), .slf_op(net_6892[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_7004[0:7]),
     .bnl_op(net_6836[0:7]), .tnr_op(net_6276[0:7]),
     .tnl_op(net_6500[0:7]));
ltile4rev I_15_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7010), .lft_op(net_6500[0:7]),
     .sp12_h_l(net_6876[0:23]), .sp4_h_l(net_6877[0:47]),
     .sp4_v_b(net_6880[0:47]), .sp12_v_b(net_6990[0:23]),
     .sp12_h_r(net_7016[0:23]), .sp4_h_r(net_7017[0:47]),
     .sp12_v_t(net_7018[0:23]), .sp4_v_t(net_6404[0:47]),
     .sp4_r_v_b(net_7020[0:47]), .wl(wl[143:128]),
     .top_op(net_6444[0:7]), .rgt_op(net_6276[0:7]),
     .bot_op(net_6892[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_6982), .purst(purst), .slf_op(net_6416[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_7032[0:7]),
     .bnl_op(net_6864[0:7]), .tnr_op(net_6304[0:7]),
     .tnl_op(net_6472[0:7]));
ltile4rev I_16_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7038), .lft_op(net_6416[0:7]),
     .sp12_h_l(net_7016[0:23]), .sp4_h_l(net_7017[0:47]),
     .sp4_v_b(net_7020[0:47]), .sp12_v_b(net_7074[0:23]),
     .sp12_h_r(net_7044[0:23]), .sp4_h_r(net_7045[0:47]),
     .sp12_v_t(net_7046[0:23]), .sp4_v_t(net_6264[0:47]),
     .sp4_r_v_b(net_7048[0:47]), .wl(wl[143:128]),
     .top_op(net_6304[0:7]), .rgt_op(net_6360[0:7]),
     .bot_op(net_7032[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_7066), .purst(purst), .slf_op(net_6276[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_7060[0:7]),
     .bnl_op(net_6892[0:7]), .tnr_op(net_6332[0:7]),
     .tnl_op(net_6444[0:7]));
ltile4rev I_16_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_7066), .lft_op(net_6892[0:7]),
     .sp12_h_l(net_6988[0:23]), .sp4_h_l(net_6989[0:47]),
     .sp4_v_b(net_6992[0:47]), .sp12_v_b(net_5702[0:23]),
     .sp12_h_r(net_7072[0:23]), .sp4_h_r(net_7073[0:47]),
     .sp12_v_t(net_7074[0:23]), .sp4_v_t(net_7020[0:47]),
     .sp4_r_v_b(net_7076[0:47]), .wl(wl[127:112]),
     .top_op(net_6276[0:7]), .rgt_op(net_7060[0:7]),
     .bot_op(net_7004[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_5694), .purst(purst), .slf_op(net_7032[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_7088[0:7]),
     .bnl_op(net_6920[0:7]), .tnr_op(net_6360[0:7]),
     .tnl_op(net_6416[0:7]));
ltile4rev I_18_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7094), .lft_op(net_6360[0:7]),
     .sp12_h_l(net_6960[0:23]), .sp4_h_l(net_6961[0:47]),
     .sp4_v_b(net_6964[0:47]), .sp12_v_b(net_7130[0:23]),
     .sp12_h_r(net_7100[0:23]), .sp4_h_r(net_7101[0:47]),
     .sp12_v_t(net_7102[0:23]), .sp4_v_t(net_6208[0:47]),
     .sp4_r_v_b(net_7104[0:47]), .wl(wl[143:128]),
     .top_op(net_6248[0:7]), .rgt_op(net_6528[0:7]),
     .bot_op(net_6976[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_7122), .purst(purst), .slf_op(net_6220[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_4953[0:7]),
     .bnl_op(net_7060[0:7]), .tnr_op(net_7118[0:7]),
     .tnl_op(net_6332[0:7]));
ltile4rev I_18_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_7122), .lft_op(net_7060[0:7]),
     .sp12_h_l(net_6932[0:23]), .sp4_h_l(net_6933[0:47]),
     .sp4_v_b(net_6936[0:47]), .sp12_v_b(net_5758[0:23]),
     .sp12_h_r(net_7128[0:23]), .sp4_h_r(net_7129[0:47]),
     .sp12_v_t(net_7130[0:23]), .sp4_v_t(net_6964[0:47]),
     .sp4_r_v_b(net_7132[0:47]), .wl(wl[127:112]),
     .top_op(net_6220[0:7]), .rgt_op(net_4953[0:7]),
     .bot_op(net_6948[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_5750), .purst(purst), .slf_op(net_6976[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_7144[0:7]),
     .bnl_op(net_7088[0:7]), .tnr_op(net_6528[0:7]),
     .tnl_op(net_6360[0:7]));
ltile4rev I_20_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_7150), .lft_op(net_4953[0:7]),
     .sp12_h_l(net_4939[0:23]), .sp4_h_l(net_4940[0:47]),
     .sp4_v_b(net_4944[0:47]), .sp12_v_b(net_5954[0:23]),
     .sp12_h_r(net_7156[0:23]), .sp4_h_r(net_7157[0:47]),
     .sp12_v_t(net_7158[0:23]), .sp4_v_t(net_4943[0:47]),
     .sp4_r_v_b(net_7160[0:47]), .wl(wl[127:112]),
     .top_op(net_5094[0:7]), .rgt_op(net_7200[0:7]),
     .bot_op(net_4945[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_5946), .purst(purst), .slf_op(net_5958[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_7172[0:7]),
     .bnl_op(net_7144[0:7]), .tnr_op(net_6556[0:7]),
     .tnl_op(net_6528[0:7]));
ltile4rev I_20_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7178), .lft_op(net_6528[0:7]),
     .sp12_h_l(net_4938[0:23]), .sp4_h_l(net_4941[0:47]),
     .sp4_v_b(net_4943[0:47]), .sp12_v_b(net_7158[0:23]),
     .sp12_h_r(net_7184[0:23]), .sp4_h_r(net_7185[0:47]),
     .sp12_v_t(net_7186[0:23]), .sp4_v_t(net_5108[0:47]),
     .sp4_r_v_b(net_7188[0:47]), .wl(wl[143:128]),
     .top_op(net_4936[0:7]), .rgt_op(net_6556[0:7]),
     .bot_op(net_5958[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_7150), .purst(purst), .slf_op(net_5094[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_7200[0:7]),
     .bnl_op(net_4953[0:7]), .tnr_op(net_6584[0:7]),
     .tnl_op(net_7118[0:7]));
ltile4rev I_21_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7206), .lft_op(net_5094[0:7]),
     .sp12_h_l(net_7184[0:23]), .sp4_h_l(net_7185[0:47]),
     .sp4_v_b(net_7188[0:47]), .sp12_v_b(net_7242[0:23]),
     .sp12_h_r(net_7212[0:23]), .sp4_h_r(net_7213[0:47]),
     .sp12_v_t(net_7214[0:23]), .sp4_v_t(net_6544[0:47]),
     .sp4_r_v_b(net_7216[0:47]), .wl(wl[143:128]),
     .top_op(net_6584[0:7]), .rgt_op(net_6640[0:7]),
     .bot_op(net_7200[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_7234), .purst(purst), .slf_op(net_6556[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_7228[0:7]),
     .bnl_op(net_5958[0:7]), .tnr_op(net_6612[0:7]),
     .tnl_op(net_4936[0:7]));
ltile4rev I_21_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_7234), .lft_op(net_5958[0:7]),
     .sp12_h_l(net_7156[0:23]), .sp4_h_l(net_7157[0:47]),
     .sp4_v_b(net_7160[0:47]), .sp12_v_b(net_5982[0:23]),
     .sp12_h_r(net_7240[0:23]), .sp4_h_r(net_7241[0:47]),
     .sp12_v_t(net_7242[0:23]), .sp4_v_t(net_7188[0:47]),
     .sp4_r_v_b(net_7244[0:47]), .wl(wl[127:112]),
     .top_op(net_6556[0:7]), .rgt_op(net_7228[0:7]),
     .bot_op(net_7172[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_5974), .purst(purst), .slf_op(net_7200[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_7256[0:7]),
     .bnl_op(net_4945[0:7]), .tnr_op(net_6640[0:7]),
     .tnl_op(net_5094[0:7]));
ltile4rev I_23_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_7262), .lft_op(net_7228[0:7]),
     .sp12_h_l(net_7324[0:23]), .sp4_h_l(net_7325[0:47]),
     .sp4_v_b(net_7328[0:47]), .sp12_v_b(net_6178[0:23]),
     .sp12_h_r(net_7268[0:23]), .sp4_h_r(net_7269[0:47]),
     .sp12_v_t(net_7270[0:23]), .sp4_v_t(net_7356[0:47]),
     .sp4_r_v_b(net_7272[0:47]), .wl(wl[127:112]),
     .top_op(net_6724[0:7]), .rgt_op(net_7424[0:7]),
     .bot_op(net_7340[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_6170), .purst(purst), .slf_op(net_7368[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_7284[0:7]),
     .bnl_op(net_7256[0:7]), .tnr_op(net_6668[0:7]),
     .tnl_op(net_6640[0:7]));
ltile4rev I_24_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7290), .lft_op(net_6724[0:7]),
     .sp12_h_l(net_7408[0:23]), .sp4_h_l(net_7409[0:47]),
     .sp4_v_b(net_7412[0:47]), .sp12_v_b(net_7382[0:23]),
     .sp12_h_r(net_7296[0:23]), .sp4_h_r(net_7297[0:47]),
     .sp12_v_t(net_7298[0:23]), .sp4_v_t(net_6656[0:47]),
     .sp4_r_v_b(net_7300[0:47]), .wl(wl[143:128]),
     .top_op(net_6808[0:7]), .rgt_op({io_r_07[3], io_r_07[2],
     io_r_07[1], io_r_07[0], io_r_07[3], io_r_07[2], io_r_07[1],
     io_r_07[0]}), .bot_op(net_7424[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_7374), .purst(purst), .slf_op(net_6668[0:7]),
     .pgate(pgate[143:128]), .bnr_op({io_r_06[3], io_r_06[2],
     io_r_06[1], io_r_06[0], io_r_06[3], io_r_06[2], io_r_06[1],
     io_r_06[0]}), .bnl_op(net_7368[0:7]), .tnr_op({io_r_08[3],
     io_r_08[2], io_r_08[1], io_r_08[0], io_r_08[3], io_r_08[2],
     io_r_08[1], io_r_08[0]}), .tnl_op(net_6752[0:7]));
ltile4rev I_22_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_7318), .lft_op(net_7200[0:7]),
     .sp12_h_l(net_7240[0:23]), .sp4_h_l(net_7241[0:47]),
     .sp4_v_b(net_7244[0:47]), .sp12_v_b(net_6122[0:23]),
     .sp12_h_r(net_7324[0:23]), .sp4_h_r(net_7325[0:47]),
     .sp12_v_t(net_7326[0:23]), .sp4_v_t(net_7216[0:47]),
     .sp4_r_v_b(net_7328[0:47]), .wl(wl[127:112]),
     .top_op(net_6640[0:7]), .rgt_op(net_7368[0:7]),
     .bot_op(net_7256[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_6114), .purst(purst), .slf_op(net_7228[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net_7340[0:7]),
     .bnl_op(net_7172[0:7]), .tnr_op(net_6724[0:7]),
     .tnl_op(net_6556[0:7]));
ltile4rev I_22_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7346), .lft_op(net_6556[0:7]),
     .sp12_h_l(net_7212[0:23]), .sp4_h_l(net_7213[0:47]),
     .sp4_v_b(net_7216[0:47]), .sp12_v_b(net_7326[0:23]),
     .sp12_h_r(net_7352[0:23]), .sp4_h_r(net_7353[0:47]),
     .sp12_v_t(net_7354[0:23]), .sp4_v_t(net_6628[0:47]),
     .sp4_r_v_b(net_7356[0:47]), .wl(wl[143:128]),
     .top_op(net_6612[0:7]), .rgt_op(net_6724[0:7]),
     .bot_op(net_7228[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_7318), .purst(purst), .slf_op(net_6640[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_7368[0:7]),
     .bnl_op(net_7200[0:7]), .tnr_op(net_6752[0:7]),
     .tnl_op(net_6584[0:7]));
ltile4rev I_24_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net_7374), .lft_op(net_7368[0:7]),
     .sp12_h_l(net_7268[0:23]), .sp4_h_l(net_7269[0:47]),
     .sp4_v_b(net_7272[0:47]), .sp12_v_b(net_6066[0:23]),
     .sp12_h_r(net_7380[0:23]), .sp4_h_r(net_7381[0:47]),
     .sp12_v_t(net_7382[0:23]), .sp4_v_t(net_7412[0:47]),
     .sp4_r_v_b(net_7384[0:47]), .wl(wl[127:112]),
     .top_op(net_6668[0:7]), .rgt_op({io_r_06[3], io_r_06[2],
     io_r_06[1], io_r_06[0], io_r_06[3], io_r_06[2], io_r_06[1],
     io_r_06[0]}), .bot_op(net_7284[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_6058), .purst(purst), .slf_op(net_7424[0:7]),
     .pgate(pgate[127:112]), .bnr_op({io_r_05[3], io_r_05[2],
     io_r_05[1], io_r_05[0], io_r_05[3], io_r_05[2], io_r_05[1],
     io_r_05[0]}), .bnl_op(net_7340[0:7]), .tnr_op({io_r_07[3],
     io_r_07[2], io_r_07[1], io_r_07[0], io_r_07[3], io_r_07[2],
     io_r_07[1], io_r_07[0]}), .tnl_op(net_6724[0:7]));
ltile4rev I_23_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net_7402), .lft_op(net_6640[0:7]),
     .sp12_h_l(net_7352[0:23]), .sp4_h_l(net_7353[0:47]),
     .sp4_v_b(net_7356[0:47]), .sp12_v_b(net_7270[0:23]),
     .sp12_h_r(net_7408[0:23]), .sp4_h_r(net_7409[0:47]),
     .sp12_v_t(net_7410[0:23]), .sp4_v_t(net_6712[0:47]),
     .sp4_r_v_b(net_7412[0:47]), .wl(wl[143:128]),
     .top_op(net_6752[0:7]), .rgt_op(net_6668[0:7]),
     .bot_op(net_7368[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_7262), .purst(purst), .slf_op(net_6724[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net_7424[0:7]),
     .bnl_op(net_7228[0:7]), .tnr_op(net_6808[0:7]),
     .tnl_op(net_6612[0:7]));
ltile4rev I_23_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_7430), .lft_op(net_5548[0:7]),
     .sp12_h_l(net_7492[0:23]), .sp4_h_l(net_7493[0:47]),
     .sp4_v_b(net_7496[0:47]), .sp12_v_b(net_4369[0:23]),
     .sp12_h_r(net_7436[0:23]), .sp4_h_r(net_7437[0:47]),
     .sp12_v_t(net_7438[0:23]), .sp4_v_t(net_7524[0:47]),
     .sp4_r_v_b(net_7440[0:47]), .wl(wl[31:16]),
     .top_op(net_8124[0:7]), .rgt_op(net_7592[0:7]),
     .bot_op({io_b_44[3], io_b_44[2], io_b_44[1], io_b_44[0],
     io_b_44[3], io_b_44[2], io_b_44[1], io_b_44[0]}),
     .bl(bl[1239:1186]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_23[7:0]), .carry_in(net_8259), .purst(purst),
     .slf_op(net_7536[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_46[3],
     io_b_46[2], io_b_46[1], io_b_46[0], io_b_46[3], io_b_46[2],
     io_b_46[1], io_b_46[0]}), .bnl_op({io_b_42[3], io_b_42[2],
     io_b_42[1], io_b_42[0], io_b_42[3], io_b_42[2], io_b_42[1],
     io_b_42[0]}), .tnr_op(net_8068[0:7]), .tnl_op(net_8040[0:7]));
ltile4rev I_24_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_7458), .lft_op(net_8124[0:7]),
     .sp12_h_l(net_7576[0:23]), .sp4_h_l(net_7577[0:47]),
     .sp4_v_b(net_7580[0:47]), .sp12_v_b(net_7550[0:23]),
     .sp12_h_r(net_7464[0:23]), .sp4_h_r(net_7465[0:47]),
     .sp12_v_t(net_7466[0:23]), .sp4_v_t(net_8056[0:47]),
     .sp4_r_v_b(net_7468[0:47]), .wl(wl[47:32]),
     .top_op(net_8208[0:7]), .rgt_op({io_r_01[3], io_r_01[2],
     io_r_01[1], io_r_01[0], io_r_01[3], io_r_01[2], io_r_01[1],
     io_r_01[0]}), .bot_op(net_7592[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_7542), .purst(purst), .slf_op(net_8068[0:7]),
     .pgate(pgate[47:32]), .bnr_op({io_r_00[3], io_r_00[2], io_r_00[1],
     io_r_00[0], io_r_00[3], io_r_00[2], io_r_00[1], io_r_00[0]}),
     .bnl_op(net_7536[0:7]), .tnr_op({io_r_02[3], io_r_02[2],
     io_r_02[1], io_r_02[0], io_r_02[3], io_r_02[2], io_r_02[1],
     io_r_02[0]}), .tnl_op(net_8152[0:7]));
ltile4rev I_22_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_7486), .lft_op(net_5520[0:7]),
     .sp12_h_l(net_5560[0:23]), .sp4_h_l(net_5561[0:47]),
     .sp4_v_b(net_5564[0:47]), .sp12_v_b(net_4403[0:23]),
     .sp12_h_r(net_7492[0:23]), .sp4_h_r(net_7493[0:47]),
     .sp12_v_t(net_7494[0:23]), .sp4_v_t(net_5536[0:47]),
     .sp4_r_v_b(net_7496[0:47]), .wl(wl[31:16]),
     .top_op(net_8040[0:7]), .rgt_op(net_7536[0:7]),
     .bot_op({io_b_42[3], io_b_42[2], io_b_42[1], io_b_42[0],
     io_b_42[3], io_b_42[2], io_b_42[1], io_b_42[0]}),
     .bl(bl[1185:1132]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_22[7:0]), .carry_in(net_7504), .purst(purst),
     .slf_op(net_5548[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_44[3],
     io_b_44[2], io_b_44[1], io_b_44[0], io_b_44[3], io_b_44[2],
     io_b_44[1], io_b_44[0]}), .bnl_op({io_b_40[3], io_b_40[2],
     io_b_40[1], io_b_40[0], io_b_40[3], io_b_40[2], io_b_40[1],
     io_b_40[0]}), .tnr_op(net_8124[0:7]), .tnl_op(net_7956[0:7]));
ltile4rev I_22_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_7514), .lft_op(net_7956[0:7]),
     .sp12_h_l(net_5532[0:23]), .sp4_h_l(net_5533[0:47]),
     .sp4_v_b(net_5536[0:47]), .sp12_v_b(net_7494[0:23]),
     .sp12_h_r(net_7520[0:23]), .sp4_h_r(net_7521[0:47]),
     .sp12_v_t(net_7522[0:23]), .sp4_v_t(net_8028[0:47]),
     .sp4_r_v_b(net_7524[0:47]), .wl(wl[47:32]),
     .top_op(net_8012[0:7]), .rgt_op(net_8124[0:7]),
     .bot_op(net_5548[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_7486), .purst(purst), .slf_op(net_8040[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_7536[0:7]),
     .bnl_op(net_5520[0:7]), .tnr_op(net_8152[0:7]),
     .tnl_op(net_7984[0:7]));
ltile4rev I_24_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net_7542), .lft_op(net_7536[0:7]),
     .sp12_h_l(net_7436[0:23]), .sp4_h_l(net_7437[0:47]),
     .sp4_v_b(net_7440[0:47]), .sp12_v_b(net_4709[0:23]),
     .sp12_h_r(net_7548[0:23]), .sp4_h_r(net_7549[0:47]),
     .sp12_v_t(net_7550[0:23]), .sp4_v_t(net_7580[0:47]),
     .sp4_r_v_b(net_7552[0:47]), .wl(wl[31:16]),
     .top_op(net_8068[0:7]), .rgt_op({io_r_00[3], io_r_00[2],
     io_r_00[1], io_r_00[0], io_r_00[3], io_r_00[2], io_r_00[1],
     io_r_00[0]}), .bot_op({io_b_46[3], io_b_46[2], io_b_46[1],
     io_b_46[0], io_b_46[3], io_b_46[2], io_b_46[1], io_b_46[0]}),
     .bl(bl[1293:1240]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_24[7:0]), .carry_in(net_7560), .purst(purst),
     .slf_op(net_7592[0:7]), .pgate(pgate[31:16]), .bnr_op({tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .bnl_op({io_b_44[3], io_b_44[2], io_b_44[1], io_b_44[0],
     io_b_44[3], io_b_44[2], io_b_44[1], io_b_44[0]}),
     .tnr_op({io_r_01[3], io_r_01[2], io_r_01[1], io_r_01[0],
     io_r_01[3], io_r_01[2], io_r_01[1], io_r_01[0]}),
     .tnl_op(net_8124[0:7]));
ltile4rev I_23_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net_7570), .lft_op(net_8040[0:7]),
     .sp12_h_l(net_7520[0:23]), .sp4_h_l(net_7521[0:47]),
     .sp4_v_b(net_7524[0:47]), .sp12_v_b(net_7438[0:23]),
     .sp12_h_r(net_7576[0:23]), .sp4_h_r(net_7577[0:47]),
     .sp12_v_t(net_7578[0:23]), .sp4_v_t(net_8112[0:47]),
     .sp4_r_v_b(net_7580[0:47]), .wl(wl[47:32]),
     .top_op(net_8152[0:7]), .rgt_op(net_8068[0:7]),
     .bot_op(net_7536[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_7430), .purst(purst), .slf_op(net_8124[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net_7592[0:7]),
     .bnl_op(net_5548[0:7]), .tnr_op(net_8208[0:7]),
     .tnl_op(net_8012[0:7]));
ltile4rev I_13_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_7598), .lft_op(lft_op_13_03[7:0]),
     .sp12_h_l(sp12_h_l_13_03[23:0]), .sp4_h_l(sp4_h_l_13_03[47:0]),
     .sp4_v_b(sp4_v_b_13_03[47:0]), .sp12_v_b(net_5394[0:23]),
     .sp12_h_r(net_7604[0:23]), .sp4_h_r(net_7605[0:47]),
     .sp12_v_t(net_7606[0:23]), .sp4_v_t(sp4_v_b_13_04[47:0]),
     .sp4_r_v_b(net_7608[0:47]), .wl(wl[63:48]),
     .top_op(slf_op_13_04[7:0]), .rgt_op(net_7648[0:7]),
     .bot_op(slf_op_13_02[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5386), .purst(purst), .slf_op(slf_op_13_03[7:0]),
     .pgate(pgate[63:48]), .bnr_op(net_7620[0:7]),
     .bnl_op(lft_op_13_02[7:0]), .tnr_op(net_5884[0:7]),
     .tnl_op(lft_op_13_04[7:0]));
ltile4rev I_13_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7626), .lft_op(lft_op_13_04[7:0]),
     .sp12_h_l(sp12_h_l_13_04[23:0]), .sp4_h_l(sp4_h_l_13_04[47:0]),
     .sp4_v_b(sp4_v_b_13_04[47:0]), .sp12_v_b(net_7606[0:23]),
     .sp12_h_r(net_7632[0:23]), .sp4_h_r(net_7633[0:47]),
     .sp12_v_t(net_7634[0:23]), .sp4_v_t(sp4_v_b_13_05[47:0]),
     .sp4_r_v_b(net_7636[0:47]), .wl(wl[79:64]),
     .top_op(slf_op_13_05[7:0]), .rgt_op(net_5884[0:7]),
     .bot_op(slf_op_13_03[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_7598), .purst(purst), .slf_op(slf_op_13_04[7:0]),
     .pgate(pgate[79:64]), .bnr_op(net_7648[0:7]),
     .bnl_op(lft_op_13_03[7:0]), .tnr_op(net_5856[0:7]),
     .tnl_op(lft_op_13_05[7:0]));
ltile4rev I_14_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7654), .lft_op(slf_op_13_04[7:0]),
     .sp12_h_l(net_7632[0:23]), .sp4_h_l(net_7633[0:47]),
     .sp4_v_b(net_7636[0:47]), .sp12_v_b(net_7690[0:23]),
     .sp12_h_r(net_7660[0:23]), .sp4_h_r(net_7661[0:47]),
     .sp12_v_t(net_7662[0:23]), .sp4_v_t(net_5872[0:47]),
     .sp4_r_v_b(net_7664[0:47]), .wl(wl[79:64]),
     .top_op(net_5856[0:7]), .rgt_op(net_5800[0:7]),
     .bot_op(net_7648[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_7682), .purst(purst), .slf_op(net_5884[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_7676[0:7]),
     .bnl_op(slf_op_13_03[7:0]), .tnr_op(net_5828[0:7]),
     .tnl_op(slf_op_13_05[7:0]));
ltile4rev I_14_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_7682), .lft_op(slf_op_13_03[7:0]),
     .sp12_h_l(net_7604[0:23]), .sp4_h_l(net_7605[0:47]),
     .sp4_v_b(net_7608[0:47]), .sp12_v_b(net_5366[0:23]),
     .sp12_h_r(net_7688[0:23]), .sp4_h_r(net_7689[0:47]),
     .sp12_v_t(net_7690[0:23]), .sp4_v_t(net_7636[0:47]),
     .sp4_r_v_b(net_7692[0:47]), .wl(wl[63:48]),
     .top_op(net_5884[0:7]), .rgt_op(net_7676[0:7]),
     .bot_op(net_7620[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_5358), .purst(purst), .slf_op(net_7648[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_7704[0:7]),
     .bnl_op(slf_op_13_02[7:0]), .tnr_op(net_5800[0:7]),
     .tnl_op(slf_op_13_04[7:0]));
ltile4rev I_17_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_7710), .lft_op(net_7816[0:7]),
     .sp12_h_l(net_7856[0:23]), .sp4_h_l(net_7857[0:47]),
     .sp4_v_b(net_7860[0:47]), .sp12_v_b(net_5170[0:23]),
     .sp12_h_r(net_7716[0:23]), .sp4_h_r(net_7717[0:47]),
     .sp12_v_t(net_7718[0:23]), .sp4_v_t(net_7832[0:47]),
     .sp4_r_v_b(net_7720[0:47]), .wl(wl[63:48]),
     .top_op(net_5744[0:7]), .rgt_op(net_7760[0:7]),
     .bot_op(net_7872[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_5162), .purst(purst), .slf_op(net_7844[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_7732[0:7]),
     .bnl_op(net_7788[0:7]), .tnr_op(net_5604[0:7]),
     .tnl_op(net_5660[0:7]));
ltile4rev I_17_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7738), .lft_op(net_5660[0:7]),
     .sp12_h_l(net_7828[0:23]), .sp4_h_l(net_7829[0:47]),
     .sp4_v_b(net_7832[0:47]), .sp12_v_b(net_7718[0:23]),
     .sp12_h_r(net_7744[0:23]), .sp4_h_r(net_7745[0:47]),
     .sp12_v_t(net_7746[0:23]), .sp4_v_t(net_5732[0:47]),
     .sp4_r_v_b(net_7748[0:47]), .wl(wl[79:64]),
     .top_op(net_5716[0:7]), .rgt_op(net_5604[0:7]),
     .bot_op(net_7844[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_7710), .purst(purst), .slf_op(net_5744[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_7760[0:7]),
     .bnl_op(net_7816[0:7]), .tnr_op(net_5632[0:7]),
     .tnl_op(net_5688[0:7]));
ltile4rev I_15_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_7766), .lft_op(net_7648[0:7]),
     .sp12_h_l(net_7688[0:23]), .sp4_h_l(net_7689[0:47]),
     .sp4_v_b(net_7692[0:47]), .sp12_v_b(net_5226[0:23]),
     .sp12_h_r(net_7772[0:23]), .sp4_h_r(net_7773[0:47]),
     .sp12_v_t(net_7774[0:23]), .sp4_v_t(net_7664[0:47]),
     .sp4_r_v_b(net_7776[0:47]), .wl(wl[63:48]),
     .top_op(net_5800[0:7]), .rgt_op(net_7816[0:7]),
     .bot_op(net_7704[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_5218), .purst(purst), .slf_op(net_7676[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_7788[0:7]),
     .bnl_op(net_7620[0:7]), .tnr_op(net_5660[0:7]),
     .tnl_op(net_5884[0:7]));
ltile4rev I_15_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7794), .lft_op(net_5884[0:7]),
     .sp12_h_l(net_7660[0:23]), .sp4_h_l(net_7661[0:47]),
     .sp4_v_b(net_7664[0:47]), .sp12_v_b(net_7774[0:23]),
     .sp12_h_r(net_7800[0:23]), .sp4_h_r(net_7801[0:47]),
     .sp12_v_t(net_7802[0:23]), .sp4_v_t(net_5788[0:47]),
     .sp4_r_v_b(net_7804[0:47]), .wl(wl[79:64]),
     .top_op(net_5828[0:7]), .rgt_op(net_5660[0:7]),
     .bot_op(net_7676[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_7766), .purst(purst), .slf_op(net_5800[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_7816[0:7]),
     .bnl_op(net_7648[0:7]), .tnr_op(net_5688[0:7]),
     .tnl_op(net_5856[0:7]));
ltile4rev I_16_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7822), .lft_op(net_5800[0:7]),
     .sp12_h_l(net_7800[0:23]), .sp4_h_l(net_7801[0:47]),
     .sp4_v_b(net_7804[0:47]), .sp12_v_b(net_7858[0:23]),
     .sp12_h_r(net_7828[0:23]), .sp4_h_r(net_7829[0:47]),
     .sp12_v_t(net_7830[0:23]), .sp4_v_t(net_5648[0:47]),
     .sp4_r_v_b(net_7832[0:47]), .wl(wl[79:64]),
     .top_op(net_5688[0:7]), .rgt_op(net_5744[0:7]),
     .bot_op(net_7816[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_7850), .purst(purst), .slf_op(net_5660[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_7844[0:7]),
     .bnl_op(net_7676[0:7]), .tnr_op(net_5716[0:7]),
     .tnl_op(net_5828[0:7]));
ltile4rev I_16_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_7850), .lft_op(net_7676[0:7]),
     .sp12_h_l(net_7772[0:23]), .sp4_h_l(net_7773[0:47]),
     .sp4_v_b(net_7776[0:47]), .sp12_v_b(net_5254[0:23]),
     .sp12_h_r(net_7856[0:23]), .sp4_h_r(net_7857[0:47]),
     .sp12_v_t(net_7858[0:23]), .sp4_v_t(net_7804[0:47]),
     .sp4_r_v_b(net_7860[0:47]), .wl(wl[63:48]),
     .top_op(net_5660[0:7]), .rgt_op(net_7844[0:7]),
     .bot_op(net_7788[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_5246), .purst(purst), .slf_op(net_7816[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_7872[0:7]),
     .bnl_op(net_7704[0:7]), .tnr_op(net_5744[0:7]),
     .tnl_op(net_5800[0:7]));
ltile4rev I_18_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7878), .lft_op(net_5744[0:7]),
     .sp12_h_l(net_7744[0:23]), .sp4_h_l(net_7745[0:47]),
     .sp4_v_b(net_7748[0:47]), .sp12_v_b(net_7914[0:23]),
     .sp12_h_r(net_7884[0:23]), .sp4_h_r(net_7885[0:47]),
     .sp12_v_t(net_7886[0:23]), .sp4_v_t(net_5592[0:47]),
     .sp4_r_v_b(net_7888[0:47]), .wl(wl[79:64]),
     .top_op(net_5632[0:7]), .rgt_op(net_5912[0:7]),
     .bot_op(net_7760[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_7906), .purst(purst), .slf_op(net_5604[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_4829[0:7]),
     .bnl_op(net_7844[0:7]), .tnr_op(net_7902[0:7]),
     .tnl_op(net_5716[0:7]));
ltile4rev I_18_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_7906), .lft_op(net_7844[0:7]),
     .sp12_h_l(net_7716[0:23]), .sp4_h_l(net_7717[0:47]),
     .sp4_v_b(net_7720[0:47]), .sp12_v_b(net_5310[0:23]),
     .sp12_h_r(net_7912[0:23]), .sp4_h_r(net_7913[0:47]),
     .sp12_v_t(net_7914[0:23]), .sp4_v_t(net_7748[0:47]),
     .sp4_r_v_b(net_7916[0:47]), .wl(wl[63:48]),
     .top_op(net_5604[0:7]), .rgt_op(net_4829[0:7]),
     .bot_op(net_7732[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_5302), .purst(purst), .slf_op(net_7760[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_5466[0:7]),
     .bnl_op(net_7872[0:7]), .tnr_op(net_5912[0:7]),
     .tnl_op(net_5744[0:7]));
ltile4rev I_20_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_7934), .lft_op(net_4829[0:7]),
     .sp12_h_l(net_5016[0:23]), .sp4_h_l(net_5017[0:47]),
     .sp4_v_b(net_5021[0:47]), .sp12_v_b(net_5506[0:23]),
     .sp12_h_r(net_7940[0:23]), .sp4_h_r(net_7941[0:47]),
     .sp12_v_t(net_7942[0:23]), .sp4_v_t(net_5020[0:47]),
     .sp4_r_v_b(net_7944[0:47]), .wl(wl[63:48]),
     .top_op(net_4970[0:7]), .rgt_op(net_7984[0:7]),
     .bot_op(net_5022[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_5498), .purst(purst), .slf_op(net_5510[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_7956[0:7]),
     .bnl_op(net_5466[0:7]), .tnr_op(net_5940[0:7]),
     .tnl_op(net_5912[0:7]));
ltile4rev I_20_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7962), .lft_op(net_5912[0:7]),
     .sp12_h_l(net_5015[0:23]), .sp4_h_l(net_5018[0:47]),
     .sp4_v_b(net_5020[0:47]), .sp12_v_b(net_7942[0:23]),
     .sp12_h_r(net_7968[0:23]), .sp4_h_r(net_7969[0:47]),
     .sp12_v_t(net_7970[0:23]), .sp4_v_t(net_4984[0:47]),
     .sp4_r_v_b(net_7972[0:47]), .wl(wl[79:64]),
     .top_op(net_5013[0:7]), .rgt_op(net_5940[0:7]),
     .bot_op(net_5510[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_7934), .purst(purst), .slf_op(net_4970[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_7984[0:7]),
     .bnl_op(net_4829[0:7]), .tnr_op(net_5968[0:7]),
     .tnl_op(net_7902[0:7]));
ltile4rev I_21_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_7990), .lft_op(net_4970[0:7]),
     .sp12_h_l(net_7968[0:23]), .sp4_h_l(net_7969[0:47]),
     .sp4_v_b(net_7972[0:47]), .sp12_v_b(net_8026[0:23]),
     .sp12_h_r(net_7996[0:23]), .sp4_h_r(net_7997[0:47]),
     .sp12_v_t(net_7998[0:23]), .sp4_v_t(net_5928[0:47]),
     .sp4_r_v_b(net_8000[0:47]), .wl(wl[79:64]),
     .top_op(net_5968[0:7]), .rgt_op(net_6024[0:7]),
     .bot_op(net_7984[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_8018), .purst(purst), .slf_op(net_5940[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_8012[0:7]),
     .bnl_op(net_5510[0:7]), .tnr_op(net_5996[0:7]),
     .tnl_op(net_5013[0:7]));
ltile4rev I_21_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_8018), .lft_op(net_5510[0:7]),
     .sp12_h_l(net_7940[0:23]), .sp4_h_l(net_7941[0:47]),
     .sp4_v_b(net_7944[0:47]), .sp12_v_b(net_5534[0:23]),
     .sp12_h_r(net_8024[0:23]), .sp4_h_r(net_8025[0:47]),
     .sp12_v_t(net_8026[0:23]), .sp4_v_t(net_7972[0:47]),
     .sp4_r_v_b(net_8028[0:47]), .wl(wl[63:48]),
     .top_op(net_5940[0:7]), .rgt_op(net_8012[0:7]),
     .bot_op(net_7956[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_5526), .purst(purst), .slf_op(net_7984[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_8040[0:7]),
     .bnl_op(net_5022[0:7]), .tnr_op(net_6024[0:7]),
     .tnl_op(net_4970[0:7]));
ltile4rev I_23_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_8046), .lft_op(net_8012[0:7]),
     .sp12_h_l(net_8108[0:23]), .sp4_h_l(net_8109[0:47]),
     .sp4_v_b(net_8112[0:47]), .sp12_v_b(net_7578[0:23]),
     .sp12_h_r(net_8052[0:23]), .sp4_h_r(net_8053[0:47]),
     .sp12_v_t(net_8054[0:23]), .sp4_v_t(net_8140[0:47]),
     .sp4_r_v_b(net_8056[0:47]), .wl(wl[63:48]),
     .top_op(net_6108[0:7]), .rgt_op(net_8208[0:7]),
     .bot_op(net_8124[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_7570), .purst(purst), .slf_op(net_8152[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_8068[0:7]),
     .bnl_op(net_8040[0:7]), .tnr_op(net_6052[0:7]),
     .tnl_op(net_6024[0:7]));
ltile4rev I_24_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_8074), .lft_op(net_6108[0:7]),
     .sp12_h_l(net_8192[0:23]), .sp4_h_l(net_8193[0:47]),
     .sp4_v_b(net_8196[0:47]), .sp12_v_b(net_8166[0:23]),
     .sp12_h_r(net_8080[0:23]), .sp4_h_r(net_8081[0:47]),
     .sp12_v_t(net_8082[0:23]), .sp4_v_t(net_6040[0:47]),
     .sp4_r_v_b(net_8084[0:47]), .wl(wl[79:64]),
     .top_op(net_6192[0:7]), .rgt_op({io_r_03[3], io_r_03[2],
     io_r_03[1], io_r_03[0], io_r_03[3], io_r_03[2], io_r_03[1],
     io_r_03[0]}), .bot_op(net_8208[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_8158), .purst(purst), .slf_op(net_6052[0:7]),
     .pgate(pgate[79:64]), .bnr_op({io_r_02[3], io_r_02[2], io_r_02[1],
     io_r_02[0], io_r_02[3], io_r_02[2], io_r_02[1], io_r_02[0]}),
     .bnl_op(net_8152[0:7]), .tnr_op({io_r_04[3], io_r_04[2],
     io_r_04[1], io_r_04[0], io_r_04[3], io_r_04[2], io_r_04[1],
     io_r_04[0]}), .tnl_op(net_6136[0:7]));
ltile4rev I_22_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_8102), .lft_op(net_7984[0:7]),
     .sp12_h_l(net_8024[0:23]), .sp4_h_l(net_8025[0:47]),
     .sp4_v_b(net_8028[0:47]), .sp12_v_b(net_7522[0:23]),
     .sp12_h_r(net_8108[0:23]), .sp4_h_r(net_8109[0:47]),
     .sp12_v_t(net_8110[0:23]), .sp4_v_t(net_8000[0:47]),
     .sp4_r_v_b(net_8112[0:47]), .wl(wl[63:48]),
     .top_op(net_6024[0:7]), .rgt_op(net_8152[0:7]),
     .bot_op(net_8040[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_7514), .purst(purst), .slf_op(net_8012[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net_8124[0:7]),
     .bnl_op(net_7956[0:7]), .tnr_op(net_6108[0:7]),
     .tnl_op(net_5940[0:7]));
ltile4rev I_22_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_8130), .lft_op(net_5940[0:7]),
     .sp12_h_l(net_7996[0:23]), .sp4_h_l(net_7997[0:47]),
     .sp4_v_b(net_8000[0:47]), .sp12_v_b(net_8110[0:23]),
     .sp12_h_r(net_8136[0:23]), .sp4_h_r(net_8137[0:47]),
     .sp12_v_t(net_8138[0:23]), .sp4_v_t(net_6012[0:47]),
     .sp4_r_v_b(net_8140[0:47]), .wl(wl[79:64]),
     .top_op(net_5996[0:7]), .rgt_op(net_6108[0:7]),
     .bot_op(net_8012[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_8102), .purst(purst), .slf_op(net_6024[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_8152[0:7]),
     .bnl_op(net_7984[0:7]), .tnr_op(net_6136[0:7]),
     .tnl_op(net_5968[0:7]));
ltile4rev I_24_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net_8158), .lft_op(net_8152[0:7]),
     .sp12_h_l(net_8052[0:23]), .sp4_h_l(net_8053[0:47]),
     .sp4_v_b(net_8056[0:47]), .sp12_v_b(net_7466[0:23]),
     .sp12_h_r(net_8164[0:23]), .sp4_h_r(net_8165[0:47]),
     .sp12_v_t(net_8166[0:23]), .sp4_v_t(net_8196[0:47]),
     .sp4_r_v_b(net_8168[0:47]), .wl(wl[63:48]),
     .top_op(net_6052[0:7]), .rgt_op({io_r_02[3], io_r_02[2],
     io_r_02[1], io_r_02[0], io_r_02[3], io_r_02[2], io_r_02[1],
     io_r_02[0]}), .bot_op(net_8068[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_7458), .purst(purst), .slf_op(net_8208[0:7]),
     .pgate(pgate[63:48]), .bnr_op({io_r_01[3], io_r_01[2], io_r_01[1],
     io_r_01[0], io_r_01[3], io_r_01[2], io_r_01[1], io_r_01[0]}),
     .bnl_op(net_8124[0:7]), .tnr_op({io_r_03[3], io_r_03[2],
     io_r_03[1], io_r_03[0], io_r_03[3], io_r_03[2], io_r_03[1],
     io_r_03[0]}), .tnl_op(net_6108[0:7]));
ltile4rev I_23_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net_8186), .lft_op(net_6024[0:7]),
     .sp12_h_l(net_8136[0:23]), .sp4_h_l(net_8137[0:47]),
     .sp4_v_b(net_8140[0:47]), .sp12_v_b(net_8054[0:23]),
     .sp12_h_r(net_8192[0:23]), .sp4_h_r(net_8193[0:47]),
     .sp12_v_t(net_8194[0:23]), .sp4_v_t(net_6096[0:47]),
     .sp4_r_v_b(net_8196[0:47]), .wl(wl[79:64]),
     .top_op(net_6136[0:7]), .rgt_op(net_6052[0:7]),
     .bot_op(net_8152[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_8046), .purst(purst), .slf_op(net_6108[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net_8208[0:7]),
     .bnl_op(net_8012[0:7]), .tnr_op(net_6192[0:7]),
     .tnl_op(net_5996[0:7]));
clk_colbufx8 I785 ( .clko(glb_netwk_13[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I786 ( .clko(glb_netwk_14[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I787 ( .clko(glb_netwk_16[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I788 ( .clko(glb_netwk_15[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I789 ( .clko(glb_netwk_19[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I790 ( .clko(glb_netwk_20[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I791 ( .clko(glb_netwk_18[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I792 ( .clko(glb_netwk_17[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I793 ( .clko(glb_netwk_io_r[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I797 ( .clko(glb_netwk_23[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I798 ( .clko(glb_netwk_24[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I799 ( .clko(glb_netwk_22[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I800 ( .clko(glb_netwk_21[7:0]),
     .clki(net2col_drivers[7:0]));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbankin_pbuffer_top, View -
//schematic
// LAST TIME SAVED: Aug 24 17:33:59 2007
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module bram_4kbankin_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [7:0]  bm_sa_i;
input [7:0]  bm_ab;
input [7:0]  bm_aa;
input [15:0]  bm_d;
input [15:0]  bm_bweb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankin I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbankin, View - schematic
// LAST TIME SAVED: Aug 22 17:37:06 2007
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module bram_4kprouting_tbankin ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [47:0]  sp4_h_l_top;
inout [23:0]  sp12_h_l_top;
inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_bot;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_r_v_b_bot;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_v_b_top;

input [7:0]  rgt_op_bot;
input [7:0]  bot_op_bot;
input [7:0]  top_op_top;
input [7:0]  bnr_op_bot;
input [15:0]  reset_b_top;
input [7:0]  bnr_op_top;
input [15:0]  pgate_bot;
input [15:0]  pgate_top;
input [15:0]  wl_top;
input [15:0]  vdd_cntl_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  lft_op_bot;
input [7:0]  tnr_op_bot;
input [7:0]  bnl_op_top;
input [7:0]  tnl_op_top;
input [7:0]  rgt_op_top;
input [7:0]  tnl_op_bot;
input [15:0]  wl_bot;
input [7:0]  bnl_op_bot;
input [7:0]  tnr_op_top;
input [7:0]  bm_sa_i;
input [7:0]  glb_netwk;
input [7:0]  lft_op_top;
input [15:0]  reset_b_bot;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net208;

wire  [0:7]  net210;

wire  [0:7]  net242;

wire  [0:7]  net316;

wire  [0:7]  net243;

wire  [0:7]  net240;

wire  [0:7]  net295;

wire  [0:7]  net241;

wire  [0:7]  net211;

wire  [0:7]  net209;



bram_4kbankin_pbuffer_top I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net245), .bm_wen(net213),
     .bm_d(bm_d[15:0]), .bm_clkr(net244), .bm_clkw(net212),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sdo_i(bm_sdo_i),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(bm_sdi_o),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net295[0:7]),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl(vdd_cntl_bot[15:0]), .bl(bl[15:0]),
     .wl(wl_bot[15:0]), .reset_b(reset_b_bot[15:0]), .prog(prog),
     .pgate(pgate_bot[15:0]), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net295[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl(vdd_cntl_top[15:0]), .bl(bl[15:0]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl(wl_top[15:0]), .reset_b(reset_b_top[15:0]), .prog(prog),
     .pgate(pgate_top[15:0]), .op(slf_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net316[0:7]));
tielo I14 ( .tielo(net0226));
tielo I15 ( .tielo(net0227));
bram_routing_tracks4rev I5 ( .vdd_cntl(vdd_cntl_bot[15:0]),
     .s_r(net213), .wl(wl_bot[15:0]), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b(reset_b_bot[15:0]), .prog(prog), .pgate(pgate_bot[15:0]),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net0227), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[41:16]));
bram_routing_tracks4rev I3 ( .vdd_cntl(vdd_cntl_top[15:0]),
     .s_r(net245), .wl(wl_top[15:0]), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b(reset_b_top[15:0]), .prog(prog), .pgate(pgate_top[15:0]),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net0226), .bot_op(slf_op_bot[7:0]),
     .bnr_op(bnr_op_top[7:0]), .bnl_op(bnl_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[41:16]));

endmodule
// Library - ice4chip, Cell - CHIP_route_right0smc, View - schematic
// LAST TIME SAVED: Aug 28 14:38:45 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module CHIP_route_right0smc ( cm_banksel_blbrd_2_, cm_banksel_bldld,
     cm_banksel_bltrd1_3_, cm_clk_blbrd, cm_clk_bltrd1, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2d, cm_sdi_u3d2, cm_sdo_u3d1, cnt_podt_out,
     core_por_b0, core_por_b1, core_por_b_rowu2, core_por_b_rowu3,
     core_por_bb, cram_pgateoff, cram_prec, cram_prec_blbrd,
     cram_prec_bltrd1, cram_pullup_b,
     .cram_pullup_b_blbrd(cram_pullup_b_bldrd), cram_pullup_b_bltrd1,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, cram_write_blbrd,
     cram_write_bltrd1, data_muxsel1_blbrd, data_muxsel1_bltrd1,
     data_muxsel_blbrd, data_muxsel_bltrd1,
     .en_8bcibfig_b_bltrd1(en_8bconfig_b_bltrd1), en_8bconfig_b_blbrd,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, last_rsr,
     monitor_celldd, osc_clk, pgate_r, reset_b_r, smc_clk_out,
     smc_por_b0, smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd,
     smc_wdis_dclk_bltrd1, spi_ss_in_rd, vdd_cntl_r, wl_r, cf_r,
     cm_banksel, cm_sdi_u2, cm_sdi_u3, cm_sdo_u3, crst_filterout,
     data_muxsel, data_muxsel1, en_8bconfig_b, j_rst_b, j_tck,
     row_test0, smc_clk, smc_core_por_bottom1, smc_core_por_bottom2,
     smc_osco_fsel, smc_oscoff_b, smc_podt_off, smc_podt_rst, smc_read,
     smc_row_inc_fromsmc, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rsr_rst_fromsmc, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_wdis_dclk, smc_write, smc_write0, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en, spi_ss_in_r,
     u0_in, u1_in, vddio_rightbank );
output  cm_banksel_blbrd_2_, cm_banksel_bltrd1_3_, cm_clk_blbrd,
     cm_clk_bltrd1, cnt_podt_out, core_por_b0, core_por_b1,
     core_por_b_rowu2, core_por_b_rowu3, core_por_bb, cram_pgateoff,
     cram_prec, cram_prec_blbrd, cram_prec_bltrd1, cram_pullup_b,
     cram_pullup_b_bldrd, cram_pullup_b_bltrd1, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, cram_write_blbrd, cram_write_bltrd1,
     data_muxsel1_blbrd, data_muxsel1_bltrd1, data_muxsel_blbrd,
     data_muxsel_bltrd1, en_8bconfig_b_bltrd1, en_8bconfig_b_blbrd,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, osc_clk,
     smc_clk_out, smc_por_b0, smc_row_inc, smc_rsr_rst,
     smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1;

input  crst_filterout, data_muxsel, data_muxsel1, en_8bconfig_b,
     j_rst_b, j_tck, row_test0, smc_clk, smc_core_por_bottom1,
     smc_core_por_bottom2, smc_oscoff_b, smc_podt_off, smc_podt_rst,
     smc_read, smc_row_inc_fromsmc, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rsr_rst_fromsmc, smc_rwl_en, smc_seq_rst,
     smc_wcram_rst, smc_wdis_dclk, smc_write, smc_write0,
     smc_wset_prec, smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en,
     vddio_rightbank;

output [3:2]  monitor_celldd;
output [1:0]  cm_banksel_bldld;
output [1:0]  cm_sdi_u2d;
output [1:0]  cm_sdo_u3d1;
output [351:0]  wl_r;
output [1:0]  cm_sdi_u3d2;
output [7:1]  spi_ss_in_rd;
output [1:0]  cm_sdi_u1;
output [1:0]  last_rsr;
output [351:0]  reset_b_r;
output [351:0]  vdd_cntl_r;
output [351:0]  pgate_r;
output [1:0]  cm_sdi_u0;

input [1:0]  cm_sdo_u3;
input [7:1]  spi_ss_in_r;
input [1:0]  cm_sdi_u3;
input [3:0]  cm_banksel;
input [1:0]  u1_in;
input [1:0]  smc_osco_fsel;
input [1:0]  cm_sdi_u2;
input [1:0]  cf_r;
input [1:0]  u0_in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net0188;

wire  [1:0]  dff_out_top;

wire  [0:1]  net0187;

wire  [1:0]  cm_sdi_u3d0;

wire  [3:3]  monitor_celld2;

wire  [3:3]  cm_banksel_bltrd0;

wire  [1:0]  dff_out_bot;

wire  [3:3]  cm_banksel_bltrd;

wire  [1:0]  cm_sdo_u3d;

wire  [1:0]  cm_sdo_u3d0;

wire  [1:0]  cm_sdo_u3dd;

wire  [2:3]  monitor_celld;

wire  [3:3]  monitor_celld1;

wire  [1:0]  cm_sdi_u3d;



tielo I462_1_ ( .tielo(net0187[0]));
tielo I462_0_ ( .tielo(net0187[1]));
tielo I463_1_ ( .tielo(net0188[0]));
tielo I463_0_ ( .tielo(net0188[1]));
sg_bufx10 I460_1_ ( .in(cm_banksel[1]), .out(cm_banksel_bldld[1]));
sg_bufx10 I460_0_ ( .in(cm_banksel[0]), .out(cm_banksel_bldld[0]));
sg_bufx10 I307 ( .in(cram_pgateoff), .out(cram_pgateoffr0));
sg_bufx10 I208 ( .in(cm_banksel[3]), .out(cm_banksel_bltrd[3]));
sg_bufx10 I308 ( .in(cram_rst), .out(cram_rstr0));
sg_bufx10 I309 ( .in(cram_vddoff), .out(cram_vddoffr0));
sg_bufx10 I310 ( .in(cram_wl_en), .out(cram_wl_enr0));
sg_bufx10 I311 ( .in(smc_row_inc), .out(smc_row_incr0));
sg_bufx10 I151 ( .in(cram_prec), .out(cram_prec_blbrd));
sg_bufx10 I312 ( .in(smc_write0), .out(smc_writer0));
sg_bufx10 I315 ( .in(cram_pgateoffr0), .out(cram_pgateoffr1));
sg_bufx10 I201 ( .in(cm_banksel_bltrd[3]), .out(cm_banksel_bltrd0[3]));
sg_bufx10 I157 ( .in(smc_wdis_dclk), .out(smc_wdis_dclk_blbrd));
sg_bufx10 I431 ( .in(monitor_celld[3]), .out(monitor_celld1[3]));
sg_bufx10 I282_1_ ( .in(cm_sdi_u3d[1]), .out(cm_sdi_u3d0[1]));
sg_bufx10 I282_0_ ( .in(cm_sdi_u3d[0]), .out(cm_sdi_u3d0[0]));
sg_bufx10 I320 ( .in(smc_writer0), .out(smc_writer1));
sg_bufx10 I322 ( .in(tck_padr0), .out(tck_padr1));
sg_bufx10 I317 ( .in(cram_vddoffr0), .out(cram_vddoffr1));
sg_bufx10 I432 ( .in(cf_r[0]), .out(monitor_celld[2]));
sg_bufx10 I323 ( .in(row_test1), .out(row_testr1));
sg_bufx10 I455_1_ ( .in(dff_out_bot[1]), .out(cm_sdo_u3d0[1]));
sg_bufx10 I455_0_ ( .in(dff_out_bot[0]), .out(cm_sdo_u3d0[0]));
sg_bufx10 I207 ( .in(en_8bconfig_b_blbrd), .out(en_8bconfig_b_bltrd0));
sg_bufx10 I434_1_ ( .in(monitor_celld2[3]), .out(monitor_celldd[3]));
sg_bufx10 I434_0_ ( .in(monitor_celld[2]), .out(monitor_celldd[2]));
sg_bufx10 I210 ( .in(cram_write_bltrd0), .out(cram_write_bltrd1));
sg_bufx10 I205 ( .in(data_muxsel_blbrd), .out(data_muxsel_bltrd0));
sg_bufx10 I206 ( .in(cram_write_blbrd), .out(cram_write_bltrd0));
sg_bufx10 I153 ( .in(data_muxsel), .out(data_muxsel_blbrd));
sg_bufx10 I458_1_ ( .in(u0_in[1]), .out(cm_sdi_u0[1]));
sg_bufx10 I458_0_ ( .in(u0_in[0]), .out(cm_sdi_u0[0]));
sg_bufx10 I433 ( .in(monitor_celld1[3]), .out(monitor_celld2[3]));
sg_bufx10 I152 ( .in(cram_write), .out(cram_write_blbrd));
sg_bufx10 I304 ( .in(j_tck), .out(tck_padr0));
sg_bufx10 I319 ( .in(smc_row_incr0), .out(smc_row_incr1));
sg_bufx10 I457 ( .in(smc_rsr_rst_fromsmc), .out(smc_rsr_rst));
sg_bufx10 I454_1_ ( .in(dff_out_top[1]), .out(cm_sdo_u3dd[1]));
sg_bufx10 I454_0_ ( .in(dff_out_top[0]), .out(cm_sdo_u3dd[0]));
sg_bufx10 I198 ( .in(cram_pullup_b), .out(cram_pullup_b_bldrd));
sg_bufx10 I156 ( .in(smc_clk_out), .out(cm_clk_blbrd));
sg_bufx10 I150 ( .in(cm_banksel[2]), .out(cm_banksel_blbrd_2_));
sg_bufx10 I288_1_ ( .in(cm_sdo_u3d0[1]), .out(cm_sdo_u3d1[1]));
sg_bufx10 I288_0_ ( .in(cm_sdo_u3d0[0]), .out(cm_sdo_u3d1[0]));
sg_bufx10 I155 ( .in(en_8bconfig_b), .out(en_8bconfig_b_blbrd));
sg_bufx10 I115_1_ ( .in(cm_sdi_u2[1]), .out(cm_sdi_u2d[1]));
sg_bufx10 I115_0_ ( .in(cm_sdi_u2[0]), .out(cm_sdi_u2d[0]));
sg_bufx10 I116_1_ ( .in(cm_sdi_u3[1]), .out(cm_sdi_u3d[1]));
sg_bufx10 I116_0_ ( .in(cm_sdi_u3[0]), .out(cm_sdi_u3d[0]));
sg_bufx10 I154 ( .in(data_muxsel1), .out(data_muxsel1_blbrd));
sg_bufx10 I324 ( .in(smc_rsr_rstr0), .out(smc_rsr_rstr1));
sg_bufx10 I202 ( .in(cm_clk_blbrd), .out(cm_clk_bltrd0));
sg_bufx10 I459_1_ ( .in(u1_in[1]), .out(cm_sdi_u1[1]));
sg_bufx10 I459_0_ ( .in(u1_in[0]), .out(cm_sdi_u1[0]));
sg_bufx10 I203 ( .in(data_muxsel1_blbrd), .out(data_muxsel1_bltrd0));
sg_bufx10 I325 ( .in(core_por_bbr0), .out(core_por_b_rowu3));
sg_bufx10 I456 ( .in(smc_row_inc_fromsmc), .out(smc_row_inc));
sg_bufx10 I215 ( .in(cm_banksel_bltrd0[3]),
     .out(cm_banksel_bltrd1_3_));
sg_bufx10 I443 ( .in(j_rst_br0), .out(j_rst_br1));
sg_bufx10 I306 ( .in(row_test0), .out(row_test1));
sg_bufx10 I212 ( .in(smc_wdis_dclk_bltrd0),
     .out(smc_wdis_dclk_bltrd1));
sg_bufx10 I209 ( .in(en_8bconfig_b_bltrd0),
     .out(en_8bconfig_b_bltrd1));
sg_bufx10 I213 ( .in(data_muxsel1_bltrd0), .out(data_muxsel1_bltrd1));
sg_bufx10 I204 ( .in(smc_wdis_dclk_blbrd), .out(smc_wdis_dclk_bltrd0));
sg_bufx10 I200 ( .in(cram_prec_blbrd), .out(cram_prec_bltrd0));
sg_bufx10 I199 ( .in(cram_pullup_b_bldrd), .out(cram_pullup_b_bltrd0));
sg_bufx10 I211 ( .in(data_muxsel_bltrd0), .out(data_muxsel_bltrd1));
sg_bufx10 I217 ( .in(cram_pullup_b_bltrd0),
     .out(cram_pullup_b_bltrd1));
sg_bufx10 I440 ( .in(j_rst_b), .out(j_rst_br0));
sg_bufx10 I214 ( .in(cm_clk_bltrd0), .out(cm_clk_bltrd1));
sg_bufx10 I216 ( .in(cram_prec_bltrd0), .out(cram_prec_bltrd1));
sg_bufx10 I305 ( .in(smc_rsr_rst), .out(smc_rsr_rstr0));
sg_bufx10 I285_1_ ( .in(cm_sdo_u3[1]), .out(cm_sdo_u3d[1]));
sg_bufx10 I285_0_ ( .in(cm_sdo_u3[0]), .out(cm_sdo_u3d[0]));
sg_bufx10 I318 ( .in(cram_wl_enr0), .out(cram_wl_enr1));
sg_bufx10 I283_1_ ( .in(cm_sdi_u3d0[1]), .out(cm_sdi_u3d2[1]));
sg_bufx10 I283_0_ ( .in(cm_sdi_u3d0[0]), .out(cm_sdi_u3d2[0]));
sg_bufx10 I314 ( .in(core_por_bb), .out(core_por_bbr0));
sg_bufx10 I316 ( .in(cram_rstr0), .out(cram_rstr1));
sg_bufx10 I430 ( .in(cf_r[1]), .out(monitor_celld[3]));
inv_hvt I136 ( .A(core_por_b0), .Y(core_por_bb));
ml_osc_top Iml_osc ( .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]), .por_b(core_por_b0),
     .crst_b(crst_filterout), .smc_clk(osc_clk),
     .cnt_podt_out(cnt_podt_out));
ml_rowdrv_bank Irowur ( .smc_write(smc_write_rowu3),
     .smc_rsr_inc(smc_row_inc_rowu3), .rsr_rst(smc_rsr_rst_rowu3),
     .por_rst(core_por_b_rowu3), .cram_wl_en(cram_wl_en_rowu3),
     .cram_vddoff(cram_vddoff_rowu3), .cram_rst(cram_rst_rowu3),
     .cram_pgateoff(cram_pgateoff_rowu3),
     .banksel(cm_banksel_bltrd0[3]), .vddctrl(vdd_cntl_r[351:176]),
     .last_rsr(last_rsr[1]), .reset(reset_b_r[351:176]),
     .pgate(pgate_r[351:176]), .trst_b(j_rst_b_rowu3),
     .jtag_rowtest_rst(row_test_rowu3), .jtag_clk(tck_pad_rowu3),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu3_b),
     .wl(wl_r[351:176]));
ml_rowdrv_bank Irowlr ( .smc_write(smc_write_rowu2),
     .smc_rsr_inc(smc_row_inc_rowu2), .rsr_rst(smc_rsr_rst_rowu2),
     .por_rst(core_por_b_rowu2), .cram_wl_en(cram_wl_en_rowu2),
     .cram_vddoff(cram_vddoff_rowu2), .cram_rst(cram_rst_rowu2),
     .cram_pgateoff(cram_pgateoff_rowu2),
     .banksel(cm_banksel_blbrd_2_), .vddctrl(vdd_cntl_r[175:0]),
     .last_rsr(last_rsr[0]), .reset(reset_b_r[175:0]),
     .pgate(pgate_r[175:0]), .trst_b(j_rst_b_rowu2),
     .jtag_rowtest_rst(row_test_rowu2), .jtag_clk(tck_pad_rowu2),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu2_b),
     .wl(wl_r[175:0]));
sg_dffbuf I286_1_ ( .r(net0187[0]), .d(cm_sdo_u3d[1]), .clk(net373),
     .dffout(dff_out_top[1]));
sg_dffbuf I286_0_ ( .r(net0187[1]), .d(cm_sdo_u3d[0]), .clk(net373),
     .dffout(dff_out_top[0]));
sg_dffbuf I453_1_ ( .r(net0188[0]), .d(cm_sdo_u3dd[1]), .clk(net375),
     .dffout(dff_out_bot[1]));
sg_dffbuf I453_0_ ( .r(net0188[1]), .d(cm_sdo_u3dd[0]), .clk(net375),
     .dffout(dff_out_bot[0]));
bram_bufferx16 I407 ( .in(cram_wl_enr0), .out(cram_wl_en_rowu2));
bram_bufferx16 I416 ( .in(cram_rstr1), .out(cram_rst_rowu3));
bram_bufferx16 I185 ( .in(core_por_b0), .out(core_por_b1));
bram_bufferx16 I442 ( .in(j_rst_br1), .out(j_rst_b_rowu3));
bram_bufferx16 I441 ( .in(j_rst_br0), .out(j_rst_b_rowu2));
bram_bufferx16 I409 ( .in(smc_writer0), .out(smc_write_rowu2));
bram_bufferx16 I287 ( .in(cm_clk_bltrd0), .out(net373));
bram_bufferx16 I452 ( .in(smc_clk_out), .out(net375));
bram_bufferx16 I451_6_ ( .in(spi_ss_in_r[7]), .out(spi_ss_in_rd[7]));
bram_bufferx16 I451_5_ ( .in(spi_ss_in_r[6]), .out(spi_ss_in_rd[6]));
bram_bufferx16 I451_4_ ( .in(spi_ss_in_r[5]), .out(spi_ss_in_rd[5]));
bram_bufferx16 I451_3_ ( .in(spi_ss_in_r[4]), .out(spi_ss_in_rd[4]));
bram_bufferx16 I451_2_ ( .in(spi_ss_in_r[3]), .out(spi_ss_in_rd[3]));
bram_bufferx16 I451_1_ ( .in(spi_ss_in_r[2]), .out(spi_ss_in_rd[2]));
bram_bufferx16 I451_0_ ( .in(spi_ss_in_r[1]), .out(spi_ss_in_rd[1]));
bram_bufferx16 I402 ( .in(smc_rsr_rstr0), .out(smc_rsr_rst_rowu2));
bram_bufferx16 I410 ( .in(core_por_bbr0), .out(core_por_b_rowu2));
bram_bufferx16 I406 ( .in(cram_vddoffr0), .out(cram_vddoff_rowu2));
bram_bufferx16 I405 ( .in(cram_rstr0), .out(cram_rst_rowu2));
bram_bufferx16 I401 ( .in(tck_padr0), .out(tck_pad_rowu2));
bram_bufferx16 I403 ( .in(row_test1), .out(row_test_rowu2));
bram_bufferx16 I420 ( .in(tck_padr1), .out(tck_pad_rowu3));
bram_bufferx16 I418 ( .in(row_testr1), .out(row_test_rowu3));
bram_bufferx16 I408 ( .in(smc_row_incr0), .out(smc_row_inc_rowu2));
bram_bufferx16 I404 ( .in(cram_pgateoffr0), .out(cram_pgateoff_rowu2));
bram_bufferx16 I412 ( .in(smc_writer1), .out(smc_write_rowu3));
bram_bufferx16 I414 ( .in(cram_wl_enr1), .out(cram_wl_en_rowu3));
bram_bufferx16 I413 ( .in(smc_row_incr1), .out(smc_row_inc_rowu3));
bram_bufferx16 I417 ( .in(cram_pgateoffr1), .out(cram_pgateoff_rowu3));
bram_bufferx16 I419 ( .in(smc_rsr_rstr1), .out(smc_rsr_rst_rowu3));
bram_bufferx16 I415 ( .in(cram_vddoffr1), .out(cram_vddoff_rowu3));
ml_cram_logic Iml_cram_logic ( .smc_wwlwrt_en(smc_wwlwrt_en),
     .smc_wset_precgnd(smc_wset_precgnd), .smc_write(smc_write),
     .cram_pgateoff(cram_pgateoff), .smc_wcram_rst(smc_wcram_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rrst_pullwlen(smc_rrst_pullwlen),
     .smc_rpull_b(smc_rpull_b), .smc_rprec(smc_rprec),
     .smc_read(smc_read), .smc_clk(smc_clk), .por(core_por_bb),
     .cram_write(cram_write), .cram_wl_en(cram_wl_en),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_vddoff(cram_vddoff),
     .smc_seq_rst(smc_seq_rst), .smc_clk_out(smc_clk_out),
     .smc_wwlwrt_dis(smc_wwlwrt_dis), .smc_wset_prec(smc_wset_prec));
SMC_CORE_POR_right I450 ( .vddio_rightbank(vddio_rightbank),
     .smc_por_b(smc_por_b0), .core_por_b(core_por_b0),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbank_pbuffer_top, View -
//schematic
// LAST TIME SAVED: Aug 24 17:33:08 2007
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [7:0]  bm_sa_o;

input [15:0]  bm_bweb;
input [7:0]  bm_aa;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbank, View - schematic
// LAST TIME SAVED: Aug 22 17:36:22 2007
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module bram_4kprouting_tbank ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_bot;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_v_t_top;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_h_r_top;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_r_v_b_bot;

input [15:0]  wl_top;
input [7:0]  lft_op_top;
input [15:0]  pgate_top;
input [7:0]  bnl_op_top;
input [7:0]  rgt_op_bot;
input [7:0]  bnr_op_top;
input [7:0]  rgt_op_top;
input [7:0]  bnl_op_bot;
input [7:0]  lft_op_bot;
input [7:0]  tnr_op_top;
input [7:0]  top_op_top;
input [15:0]  pgate_bot;
input [7:0]  tnl_op_top;
input [7:0]  bot_op_bot;
input [7:0]  tnr_op_bot;
input [15:0]  vdd_cntl_top;
input [15:0]  vdd_cntl_bot;
input [7:0]  glb_netwk;
input [15:0]  wl_bot;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_bot;
input [7:0]  bnr_op_bot;
input [15:0]  reset_b_top;
input [15:0]  reset_b_bot;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net208;

wire  [0:7]  net316;

wire  [0:7]  net242;

wire  [0:7]  net241;

wire  [0:7]  net243;

wire  [0:7]  net240;

wire  [0:7]  net295;

wire  [0:7]  net211;

wire  [0:7]  net210;

wire  [0:7]  net209;



bram_4kbank_pbuffer_top I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net245), .bm_wen(net213),
     .bm_d(bm_d[15:0]), .bm_clkr(net244), .bm_clkw(net212),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sdo_i(bm_sdo_i),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(bm_sdi_o),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net295[0:7]),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl(vdd_cntl_bot[15:0]), .bl(bl[15:0]),
     .wl(wl_bot[15:0]), .reset_b(reset_b_bot[15:0]), .prog(prog),
     .pgate(pgate_bot[15:0]), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net295[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl(vdd_cntl_top[15:0]), .bl(bl[15:0]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl(wl_top[15:0]), .reset_b(reset_b_top[15:0]), .prog(prog),
     .pgate(pgate_top[15:0]), .op(slf_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net316[0:7]));
tielo I14 ( .tielo(net0226));
tielo I15 ( .tielo(net0227));
bram_routing_tracks4rev I5 ( .vdd_cntl(vdd_cntl_bot[15:0]),
     .s_r(net213), .wl(wl_bot[15:0]), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b(reset_b_bot[15:0]), .prog(prog), .pgate(pgate_bot[15:0]),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net0227), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[41:16]));
bram_routing_tracks4rev I3 ( .vdd_cntl(vdd_cntl_top[15:0]),
     .s_r(net245), .wl(wl_top[15:0]), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b(reset_b_top[15:0]), .prog(prog), .pgate(pgate_top[15:0]),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net0226), .bot_op(slf_op_bot[7:0]),
     .bnr_op(bnr_op_top[7:0]), .bnl_op(bnl_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[41:16]));

endmodule
// Library - BRAM_WRAPPER, Cell - bram_4kbankout_pbuffer_top, View -
//schematic
// LAST TIME SAVED: Aug 24 17:34:59 2007
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module bram_4kbankout_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_aa;
input [7:0]  bm_sa_i;
input [7:0]  bm_ab;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_bankout I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbankout, View -
//schematic
// LAST TIME SAVED: Aug 22 17:39:11 2007
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module bram_4kprouting_tbankout ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_bot;
inout [41:0]  bl;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_r_top;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [23:0]  sp12_h_l_top;

input [15:0]  reset_b_top;
input [15:0]  pgate_top;
input [7:0]  bnr_op_top;
input [15:0]  vdd_cntl_top;
input [7:0]  rgt_op_bot;
input [15:0]  pgate_bot;
input [7:0]  lft_op_top;
input [7:0]  glb_netwk;
input [15:0]  vdd_cntl_bot;
input [7:0]  tnr_op_top;
input [7:0]  rgt_op_top;
input [7:0]  top_op_top;
input [7:0]  tnr_op_bot;
input [7:0]  bot_op_bot;
input [7:0]  bnl_op_top;
input [7:0]  bnr_op_bot;
input [7:0]  bnl_op_bot;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_bot;
input [15:0]  reset_b_bot;
input [7:0]  lft_op_bot;
input [7:0]  tnl_op_top;
input [15:0]  wl_bot;
input [15:0]  wl_top;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net208;

wire  [0:7]  net316;

wire  [0:7]  net242;

wire  [0:7]  net241;

wire  [0:7]  net243;

wire  [0:7]  net240;

wire  [0:7]  net295;

wire  [0:7]  net210;

wire  [0:7]  net211;

wire  [0:7]  net209;



bram_4kbankout_pbuffer_top I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net245), .bm_wen(net213),
     .bm_d(bm_d[15:0]), .bm_clkr(net244), .bm_clkw(net212),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sdo_i(bm_sdo_i),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(bm_sdi_o),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net295[0:7]),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl(vdd_cntl_bot[15:0]), .bl(bl[15:0]),
     .wl(wl_bot[15:0]), .reset_b(reset_b_bot[15:0]), .prog(prog),
     .pgate(pgate_bot[15:0]), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net295[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl(vdd_cntl_top[15:0]), .bl(bl[15:0]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl(wl_top[15:0]), .reset_b(reset_b_top[15:0]), .prog(prog),
     .pgate(pgate_top[15:0]), .op(slf_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net316[0:7]));
tielo I14 ( .tielo(net0226));
tielo I15 ( .tielo(net0227));
bram_routing_tracks4rev I5 ( .vdd_cntl(vdd_cntl_bot[15:0]),
     .s_r(net213), .wl(wl_bot[15:0]), .top_op(slf_op_top[7:0]),
     .tnr_op(tnr_op_bot[7:0]), .tnl_op(tnl_op_bot[7:0]),
     .slf_op(slf_op_bot[7:0]), .rgt_op(rgt_op_bot[7:0]),
     .reset_b(reset_b_bot[15:0]), .prog(prog), .pgate(pgate_bot[15:0]),
     .lft_op(lft_op_bot[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net0227), .bot_op(bot_op_bot[7:0]),
     .bnr_op(bnr_op_bot[7:0]), .bnl_op(bnl_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[41:16]));
bram_routing_tracks4rev I3 ( .vdd_cntl(vdd_cntl_top[15:0]),
     .s_r(net245), .wl(wl_top[15:0]), .top_op(top_op_top[7:0]),
     .tnr_op(tnr_op_top[7:0]), .tnl_op(tnl_op_top[7:0]),
     .slf_op(slf_op_top[7:0]), .rgt_op(rgt_op_top[7:0]),
     .reset_b(reset_b_top[15:0]), .prog(prog), .pgate(pgate_top[15:0]),
     .lft_op(lft_op_top[7:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net0226), .bot_op(slf_op_bot[7:0]),
     .bnr_op(bnr_op_top[7:0]), .bnl_op(bnl_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[41:16]));

endmodule
// Library - io, Cell - io_col4, View - schematic
// LAST TIME SAVED: Feb  8 13:37:35 2008
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module io_col4 ( cf, fabric_out, padeb, pado, sdo, slf_op, spi_ss_in_b,
     bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op, bs_en, cdone_in,
     ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin, pgate, prog, r,
     reset, sdi, shift, spioeb, spiout, tclk, tnl_op, update, vdd_cntl,
     wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  spi_ss_in_b;
output [1:0]  pado;
output [1:0]  padeb;
output [23:0]  cf;
output [3:0]  slf_op;

inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;

input [1:0]  padin;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [1:0]  spioeb;
input [15:0]  wl;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [7:0]  lft_op;
input [1:0]  spiout;
input [15:0]  reset;
input [7:0]  glb_netwk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



rm6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[17:14],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, pgate[15:0], prog, reset[15:0], vdd_cntl[15:0],
     wl[15:0]);
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl(vdd_cntl[15:0]),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[13:8]), .wl(wl[15:0]),
     .reset(reset[15:0]), .pgate(pgate[15:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(prog),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl(vdd_cntl[15:0]), .outclk(outclk),
     .fabric_out(fabric_out), .min6({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .inclk_in({lc_trk_g1[3],
     lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0], glb_netwk[7:0]}),
     .ceb_in({lc_trk_g1[5], lc_trk_g1[2], lc_trk_g0[5], lc_trk_g0[2],
     glb_netwk[6], glb_netwk[4], glb_netwk[2], glb_netwk[0]}),
     .clk_in({lc_trk_g1[4], lc_trk_g1[1], lc_trk_g0[4], lc_trk_g0[1],
     glb_netwk[7:0]}), .update(update), .spiout(spiout[1:0]),
     .spioeb(spioeb[1:0]), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[7:2]), .inclk(inclk), .wl(wl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]), .prog(prog));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl(vdd_cntl[15:0]),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl(wl[15:0]), .reset(reset[15:0]), .pgate(pgate[15:0]),
     .hiz_b(hiz_b), .update(enable_update), .ti(ti[5:0]), .tclk(tclk),
     .shift(shift), .sdi(sdi), .prog(prog), .padin(padin[1:0]),
     .mode(mode), .inclk(inclk), .bs_en(bs_en),
     .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo), .pado(om[1:0]),
     .padeb(oenm[1:0]), .bl(bl[1:0]));

endmodule
// Library - leafcell, Cell - QUAD_TR, View - schematic
// LAST TIME SAVED: Sep 15 14:06:50 2008
// NETLIST TIME: Nov 14 16:12:03 2008
`timescale 1ns / 1ns 

module QUAD_TR ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, ceb_o, cf_r, cf_t, fabric_out_163,
     fabric_out_168, fabric_out_223, hiz_b_o, io_r_00_24_11, mode_o,
     padeb_r, padeb_t, padin_163, padin_223, pado_r, pado_t, r_o, sdo,
     shift_o, slf_op_13_02, slf_op_13_03, slf_op_13_04, slf_op_13_05,
     slf_op_13_06, slf_op_13_07, slf_op_13_08, slf_op_13_09,
     slf_op_13_10, slf_op_13_11, slf_op_13_21, slf_op_14_11,
     slf_op_15_11, slf_op_16_11, slf_op_17_11, slf_op_18_11,
     slf_op_19_11, slf_op_20_11, slf_op_21_11, slf_op_22_11,
     slf_op_23_11, slf_op_24_11, spi_ss_in_r, tclk_o, update_o, bl,
     sp4_h_l_13_01, sp4_h_l_13_02, sp4_h_l_13_03, sp4_h_l_13_04,
     sp4_h_l_13_05, sp4_h_l_13_06, sp4_h_l_13_07, sp4_h_l_13_08,
     sp4_h_l_13_09, sp4_h_l_13_10, sp4_h_l_13_21, sp4_v_b_13_02,
     sp4_v_b_13_03, sp4_v_b_13_04, sp4_v_b_13_05, sp4_v_b_13_06,
     sp4_v_b_13_07, sp4_v_b_13_08, sp4_v_b_13_09, sp4_v_b_13_10,
     sp4_v_b_13_11, sp4_v_b_14_11, sp4_v_b_15_11, sp4_v_b_16_11,
     sp4_v_b_17_11, sp4_v_b_18_11, sp4_v_b_19_11, sp4_v_b_20_11,
     sp4_v_b_21_11, sp4_v_b_22_11, sp4_v_b_23_11, sp4_v_b_24_11,
     sp4_v_b_25_11, sp12_h_l_13_01, sp12_h_l_13_02, sp12_h_l_13_03,
     sp12_h_l_13_04, sp12_h_l_13_05, sp12_h_l_13_06, sp12_h_l_13_07,
     sp12_h_l_13_08, sp12_h_l_13_09, sp12_h_l_13_10, sp12_v_b_13_11,
     sp12_v_b_14_11, sp12_v_b_15_11, sp12_v_b_16_11, sp12_v_b_17_11,
     sp12_v_b_18_11, sp12_v_b_19_11, sp12_v_b_20_11, sp12_v_b_21_11,
     sp12_v_b_22_11, sp12_v_b_23_11, sp12_v_b_24_11, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_13_11,
     bnl_op_14_11, bnl_op_15_11, bnl_op_16_11, bnl_op_17_11,
     bnl_op_18_11, bnl_op_19_11, bnl_op_20_11, bnl_op_21_11,
     bnl_op_22_11, bnl_op_23_11, bnl_op_24_11, bnl_op_25_11,
     bnr_op_13_11, bnr_op_14_11, bnr_op_15_11, bnr_op_16_11,
     bnr_op_17_11, bnr_op_18_11, bnr_op_19_11, bnr_op_20_11,
     bnr_op_21_11, bnr_op_22_11, bnr_op_23_11, bnr_op_24_11,
     bot_op_13_11, bot_op_14_11, bot_op_15_11, bot_op_16_11,
     bot_op_17_11, bot_op_18_11, bot_op_19_11, bot_op_20_11,
     bot_op_21_11, bot_op_22_11, bot_op_23_11, bot_op_24_11, bs_en_i,
     carry_in_13_11, carry_in_14_11, carry_in_15_11, carry_in_16_11,
     carry_in_17_11, carry_in_18_11, carry_in_20_11, carry_in_21_11,
     carry_in_22_11, carry_in_23_11, carry_in_24_11, ceb_i,
     end_of_startup_r, end_of_startup_top_r, glb_in, hiz_b_i, hold_r_t,
     hold_t_r, lft_op_13_01, lft_op_13_02, lft_op_13_03, lft_op_13_04,
     lft_op_13_05, lft_op_13_06, lft_op_13_07, lft_op_13_08,
     lft_op_13_09, lft_op_13_10, mode_i, padin_r, padin_t, pgate, prog,
     purst, r_i, reset_b, sdi, shift_i, tclk_i, tiegnd, tievdd,
     tnl_op_13_20, update_i, vdd_cntl, wl );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bs_en_o, ceb_o,
     fabric_out_163, fabric_out_168, fabric_out_223, hiz_b_o, mode_o,
     padin_163, padin_223, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en_i,
     carry_in_13_11, carry_in_14_11, carry_in_15_11, carry_in_16_11,
     carry_in_17_11, carry_in_18_11, carry_in_20_11, carry_in_21_11,
     carry_in_22_11, carry_in_23_11, carry_in_24_11, ceb_i, hiz_b_i,
     hold_r_t, hold_t_r, mode_i, prog, purst, r_i, sdi, shift_i,
     tclk_i, tiegnd, tievdd, update_i;

output [7:0]  slf_op_13_10;
output [7:0]  slf_op_14_11;
output [7:0]  slf_op_20_11;
output [7:0]  slf_op_13_06;
output [7:0]  slf_op_13_08;
output [7:0]  slf_op_23_11;
output [7:0]  slf_op_22_11;
output [7:0]  slf_op_13_04;
output [7:0]  slf_op_13_03;
output [7:0]  slf_op_13_05;
output [7:0]  slf_op_24_11;
output [3:0]  io_r_00_24_11;
output [7:0]  bm_sa_o;
output [39:20]  padeb_r;
output [7:0]  slf_op_21_11;
output [47:24]  padeb_t;
output [575:288]  cf_t;
output [47:24]  pado_t;
output [7:0]  slf_op_13_07;
output [39:20]  spi_ss_in_r;
output [479:240]  cf_r;
output [3:0]  slf_op_13_21;
output [39:20]  pado_r;
output [7:0]  slf_op_18_11;
output [7:0]  slf_op_13_11;
output [7:0]  slf_op_13_02;
output [7:0]  slf_op_19_11;
output [7:0]  slf_op_15_11;
output [7:0]  slf_op_13_09;
output [7:0]  slf_op_16_11;
output [7:0]  slf_op_17_11;

inout [47:0]  sp4_v_b_13_03;
inout [47:0]  sp4_v_b_13_02;
inout [23:0]  sp12_h_l_13_03;
inout [23:0]  sp12_v_b_22_11;
inout [23:0]  sp12_h_l_13_06;
inout [23:0]  sp12_h_l_13_02;
inout [23:0]  sp12_h_l_13_10;
inout [23:0]  sp12_h_l_13_09;
inout [47:0]  sp4_h_l_13_06;
inout [47:0]  sp4_v_b_20_11;
inout [23:0]  sp12_h_l_13_05;
inout [23:0]  sp12_h_l_13_07;
inout [23:0]  sp12_v_b_23_11;
inout [47:0]  sp4_h_l_13_10;
inout [15:0]  sp4_v_b_25_11;
inout [47:0]  sp4_v_b_15_11;
inout [47:0]  sp4_v_b_18_11;
inout [47:0]  sp4_v_b_14_11;
inout [23:0]  sp12_v_b_16_11;
inout [47:0]  sp4_v_b_13_10;
inout [47:0]  sp4_v_b_13_06;
inout [23:0]  sp12_v_b_13_11;
inout [47:0]  sp4_h_l_13_04;
inout [47:0]  sp4_v_b_23_11;
inout [47:0]  sp4_v_b_13_04;
inout [47:0]  sp4_v_b_13_07;
inout [47:0]  sp4_v_b_17_11;
inout [15:0]  sp4_h_l_13_21;
inout [23:0]  sp12_v_b_24_11;
inout [47:0]  sp4_h_l_13_09;
inout [23:0]  sp12_v_b_20_11;
inout [23:0]  sp12_h_l_13_08;
inout [47:0]  sp4_v_b_13_11;
inout [47:0]  sp4_v_b_16_11;
inout [47:0]  sp4_h_l_13_02;
inout [47:0]  sp4_v_b_13_09;
inout [1311:658]  bl;
inout [23:0]  sp12_h_l_13_04;
inout [47:0]  sp4_v_b_13_05;
inout [47:0]  sp4_v_b_19_11;
inout [47:0]  sp4_v_b_24_11;
inout [23:0]  sp12_v_b_21_11;
inout [47:0]  sp4_h_l_13_08;
inout [47:0]  sp4_h_l_13_03;
inout [47:0]  sp4_v_b_22_11;
inout [23:0]  sp12_v_b_15_11;
inout [23:0]  sp12_v_b_14_11;
inout [47:0]  sp4_h_l_13_07;
inout [23:0]  sp12_h_l_13_01;
inout [47:0]  sp4_v_b_13_08;
inout [23:0]  sp12_v_b_19_11;
inout [23:0]  sp12_v_b_18_11;
inout [47:0]  sp4_h_l_13_05;
inout [23:0]  sp12_v_b_17_11;
inout [47:0]  sp4_h_l_13_01;
inout [47:0]  sp4_v_b_21_11;

input [7:0]  lft_op_13_07;
input [7:0]  bnl_op_24_11;
input [7:0]  bnr_op_21_11;
input [7:0]  bnr_op_14_11;
input [7:0]  lft_op_13_03;
input [7:0]  bot_op_24_11;
input [7:0]  lft_op_13_08;
input [7:0]  bnl_op_20_11;
input [7:0]  bot_op_18_11;
input [7:0]  bnr_op_18_11;
input [7:0]  lft_op_13_10;
input [7:0]  lft_op_13_05;
input [7:0]  bm_sa_i;
input [7:0]  bnl_op_14_11;
input [7:0]  bnr_op_13_11;
input [9:0]  end_of_startup_r;
input [7:0]  bnl_op_16_11;
input [7:0]  bnr_op_24_11;
input [7:0]  lft_op_13_09;
input [7:0]  bnl_op_25_11;
input [7:0]  bot_op_20_11;
input [7:0]  bnr_op_16_11;
input [3:0]  tnl_op_13_20;
input [7:0]  bot_op_15_11;
input [7:0]  bot_op_19_11;
input [7:0]  lft_op_13_06;
input [7:0]  lft_op_13_02;
input [351:176]  pgate;
input [351:176]  vdd_cntl;
input [351:176]  wl;
input [7:0]  bnr_op_17_11;
input [7:0]  bnr_op_22_11;
input [7:0]  bot_op_14_11;
input [47:24]  padin_t;
input [7:0]  bot_op_13_11;
input [7:0]  lft_op_13_01;
input [7:0]  bnl_op_23_11;
input [351:176]  reset_b;
input [7:0]  bnl_op_15_11;
input [7:0]  bnl_op_21_11;
input [7:0]  bnr_op_23_11;
input [7:0]  bnr_op_19_11;
input [7:0]  bnl_op_13_11;
input [7:0]  glb_in;
input [7:0]  bot_op_21_11;
input [24:13]  end_of_startup_top_r;
input [7:0]  bnr_op_20_11;
input [7:0]  bnl_op_18_11;
input [7:0]  bot_op_23_11;
input [7:0]  bot_op_22_11;
input [7:0]  bnl_op_17_11;
input [7:0]  bnr_op_15_11;
input [7:0]  lft_op_13_04;
input [7:0]  bnl_op_19_11;
input [39:20]  padin_r;
input [7:0]  bot_op_17_11;
input [7:0]  bot_op_16_11;
input [7:0]  bnl_op_22_11;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:47]  net_5331;

wire  [0:23]  net_6027;

wire  [0:7]  net_4031;

wire  [0:23]  net_4601;

wire  [0:7]  net_8055;

wire  [3:0]  io_t_24;

wire  [3:0]  slf_op_25_10;

wire  [3:0]  io_r_07;

wire  [0:1]  net_7542;

wire  [3:0]  io_t_23;

wire  [0:23]  net_6727;

wire  [0:47]  net_4320;

wire  [0:23]  net_6559;

wire  [0:23]  net_5635;

wire  [3:0]  io_r_08;

wire  [0:23]  net_4627;

wire  [0:15]  net_7820;

wire  [0:23]  net_4937;

wire  [0:7]  net_4783;

wire  [0:7]  net_4729;

wire  [0:47]  net_6336;

wire  [3:0]  io_r_06;

wire  [0:47]  net_4294;

wire  [3:0]  io_t_22;

wire  [3:0]  io_t_21;

wire  [3:0]  io_r_03;

wire  [3:0]  io_r_05;

wire  [3:0]  io_r_01;

wire  [3:0]  io_r_02;

wire  [3:0]  io_r_04;

wire  [3:0]  io_t_17;

wire  [3:0]  io_t_20;

wire  [3:0]  io_t_15;

wire  [3:0]  io_t_19;

wire  [3:0]  io_t_14;

wire  [3:0]  io_t_16;

wire  [7:0]  net2col_drivers;

wire  [7:0]  glb_netwk_13;

wire  [7:0]  glb_netwk_14;

wire  [7:0]  glb_netwk_15;

wire  [7:0]  glb_netwk_16;

wire  [7:0]  glb_netwk_17;

wire  [7:0]  glb_netwk_18;

wire  [7:0]  glb_netwk_19;

wire  [7:0]  glb_netwk_20;

wire  [7:0]  glb_netwk_21;

wire  [7:0]  glb_netwk_22;

wire  [7:0]  glb_netwk_23;

wire  [7:0]  glb_netwk_24;

wire  [7:0]  glb_netwk_io_r;

wire  [3:0]  io_t_18;

wire  [0:7]  net_6239;

wire  [0:47]  net_5303;

wire  [0:47]  net_7263;

wire  [0:7]  net_5931;

wire  [0:7]  net_8157;

wire  [0:23]  net_5215;

wire  [0:23]  net_6307;

wire  [0:47]  net_4202;

wire  [0:47]  net_5300;

wire  [0:23]  net_5887;

wire  [0:7]  net_5427;

wire  [0:23]  net_4741;

wire  [0:1]  net_7610;

wire  [0:47]  net_5415;

wire  [0:15]  net_8082;

wire  [0:23]  net_6225;

wire  [0:23]  net_6505;

wire  [0:47]  net_6140;

wire  [0:23]  net_5271;

wire  [0:47]  net_6115;

wire  [0:47]  net_4883;

wire  [0:7]  net_4689;

wire  [0:47]  net_7375;

wire  [0:7]  net_6015;

wire  [0:23]  net_6001;

wire  [0:23]  net_5917;

wire  [0:23]  net_5859;

wire  [0:47]  net_4908;

wire  [0:47]  net_6367;

wire  [0:47]  net_6252;

wire  [0:47]  net_7092;

wire  [0:47]  net_7067;

wire  [0:23]  net_4405;

wire  [0:15]  net_7572;

wire  [0:47]  net_5443;

wire  [0:23]  net_5133;

wire  [0:47]  net_6395;

wire  [0:23]  net_4851;

wire  [0:47]  net_5023;

wire  [0:23]  net_5159;

wire  [0:47]  net_5580;

wire  [0:47]  net_5916;

wire  [0:7]  net_6267;

wire  [0:7]  net_4839;

wire  [0:23]  net_4823;

wire  [0:7]  net_5651;

wire  [0:23]  net_6113;

wire  [0:47]  net_6672;

wire  [0:23]  net_5663;

wire  [0:47]  net_6644;

wire  [0:23]  net_5915;

wire  [0:7]  net_5007;

wire  [0:47]  net_6952;

wire  [0:47]  net_4348;

wire  [0:47]  net_6535;

wire  [0:47]  net_4575;

wire  [0:23]  net_6897;

wire  [0:47]  net_4120;

wire  [0:7]  net_4138;

wire  [0:23]  net_4515;

wire  [0:7]  net_4867;

wire  [0:47]  net_6392;

wire  [0:23]  net_4116;

wire  [0:23]  net_7091;

wire  [0:23]  net_5553;

wire  [0:47]  net_4936;

wire  [0:7]  net_6043;

wire  [0:15]  net_7878;

wire  [0:47]  net_5751;

wire  [0:23]  net_6419;

wire  [0:47]  net_4827;

wire  [0:23]  net_4713;

wire  [0:23]  net_4881;

wire  [0:7]  net_6435;

wire  [0:23]  net_4200;

wire  [0:23]  net_7231;

wire  [0:47]  net_4771;

wire  [0:23]  net_5327;

wire  [0:47]  net_4295;

wire  [0:23]  net_6925;

wire  [0:23]  net_5469;

wire  [0:23]  net_4573;

wire  [0:23]  net_7147;

wire  [0:23]  net_6055;

wire  [0:23]  net_6279;

wire  [0:47]  net_5359;

wire  [0:23]  net_4935;

wire  [0:7]  net_6351;

wire  [0:47]  net_5807;

wire  [0:23]  net_4034;

wire  [0:47]  net_4687;

wire  [0:47]  net_7811;

wire  [0:47]  net_4992;

wire  [0:47]  net_7291;

wire  [0:47]  net_4852;

wire  [0:47]  net_5048;

wire  [0:7]  net_5763;

wire  [0:23]  net_5637;

wire  [0:47]  net_5244;

wire  [0:47]  net_5160;

wire  [0:47]  net_7471;

wire  [0:47]  net_6616;

wire  [0:47]  net_4712;

wire  [0:47]  net_5387;

wire  [0:7]  net_6463;

wire  [0:7]  net_6183;

wire  [0:7]  net_4113;

wire  [0:7]  net_6071;

wire  [0:15]  net_8014;

wire  [0:47]  net_6924;

wire  [0:23]  net_4161;

wire  [0:47]  net_7319;

wire  [0:7]  net_5679;

wire  [0:23]  net_5775;

wire  [0:15]  net_7752;

wire  [0:23]  net_6671;

wire  [0:23]  net_4038;

wire  [0:47]  net_6532;

wire  [0:23]  net_5131;

wire  [0:1]  net_7508;

wire  [0:23]  net_6841;

wire  [0:23]  net_6643;

wire  [0:7]  net_6407;

wire  [0:47]  net_5639;

wire  [0:7]  net_7715;

wire  [0:23]  net_7315;

wire  [0:7]  net_5735;

wire  [0:47]  net_6087;

wire  [0:47]  net_6003;

wire  [0:47]  net_5611;

wire  [0:47]  net_5524;

wire  [0:7]  net_5177;

wire  [0:23]  net_5609;

wire  [0:23]  net_4461;

wire  [0:7]  net_7511;

wire  [0:7]  net_5035;

wire  [0:23]  net_7259;

wire  [0:23]  net_5441;

wire  [0:7]  net_5707;

wire  [0:7]  net_4155;

wire  [0:23]  net_7345;

wire  [0:23]  net_4226;

wire  [0:23]  net_5665;

wire  [0:23]  net_6169;

wire  [0:7]  net_4122;

wire  [0:23]  net_7009;

wire  [0:47]  net_5552;

wire  [0:23]  net_4158;

wire  [0:23]  net_6867;

wire  [0:23]  net_5383;

wire  [0:47]  net_5440;

wire  [0:47]  net_5748;

wire  [0:23]  net_4489;

wire  [0:23]  net_5551;

wire  [0:23]  net_4487;

wire  [0:47]  net_7095;

wire  [0:7]  net_7545;

wire  [0:23]  net_5161;

wire  [0:47]  net_5275;

wire  [0:23]  net_4545;

wire  [0:7]  net_5595;

wire  [0:7]  net_5903;

wire  [0:23]  net_5439;

wire  [0:15]  net_8116;

wire  [0:47]  net_7179;

wire  [0:23]  net_4739;

wire  [0:23]  net_4282;

wire  [0:47]  net_7176;

wire  [0:47]  net_7777;

wire  [0:47]  net_4171;

wire  [0:7]  net_5137;

wire  [0:7]  net_7331;

wire  [0:47]  net_4684;

wire  [0:23]  net_7149;

wire  [0:47]  net_6840;

wire  [0:23]  net_7205;

wire  [0:23]  net_6785;

wire  [0:47]  net_6056;

wire  [0:47]  net_4170;

wire  [0:23]  net_4162;

wire  [0:47]  net_6311;

wire  [0:7]  net_7219;

wire  [0:47]  net_7011;

wire  [0:47]  net_4404;

wire  [0:47]  net_5608;

wire  [0:23]  net_4769;

wire  [0:7]  net_4198;

wire  [0:23]  net_6811;

wire  [0:47]  net_6227;

wire  [0:23]  net_7343;

wire  [0:47]  net_4572;

wire  [0:47]  net_4656;

wire  [0:47]  net_5667;

wire  [0:23]  net_7093;

wire  [0:47]  net_5944;

wire  [0:23]  net_4431;

wire  [0:23]  net_4909;

wire  [0:23]  net_4683;

wire  [0:47]  net_6143;

wire  [0:23]  net_6755;

wire  [0:47]  net_7505;

wire  [0:23]  net_6645;

wire  [0:47]  net_4121;

wire  [0:47]  net_5020;

wire  [0:47]  net_4600;

wire  [0:23]  net_5467;

wire  [0:47]  net_6479;

wire  [0:47]  net_6168;

wire  [0:23]  net_6253;

wire  [0:47]  net_5664;

wire  [0:23]  net_4201;

wire  [0:47]  net_5832;

wire  [0:15]  net_7912;

wire  [0:23]  net_4285;

wire  [0:7]  net_5511;

wire  [0:47]  net_4046;

wire  [0:23]  net_5047;

wire  [0:47]  net_6843;

wire  [0:1]  net_7712;

wire  [0:23]  net_6197;

wire  [0:47]  net_5947;

wire  [0:23]  net_4767;

wire  [0:47]  net_6280;

wire  [0:23]  net_4403;

wire  [0:23]  net_7233;

wire  [0:23]  net_4090;

wire  [0:47]  net_6868;

wire  [0:47]  net_6423;

wire  [0:1]  net_8052;

wire  [0:15]  net_8058;

wire  [0:23]  net_4853;

wire  [0:47]  net_6339;

wire  [0:7]  net_6855;

wire  [0:23]  net_5693;

wire  [0:23]  net_4685;

wire  [0:47]  net_6476;

wire  [0:47]  net_6560;

wire  [0:23]  net_5943;

wire  [0:23]  net_4993;

wire  [0:47]  net_5216;

wire  [0:15]  net_7844;

wire  [0:1]  net_7746;

wire  [0:7]  net_6603;

wire  [0:23]  net_6869;

wire  [0:23]  net_6449;

wire  [0:15]  net_7548;

wire  [0:47]  net_6980;

wire  [0:47]  net_6031;

wire  [0:47]  net_5583;

wire  [0:23]  net_6083;

wire  [0:23]  net_5999;

wire  [0:47]  net_4044;

wire  [0:15]  net_7786;

wire  [0:23]  net_4655;

wire  [0:47]  net_6871;

wire  [0:7]  net_5539;

wire  [0:7]  net_6967;

wire  [0:7]  net_7135;

wire  [0:7]  net_6799;

wire  [0:7]  net_5231;

wire  [0:7]  net_7613;

wire  [0:7]  net_6099;

wire  [0:47]  net_5076;

wire  [0:23]  net_6029;

wire  [0:47]  net_6504;

wire  [0:23]  net_6195;

wire  [0:47]  net_4796;

wire  [0:47]  net_4432;

wire  [0:23]  net_5075;

wire  [0:47]  net_4544;

wire  [0:7]  net_7051;

wire  [0:47]  net_7235;

wire  [0:23]  net_6839;

wire  [0:47]  net_4407;

wire  [0:47]  net_6647;

wire  [0:23]  net_6953;

wire  [0:7]  net_4811;

wire  [0:47]  net_4824;

wire  [0:47]  net_7039;

wire  [0:47]  net_5188;

wire  [0:47]  net_4292;

wire  [0:47]  net_4547;

wire  [0:7]  net_6127;

wire  [0:23]  net_5019;

wire  [0:47]  net_5079;

wire  [0:15]  net_7980;

wire  [0:7]  net_7387;

wire  [0:47]  net_7344;

wire  [0:47]  net_5219;

wire  [0:47]  net_7123;

wire  [0:47]  net_5835;

wire  [0:47]  net_7316;

wire  [0:47]  net_6815;

wire  [0:23]  net_5021;

wire  [0:23]  net_6729;

wire  [0:47]  net_6756;

wire  [0:23]  net_7317;

wire  [0:23]  net_6951;

wire  [0:23]  net_5413;

wire  [0:23]  net_6699;

wire  [0:15]  net_7514;

wire  [0:47]  net_4880;

wire  [0:47]  net_6703;

wire  [0:47]  net_5471;

wire  [0:23]  net_4459;

wire  [0:23]  net_7261;

wire  [0:1]  net_7814;

wire  [0:47]  net_5972;

wire  [0:47]  net_5384;

wire  [0:47]  net_4911;

wire  [0:23]  net_6533;

wire  [0:23]  net_5971;

wire  [0:47]  net_5051;

wire  [0:23]  net_6757;

wire  [0:23]  net_4657;

wire  [0:47]  net_6927;

wire  [0:7]  net_8170;

wire  [0:23]  net_6561;

wire  [0:47]  net_4460;

wire  [0:23]  net_4433;

wire  [0:7]  net_7247;

wire  [0:47]  net_7036;

wire  [0:1]  net_7678;

wire  [0:23]  net_6981;

wire  [0:47]  net_4491;

wire  [0:47]  net_5104;

wire  [0:47]  net_5776;

wire  [0:47]  net_5247;

wire  [0:7]  net_6547;

wire  [0:7]  net_5119;

wire  [0:15]  net_8160;

wire  [0:23]  net_6393;

wire  [0:47]  net_7539;

wire  [0:23]  net_4517;

wire  [0:23]  net_7373;

wire  [0:23]  net_5301;

wire  [0:47]  net_4205;

wire  [0:47]  net_5695;

wire  [0:7]  net_7193;

wire  [0:23]  net_5719;

wire  [0:23]  net_5245;

wire  [0:23]  net_5187;

wire  [0:23]  net_4115;

wire  [0:47]  net_6731;

wire  [0:47]  net_4995;

wire  [0:47]  net_5863;

wire  [0:23]  net_7007;

wire  [0:47]  net_4488;

wire  [0:23]  net_7371;

wire  [0:23]  net_6615;

wire  [0:7]  net_5091;

wire  [0:23]  net_6335;

wire  [0:47]  net_5272;

wire  [0:23]  net_5243;

wire  [0:23]  net_6503;

wire  [0:23]  net_6363;

wire  [0:47]  net_4045;

wire  [0:7]  net_6827;

wire  [0:7]  net_5987;

wire  [0:23]  net_6281;

wire  [0:23]  net_5355;

wire  [0:47]  net_5723;

wire  [0:47]  net_7064;

wire  [0:47]  net_6591;

wire  [0:47]  net_4117;

wire  [0:7]  net_7681;

wire  [0:23]  net_7119;

wire  [0:47]  net_6420;

wire  [0:23]  net_4795;

wire  [0:23]  net_4825;

wire  [0:7]  net_4262;

wire  [0:23]  net_4375;

wire  [0:23]  net_5749;

wire  [0:23]  net_5777;

wire  [0:47]  net_5468;

wire  [0:7]  net_5287;

wire  [0:7]  net_4645;

wire  [0:47]  net_5555;

wire  [0:23]  net_5329;

wire  [0:47]  net_4740;

wire  [0:47]  net_7232;

wire  [0:23]  net_5831;

wire  [0:7]  net_4107;

wire  [0:23]  net_6531;

wire  [0:47]  net_7204;

wire  [0:7]  net_6519;

wire  [0:7]  net_7303;

wire  [0:23]  net_7037;

wire  [0:23]  net_5217;

wire  [0:7]  net_4305;

wire  [0:23]  net_4797;

wire  [0:47]  net_5720;

wire  [0:23]  net_5803;

wire  [0:23]  net_6167;

wire  [0:7]  net_6211;

wire  [0:47]  net_4967;

wire  [0:47]  net_6255;

wire  [0:7]  net_5455;

wire  [0:23]  net_5861;

wire  [0:47]  net_4351;

wire  [0:47]  net_4118;

wire  [0:47]  net_6896;

wire  [0:23]  net_4037;

wire  [0:23]  net_5889;

wire  [0:23]  net_5747;

wire  [0:23]  net_6057;

wire  [0:47]  net_5163;

wire  [0:23]  net_4571;

wire  [0:15]  net_7718;

wire  [0:23]  net_4377;

wire  [0:47]  net_6224;

wire  [0:23]  net_5523;

wire  [0:47]  net_6364;

wire  [0:47]  net_6000;

wire  [0:47]  net_6283;

wire  [0:23]  net_7287;

wire  [0:15]  net_7480;

wire  [0:7]  net_6883;

wire  [0:23]  net_4991;

wire  [0:47]  net_6196;

wire  [0:47]  net_6955;

wire  [0:7]  net_6155;

wire  [0:23]  net_5945;

wire  [0:23]  net_4711;

wire  [0:7]  net_7443;

wire  [0:23]  net_6477;

wire  [0:7]  net_7081;

wire  [0:47]  net_6507;

wire  [0:23]  net_5833;

wire  [0:47]  net_6588;

wire  [0:23]  net_5077;

wire  [0:23]  net_6979;

wire  [0:47]  net_7347;

wire  [0:47]  net_4435;

wire  [0:47]  net_6784;

wire  [0:47]  net_6199;

wire  [0:23]  net_7289;

wire  [0:47]  net_5107;

wire  [0:23]  net_6391;

wire  [0:7]  net_5483;

wire  [0:23]  net_4629;

wire  [0:23]  net_5357;

wire  [0:23]  net_6309;

wire  [0:7]  net_6323;

wire  [0:23]  net_4543;

wire  [0:7]  net_7783;

wire  [0:47]  net_6171;

wire  [0:23]  net_6617;

wire  [0:7]  net_4979;

wire  [0:23]  net_5385;

wire  [0:47]  net_6728;

wire  [0:47]  net_4799;

wire  [0:7]  net_5371;

wire  [0:7]  net_4923;

wire  [0:23]  net_6421;

wire  [0:23]  net_6139;

wire  [0:47]  net_5779;

wire  [0:23]  net_4879;

wire  [0:47]  net_6787;

wire  [0:23]  net_7203;

wire  [0:7]  net_7163;

wire  [0:23]  net_6475;

wire  [0:23]  net_4965;

wire  [0:23]  net_7065;

wire  [0:47]  net_6983;

wire  [0:23]  net_6337;

wire  [0:47]  net_6084;

wire  [0:47]  net_4715;

wire  [0:7]  net_4243;

wire  [0:23]  net_6589;

wire  [0:7]  net_5315;

wire  [0:47]  net_4169;

wire  [0:47]  net_6563;

wire  [0:23]  net_5273;

wire  [0:23]  net_6223;

wire  [0:23]  net_6141;

wire  [0:47]  net_5135;

wire  [0:47]  net_7675;

wire  [0:23]  net_5525;

wire  [0:23]  net_5497;

wire  [0:1]  net_7440;

wire  [0:47]  net_5636;

wire  [0:7]  net_5847;

wire  [0:7]  net_6995;

wire  [0:47]  net_4768;

wire  [0:47]  net_4047;

wire  [0:47]  net_7120;

wire  [0:23]  net_6251;

wire  [0:23]  net_7177;

wire  [0:23]  net_4319;

wire  [0:23]  net_4286;

wire  [0:7]  net_7477;

wire  [0:47]  net_8049;

wire  [0:15]  net_7446;

wire  [0:7]  net_6297;

wire  [0:23]  net_4349;

wire  [0:1]  net_7780;

wire  [0:47]  net_7288;

wire  [0:47]  net_5891;

wire  [0:47]  net_6899;

wire  [0:47]  net_5527;

wire  [0:47]  net_5356;

wire  [0:47]  net_6700;

wire  [0:47]  net_7148;

wire  [0:47]  net_6112;

wire  [0:47]  net_7372;

wire  [0:23]  net_5805;

wire  [0:15]  net_7684;

wire  [0:23]  net_6111;

wire  [0:47]  net_7207;

wire  [0:47]  net_4939;

wire  [0:7]  net_7749;

wire  [0:7]  net_4181;

wire  [0:23]  net_4347;

wire  [0:7]  net_7191;

wire  [0:23]  net_5299;

wire  [0:7]  net_6409;

wire  [0:23]  net_6895;

wire  [0:7]  net_5147;

wire  [0:7]  net_6379;

wire  [0:47]  net_6759;

wire  [0:23]  net_4907;

wire  [0:47]  net_5975;

wire  [0:7]  net_6911;

wire  [0:47]  net_4206;

wire  [0:15]  net_7640;

wire  [0:23]  net_6365;

wire  [0:15]  net_7616;

wire  [0:47]  net_4964;

wire  [0:47]  net_7151;

wire  [0:47]  net_5328;

wire  [0:47]  net_7008;

wire  [0:7]  net_4895;

wire  [0:47]  net_7437;

wire  [0:47]  net_6448;

wire  [0:47]  net_5554;

wire  [0:47]  net_4168;

wire  [0:47]  net_5888;

wire  [0:47]  net_4516;

wire  [0:47]  net_4203;

wire  [0:23]  net_5189;

wire  [0:23]  net_7121;

wire  [0:1]  net_7474;

wire  [0:23]  net_7175;

wire  [0:47]  net_6028;

wire  [0:47]  net_4628;

wire  [0:23]  net_5495;

wire  [0:23]  net_6813;

wire  [0:23]  net_7035;

wire  [0:47]  net_5804;

wire  [0:23]  net_5721;

wire  [0:23]  net_4963;

wire  [0:23]  net_6923;

wire  [0:23]  net_5973;

wire  [0:47]  net_4855;

wire  [0:47]  net_7607;

wire  [0:47]  net_6812;

wire  [0:47]  net_5860;

wire  [0:23]  net_4599;

wire  [0:23]  net_5579;

wire  [0:23]  net_6673;

wire  [0:23]  net_5049;

wire  [0:23]  net_7063;

wire  [0:7]  net_7023;

wire  [0:47]  net_5919;

wire  [0:1]  net_8154;

wire  [0:23]  net_6783;

wire  [0:47]  net_7743;

wire  [0:23]  net_5581;

wire  [0:23]  net_5103;

wire  [0:47]  net_7260;

wire  [0:23]  net_6447;

wire  [0:47]  net_7709;

wire  [0:23]  net_6085;

wire  [0:47]  net_5496;

wire  [0:47]  net_5191;

wire  [0:23]  net_6587;

wire  [0:7]  net_5623;

wire  [0:23]  net_5607;

wire  [0:23]  net_4321;

wire  [0:47]  net_6059;

wire  [0:47]  net_6451;

wire  [0:23]  net_5691;

wire  [0:7]  net_5399;

wire  [0:47]  net_6308;

wire  [0:23]  net_5105;

wire  [0:47]  net_5132;

wire  [0:47]  net_5412;

wire  [0:47]  net_5692;

wire  [0:47]  net_4376;

wire  [0:7]  net_5063;

wire  [0:47]  net_5499;

wire  [0:7]  net_6939;

wire  [0:7]  net_4207;

wire  [0:23]  net_5411;

wire  [0:23]  net_6701;



bram_bufferx4x6 I904 ( .in(sdi), .out(net_03985));
bram_bufferx4x6 I905 ( .in(net_7931), .out(net_03983));
lowla_modified I896 ( .clk(tclk_i), .min(net_03985), .lao(net_3948));
lowla_modified I1083 ( .clk(net_03953), .min(net_03983),
     .lao(net_3950));
io_col4_rowright I_25_11_ior21 ( .ceb(net_04306), .cf(cf_r[263:240]),
     .vdd_cntl(vdd_cntl[191:176]), .hold(hold_r_t),
     .fabric_out(net_7556), .sdo(net_7557), .sdi(net_3948),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[0]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[21:20]),
     .pado(pado_r[21:20]), .padeb(padeb_r[21:20]),
     .sp4_v_t(net_7572[0:15]), .sp4_h_l(net_6728[0:47]),
     .sp12_h_l(net_6727[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[21:20]), .tnl_op(net_7247[0:7]),
     .lft_op(slf_op_24_11[7:0]), .bnl_op(bnl_op_25_11[7:0]),
     .pgate(pgate[191:176]), .reset(reset_b[191:176]),
     .sp4_v_b(sp4_v_b_25_11[15:0]), .wl(wl[191:176]),
     .bl(bl[1311:1294]), .slf_op(io_r_00_24_11[3:0]),
     .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_12_ior23 ( .ceb(net_04306), .cf(cf_r[287:264]),
     .vdd_cntl(vdd_cntl[207:192]), .hold(hold_r_t),
     .fabric_out(net_7624), .sdo(net_8068), .sdi(net_7557),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[1]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[23:22]),
     .pado(pado_r[23:22]), .padeb(padeb_r[23:22]),
     .sp4_v_t(net_7640[0:15]), .sp4_h_l(net_6644[0:47]),
     .sp12_h_l(net_6643[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[23:22]), .tnl_op(net_7387[0:7]),
     .lft_op(net_7247[0:7]), .bnl_op(slf_op_24_11[7:0]),
     .pgate(pgate[207:192]), .reset(reset_b[207:192]),
     .sp4_v_b(net_7572[0:15]), .wl(wl[207:192]), .bl(bl[1311:1294]),
     .slf_op(io_r_01[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_15_ior29 ( .ceb(net_04306), .cf(cf_r[359:336]),
     .vdd_cntl(vdd_cntl[255:240]), .hold(hold_r_t),
     .fabric_out(net_7828), .sdo(net_7829), .sdi(net_8101),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[4]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[29:28]),
     .pado(pado_r[29:28]), .padeb(padeb_r[29:28]),
     .sp4_v_t(net_7844[0:15]), .sp4_h_l(net_5328[0:47]),
     .sp12_h_l(net_5327[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[29:28]), .tnl_op(net_6463[0:7]),
     .lft_op(net_5371[0:7]), .bnl_op(net_5231[0:7]),
     .pgate(pgate[255:240]), .reset(reset_b[255:240]),
     .sp4_v_b(net_8116[0:15]), .wl(wl[255:240]), .bl(bl[1311:1294]),
     .slf_op(io_r_04[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_16_ior31 ( .ceb(net_04306), .cf(cf_r[383:360]),
     .vdd_cntl(vdd_cntl[271:256]), .hold(hold_r_t),
     .fabric_out(net_7862), .sdo(net_7863), .sdi(net_7829),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[5]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[31:30]),
     .pado(pado_r[31:30]), .padeb(padeb_r[31:30]),
     .sp4_v_t(net_7878[0:15]), .sp4_h_l(net_5244[0:47]),
     .sp12_h_l(net_5243[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[31:30]), .tnl_op(net_6603[0:7]),
     .lft_op(net_6463[0:7]), .bnl_op(net_5371[0:7]),
     .pgate(pgate[271:256]), .reset(reset_b[271:256]),
     .sp4_v_b(net_7844[0:15]), .wl(wl[271:256]), .bl(bl[1311:1294]),
     .slf_op(io_r_05[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_19_ior37 ( .ceb(net_04306), .cf(cf_r[455:432]),
     .vdd_cntl(vdd_cntl[319:304]), .hold(hold_r_t),
     .fabric_out(net_7896), .sdo(net_7897), .sdi(net_7999),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[8]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[37:36]),
     .pado(pado_r[37:36]), .padeb(padeb_r[37:36]),
     .sp4_v_t(net_7912[0:15]), .sp4_h_l(net_5944[0:47]),
     .sp12_h_l(net_5943[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[37:36]), .tnl_op(net_7783[0:7]),
     .lft_op(net_5987[0:7]), .bnl_op(net_5847[0:7]),
     .pgate(pgate[319:304]), .reset(reset_b[319:304]),
     .sp4_v_b(net_8014[0:15]), .wl(wl[319:304]), .bl(bl[1311:1294]),
     .slf_op(io_r_08[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_20_ior39 ( .ceb(net_04306), .cf(cf_r[479:456]),
     .vdd_cntl(vdd_cntl[335:320]), .hold(hold_r_t),
     .fabric_out(net_7930), .sdo(net_7931), .sdi(net_7897),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[9]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[39:38]),
     .pado(pado_r[39:38]), .padeb(padeb_r[39:38]),
     .sp4_v_t(net_7820[0:15]), .sp4_h_l(net_5860[0:47]),
     .sp12_h_l(net_5859[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[39:38]), .tnl_op({io_t_24[3], io_t_24[2],
     io_t_24[1], io_t_24[0], io_t_24[3], io_t_24[2], io_t_24[1],
     io_t_24[0]}), .lft_op(net_7783[0:7]), .bnl_op(net_5987[0:7]),
     .pgate(pgate[335:320]), .reset(reset_b[335:320]),
     .sp4_v_b(net_7912[0:15]), .wl(wl[335:320]), .bl(bl[1311:1294]),
     .slf_op(slf_op_25_10[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_17_ior33 ( .ceb(net_04306), .cf(cf_r[407:384]),
     .vdd_cntl(vdd_cntl[287:272]), .hold(hold_r_t),
     .fabric_out(net_7964), .sdo(net_7965), .sdi(net_7863),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[6]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[33:32]),
     .pado(pado_r[33:32]), .padeb(padeb_r[33:32]),
     .sp4_v_t(net_7980[0:15]), .sp4_h_l(net_6560[0:47]),
     .sp12_h_l(net_6559[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[33:32]), .tnl_op(net_5847[0:7]),
     .lft_op(net_6603[0:7]), .bnl_op(net_6463[0:7]),
     .pgate(pgate[287:272]), .reset(reset_b[287:272]),
     .sp4_v_b(net_7878[0:15]), .wl(wl[287:272]), .bl(bl[1311:1294]),
     .slf_op(io_r_06[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_18_ior35 ( .ceb(net_04306), .cf(cf_r[431:408]),
     .vdd_cntl(vdd_cntl[303:288]), .hold(hold_r_t),
     .fabric_out(net_7998), .sdo(net_7999), .sdi(net_7965),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[7]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[35:34]),
     .pado(pado_r[35:34]), .padeb(padeb_r[35:34]),
     .sp4_v_t(net_8014[0:15]), .sp4_h_l(net_6476[0:47]),
     .sp12_h_l(net_6475[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[35:34]), .tnl_op(net_5987[0:7]),
     .lft_op(net_5847[0:7]), .bnl_op(net_6603[0:7]),
     .pgate(pgate[303:288]), .reset(reset_b[303:288]),
     .sp4_v_b(net_7980[0:15]), .wl(wl[303:288]), .bl(bl[1311:1294]),
     .slf_op(io_r_07[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_13_ior25 ( .ceb(net_04306), .cf(cf_r[311:288]),
     .vdd_cntl(vdd_cntl[223:208]), .hold(hold_r_t),
     .fabric_out(net_8066), .sdo(net_8067), .sdi(net_8068),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[2]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[25:24]),
     .pado(pado_r[25:24]), .padeb(padeb_r[25:24]),
     .sp4_v_t(net_8082[0:15]), .sp4_h_l(net_7344[0:47]),
     .sp12_h_l(net_7343[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[25:24]), .tnl_op(net_5231[0:7]),
     .lft_op(net_7387[0:7]), .bnl_op(net_7247[0:7]),
     .pgate(pgate[223:208]), .reset(reset_b[223:208]),
     .sp4_v_b(net_7640[0:15]), .wl(wl[223:208]), .bl(bl[1311:1294]),
     .slf_op(io_r_02[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
io_col4_rowright I_25_14_ior27 ( .ceb(net_04306), .cf(cf_r[335:312]),
     .vdd_cntl(vdd_cntl[239:224]), .hold(hold_r_t),
     .fabric_out(net_8100), .sdo(net_8101), .sdi(net_8067),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_r[3]),
     .spioeb({tievdd, tievdd}), .mode(net_3953), .shift(net_3973),
     .hiz_b(net_7564), .r(net_7565), .bs_en(net_7566),
     .tclk(net_03953), .update(net_3955), .padin(padin_r[27:26]),
     .pado(pado_r[27:26]), .padeb(padeb_r[27:26]),
     .sp4_v_t(net_8116[0:15]), .sp4_h_l(net_7260[0:47]),
     .sp12_h_l(net_7259[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_r[27:26]), .tnl_op(net_5371[0:7]),
     .lft_op(net_5231[0:7]), .bnl_op(net_7387[0:7]),
     .pgate(pgate[239:224]), .reset(reset_b[239:224]),
     .sp4_v_b(net_8082[0:15]), .wl(wl[239:224]), .bl(bl[1311:1294]),
     .slf_op(io_r_03[3:0]), .glb_netwk(glb_netwk_io_r[7:0]));
bram_bufferx4 I903 ( .in(net_04306), .out(ceb_o));
bram_bufferx4 I889 ( .in(mode_i), .out(net_3953));
bram_bufferx4 I902 ( .in(ceb_i), .out(net_04306));
bram_bufferx4 I1076 ( .in(net_3953), .out(mode_o));
bram_bufferx4 I1082 ( .in(net_3955), .out(update_o));
bram_bufferx4 I895 ( .in(hiz_b_i), .out(net_7564));
bram_bufferx4 I894 ( .in(r_i), .out(net_7565));
bram_bufferx4 I893 ( .in(shift_i), .out(net_3973));
bram_bufferx4 I890 ( .in(update_i), .out(net_3955));
bram_bufferx4 I892 ( .in(bs_en_i), .out(net_7566));
bram_bufferx4 I891 ( .in(tclk_i), .out(net_03953));
bram_bufferx4 I1077 ( .in(net_03953), .out(tclk_o));
bram_bufferx4 I1079 ( .in(net_7566), .out(bs_en_o));
bram_bufferx4 I1078 ( .in(net_3973), .out(shift_o));
bram_bufferx4 I1080 ( .in(net_7565), .out(r_o));
bram_bufferx4 I1081 ( .in(net_7564), .out(hiz_b_o));
inv_hvt I1017 ( .A(net_3979), .Y(padin_223));
inv_hvt I1018 ( .A(padin_t[24]), .Y(net_3979));
inv_hvt I855 ( .A(padin_r[20]), .Y(net_3984));
inv_hvt I856 ( .A(net_3984), .Y(padin_163));
inv_hvt I859 ( .A(net_7624), .Y(net_3988));
inv_hvt I860 ( .A(net_3988), .Y(fabric_out_168));
inv_hvt I857 ( .A(net_3991), .Y(fabric_out_223));
inv_hvt I862 ( .A(net_3996), .Y(fabric_out_163));
inv_hvt I861 ( .A(net_7556), .Y(net_3996));
inv_hvt I858 ( .A(net_3997), .Y(net_3991));
bram_4kprouting_tbankin I_bram1919 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_bot(vdd_cntl[319:304]),
     .vdd_cntl_top(vdd_cntl[335:320]), .bm_sdo_o(net_4067),
     .bm_sdi_i(net_4069), .bm_sclkrw_i(net_4070), .bm_sdo_i(bm_sdo_i),
     .bm_sweb_i(net_4071), .bm_sdi_o(bm_sdi_o),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_sweb_o(bm_sweb_o),
     .slf_op_top(net_8157[0:7]), .slf_op_bot(net_6297[0:7]),
     .wl_top(wl[335:320]), .wl_bot(wl[319:304]),
     .top_op_top({io_t_19[3], io_t_19[2], io_t_19[1], io_t_19[0],
     io_t_19[3], io_t_19[2], io_t_19[1], io_t_19[0]}),
     .tnr_op_top({io_t_20[3], io_t_20[2], io_t_20[1], io_t_20[0],
     io_t_20[3], io_t_20[2], io_t_20[1], io_t_20[0]}),
     .tnr_op_bot(net_7613[0:7]), .tnl_op_top({io_t_18[3], io_t_18[2],
     io_t_18[1], io_t_18[0], io_t_18[3], io_t_18[2], io_t_18[1],
     io_t_18[0]}), .tnl_op_bot(net_7545[0:7]),
     .rgt_op_top(net_7613[0:7]), .rgt_op_bot(net_4113[0:7]),
     .reset_b_top(reset_b[335:320]), .reset_b_bot(reset_b[319:304]),
     .prog(prog), .pgate_top(pgate[335:320]),
     .pgate_bot(pgate[319:304]), .lft_op_top(net_7545[0:7]),
     .lft_op_bot(net_5427[0:7]), .bm_wdummymux_en_i(net_4110),
     .bot_op_bot(net_5707[0:7]), .bnr_op_top(net_4113[0:7]),
     .bnr_op_bot(net_4031[0:7]), .bnl_op_top(net_5427[0:7]),
     .bnl_op_bot(net_5399[0:7]), .sp12_v_t_top(net_4034[0:23]),
     .sp12_v_b_bot(net_4090[0:23]), .bm_init_i(net_4106),
     .sp12_h_r_top(net_4037[0:23]), .sp12_h_r_bot(net_4038[0:23]),
     .sp12_h_l_top(net_5551[0:23]), .sp12_h_l_bot(net_5691[0:23]),
     .sp4_v_t_top(net_7607[0:47]), .sp4_v_b_top(net_5555[0:47]),
     .sp4_v_b_bot(net_5695[0:47]), .sp4_r_v_b_top(net_4044[0:47]),
     .sp4_r_v_b_bot(net_4045[0:47]), .sp4_h_r_top(net_4046[0:47]),
     .sp4_h_r_bot(net_4047[0:47]), .sp4_h_l_top(net_5552[0:47]),
     .sp4_h_l_bot(net_5692[0:47]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(net_4105), .bm_sa_i(net_4107[0:7]),
     .bm_sclk_i(net_4108), .bm_sreb_i(net_4109),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4kprouting_tbank I_bram1917 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_bot(vdd_cntl[287:272]),
     .vdd_cntl_top(vdd_cntl[303:288]), .bm_sdo_o(net_4129),
     .bm_sdi_i(net_4131), .bm_sclkrw_i(net_4132), .bm_sdo_i(net_4067),
     .bm_sweb_i(net_4133), .bm_sdi_o(net_4069), .bm_sclkrw_o(net_4070),
     .bm_sweb_o(net_4071), .slf_op_top(net_5707[0:7]),
     .slf_op_bot(net_4138[0:7]), .wl_top(wl[303:288]),
     .wl_bot(wl[287:272]), .top_op_top(net_6297[0:7]),
     .tnl_op_top(net_5427[0:7]), .tnl_op_bot(net_5399[0:7]),
     .reset_b_top(reset_b[303:288]), .reset_b_bot(reset_b[287:272]),
     .prog(prog), .pgate_top(pgate[303:288]),
     .pgate_bot(pgate[287:272]), .lft_op_top(net_5399[0:7]),
     .lft_op_bot(net_6155[0:7]), .bm_wdummymux_en_i(net_4184),
     .bot_op_bot(net_6323[0:7]), .bnl_op_top(net_6155[0:7]),
     .bnl_op_bot(net_6127[0:7]), .sp12_v_t_top(net_4090[0:23]),
     .sp12_v_b_bot(net_4158[0:23]), .bm_init_i(net_4180),
     .sp12_h_l_top(net_6279[0:23]), .sp12_h_l_bot(net_6307[0:23]),
     .sp4_v_t_top(net_5695[0:47]), .sp4_v_b_top(net_6283[0:47]),
     .sp4_v_b_bot(net_6311[0:47]), .sp4_h_l_top(net_6280[0:47]),
     .sp4_h_l_bot(net_6308[0:47]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(net_4179), .bm_sa_i(net_4181[0:7]),
     .bm_sclk_i(net_4182), .bm_sreb_i(net_4183),
     .bm_rcapmux_en_o(net_4105), .bm_init_o(net_4106),
     .bm_sa_o(net_4107[0:7]), .bm_sclk_o(net_4108),
     .bm_sreb_o(net_4109), .bm_wdummymux_en_o(net_4110),
     .bnr_op_top(net_5137[0:7]), .rgt_op_top(net_4031[0:7]),
     .tnr_op_top(net_4113[0:7]), .tnr_op_bot(net_4031[0:7]),
     .sp12_h_r_top(net_4115[0:23]), .sp12_h_r_bot(net_4116[0:23]),
     .sp4_h_r_bot(net_4117[0:47]), .sp4_h_r_top(net_4118[0:47]),
     .rgt_op_bot(net_5137[0:7]), .sp4_r_v_b_top(net_4120[0:47]),
     .sp4_r_v_b_bot(net_4121[0:47]), .bnr_op_bot(net_4122[0:7]));
bram_4kprouting_tbank I_bram1915 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_bot(vdd_cntl[255:240]),
     .vdd_cntl_top(vdd_cntl[271:256]), .bm_sdo_o(net_4191),
     .bm_sdi_i(net_4193), .bm_sclkrw_i(net_4194), .bm_sdo_i(net_4129),
     .bm_sweb_i(net_4195), .bm_sdi_o(net_4131), .bm_sclkrw_o(net_4132),
     .bm_sweb_o(net_4133), .slf_op_top(net_6323[0:7]),
     .slf_op_bot(net_7081[0:7]), .wl_top(wl[271:256]),
     .wl_bot(wl[255:240]), .top_op_top(net_4138[0:7]),
     .tnr_op_top(net_5137[0:7]), .tnr_op_bot(net_4122[0:7]),
     .tnl_op_top(net_6155[0:7]), .tnl_op_bot(net_6127[0:7]),
     .rgt_op_top(net_4122[0:7]), .rgt_op_bot(net_4198[0:7]),
     .reset_b_top(reset_b[271:256]), .reset_b_bot(reset_b[255:240]),
     .prog(prog), .pgate_top(pgate[271:256]),
     .pgate_bot(pgate[255:240]), .lft_op_top(net_6127[0:7]),
     .lft_op_bot(net_4811[0:7]), .bm_wdummymux_en_i(net_4246),
     .bot_op_bot(net_5091[0:7]), .bnr_op_top(net_4198[0:7]),
     .bnr_op_bot(net_4155[0:7]), .bnl_op_top(net_4811[0:7]),
     .bnl_op_bot(net_4783[0:7]), .sp12_v_t_top(net_4158[0:23]),
     .sp12_v_b_bot(net_4226[0:23]), .bm_init_i(net_4242),
     .sp12_h_r_top(net_4161[0:23]), .sp12_h_r_bot(net_4162[0:23]),
     .sp12_h_l_top(net_4935[0:23]), .sp12_h_l_bot(net_5075[0:23]),
     .sp4_v_t_top(net_6311[0:47]), .sp4_v_b_top(net_4939[0:47]),
     .sp4_v_b_bot(net_5079[0:47]), .sp4_r_v_b_top(net_4168[0:47]),
     .sp4_r_v_b_bot(net_4169[0:47]), .sp4_h_r_top(net_4170[0:47]),
     .sp4_h_r_bot(net_4171[0:47]), .sp4_h_l_top(net_4936[0:47]),
     .sp4_h_l_bot(net_5076[0:47]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(net_4241), .bm_sa_i(net_4243[0:7]),
     .bm_sclk_i(net_4244), .bm_sreb_i(net_4245),
     .bm_rcapmux_en_o(net_4179), .bm_init_o(net_4180),
     .bm_sa_o(net_4181[0:7]), .bm_sclk_o(net_4182),
     .bm_sreb_o(net_4183), .bm_wdummymux_en_o(net_4184));
bram_4kprouting_tbank I_bram1913 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_bot(vdd_cntl[223:208]),
     .vdd_cntl_top(vdd_cntl[239:224]), .bm_sdo_o(net_4253),
     .bm_sdi_i(net_4255), .bm_sclkrw_i(net_4256), .bm_sdo_i(net_4191),
     .bm_sweb_i(net_4257), .bm_sdi_o(net_4193), .bm_sclkrw_o(net_4194),
     .bm_sweb_o(net_4195), .bnr_op_top(net_4689[0:7]),
     .rgt_op_top(net_4155[0:7]), .tnr_op_top(net_4198[0:7]),
     .tnr_op_bot(net_4155[0:7]), .sp12_h_r_top(net_4200[0:23]),
     .sp12_h_r_bot(net_4201[0:23]), .sp4_h_r_bot(net_4202[0:47]),
     .sp4_h_r_top(net_4203[0:47]), .rgt_op_bot(net_4689[0:7]),
     .sp4_r_v_b_top(net_4205[0:47]), .sp4_r_v_b_bot(net_4206[0:47]),
     .bnr_op_bot(net_4207[0:7]), .slf_op_top(net_5091[0:7]),
     .slf_op_bot(net_4262[0:7]), .wl_top(wl[239:224]),
     .wl_bot(wl[223:208]), .top_op_top(net_7081[0:7]),
     .tnl_op_top(net_4811[0:7]), .tnl_op_bot(net_4783[0:7]),
     .reset_b_top(reset_b[239:224]), .reset_b_bot(reset_b[223:208]),
     .prog(prog), .pgate_top(pgate[239:224]),
     .pgate_bot(pgate[223:208]), .lft_op_top(net_4783[0:7]),
     .lft_op_bot(net_6939[0:7]), .bm_wdummymux_en_i(net_4308),
     .bot_op_bot(net_4645[0:7]), .bnl_op_top(net_6939[0:7]),
     .bnl_op_bot(net_6911[0:7]), .sp12_v_t_top(net_4226[0:23]),
     .sp12_v_b_bot(net_4282[0:23]), .bm_init_i(net_4304),
     .sp12_h_l_top(net_7063[0:23]), .sp12_h_l_bot(net_7091[0:23]),
     .sp4_v_t_top(net_5079[0:47]), .sp4_v_b_top(net_7067[0:47]),
     .sp4_v_b_bot(net_7095[0:47]), .sp4_h_l_top(net_7064[0:47]),
     .sp4_h_l_bot(net_7092[0:47]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(net_4303), .bm_sa_i(net_4305[0:7]),
     .bm_sclk_i(net_4306), .bm_sreb_i(net_4307),
     .bm_rcapmux_en_o(net_4241), .bm_init_o(net_4242),
     .bm_sa_o(net_4243[0:7]), .bm_sclk_o(net_4244),
     .bm_sreb_o(net_4245), .bm_wdummymux_en_o(net_4246));
bram_4kprouting_tbankout I_bram1911 ( .glb_netwk(glb_netwk_19[7:0]),
     .vdd_cntl_bot(vdd_cntl[191:176]),
     .vdd_cntl_top(vdd_cntl[207:192]), .bm_sdo_o(bm_sdo_o),
     .bm_sdi_i(bm_sdi_i), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sdo_i(net_4253), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(net_4255),
     .bm_sclkrw_o(net_4256), .bm_sweb_o(net_4257),
     .slf_op_top(net_4645[0:7]), .slf_op_bot(slf_op_19_11[7:0]),
     .wl_top(wl[207:192]), .wl_bot(wl[191:176]),
     .top_op_top(net_4262[0:7]), .tnr_op_top(net_4689[0:7]),
     .tnr_op_bot(net_4207[0:7]), .tnl_op_top(net_6939[0:7]),
     .tnl_op_bot(net_6911[0:7]), .rgt_op_top(net_4207[0:7]),
     .rgt_op_bot(slf_op_20_11[7:0]), .reset_b_top(reset_b[207:192]),
     .reset_b_bot(reset_b[191:176]), .prog(prog),
     .pgate_top(pgate[207:192]), .pgate_bot(pgate[191:176]),
     .lft_op_top(net_6911[0:7]), .lft_op_bot(slf_op_18_11[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_19_11[7:0]), .bnr_op_top(slf_op_20_11[7:0]),
     .bnr_op_bot(bnr_op_19_11[7:0]), .bnl_op_top(slf_op_18_11[7:0]),
     .bnl_op_bot(bnl_op_19_11[7:0]), .sp12_v_t_top(net_4282[0:23]),
     .sp12_v_b_bot(sp12_v_b_19_11[23:0]), .bm_init_i(bm_init_i),
     .sp12_h_r_top(net_4285[0:23]), .sp12_h_r_bot(net_4286[0:23]),
     .sp12_h_l_top(net_4487[0:23]), .sp12_h_l_bot(net_4627[0:23]),
     .sp4_v_t_top(net_7095[0:47]), .sp4_v_b_top(net_4491[0:47]),
     .sp4_v_b_bot(sp4_v_b_19_11[47:0]), .sp4_r_v_b_top(net_4292[0:47]),
     .sp4_r_v_b_bot(sp4_v_b_20_11[47:0]), .sp4_h_r_top(net_4294[0:47]),
     .sp4_h_r_bot(net_4295[0:47]), .sp4_h_l_top(net_4488[0:47]),
     .sp4_h_l_bot(net_4628[0:47]), .bl(bl[1023:982]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(net_4303), .bm_init_o(net_4304),
     .bm_sa_o(net_4305[0:7]), .bm_sclk_o(net_4306),
     .bm_sreb_o(net_4307), .bm_wdummymux_en_o(net_4308));
clk_quad_bufx8 I_quad_driver ( .clko(net2col_drivers[7:0]),
     .clki(glb_in[7:0]));
ltile4rev I_17_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4313), .lft_op(slf_op_16_11[7:0]),
     .sp12_h_l(net_4459[0:23]), .sp4_h_l(net_4460[0:47]),
     .sp4_v_b(sp4_v_b_17_11[47:0]), .sp12_v_b(sp12_v_b_17_11[23:0]),
     .sp12_h_r(net_4319[0:23]), .sp4_h_r(net_4320[0:47]),
     .sp12_v_t(net_4321[0:23]), .sp4_v_t(net_4435[0:47]),
     .sp4_r_v_b(sp4_v_b_18_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7051[0:7]), .rgt_op(slf_op_18_11[7:0]),
     .bot_op(bot_op_17_11[7:0]), .bl(bl[927:874]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(carry_in_17_11), .purst(purst),
     .slf_op(slf_op_17_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_17_11[7:0]), .bnl_op(bnl_op_17_11[7:0]),
     .tnr_op(net_6911[0:7]), .tnl_op(net_6967[0:7]));
ltile4rev I_17_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4341), .lft_op(net_6967[0:7]),
     .sp12_h_l(net_4431[0:23]), .sp4_h_l(net_4432[0:47]),
     .sp4_v_b(net_4435[0:47]), .sp12_v_b(net_4321[0:23]),
     .sp12_h_r(net_4347[0:23]), .sp4_h_r(net_4348[0:47]),
     .sp12_v_t(net_4349[0:23]), .sp4_v_t(net_7039[0:47]),
     .sp4_r_v_b(net_4351[0:47]), .wl(wl[207:192]),
     .top_op(net_7023[0:7]), .rgt_op(net_6911[0:7]),
     .bot_op(slf_op_17_11[7:0]), .bl(bl[927:874]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_4313), .purst(purst), .slf_op(net_7051[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_18_11[7:0]),
     .bnl_op(slf_op_16_11[7:0]), .tnr_op(net_6939[0:7]),
     .tnl_op(net_6995[0:7]));
ltile4rev I_15_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4369), .lft_op(slf_op_14_11[7:0]),
     .sp12_h_l(net_4515[0:23]), .sp4_h_l(net_4516[0:47]),
     .sp4_v_b(sp4_v_b_15_11[47:0]), .sp12_v_b(sp12_v_b_15_11[23:0]),
     .sp12_h_r(net_4375[0:23]), .sp4_h_r(net_4376[0:47]),
     .sp12_v_t(net_4377[0:23]), .sp4_v_t(net_4547[0:47]),
     .sp4_r_v_b(sp4_v_b_16_11[47:0]), .wl(wl[191:176]),
     .top_op(net_6883[0:7]), .rgt_op(slf_op_16_11[7:0]),
     .bot_op(bot_op_15_11[7:0]), .bl(bl[819:766]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(carry_in_15_11), .purst(purst),
     .slf_op(slf_op_15_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_15_11[7:0]), .bnl_op(bnl_op_15_11[7:0]),
     .tnr_op(net_6967[0:7]), .tnl_op(net_6799[0:7]));
ltile4rev I_15_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4397), .lft_op(net_6799[0:7]),
     .sp12_h_l(net_4543[0:23]), .sp4_h_l(net_4544[0:47]),
     .sp4_v_b(net_4547[0:47]), .sp12_v_b(net_4377[0:23]),
     .sp12_h_r(net_4403[0:23]), .sp4_h_r(net_4404[0:47]),
     .sp12_v_t(net_4405[0:23]), .sp4_v_t(net_6871[0:47]),
     .sp4_r_v_b(net_4407[0:47]), .wl(wl[207:192]),
     .top_op(net_6855[0:7]), .rgt_op(net_6967[0:7]),
     .bot_op(slf_op_15_11[7:0]), .bl(bl[819:766]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_4369), .purst(purst), .slf_op(net_6883[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_16_11[7:0]),
     .bnl_op(slf_op_14_11[7:0]), .tnr_op(net_6995[0:7]),
     .tnl_op(net_6827[0:7]));
ltile4rev I_16_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4425), .lft_op(net_6883[0:7]),
     .sp12_h_l(net_4403[0:23]), .sp4_h_l(net_4404[0:47]),
     .sp4_v_b(net_4407[0:47]), .sp12_v_b(net_4461[0:23]),
     .sp12_h_r(net_4431[0:23]), .sp4_h_r(net_4432[0:47]),
     .sp12_v_t(net_4433[0:23]), .sp4_v_t(net_6955[0:47]),
     .sp4_r_v_b(net_4435[0:47]), .wl(wl[207:192]),
     .top_op(net_6995[0:7]), .rgt_op(net_7051[0:7]),
     .bot_op(slf_op_16_11[7:0]), .bl(bl[873:820]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_4453), .purst(purst), .slf_op(net_6967[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_17_11[7:0]),
     .bnl_op(slf_op_15_11[7:0]), .tnr_op(net_7023[0:7]),
     .tnl_op(net_6855[0:7]));
ltile4rev I_16_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4453), .lft_op(slf_op_15_11[7:0]),
     .sp12_h_l(net_4375[0:23]), .sp4_h_l(net_4376[0:47]),
     .sp4_v_b(sp4_v_b_16_11[47:0]), .sp12_v_b(sp12_v_b_16_11[23:0]),
     .sp12_h_r(net_4459[0:23]), .sp4_h_r(net_4460[0:47]),
     .sp12_v_t(net_4461[0:23]), .sp4_v_t(net_4407[0:47]),
     .sp4_r_v_b(sp4_v_b_17_11[47:0]), .wl(wl[191:176]),
     .top_op(net_6967[0:7]), .rgt_op(slf_op_17_11[7:0]),
     .bot_op(bot_op_16_11[7:0]), .bl(bl[873:820]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(carry_in_16_11), .purst(purst),
     .slf_op(slf_op_16_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_16_11[7:0]), .bnl_op(bnl_op_16_11[7:0]),
     .tnr_op(net_7051[0:7]), .tnl_op(net_6883[0:7]));
ltile4rev I_18_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4481), .lft_op(net_7051[0:7]),
     .sp12_h_l(net_4347[0:23]), .sp4_h_l(net_4348[0:47]),
     .sp4_v_b(net_4351[0:47]), .sp12_v_b(net_4629[0:23]),
     .sp12_h_r(net_4487[0:23]), .sp4_h_r(net_4488[0:47]),
     .sp12_v_t(net_4489[0:23]), .sp4_v_t(net_6899[0:47]),
     .sp4_r_v_b(net_4491[0:47]), .wl(wl[207:192]),
     .top_op(net_6939[0:7]), .rgt_op(net_4645[0:7]),
     .bot_op(slf_op_18_11[7:0]), .bl(bl[981:928]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_4621), .purst(purst), .slf_op(net_6911[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_19_11[7:0]),
     .bnl_op(slf_op_17_11[7:0]), .tnr_op(net_4262[0:7]),
     .tnl_op(net_7023[0:7]));
ltile4rev I_14_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4509), .lft_op(slf_op_13_11[7:0]),
     .sp12_h_l(net_4599[0:23]), .sp4_h_l(net_4600[0:47]),
     .sp4_v_b(sp4_v_b_14_11[47:0]), .sp12_v_b(sp12_v_b_14_11[23:0]),
     .sp12_h_r(net_4515[0:23]), .sp4_h_r(net_4516[0:47]),
     .sp12_v_t(net_4517[0:23]), .sp4_v_t(net_4575[0:47]),
     .sp4_r_v_b(sp4_v_b_15_11[47:0]), .wl(wl[191:176]),
     .top_op(net_6799[0:7]), .rgt_op(slf_op_15_11[7:0]),
     .bot_op(bot_op_14_11[7:0]), .bl(bl[765:712]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(carry_in_14_11), .purst(purst),
     .slf_op(slf_op_14_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_14_11[7:0]), .bnl_op(bnl_op_14_11[7:0]),
     .tnr_op(net_6883[0:7]), .tnl_op(slf_op_13_02[7:0]));
ltile4rev I_14_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4537), .lft_op(slf_op_13_02[7:0]),
     .sp12_h_l(net_4571[0:23]), .sp4_h_l(net_4572[0:47]),
     .sp4_v_b(net_4575[0:47]), .sp12_v_b(net_4517[0:23]),
     .sp12_h_r(net_4543[0:23]), .sp4_h_r(net_4544[0:47]),
     .sp12_v_t(net_4545[0:23]), .sp4_v_t(net_6787[0:47]),
     .sp4_r_v_b(net_4547[0:47]), .wl(wl[207:192]),
     .top_op(net_6827[0:7]), .rgt_op(net_6883[0:7]),
     .bot_op(slf_op_14_11[7:0]), .bl(bl[765:712]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_4509), .purst(purst), .slf_op(net_6799[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_15_11[7:0]),
     .bnl_op(slf_op_13_11[7:0]), .tnr_op(net_6855[0:7]),
     .tnl_op(slf_op_13_03[7:0]));
ltile4rev I_13_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4565), .lft_op(lft_op_13_02[7:0]),
     .sp12_h_l(sp12_h_l_13_02[23:0]), .sp4_h_l(sp4_h_l_13_02[47:0]),
     .sp4_v_b(sp4_v_b_13_02[47:0]), .sp12_v_b(net_4601[0:23]),
     .sp12_h_r(net_4571[0:23]), .sp4_h_r(net_4572[0:47]),
     .sp12_v_t(net_4573[0:23]), .sp4_v_t(sp4_v_b_13_03[47:0]),
     .sp4_r_v_b(net_4575[0:47]), .wl(wl[207:192]),
     .top_op(slf_op_13_03[7:0]), .rgt_op(net_6799[0:7]),
     .bot_op(slf_op_13_11[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_4593), .purst(purst), .slf_op(slf_op_13_02[7:0]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_14_11[7:0]),
     .bnl_op(lft_op_13_01[7:0]), .tnr_op(net_6827[0:7]),
     .tnl_op(lft_op_13_03[7:0]));
ltile4rev I_13_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4593), .lft_op(lft_op_13_01[7:0]),
     .sp12_h_l(sp12_h_l_13_01[23:0]), .sp4_h_l(sp4_h_l_13_01[47:0]),
     .sp4_v_b(sp4_v_b_13_11[47:0]), .sp12_v_b(sp12_v_b_13_11[23:0]),
     .sp12_h_r(net_4599[0:23]), .sp4_h_r(net_4600[0:47]),
     .sp12_v_t(net_4601[0:23]), .sp4_v_t(sp4_v_b_13_02[47:0]),
     .sp4_r_v_b(sp4_v_b_14_11[47:0]), .wl(wl[191:176]),
     .top_op(slf_op_13_02[7:0]), .rgt_op(slf_op_14_11[7:0]),
     .bot_op(bot_op_13_11[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(carry_in_13_11), .purst(purst),
     .slf_op(slf_op_13_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_13_11[7:0]), .bnl_op(bnl_op_13_11[7:0]),
     .tnr_op(net_6799[0:7]), .tnl_op(lft_op_13_02[7:0]));
ltile4rev I_18_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4621), .lft_op(slf_op_17_11[7:0]),
     .sp12_h_l(net_4319[0:23]), .sp4_h_l(net_4320[0:47]),
     .sp4_v_b(sp4_v_b_18_11[47:0]), .sp12_v_b(sp12_v_b_18_11[23:0]),
     .sp12_h_r(net_4627[0:23]), .sp4_h_r(net_4628[0:47]),
     .sp12_v_t(net_4629[0:23]), .sp4_v_t(net_4351[0:47]),
     .sp4_r_v_b(sp4_v_b_19_11[47:0]), .wl(wl[191:176]),
     .top_op(net_6911[0:7]), .rgt_op(slf_op_19_11[7:0]),
     .bot_op(bot_op_18_11[7:0]), .bl(bl[981:928]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(carry_in_18_11), .purst(purst),
     .slf_op(slf_op_18_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_18_11[7:0]), .bnl_op(bnl_op_18_11[7:0]),
     .tnr_op(net_4645[0:7]), .tnl_op(net_7051[0:7]));
ltile4rev I_20_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4649), .lft_op(slf_op_19_11[7:0]),
     .sp12_h_l(net_4286[0:23]), .sp4_h_l(net_4295[0:47]),
     .sp4_v_b(sp4_v_b_20_11[47:0]), .sp12_v_b(sp12_v_b_20_11[23:0]),
     .sp12_h_r(net_4655[0:23]), .sp4_h_r(net_4656[0:47]),
     .sp12_v_t(net_4657[0:23]), .sp4_v_t(net_4292[0:47]),
     .sp4_r_v_b(sp4_v_b_21_11[47:0]), .wl(wl[191:176]),
     .top_op(net_4207[0:7]), .rgt_op(slf_op_21_11[7:0]),
     .bot_op(bot_op_20_11[7:0]), .bl(bl[1077:1024]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(carry_in_20_11), .purst(purst),
     .slf_op(slf_op_20_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_20_11[7:0]), .bnl_op(bnl_op_20_11[7:0]),
     .tnr_op(net_7135[0:7]), .tnl_op(net_4645[0:7]));
ltile4rev I_20_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4677), .lft_op(net_4645[0:7]),
     .sp12_h_l(net_4285[0:23]), .sp4_h_l(net_4294[0:47]),
     .sp4_v_b(net_4292[0:47]), .sp12_v_b(net_4657[0:23]),
     .sp12_h_r(net_4683[0:23]), .sp4_h_r(net_4684[0:47]),
     .sp12_v_t(net_4685[0:23]), .sp4_v_t(net_4206[0:47]),
     .sp4_r_v_b(net_4687[0:47]), .wl(wl[207:192]),
     .top_op(net_4689[0:7]), .rgt_op(net_7135[0:7]),
     .bot_op(slf_op_20_11[7:0]), .bl(bl[1077:1024]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_4649), .purst(purst), .slf_op(net_4207[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_21_11[7:0]),
     .bnl_op(slf_op_19_11[7:0]), .tnr_op(net_7163[0:7]),
     .tnl_op(net_4262[0:7]));
ltile4rev I_21_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4705), .lft_op(net_4207[0:7]),
     .sp12_h_l(net_4683[0:23]), .sp4_h_l(net_4684[0:47]),
     .sp4_v_b(net_4687[0:47]), .sp12_v_b(net_4741[0:23]),
     .sp12_h_r(net_4711[0:23]), .sp4_h_r(net_4712[0:47]),
     .sp12_v_t(net_4713[0:23]), .sp4_v_t(net_7123[0:47]),
     .sp4_r_v_b(net_4715[0:47]), .wl(wl[207:192]),
     .top_op(net_7163[0:7]), .rgt_op(net_7219[0:7]),
     .bot_op(slf_op_21_11[7:0]), .bl(bl[1131:1078]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_4733), .purst(purst), .slf_op(net_7135[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_22_11[7:0]),
     .bnl_op(slf_op_20_11[7:0]), .tnr_op(net_4729[0:7]),
     .tnl_op(net_4689[0:7]));
ltile4rev I_21_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4733), .lft_op(slf_op_20_11[7:0]),
     .sp12_h_l(net_4655[0:23]), .sp4_h_l(net_4656[0:47]),
     .sp4_v_b(sp4_v_b_21_11[47:0]), .sp12_v_b(sp12_v_b_21_11[23:0]),
     .sp12_h_r(net_4739[0:23]), .sp4_h_r(net_4740[0:47]),
     .sp12_v_t(net_4741[0:23]), .sp4_v_t(net_4687[0:47]),
     .sp4_r_v_b(sp4_v_b_22_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7135[0:7]), .rgt_op(slf_op_22_11[7:0]),
     .bot_op(bot_op_21_11[7:0]), .bl(bl[1131:1078]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(carry_in_21_11), .purst(purst),
     .slf_op(slf_op_21_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_21_11[7:0]), .bnl_op(bnl_op_21_11[7:0]),
     .tnr_op(net_7219[0:7]), .tnl_op(net_4207[0:7]));
ltile4rev I_17_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_4761), .lft_op(net_4867[0:7]),
     .sp12_h_l(net_4907[0:23]), .sp4_h_l(net_4908[0:47]),
     .sp4_v_b(net_4911[0:47]), .sp12_v_b(net_6925[0:23]),
     .sp12_h_r(net_4767[0:23]), .sp4_h_r(net_4768[0:47]),
     .sp12_v_t(net_4769[0:23]), .sp4_v_t(net_4883[0:47]),
     .sp4_r_v_b(net_4771[0:47]), .wl(wl[255:240]),
     .top_op(net_6267[0:7]), .rgt_op(net_4811[0:7]),
     .bot_op(net_4923[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_6917), .purst(purst), .slf_op(net_4895[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_4783[0:7]),
     .bnl_op(net_4839[0:7]), .tnr_op(net_6127[0:7]),
     .tnl_op(net_6183[0:7]));
ltile4rev I_17_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4789), .lft_op(net_6183[0:7]),
     .sp12_h_l(net_4879[0:23]), .sp4_h_l(net_4880[0:47]),
     .sp4_v_b(net_4883[0:47]), .sp12_v_b(net_4769[0:23]),
     .sp12_h_r(net_4795[0:23]), .sp4_h_r(net_4796[0:47]),
     .sp12_v_t(net_4797[0:23]), .sp4_v_t(net_6255[0:47]),
     .sp4_r_v_b(net_4799[0:47]), .wl(wl[271:256]),
     .top_op(net_6239[0:7]), .rgt_op(net_6127[0:7]),
     .bot_op(net_4895[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_4761), .purst(purst), .slf_op(net_6267[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_4811[0:7]),
     .bnl_op(net_4867[0:7]), .tnr_op(net_6155[0:7]),
     .tnl_op(net_6211[0:7]));
ltile4rev I_15_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_4817), .lft_op(net_5035[0:7]),
     .sp12_h_l(net_4963[0:23]), .sp4_h_l(net_4964[0:47]),
     .sp4_v_b(net_4967[0:47]), .sp12_v_b(net_6981[0:23]),
     .sp12_h_r(net_4823[0:23]), .sp4_h_r(net_4824[0:47]),
     .sp12_v_t(net_4825[0:23]), .sp4_v_t(net_4995[0:47]),
     .sp4_r_v_b(net_4827[0:47]), .wl(wl[255:240]),
     .top_op(net_6099[0:7]), .rgt_op(net_4867[0:7]),
     .bot_op(net_4979[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_6973), .purst(purst), .slf_op(net_5007[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_4839[0:7]),
     .bnl_op(net_5063[0:7]), .tnr_op(net_6183[0:7]),
     .tnl_op(net_6015[0:7]));
ltile4rev I_15_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4845), .lft_op(net_6015[0:7]),
     .sp12_h_l(net_4991[0:23]), .sp4_h_l(net_4992[0:47]),
     .sp4_v_b(net_4995[0:47]), .sp12_v_b(net_4825[0:23]),
     .sp12_h_r(net_4851[0:23]), .sp4_h_r(net_4852[0:47]),
     .sp12_v_t(net_4853[0:23]), .sp4_v_t(net_6087[0:47]),
     .sp4_r_v_b(net_4855[0:47]), .wl(wl[271:256]),
     .top_op(net_6071[0:7]), .rgt_op(net_6183[0:7]),
     .bot_op(net_5007[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_4817), .purst(purst), .slf_op(net_6099[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_4867[0:7]),
     .bnl_op(net_5035[0:7]), .tnr_op(net_6211[0:7]),
     .tnl_op(net_6043[0:7]));
ltile4rev I_16_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4873), .lft_op(net_6099[0:7]),
     .sp12_h_l(net_4851[0:23]), .sp4_h_l(net_4852[0:47]),
     .sp4_v_b(net_4855[0:47]), .sp12_v_b(net_4909[0:23]),
     .sp12_h_r(net_4879[0:23]), .sp4_h_r(net_4880[0:47]),
     .sp12_v_t(net_4881[0:23]), .sp4_v_t(net_6171[0:47]),
     .sp4_r_v_b(net_4883[0:47]), .wl(wl[271:256]),
     .top_op(net_6211[0:7]), .rgt_op(net_6267[0:7]),
     .bot_op(net_4867[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_4901), .purst(purst), .slf_op(net_6183[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_4895[0:7]),
     .bnl_op(net_5007[0:7]), .tnr_op(net_6239[0:7]),
     .tnl_op(net_6071[0:7]));
ltile4rev I_16_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_4901), .lft_op(net_5007[0:7]),
     .sp12_h_l(net_4823[0:23]), .sp4_h_l(net_4824[0:47]),
     .sp4_v_b(net_4827[0:47]), .sp12_v_b(net_7009[0:23]),
     .sp12_h_r(net_4907[0:23]), .sp4_h_r(net_4908[0:47]),
     .sp12_v_t(net_4909[0:23]), .sp4_v_t(net_4855[0:47]),
     .sp4_r_v_b(net_4911[0:47]), .wl(wl[255:240]),
     .top_op(net_6183[0:7]), .rgt_op(net_4895[0:7]),
     .bot_op(net_4839[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_7001), .purst(purst), .slf_op(net_4867[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_4923[0:7]),
     .bnl_op(net_4979[0:7]), .tnr_op(net_6267[0:7]),
     .tnl_op(net_6099[0:7]));
ltile4rev I_18_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4929), .lft_op(net_6267[0:7]),
     .sp12_h_l(net_4795[0:23]), .sp4_h_l(net_4796[0:47]),
     .sp4_v_b(net_4799[0:47]), .sp12_v_b(net_5077[0:23]),
     .sp12_h_r(net_4935[0:23]), .sp4_h_r(net_4936[0:47]),
     .sp12_v_t(net_4937[0:23]), .sp4_v_t(net_6115[0:47]),
     .sp4_r_v_b(net_4939[0:47]), .wl(wl[271:256]),
     .top_op(net_6155[0:7]), .rgt_op(net_6323[0:7]),
     .bot_op(net_4811[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_5069), .purst(purst), .slf_op(net_6127[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_7081[0:7]),
     .bnl_op(net_4895[0:7]), .tnr_op(net_4138[0:7]),
     .tnl_op(net_6239[0:7]));
ltile4rev I_14_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_4957), .lft_op(slf_op_13_05[7:0]),
     .sp12_h_l(net_5047[0:23]), .sp4_h_l(net_5048[0:47]),
     .sp4_v_b(net_5051[0:47]), .sp12_v_b(net_6841[0:23]),
     .sp12_h_r(net_4963[0:23]), .sp4_h_r(net_4964[0:47]),
     .sp12_v_t(net_4965[0:23]), .sp4_v_t(net_5023[0:47]),
     .sp4_r_v_b(net_4967[0:47]), .wl(wl[255:240]),
     .top_op(net_6015[0:7]), .rgt_op(net_5007[0:7]),
     .bot_op(net_5063[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_6833), .purst(purst), .slf_op(net_5035[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_4979[0:7]),
     .bnl_op(slf_op_13_04[7:0]), .tnr_op(net_6099[0:7]),
     .tnl_op(slf_op_13_06[7:0]));
ltile4rev I_14_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4985), .lft_op(slf_op_13_06[7:0]),
     .sp12_h_l(net_5019[0:23]), .sp4_h_l(net_5020[0:47]),
     .sp4_v_b(net_5023[0:47]), .sp12_v_b(net_4965[0:23]),
     .sp12_h_r(net_4991[0:23]), .sp4_h_r(net_4992[0:47]),
     .sp12_v_t(net_4993[0:23]), .sp4_v_t(net_6003[0:47]),
     .sp4_r_v_b(net_4995[0:47]), .wl(wl[271:256]),
     .top_op(net_6043[0:7]), .rgt_op(net_6099[0:7]),
     .bot_op(net_5035[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_4957), .purst(purst), .slf_op(net_6015[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5007[0:7]),
     .bnl_op(slf_op_13_05[7:0]), .tnr_op(net_6071[0:7]),
     .tnl_op(slf_op_13_07[7:0]));
ltile4rev I_13_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5013), .lft_op(lft_op_13_06[7:0]),
     .sp12_h_l(sp12_h_l_13_06[23:0]), .sp4_h_l(sp4_h_l_13_06[47:0]),
     .sp4_v_b(sp4_v_b_13_06[47:0]), .sp12_v_b(net_5049[0:23]),
     .sp12_h_r(net_5019[0:23]), .sp4_h_r(net_5020[0:47]),
     .sp12_v_t(net_5021[0:23]), .sp4_v_t(sp4_v_b_13_07[47:0]),
     .sp4_r_v_b(net_5023[0:47]), .wl(wl[271:256]),
     .top_op(slf_op_13_07[7:0]), .rgt_op(net_6015[0:7]),
     .bot_op(slf_op_13_05[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5041), .purst(purst), .slf_op(slf_op_13_06[7:0]),
     .pgate(pgate[271:256]), .bnr_op(net_5035[0:7]),
     .bnl_op(lft_op_13_05[7:0]), .tnr_op(net_6043[0:7]),
     .tnl_op(lft_op_13_07[7:0]));
ltile4rev I_13_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5041), .lft_op(lft_op_13_05[7:0]),
     .sp12_h_l(sp12_h_l_13_05[23:0]), .sp4_h_l(sp4_h_l_13_05[47:0]),
     .sp4_v_b(sp4_v_b_13_05[47:0]), .sp12_v_b(net_6813[0:23]),
     .sp12_h_r(net_5047[0:23]), .sp4_h_r(net_5048[0:47]),
     .sp12_v_t(net_5049[0:23]), .sp4_v_t(sp4_v_b_13_06[47:0]),
     .sp4_r_v_b(net_5051[0:47]), .wl(wl[255:240]),
     .top_op(slf_op_13_06[7:0]), .rgt_op(net_5035[0:7]),
     .bot_op(slf_op_13_04[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_6805), .purst(purst), .slf_op(slf_op_13_05[7:0]),
     .pgate(pgate[255:240]), .bnr_op(net_5063[0:7]),
     .bnl_op(lft_op_13_04[7:0]), .tnr_op(net_6015[0:7]),
     .tnl_op(lft_op_13_06[7:0]));
ltile4rev I_18_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5069), .lft_op(net_4895[0:7]),
     .sp12_h_l(net_4767[0:23]), .sp4_h_l(net_4768[0:47]),
     .sp4_v_b(net_4771[0:47]), .sp12_v_b(net_7065[0:23]),
     .sp12_h_r(net_5075[0:23]), .sp4_h_r(net_5076[0:47]),
     .sp12_v_t(net_5077[0:23]), .sp4_v_t(net_4799[0:47]),
     .sp4_r_v_b(net_5079[0:47]), .wl(wl[255:240]),
     .top_op(net_6127[0:7]), .rgt_op(net_7081[0:7]),
     .bot_op(net_4783[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_7057), .purst(purst), .slf_op(net_4811[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5091[0:7]),
     .bnl_op(net_4923[0:7]), .tnr_op(net_6323[0:7]),
     .tnl_op(net_6267[0:7]));
ltile4rev I_20_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5097), .lft_op(net_7081[0:7]),
     .sp12_h_l(net_4162[0:23]), .sp4_h_l(net_4171[0:47]),
     .sp4_v_b(net_4169[0:47]), .sp12_v_b(net_7149[0:23]),
     .sp12_h_r(net_5103[0:23]), .sp4_h_r(net_5104[0:47]),
     .sp12_v_t(net_5105[0:23]), .sp4_v_t(net_4168[0:47]),
     .sp4_r_v_b(net_5107[0:47]), .wl(wl[255:240]),
     .top_op(net_4122[0:7]), .rgt_op(net_5147[0:7]),
     .bot_op(net_4155[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_7141), .purst(purst), .slf_op(net_4198[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5119[0:7]),
     .bnl_op(net_5091[0:7]), .tnr_op(net_6351[0:7]),
     .tnl_op(net_6323[0:7]));
ltile4rev I_20_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5125), .lft_op(net_6323[0:7]),
     .sp12_h_l(net_4161[0:23]), .sp4_h_l(net_4170[0:47]),
     .sp4_v_b(net_4168[0:47]), .sp12_v_b(net_5105[0:23]),
     .sp12_h_r(net_5131[0:23]), .sp4_h_r(net_5132[0:47]),
     .sp12_v_t(net_5133[0:23]), .sp4_v_t(net_4121[0:47]),
     .sp4_r_v_b(net_5135[0:47]), .wl(wl[271:256]),
     .top_op(net_5137[0:7]), .rgt_op(net_6351[0:7]),
     .bot_op(net_4198[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_5097), .purst(purst), .slf_op(net_4122[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5147[0:7]),
     .bnl_op(net_7081[0:7]), .tnr_op(net_6379[0:7]),
     .tnl_op(net_4138[0:7]));
ltile4rev I_21_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5153), .lft_op(net_4122[0:7]),
     .sp12_h_l(net_5131[0:23]), .sp4_h_l(net_5132[0:47]),
     .sp4_v_b(net_5135[0:47]), .sp12_v_b(net_5189[0:23]),
     .sp12_h_r(net_5159[0:23]), .sp4_h_r(net_5160[0:47]),
     .sp12_v_t(net_5161[0:23]), .sp4_v_t(net_6339[0:47]),
     .sp4_r_v_b(net_5163[0:47]), .wl(wl[271:256]),
     .top_op(net_6379[0:7]), .rgt_op(net_6435[0:7]),
     .bot_op(net_5147[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_5181), .purst(purst), .slf_op(net_6351[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_7193[0:7]),
     .bnl_op(net_4198[0:7]), .tnr_op(net_5177[0:7]),
     .tnl_op(net_5137[0:7]));
ltile4rev I_21_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5181), .lft_op(net_4198[0:7]),
     .sp12_h_l(net_5103[0:23]), .sp4_h_l(net_5104[0:47]),
     .sp4_v_b(net_5107[0:47]), .sp12_v_b(net_7177[0:23]),
     .sp12_h_r(net_5187[0:23]), .sp4_h_r(net_5188[0:47]),
     .sp12_v_t(net_5189[0:23]), .sp4_v_t(net_5135[0:47]),
     .sp4_r_v_b(net_5191[0:47]), .wl(wl[255:240]),
     .top_op(net_6351[0:7]), .rgt_op(net_7193[0:7]),
     .bot_op(net_5119[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_7169), .purst(purst), .slf_op(net_5147[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_7191[0:7]),
     .bnl_op(net_4155[0:7]), .tnr_op(net_6435[0:7]),
     .tnl_op(net_4122[0:7]));
ltile4rev I_23_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5209), .lft_op(net_7193[0:7]),
     .sp12_h_l(net_5271[0:23]), .sp4_h_l(net_5272[0:47]),
     .sp4_v_b(net_5275[0:47]), .sp12_v_b(net_7373[0:23]),
     .sp12_h_r(net_5215[0:23]), .sp4_h_r(net_5216[0:47]),
     .sp12_v_t(net_5217[0:23]), .sp4_v_t(net_5303[0:47]),
     .sp4_r_v_b(net_5219[0:47]), .wl(wl[255:240]),
     .top_op(net_6519[0:7]), .rgt_op(net_5371[0:7]),
     .bot_op(net_5287[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_7365), .purst(purst), .slf_op(net_5315[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5231[0:7]),
     .bnl_op(net_7191[0:7]), .tnr_op(net_6463[0:7]),
     .tnl_op(net_6435[0:7]));
ltile4rev I_24_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5237), .lft_op(net_6519[0:7]),
     .sp12_h_l(net_5355[0:23]), .sp4_h_l(net_5356[0:47]),
     .sp4_v_b(net_5359[0:47]), .sp12_v_b(net_5329[0:23]),
     .sp12_h_r(net_5243[0:23]), .sp4_h_r(net_5244[0:47]),
     .sp12_v_t(net_5245[0:23]), .sp4_v_t(net_6451[0:47]),
     .sp4_r_v_b(net_5247[0:47]), .wl(wl[271:256]),
     .top_op(net_6603[0:7]), .rgt_op({io_r_05[3], io_r_05[2],
     io_r_05[1], io_r_05[0], io_r_05[3], io_r_05[2], io_r_05[1],
     io_r_05[0]}), .bot_op(net_5371[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_5321), .purst(purst), .slf_op(net_6463[0:7]),
     .pgate(pgate[271:256]), .bnr_op({io_r_04[3], io_r_04[2],
     io_r_04[1], io_r_04[0], io_r_04[3], io_r_04[2], io_r_04[1],
     io_r_04[0]}), .bnl_op(net_5315[0:7]), .tnr_op({io_r_06[3],
     io_r_06[2], io_r_06[1], io_r_06[0], io_r_06[3], io_r_06[2],
     io_r_06[1], io_r_06[0]}), .tnl_op(net_6547[0:7]));
ltile4rev I_22_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5265), .lft_op(net_5147[0:7]),
     .sp12_h_l(net_5187[0:23]), .sp4_h_l(net_5188[0:47]),
     .sp4_v_b(net_5191[0:47]), .sp12_v_b(net_7317[0:23]),
     .sp12_h_r(net_5271[0:23]), .sp4_h_r(net_5272[0:47]),
     .sp12_v_t(net_5273[0:23]), .sp4_v_t(net_5163[0:47]),
     .sp4_r_v_b(net_5275[0:47]), .wl(wl[255:240]),
     .top_op(net_6435[0:7]), .rgt_op(net_5315[0:7]),
     .bot_op(net_7191[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_7309), .purst(purst), .slf_op(net_7193[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5287[0:7]),
     .bnl_op(net_5119[0:7]), .tnr_op(net_6519[0:7]),
     .tnl_op(net_6351[0:7]));
ltile4rev I_22_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5293), .lft_op(net_6351[0:7]),
     .sp12_h_l(net_5159[0:23]), .sp4_h_l(net_5160[0:47]),
     .sp4_v_b(net_5163[0:47]), .sp12_v_b(net_5273[0:23]),
     .sp12_h_r(net_5299[0:23]), .sp4_h_r(net_5300[0:47]),
     .sp12_v_t(net_5301[0:23]), .sp4_v_t(net_6423[0:47]),
     .sp4_r_v_b(net_5303[0:47]), .wl(wl[271:256]),
     .top_op(net_5177[0:7]), .rgt_op(net_6519[0:7]),
     .bot_op(net_7193[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_5265), .purst(purst), .slf_op(net_6435[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5315[0:7]),
     .bnl_op(net_5147[0:7]), .tnr_op(net_6547[0:7]),
     .tnl_op(net_6379[0:7]));
ltile4rev I_24_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5321), .lft_op(net_5315[0:7]),
     .sp12_h_l(net_5215[0:23]), .sp4_h_l(net_5216[0:47]),
     .sp4_v_b(net_5219[0:47]), .sp12_v_b(net_7261[0:23]),
     .sp12_h_r(net_5327[0:23]), .sp4_h_r(net_5328[0:47]),
     .sp12_v_t(net_5329[0:23]), .sp4_v_t(net_5359[0:47]),
     .sp4_r_v_b(net_5331[0:47]), .wl(wl[255:240]),
     .top_op(net_6463[0:7]), .rgt_op({io_r_04[3], io_r_04[2],
     io_r_04[1], io_r_04[0], io_r_04[3], io_r_04[2], io_r_04[1],
     io_r_04[0]}), .bot_op(net_5231[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_7253), .purst(purst), .slf_op(net_5371[0:7]),
     .pgate(pgate[255:240]), .bnr_op({io_r_03[3], io_r_03[2],
     io_r_03[1], io_r_03[0], io_r_03[3], io_r_03[2], io_r_03[1],
     io_r_03[0]}), .bnl_op(net_5287[0:7]), .tnr_op({io_r_05[3],
     io_r_05[2], io_r_05[1], io_r_05[0], io_r_05[3], io_r_05[2],
     io_r_05[1], io_r_05[0]}), .tnl_op(net_6519[0:7]));
ltile4rev I_23_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5349), .lft_op(net_6435[0:7]),
     .sp12_h_l(net_5299[0:23]), .sp4_h_l(net_5300[0:47]),
     .sp4_v_b(net_5303[0:47]), .sp12_v_b(net_5217[0:23]),
     .sp12_h_r(net_5355[0:23]), .sp4_h_r(net_5356[0:47]),
     .sp12_v_t(net_5357[0:23]), .sp4_v_t(net_6507[0:47]),
     .sp4_r_v_b(net_5359[0:47]), .wl(wl[271:256]),
     .top_op(net_6547[0:7]), .rgt_op(net_6463[0:7]),
     .bot_op(net_5315[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_5209), .purst(purst), .slf_op(net_6519[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5371[0:7]),
     .bnl_op(net_7193[0:7]), .tnr_op(net_6603[0:7]),
     .tnl_op(net_5177[0:7]));
ltile4rev I_17_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5377), .lft_op(net_5483[0:7]),
     .sp12_h_l(net_5523[0:23]), .sp4_h_l(net_5524[0:47]),
     .sp4_v_b(net_5527[0:47]), .sp12_v_b(net_6141[0:23]),
     .sp12_h_r(net_5383[0:23]), .sp4_h_r(net_5384[0:47]),
     .sp12_v_t(net_5385[0:23]), .sp4_v_t(net_5499[0:47]),
     .sp4_r_v_b(net_5387[0:47]), .wl(wl[319:304]),
     .top_op(net_7511[0:7]), .rgt_op(net_5427[0:7]),
     .bot_op(net_5539[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_6133), .purst(purst), .slf_op(net_5511[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5399[0:7]),
     .bnl_op(net_5455[0:7]), .tnr_op(net_7545[0:7]),
     .tnl_op(net_7477[0:7]));
ltile4rev I_17_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8226), .lft_op(net_7477[0:7]),
     .sp12_h_l(net_5495[0:23]), .sp4_h_l(net_5496[0:47]),
     .sp4_v_b(net_5499[0:47]), .sp12_v_b(net_5385[0:23]),
     .sp12_h_r(net_5411[0:23]), .sp4_h_r(net_5412[0:47]),
     .sp12_v_t(net_5413[0:23]), .sp4_v_t(net_7539[0:47]),
     .sp4_r_v_b(net_5415[0:47]), .wl(wl[335:320]), .top_op({io_t_17[3],
     io_t_17[2], io_t_17[1], io_t_17[0], io_t_17[3], io_t_17[2],
     io_t_17[1], io_t_17[0]}), .rgt_op(net_7545[0:7]),
     .bot_op(net_5511[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_5377), .purst(purst), .slf_op(net_7511[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5427[0:7]),
     .bnl_op(net_5483[0:7]), .tnr_op({io_t_18[3], io_t_18[2],
     io_t_18[1], io_t_18[0], io_t_18[3], io_t_18[2], io_t_18[1],
     io_t_18[0]}), .tnl_op({io_t_16[3], io_t_16[2], io_t_16[1],
     io_t_16[0], io_t_16[3], io_t_16[2], io_t_16[1], io_t_16[0]}));
ltile4rev I_15_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5433), .lft_op(net_5651[0:7]),
     .sp12_h_l(net_5579[0:23]), .sp4_h_l(net_5580[0:47]),
     .sp4_v_b(net_5583[0:47]), .sp12_v_b(net_6197[0:23]),
     .sp12_h_r(net_5439[0:23]), .sp4_h_r(net_5440[0:47]),
     .sp12_v_t(net_5441[0:23]), .sp4_v_t(net_5611[0:47]),
     .sp4_r_v_b(net_5443[0:47]), .wl(wl[319:304]),
     .top_op(net_7443[0:7]), .rgt_op(net_5483[0:7]),
     .bot_op(net_5595[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_6189), .purst(purst), .slf_op(net_5623[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5455[0:7]),
     .bnl_op(net_5679[0:7]), .tnr_op(net_7477[0:7]),
     .tnl_op(net_8055[0:7]));
ltile4rev I_15_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8221), .lft_op(net_8055[0:7]),
     .sp12_h_l(net_5607[0:23]), .sp4_h_l(net_5608[0:47]),
     .sp4_v_b(net_5611[0:47]), .sp12_v_b(net_5441[0:23]),
     .sp12_h_r(net_5467[0:23]), .sp4_h_r(net_5468[0:47]),
     .sp12_v_t(net_5469[0:23]), .sp4_v_t(net_7471[0:47]),
     .sp4_r_v_b(net_5471[0:47]), .wl(wl[335:320]), .top_op({io_t_15[3],
     io_t_15[2], io_t_15[1], io_t_15[0], io_t_15[3], io_t_15[2],
     io_t_15[1], io_t_15[0]}), .rgt_op(net_7477[0:7]),
     .bot_op(net_5623[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_5433), .purst(purst), .slf_op(net_7443[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5483[0:7]),
     .bnl_op(net_5651[0:7]), .tnr_op({io_t_16[3], io_t_16[2],
     io_t_16[1], io_t_16[0], io_t_16[3], io_t_16[2], io_t_16[1],
     io_t_16[0]}), .tnl_op({io_t_14[3], io_t_14[2], io_t_14[1],
     io_t_14[0], io_t_14[3], io_t_14[2], io_t_14[1], io_t_14[0]}));
ltile4rev I_16_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8224), .lft_op(net_7443[0:7]),
     .sp12_h_l(net_5467[0:23]), .sp4_h_l(net_5468[0:47]),
     .sp4_v_b(net_5471[0:47]), .sp12_v_b(net_5525[0:23]),
     .sp12_h_r(net_5495[0:23]), .sp4_h_r(net_5496[0:47]),
     .sp12_v_t(net_5497[0:23]), .sp4_v_t(net_7505[0:47]),
     .sp4_r_v_b(net_5499[0:47]), .wl(wl[335:320]), .top_op({io_t_16[3],
     io_t_16[2], io_t_16[1], io_t_16[0], io_t_16[3], io_t_16[2],
     io_t_16[1], io_t_16[0]}), .rgt_op(net_7511[0:7]),
     .bot_op(net_5483[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_5517), .purst(purst), .slf_op(net_7477[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5511[0:7]),
     .bnl_op(net_5623[0:7]), .tnr_op({io_t_17[3], io_t_17[2],
     io_t_17[1], io_t_17[0], io_t_17[3], io_t_17[2], io_t_17[1],
     io_t_17[0]}), .tnl_op({io_t_15[3], io_t_15[2], io_t_15[1],
     io_t_15[0], io_t_15[3], io_t_15[2], io_t_15[1], io_t_15[0]}));
ltile4rev I_16_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5517), .lft_op(net_5623[0:7]),
     .sp12_h_l(net_5439[0:23]), .sp4_h_l(net_5440[0:47]),
     .sp4_v_b(net_5443[0:47]), .sp12_v_b(net_6225[0:23]),
     .sp12_h_r(net_5523[0:23]), .sp4_h_r(net_5524[0:47]),
     .sp12_v_t(net_5525[0:23]), .sp4_v_t(net_5471[0:47]),
     .sp4_r_v_b(net_5527[0:47]), .wl(wl[319:304]),
     .top_op(net_7477[0:7]), .rgt_op(net_5511[0:7]),
     .bot_op(net_5455[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_6217), .purst(purst), .slf_op(net_5483[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5539[0:7]),
     .bnl_op(net_5595[0:7]), .tnr_op(net_7511[0:7]),
     .tnl_op(net_7443[0:7]));
ltile4rev I_18_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8218), .lft_op(net_7511[0:7]),
     .sp12_h_l(net_5411[0:23]), .sp4_h_l(net_5412[0:47]),
     .sp4_v_b(net_5415[0:47]), .sp12_v_b(net_5693[0:23]),
     .sp12_h_r(net_5551[0:23]), .sp4_h_r(net_5552[0:47]),
     .sp12_v_t(net_5553[0:23]), .sp4_v_t(net_5554[0:47]),
     .sp4_r_v_b(net_5555[0:47]), .wl(wl[335:320]), .top_op({io_t_18[3],
     io_t_18[2], io_t_18[1], io_t_18[0], io_t_18[3], io_t_18[2],
     io_t_18[1], io_t_18[0]}), .rgt_op(net_8157[0:7]),
     .bot_op(net_5427[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_5685), .purst(purst), .slf_op(net_7545[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_6297[0:7]),
     .bnl_op(net_5511[0:7]), .tnr_op({io_t_19[3], io_t_19[2],
     io_t_19[1], io_t_19[0], io_t_19[3], io_t_19[2], io_t_19[1],
     io_t_19[0]}), .tnl_op({io_t_17[3], io_t_17[2], io_t_17[1],
     io_t_17[0], io_t_17[3], io_t_17[2], io_t_17[1], io_t_17[0]}));
ltile4rev I_14_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5573), .lft_op(slf_op_13_09[7:0]),
     .sp12_h_l(net_5663[0:23]), .sp4_h_l(net_5664[0:47]),
     .sp4_v_b(net_5667[0:47]), .sp12_v_b(net_6057[0:23]),
     .sp12_h_r(net_5579[0:23]), .sp4_h_r(net_5580[0:47]),
     .sp12_v_t(net_5581[0:23]), .sp4_v_t(net_5639[0:47]),
     .sp4_r_v_b(net_5583[0:47]), .wl(wl[319:304]),
     .top_op(net_8055[0:7]), .rgt_op(net_5623[0:7]),
     .bot_op(net_5679[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_6049), .purst(purst), .slf_op(net_5651[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5595[0:7]),
     .bnl_op(slf_op_13_08[7:0]), .tnr_op(net_7443[0:7]),
     .tnl_op(slf_op_13_10[7:0]));
ltile4rev I_14_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8198), .lft_op(slf_op_13_10[7:0]),
     .sp12_h_l(net_5635[0:23]), .sp4_h_l(net_5636[0:47]),
     .sp4_v_b(net_5639[0:47]), .sp12_v_b(net_5581[0:23]),
     .sp12_h_r(net_5607[0:23]), .sp4_h_r(net_5608[0:47]),
     .sp12_v_t(net_5609[0:23]), .sp4_v_t(net_7437[0:47]),
     .sp4_r_v_b(net_5611[0:47]), .wl(wl[335:320]), .top_op({io_t_14[3],
     io_t_14[2], io_t_14[1], io_t_14[0], io_t_14[3], io_t_14[2],
     io_t_14[1], io_t_14[0]}), .rgt_op(net_7443[0:7]),
     .bot_op(net_5651[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_5573), .purst(purst), .slf_op(net_8055[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5623[0:7]),
     .bnl_op(slf_op_13_09[7:0]), .tnr_op({io_t_15[3], io_t_15[2],
     io_t_15[1], io_t_15[0], io_t_15[3], io_t_15[2], io_t_15[1],
     io_t_15[0]}), .tnl_op({slf_op_13_21[3], slf_op_13_21[2],
     slf_op_13_21[1], slf_op_13_21[0], slf_op_13_21[3],
     slf_op_13_21[2], slf_op_13_21[1], slf_op_13_21[0]}));
ltile4rev I_13_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8199), .lft_op(lft_op_13_10[7:0]),
     .sp12_h_l(sp12_h_l_13_10[23:0]), .sp4_h_l(sp4_h_l_13_10[47:0]),
     .sp4_v_b(sp4_v_b_13_10[47:0]), .sp12_v_b(net_5665[0:23]),
     .sp12_h_r(net_5635[0:23]), .sp4_h_r(net_5636[0:47]),
     .sp12_v_t(net_5637[0:23]), .sp4_v_t(net_8049[0:47]),
     .sp4_r_v_b(net_5639[0:47]), .wl(wl[335:320]),
     .top_op({slf_op_13_21[3], slf_op_13_21[2], slf_op_13_21[1],
     slf_op_13_21[0], slf_op_13_21[3], slf_op_13_21[2],
     slf_op_13_21[1], slf_op_13_21[0]}), .rgt_op(net_8055[0:7]),
     .bot_op(slf_op_13_09[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5657), .purst(purst), .slf_op(slf_op_13_10[7:0]),
     .pgate(pgate[335:320]), .bnr_op(net_5651[0:7]),
     .bnl_op(lft_op_13_09[7:0]), .tnr_op({io_t_14[3], io_t_14[2],
     io_t_14[1], io_t_14[0], io_t_14[3], io_t_14[2], io_t_14[1],
     io_t_14[0]}), .tnl_op({tnl_op_13_20[3], tnl_op_13_20[2],
     tnl_op_13_20[1], tnl_op_13_20[0], tnl_op_13_20[3],
     tnl_op_13_20[2], tnl_op_13_20[1], tnl_op_13_20[0]}));
ltile4rev I_13_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5657), .lft_op(lft_op_13_09[7:0]),
     .sp12_h_l(sp12_h_l_13_09[23:0]), .sp4_h_l(sp4_h_l_13_09[47:0]),
     .sp4_v_b(sp4_v_b_13_09[47:0]), .sp12_v_b(net_6029[0:23]),
     .sp12_h_r(net_5663[0:23]), .sp4_h_r(net_5664[0:47]),
     .sp12_v_t(net_5665[0:23]), .sp4_v_t(sp4_v_b_13_10[47:0]),
     .sp4_r_v_b(net_5667[0:47]), .wl(wl[319:304]),
     .top_op(slf_op_13_10[7:0]), .rgt_op(net_5651[0:7]),
     .bot_op(slf_op_13_08[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_6021), .purst(purst), .slf_op(slf_op_13_09[7:0]),
     .pgate(pgate[319:304]), .bnr_op(net_5679[0:7]),
     .bnl_op(lft_op_13_08[7:0]), .tnr_op(net_8055[0:7]),
     .tnl_op(lft_op_13_10[7:0]));
ltile4rev I_18_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5685), .lft_op(net_5511[0:7]),
     .sp12_h_l(net_5383[0:23]), .sp4_h_l(net_5384[0:47]),
     .sp4_v_b(net_5387[0:47]), .sp12_v_b(net_6281[0:23]),
     .sp12_h_r(net_5691[0:23]), .sp4_h_r(net_5692[0:47]),
     .sp12_v_t(net_5693[0:23]), .sp4_v_t(net_5415[0:47]),
     .sp4_r_v_b(net_5695[0:47]), .wl(wl[319:304]),
     .top_op(net_7545[0:7]), .rgt_op(net_6297[0:7]),
     .bot_op(net_5399[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_6273), .purst(purst), .slf_op(net_5427[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5707[0:7]),
     .bnl_op(net_5539[0:7]), .tnr_op(net_8157[0:7]),
     .tnl_op(net_7511[0:7]));
ltile4rev I_20_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5713), .lft_op(net_6297[0:7]),
     .sp12_h_l(net_4038[0:23]), .sp4_h_l(net_4047[0:47]),
     .sp4_v_b(net_4045[0:47]), .sp12_v_b(net_6365[0:23]),
     .sp12_h_r(net_5719[0:23]), .sp4_h_r(net_5720[0:47]),
     .sp12_v_t(net_5721[0:23]), .sp4_v_t(net_4044[0:47]),
     .sp4_r_v_b(net_5723[0:47]), .wl(wl[319:304]),
     .top_op(net_7613[0:7]), .rgt_op(net_5763[0:7]),
     .bot_op(net_4031[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_6357), .purst(purst), .slf_op(net_4113[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5735[0:7]),
     .bnl_op(net_5707[0:7]), .tnr_op(net_7681[0:7]),
     .tnl_op(net_8157[0:7]));
ltile4rev I_20_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8222), .lft_op(net_8157[0:7]),
     .sp12_h_l(net_4037[0:23]), .sp4_h_l(net_4046[0:47]),
     .sp4_v_b(net_4044[0:47]), .sp12_v_b(net_5721[0:23]),
     .sp12_h_r(net_5747[0:23]), .sp4_h_r(net_5748[0:47]),
     .sp12_v_t(net_5749[0:23]), .sp4_v_t(net_7675[0:47]),
     .sp4_r_v_b(net_5751[0:47]), .wl(wl[335:320]), .top_op({io_t_20[3],
     io_t_20[2], io_t_20[1], io_t_20[0], io_t_20[3], io_t_20[2],
     io_t_20[1], io_t_20[0]}), .rgt_op(net_7681[0:7]),
     .bot_op(net_4113[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_5713), .purst(purst), .slf_op(net_7613[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5763[0:7]),
     .bnl_op(net_6297[0:7]), .tnr_op({io_t_21[3], io_t_21[2],
     io_t_21[1], io_t_21[0], io_t_21[3], io_t_21[2], io_t_21[1],
     io_t_21[0]}), .tnl_op({io_t_19[3], io_t_19[2], io_t_19[1],
     io_t_19[0], io_t_19[3], io_t_19[2], io_t_19[1], io_t_19[0]}));
ltile4rev I_21_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8219), .lft_op(net_7613[0:7]),
     .sp12_h_l(net_5747[0:23]), .sp4_h_l(net_5748[0:47]),
     .sp4_v_b(net_5751[0:47]), .sp12_v_b(net_5805[0:23]),
     .sp12_h_r(net_5775[0:23]), .sp4_h_r(net_5776[0:47]),
     .sp12_v_t(net_5777[0:23]), .sp4_v_t(net_7709[0:47]),
     .sp4_r_v_b(net_5779[0:47]), .wl(wl[335:320]), .top_op({io_t_21[3],
     io_t_21[2], io_t_21[1], io_t_21[0], io_t_21[3], io_t_21[2],
     io_t_21[1], io_t_21[0]}), .rgt_op(net_7715[0:7]),
     .bot_op(net_5763[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_5797), .purst(purst), .slf_op(net_7681[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_6409[0:7]),
     .bnl_op(net_4113[0:7]), .tnr_op({io_t_22[3], io_t_22[2],
     io_t_22[1], io_t_22[0], io_t_22[3], io_t_22[2], io_t_22[1],
     io_t_22[0]}), .tnl_op({io_t_20[3], io_t_20[2], io_t_20[1],
     io_t_20[0], io_t_20[3], io_t_20[2], io_t_20[1], io_t_20[0]}));
ltile4rev I_21_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5797), .lft_op(net_4113[0:7]),
     .sp12_h_l(net_5719[0:23]), .sp4_h_l(net_5720[0:47]),
     .sp4_v_b(net_5723[0:47]), .sp12_v_b(net_6393[0:23]),
     .sp12_h_r(net_5803[0:23]), .sp4_h_r(net_5804[0:47]),
     .sp12_v_t(net_5805[0:23]), .sp4_v_t(net_5751[0:47]),
     .sp4_r_v_b(net_5807[0:47]), .wl(wl[319:304]),
     .top_op(net_7681[0:7]), .rgt_op(net_6409[0:7]),
     .bot_op(net_5735[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_6385), .purst(purst), .slf_op(net_5763[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_6407[0:7]),
     .bnl_op(net_4031[0:7]), .tnr_op(net_7715[0:7]),
     .tnl_op(net_7613[0:7]));
ltile4rev I_23_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5825), .lft_op(net_6409[0:7]),
     .sp12_h_l(net_5887[0:23]), .sp4_h_l(net_5888[0:47]),
     .sp4_v_b(net_5891[0:47]), .sp12_v_b(net_6589[0:23]),
     .sp12_h_r(net_5831[0:23]), .sp4_h_r(net_5832[0:47]),
     .sp12_v_t(net_5833[0:23]), .sp4_v_t(net_5919[0:47]),
     .sp4_r_v_b(net_5835[0:47]), .wl(wl[319:304]),
     .top_op(net_7749[0:7]), .rgt_op(net_5987[0:7]),
     .bot_op(net_5903[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_6581), .purst(purst), .slf_op(net_5931[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5847[0:7]),
     .bnl_op(net_6407[0:7]), .tnr_op(net_7783[0:7]),
     .tnl_op(net_7715[0:7]));
ltile4rev I_24_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8225), .lft_op(net_7749[0:7]),
     .sp12_h_l(net_5971[0:23]), .sp4_h_l(net_5972[0:47]),
     .sp4_v_b(net_5975[0:47]), .sp12_v_b(net_5945[0:23]),
     .sp12_h_r(net_5859[0:23]), .sp4_h_r(net_5860[0:47]),
     .sp12_v_t(net_5861[0:23]), .sp4_v_t(net_7811[0:47]),
     .sp4_r_v_b(net_5863[0:47]), .wl(wl[335:320]), .top_op({io_t_24[3],
     io_t_24[2], io_t_24[1], io_t_24[0], io_t_24[3], io_t_24[2],
     io_t_24[1], io_t_24[0]}), .rgt_op({slf_op_25_10[3],
     slf_op_25_10[2], slf_op_25_10[1], slf_op_25_10[0],
     slf_op_25_10[3], slf_op_25_10[2], slf_op_25_10[1],
     slf_op_25_10[0]}), .bot_op(net_5987[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_5937), .purst(purst), .slf_op(net_7783[0:7]),
     .pgate(pgate[335:320]), .bnr_op({io_r_08[3], io_r_08[2],
     io_r_08[1], io_r_08[0], io_r_08[3], io_r_08[2], io_r_08[1],
     io_r_08[0]}), .bnl_op(net_5931[0:7]), .tnr_op({tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .tnl_op({io_t_23[3], io_t_23[2], io_t_23[1], io_t_23[0],
     io_t_23[3], io_t_23[2], io_t_23[1], io_t_23[0]}));
ltile4rev I_22_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5881), .lft_op(net_5763[0:7]),
     .sp12_h_l(net_5803[0:23]), .sp4_h_l(net_5804[0:47]),
     .sp4_v_b(net_5807[0:47]), .sp12_v_b(net_6533[0:23]),
     .sp12_h_r(net_5887[0:23]), .sp4_h_r(net_5888[0:47]),
     .sp12_v_t(net_5889[0:23]), .sp4_v_t(net_5779[0:47]),
     .sp4_r_v_b(net_5891[0:47]), .wl(wl[319:304]),
     .top_op(net_7715[0:7]), .rgt_op(net_5931[0:7]),
     .bot_op(net_6407[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_6525), .purst(purst), .slf_op(net_6409[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5903[0:7]),
     .bnl_op(net_5735[0:7]), .tnr_op(net_7749[0:7]),
     .tnl_op(net_7681[0:7]));
ltile4rev I_22_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8223), .lft_op(net_7681[0:7]),
     .sp12_h_l(net_5775[0:23]), .sp4_h_l(net_5776[0:47]),
     .sp4_v_b(net_5779[0:47]), .sp12_v_b(net_5889[0:23]),
     .sp12_h_r(net_5915[0:23]), .sp4_h_r(net_5916[0:47]),
     .sp12_v_t(net_5917[0:23]), .sp4_v_t(net_7743[0:47]),
     .sp4_r_v_b(net_5919[0:47]), .wl(wl[335:320]), .top_op({io_t_22[3],
     io_t_22[2], io_t_22[1], io_t_22[0], io_t_22[3], io_t_22[2],
     io_t_22[1], io_t_22[0]}), .rgt_op(net_7749[0:7]),
     .bot_op(net_6409[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_5881), .purst(purst), .slf_op(net_7715[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5931[0:7]),
     .bnl_op(net_5763[0:7]), .tnr_op({io_t_23[3], io_t_23[2],
     io_t_23[1], io_t_23[0], io_t_23[3], io_t_23[2], io_t_23[1],
     io_t_23[0]}), .tnl_op({io_t_21[3], io_t_21[2], io_t_21[1],
     io_t_21[0], io_t_21[3], io_t_21[2], io_t_21[1], io_t_21[0]}));
ltile4rev I_24_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5937), .lft_op(net_5931[0:7]),
     .sp12_h_l(net_5831[0:23]), .sp4_h_l(net_5832[0:47]),
     .sp4_v_b(net_5835[0:47]), .sp12_v_b(net_6477[0:23]),
     .sp12_h_r(net_5943[0:23]), .sp4_h_r(net_5944[0:47]),
     .sp12_v_t(net_5945[0:23]), .sp4_v_t(net_5975[0:47]),
     .sp4_r_v_b(net_5947[0:47]), .wl(wl[319:304]),
     .top_op(net_7783[0:7]), .rgt_op({io_r_08[3], io_r_08[2],
     io_r_08[1], io_r_08[0], io_r_08[3], io_r_08[2], io_r_08[1],
     io_r_08[0]}), .bot_op(net_5847[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_6469), .purst(purst), .slf_op(net_5987[0:7]),
     .pgate(pgate[319:304]), .bnr_op({io_r_07[3], io_r_07[2],
     io_r_07[1], io_r_07[0], io_r_07[3], io_r_07[2], io_r_07[1],
     io_r_07[0]}), .bnl_op(net_5903[0:7]), .tnr_op({slf_op_25_10[3],
     slf_op_25_10[2], slf_op_25_10[1], slf_op_25_10[0],
     slf_op_25_10[3], slf_op_25_10[2], slf_op_25_10[1],
     slf_op_25_10[0]}), .tnl_op(net_7749[0:7]));
ltile4rev I_23_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8217), .lft_op(net_7715[0:7]),
     .sp12_h_l(net_5915[0:23]), .sp4_h_l(net_5916[0:47]),
     .sp4_v_b(net_5919[0:47]), .sp12_v_b(net_5833[0:23]),
     .sp12_h_r(net_5971[0:23]), .sp4_h_r(net_5972[0:47]),
     .sp12_v_t(net_5973[0:23]), .sp4_v_t(net_7777[0:47]),
     .sp4_r_v_b(net_5975[0:47]), .wl(wl[335:320]), .top_op({io_t_23[3],
     io_t_23[2], io_t_23[1], io_t_23[0], io_t_23[3], io_t_23[2],
     io_t_23[1], io_t_23[0]}), .rgt_op(net_7783[0:7]),
     .bot_op(net_5931[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_5825), .purst(purst), .slf_op(net_7749[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5987[0:7]),
     .bnl_op(net_6409[0:7]), .tnr_op({io_t_24[3], io_t_24[2],
     io_t_24[1], io_t_24[0], io_t_24[3], io_t_24[2], io_t_24[1],
     io_t_24[0]}), .tnl_op({io_t_22[3], io_t_22[2], io_t_22[1],
     io_t_22[0], io_t_22[3], io_t_22[2], io_t_22[1], io_t_22[0]}));
ltile4rev I_13_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_5993), .lft_op(lft_op_13_07[7:0]),
     .sp12_h_l(sp12_h_l_13_07[23:0]), .sp4_h_l(sp4_h_l_13_07[47:0]),
     .sp4_v_b(sp4_v_b_13_07[47:0]), .sp12_v_b(net_5021[0:23]),
     .sp12_h_r(net_5999[0:23]), .sp4_h_r(net_6000[0:47]),
     .sp12_v_t(net_6001[0:23]), .sp4_v_t(sp4_v_b_13_08[47:0]),
     .sp4_r_v_b(net_6003[0:47]), .wl(wl[287:272]),
     .top_op(slf_op_13_08[7:0]), .rgt_op(net_6043[0:7]),
     .bot_op(slf_op_13_06[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5013), .purst(purst), .slf_op(slf_op_13_07[7:0]),
     .pgate(pgate[287:272]), .bnr_op(net_6015[0:7]),
     .bnl_op(lft_op_13_06[7:0]), .tnr_op(net_5679[0:7]),
     .tnl_op(lft_op_13_08[7:0]));
ltile4rev I_13_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6021), .lft_op(lft_op_13_08[7:0]),
     .sp12_h_l(sp12_h_l_13_08[23:0]), .sp4_h_l(sp4_h_l_13_08[47:0]),
     .sp4_v_b(sp4_v_b_13_08[47:0]), .sp12_v_b(net_6001[0:23]),
     .sp12_h_r(net_6027[0:23]), .sp4_h_r(net_6028[0:47]),
     .sp12_v_t(net_6029[0:23]), .sp4_v_t(sp4_v_b_13_09[47:0]),
     .sp4_r_v_b(net_6031[0:47]), .wl(wl[303:288]),
     .top_op(slf_op_13_09[7:0]), .rgt_op(net_5679[0:7]),
     .bot_op(slf_op_13_07[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_5993), .purst(purst), .slf_op(slf_op_13_08[7:0]),
     .pgate(pgate[303:288]), .bnr_op(net_6043[0:7]),
     .bnl_op(lft_op_13_07[7:0]), .tnr_op(net_5651[0:7]),
     .tnl_op(lft_op_13_09[7:0]));
ltile4rev I_14_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6049), .lft_op(slf_op_13_08[7:0]),
     .sp12_h_l(net_6027[0:23]), .sp4_h_l(net_6028[0:47]),
     .sp4_v_b(net_6031[0:47]), .sp12_v_b(net_6085[0:23]),
     .sp12_h_r(net_6055[0:23]), .sp4_h_r(net_6056[0:47]),
     .sp12_v_t(net_6057[0:23]), .sp4_v_t(net_5667[0:47]),
     .sp4_r_v_b(net_6059[0:47]), .wl(wl[303:288]),
     .top_op(net_5651[0:7]), .rgt_op(net_5595[0:7]),
     .bot_op(net_6043[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_6077), .purst(purst), .slf_op(net_5679[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6071[0:7]),
     .bnl_op(slf_op_13_07[7:0]), .tnr_op(net_5623[0:7]),
     .tnl_op(slf_op_13_09[7:0]));
ltile4rev I_14_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6077), .lft_op(slf_op_13_07[7:0]),
     .sp12_h_l(net_5999[0:23]), .sp4_h_l(net_6000[0:47]),
     .sp4_v_b(net_6003[0:47]), .sp12_v_b(net_4993[0:23]),
     .sp12_h_r(net_6083[0:23]), .sp4_h_r(net_6084[0:47]),
     .sp12_v_t(net_6085[0:23]), .sp4_v_t(net_6031[0:47]),
     .sp4_r_v_b(net_6087[0:47]), .wl(wl[287:272]),
     .top_op(net_5679[0:7]), .rgt_op(net_6071[0:7]),
     .bot_op(net_6015[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_4985), .purst(purst), .slf_op(net_6043[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6099[0:7]),
     .bnl_op(slf_op_13_06[7:0]), .tnr_op(net_5595[0:7]),
     .tnl_op(slf_op_13_08[7:0]));
ltile4rev I_17_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6105), .lft_op(net_6211[0:7]),
     .sp12_h_l(net_6251[0:23]), .sp4_h_l(net_6252[0:47]),
     .sp4_v_b(net_6255[0:47]), .sp12_v_b(net_4797[0:23]),
     .sp12_h_r(net_6111[0:23]), .sp4_h_r(net_6112[0:47]),
     .sp12_v_t(net_6113[0:23]), .sp4_v_t(net_6227[0:47]),
     .sp4_r_v_b(net_6115[0:47]), .wl(wl[287:272]),
     .top_op(net_5539[0:7]), .rgt_op(net_6155[0:7]),
     .bot_op(net_6267[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_4789), .purst(purst), .slf_op(net_6239[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6127[0:7]),
     .bnl_op(net_6183[0:7]), .tnr_op(net_5399[0:7]),
     .tnl_op(net_5455[0:7]));
ltile4rev I_17_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6133), .lft_op(net_5455[0:7]),
     .sp12_h_l(net_6223[0:23]), .sp4_h_l(net_6224[0:47]),
     .sp4_v_b(net_6227[0:47]), .sp12_v_b(net_6113[0:23]),
     .sp12_h_r(net_6139[0:23]), .sp4_h_r(net_6140[0:47]),
     .sp12_v_t(net_6141[0:23]), .sp4_v_t(net_5527[0:47]),
     .sp4_r_v_b(net_6143[0:47]), .wl(wl[303:288]),
     .top_op(net_5511[0:7]), .rgt_op(net_5399[0:7]),
     .bot_op(net_6239[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_6105), .purst(purst), .slf_op(net_5539[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6155[0:7]),
     .bnl_op(net_6211[0:7]), .tnr_op(net_5427[0:7]),
     .tnl_op(net_5483[0:7]));
ltile4rev I_15_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6161), .lft_op(net_6043[0:7]),
     .sp12_h_l(net_6083[0:23]), .sp4_h_l(net_6084[0:47]),
     .sp4_v_b(net_6087[0:47]), .sp12_v_b(net_4853[0:23]),
     .sp12_h_r(net_6167[0:23]), .sp4_h_r(net_6168[0:47]),
     .sp12_v_t(net_6169[0:23]), .sp4_v_t(net_6059[0:47]),
     .sp4_r_v_b(net_6171[0:47]), .wl(wl[287:272]),
     .top_op(net_5595[0:7]), .rgt_op(net_6211[0:7]),
     .bot_op(net_6099[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_4845), .purst(purst), .slf_op(net_6071[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6183[0:7]),
     .bnl_op(net_6015[0:7]), .tnr_op(net_5455[0:7]),
     .tnl_op(net_5679[0:7]));
ltile4rev I_15_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6189), .lft_op(net_5679[0:7]),
     .sp12_h_l(net_6055[0:23]), .sp4_h_l(net_6056[0:47]),
     .sp4_v_b(net_6059[0:47]), .sp12_v_b(net_6169[0:23]),
     .sp12_h_r(net_6195[0:23]), .sp4_h_r(net_6196[0:47]),
     .sp12_v_t(net_6197[0:23]), .sp4_v_t(net_5583[0:47]),
     .sp4_r_v_b(net_6199[0:47]), .wl(wl[303:288]),
     .top_op(net_5623[0:7]), .rgt_op(net_5455[0:7]),
     .bot_op(net_6071[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_6161), .purst(purst), .slf_op(net_5595[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6211[0:7]),
     .bnl_op(net_6043[0:7]), .tnr_op(net_5483[0:7]),
     .tnl_op(net_5651[0:7]));
ltile4rev I_16_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6217), .lft_op(net_5595[0:7]),
     .sp12_h_l(net_6195[0:23]), .sp4_h_l(net_6196[0:47]),
     .sp4_v_b(net_6199[0:47]), .sp12_v_b(net_6253[0:23]),
     .sp12_h_r(net_6223[0:23]), .sp4_h_r(net_6224[0:47]),
     .sp12_v_t(net_6225[0:23]), .sp4_v_t(net_5443[0:47]),
     .sp4_r_v_b(net_6227[0:47]), .wl(wl[303:288]),
     .top_op(net_5483[0:7]), .rgt_op(net_5539[0:7]),
     .bot_op(net_6211[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_6245), .purst(purst), .slf_op(net_5455[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6239[0:7]),
     .bnl_op(net_6071[0:7]), .tnr_op(net_5511[0:7]),
     .tnl_op(net_5623[0:7]));
ltile4rev I_16_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6245), .lft_op(net_6071[0:7]),
     .sp12_h_l(net_6167[0:23]), .sp4_h_l(net_6168[0:47]),
     .sp4_v_b(net_6171[0:47]), .sp12_v_b(net_4881[0:23]),
     .sp12_h_r(net_6251[0:23]), .sp4_h_r(net_6252[0:47]),
     .sp12_v_t(net_6253[0:23]), .sp4_v_t(net_6199[0:47]),
     .sp4_r_v_b(net_6255[0:47]), .wl(wl[287:272]),
     .top_op(net_5455[0:7]), .rgt_op(net_6239[0:7]),
     .bot_op(net_6183[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_4873), .purst(purst), .slf_op(net_6211[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6267[0:7]),
     .bnl_op(net_6099[0:7]), .tnr_op(net_5539[0:7]),
     .tnl_op(net_5595[0:7]));
ltile4rev I_18_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6273), .lft_op(net_5539[0:7]),
     .sp12_h_l(net_6139[0:23]), .sp4_h_l(net_6140[0:47]),
     .sp4_v_b(net_6143[0:47]), .sp12_v_b(net_6309[0:23]),
     .sp12_h_r(net_6279[0:23]), .sp4_h_r(net_6280[0:47]),
     .sp12_v_t(net_6281[0:23]), .sp4_v_t(net_5387[0:47]),
     .sp4_r_v_b(net_6283[0:47]), .wl(wl[303:288]),
     .top_op(net_5427[0:7]), .rgt_op(net_5707[0:7]),
     .bot_op(net_6155[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_6301), .purst(purst), .slf_op(net_5399[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_4138[0:7]),
     .bnl_op(net_6239[0:7]), .tnr_op(net_6297[0:7]),
     .tnl_op(net_5511[0:7]));
ltile4rev I_18_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6301), .lft_op(net_6239[0:7]),
     .sp12_h_l(net_6111[0:23]), .sp4_h_l(net_6112[0:47]),
     .sp4_v_b(net_6115[0:47]), .sp12_v_b(net_4937[0:23]),
     .sp12_h_r(net_6307[0:23]), .sp4_h_r(net_6308[0:47]),
     .sp12_v_t(net_6309[0:23]), .sp4_v_t(net_6143[0:47]),
     .sp4_r_v_b(net_6311[0:47]), .wl(wl[287:272]),
     .top_op(net_5399[0:7]), .rgt_op(net_4138[0:7]),
     .bot_op(net_6127[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_4929), .purst(purst), .slf_op(net_6155[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6323[0:7]),
     .bnl_op(net_6267[0:7]), .tnr_op(net_5707[0:7]),
     .tnl_op(net_5539[0:7]));
ltile4rev I_20_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6329), .lft_op(net_4138[0:7]),
     .sp12_h_l(net_4116[0:23]), .sp4_h_l(net_4117[0:47]),
     .sp4_v_b(net_4121[0:47]), .sp12_v_b(net_5133[0:23]),
     .sp12_h_r(net_6335[0:23]), .sp4_h_r(net_6336[0:47]),
     .sp12_v_t(net_6337[0:23]), .sp4_v_t(net_4120[0:47]),
     .sp4_r_v_b(net_6339[0:47]), .wl(wl[287:272]),
     .top_op(net_4031[0:7]), .rgt_op(net_6379[0:7]),
     .bot_op(net_4122[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_5125), .purst(purst), .slf_op(net_5137[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6351[0:7]),
     .bnl_op(net_6323[0:7]), .tnr_op(net_5735[0:7]),
     .tnl_op(net_5707[0:7]));
ltile4rev I_20_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6357), .lft_op(net_5707[0:7]),
     .sp12_h_l(net_4115[0:23]), .sp4_h_l(net_4118[0:47]),
     .sp4_v_b(net_4120[0:47]), .sp12_v_b(net_6337[0:23]),
     .sp12_h_r(net_6363[0:23]), .sp4_h_r(net_6364[0:47]),
     .sp12_v_t(net_6365[0:23]), .sp4_v_t(net_4045[0:47]),
     .sp4_r_v_b(net_6367[0:47]), .wl(wl[303:288]),
     .top_op(net_4113[0:7]), .rgt_op(net_5735[0:7]),
     .bot_op(net_5137[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_6329), .purst(purst), .slf_op(net_4031[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6379[0:7]),
     .bnl_op(net_4138[0:7]), .tnr_op(net_5763[0:7]),
     .tnl_op(net_6297[0:7]));
ltile4rev I_21_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6385), .lft_op(net_4031[0:7]),
     .sp12_h_l(net_6363[0:23]), .sp4_h_l(net_6364[0:47]),
     .sp4_v_b(net_6367[0:47]), .sp12_v_b(net_6421[0:23]),
     .sp12_h_r(net_6391[0:23]), .sp4_h_r(net_6392[0:47]),
     .sp12_v_t(net_6393[0:23]), .sp4_v_t(net_5723[0:47]),
     .sp4_r_v_b(net_6395[0:47]), .wl(wl[303:288]),
     .top_op(net_5763[0:7]), .rgt_op(net_6407[0:7]),
     .bot_op(net_6379[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_6413), .purst(purst), .slf_op(net_5735[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_5177[0:7]),
     .bnl_op(net_5137[0:7]), .tnr_op(net_6409[0:7]),
     .tnl_op(net_4113[0:7]));
ltile4rev I_21_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6413), .lft_op(net_5137[0:7]),
     .sp12_h_l(net_6335[0:23]), .sp4_h_l(net_6336[0:47]),
     .sp4_v_b(net_6339[0:47]), .sp12_v_b(net_5161[0:23]),
     .sp12_h_r(net_6419[0:23]), .sp4_h_r(net_6420[0:47]),
     .sp12_v_t(net_6421[0:23]), .sp4_v_t(net_6367[0:47]),
     .sp4_r_v_b(net_6423[0:47]), .wl(wl[287:272]),
     .top_op(net_5735[0:7]), .rgt_op(net_5177[0:7]),
     .bot_op(net_6351[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_5153), .purst(purst), .slf_op(net_6379[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6435[0:7]),
     .bnl_op(net_4122[0:7]), .tnr_op(net_6407[0:7]),
     .tnl_op(net_4031[0:7]));
ltile4rev I_23_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6441), .lft_op(net_5177[0:7]),
     .sp12_h_l(net_6503[0:23]), .sp4_h_l(net_6504[0:47]),
     .sp4_v_b(net_6507[0:47]), .sp12_v_b(net_5357[0:23]),
     .sp12_h_r(net_6447[0:23]), .sp4_h_r(net_6448[0:47]),
     .sp12_v_t(net_6449[0:23]), .sp4_v_t(net_6535[0:47]),
     .sp4_r_v_b(net_6451[0:47]), .wl(wl[287:272]),
     .top_op(net_5903[0:7]), .rgt_op(net_6603[0:7]),
     .bot_op(net_6519[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_5349), .purst(purst), .slf_op(net_6547[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6463[0:7]),
     .bnl_op(net_6435[0:7]), .tnr_op(net_5847[0:7]),
     .tnl_op(net_6407[0:7]));
ltile4rev I_24_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6469), .lft_op(net_5903[0:7]),
     .sp12_h_l(net_6587[0:23]), .sp4_h_l(net_6588[0:47]),
     .sp4_v_b(net_6591[0:47]), .sp12_v_b(net_6561[0:23]),
     .sp12_h_r(net_6475[0:23]), .sp4_h_r(net_6476[0:47]),
     .sp12_v_t(net_6477[0:23]), .sp4_v_t(net_5835[0:47]),
     .sp4_r_v_b(net_6479[0:47]), .wl(wl[303:288]),
     .top_op(net_5987[0:7]), .rgt_op({io_r_07[3], io_r_07[2],
     io_r_07[1], io_r_07[0], io_r_07[3], io_r_07[2], io_r_07[1],
     io_r_07[0]}), .bot_op(net_6603[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_6553), .purst(purst), .slf_op(net_5847[0:7]),
     .pgate(pgate[303:288]), .bnr_op({io_r_06[3], io_r_06[2],
     io_r_06[1], io_r_06[0], io_r_06[3], io_r_06[2], io_r_06[1],
     io_r_06[0]}), .bnl_op(net_6547[0:7]), .tnr_op({io_r_08[3],
     io_r_08[2], io_r_08[1], io_r_08[0], io_r_08[3], io_r_08[2],
     io_r_08[1], io_r_08[0]}), .tnl_op(net_5931[0:7]));
ltile4rev I_22_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6497), .lft_op(net_6379[0:7]),
     .sp12_h_l(net_6419[0:23]), .sp4_h_l(net_6420[0:47]),
     .sp4_v_b(net_6423[0:47]), .sp12_v_b(net_5301[0:23]),
     .sp12_h_r(net_6503[0:23]), .sp4_h_r(net_6504[0:47]),
     .sp12_v_t(net_6505[0:23]), .sp4_v_t(net_6395[0:47]),
     .sp4_r_v_b(net_6507[0:47]), .wl(wl[287:272]),
     .top_op(net_6407[0:7]), .rgt_op(net_6547[0:7]),
     .bot_op(net_6435[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_5293), .purst(purst), .slf_op(net_5177[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6519[0:7]),
     .bnl_op(net_6351[0:7]), .tnr_op(net_5903[0:7]),
     .tnl_op(net_5735[0:7]));
ltile4rev I_22_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6525), .lft_op(net_5735[0:7]),
     .sp12_h_l(net_6391[0:23]), .sp4_h_l(net_6392[0:47]),
     .sp4_v_b(net_6395[0:47]), .sp12_v_b(net_6505[0:23]),
     .sp12_h_r(net_6531[0:23]), .sp4_h_r(net_6532[0:47]),
     .sp12_v_t(net_6533[0:23]), .sp4_v_t(net_5807[0:47]),
     .sp4_r_v_b(net_6535[0:47]), .wl(wl[303:288]),
     .top_op(net_6409[0:7]), .rgt_op(net_5903[0:7]),
     .bot_op(net_5177[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_6497), .purst(purst), .slf_op(net_6407[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6547[0:7]),
     .bnl_op(net_6379[0:7]), .tnr_op(net_5931[0:7]),
     .tnl_op(net_5763[0:7]));
ltile4rev I_24_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6553), .lft_op(net_6547[0:7]),
     .sp12_h_l(net_6447[0:23]), .sp4_h_l(net_6448[0:47]),
     .sp4_v_b(net_6451[0:47]), .sp12_v_b(net_5245[0:23]),
     .sp12_h_r(net_6559[0:23]), .sp4_h_r(net_6560[0:47]),
     .sp12_v_t(net_6561[0:23]), .sp4_v_t(net_6591[0:47]),
     .sp4_r_v_b(net_6563[0:47]), .wl(wl[287:272]),
     .top_op(net_5847[0:7]), .rgt_op({io_r_06[3], io_r_06[2],
     io_r_06[1], io_r_06[0], io_r_06[3], io_r_06[2], io_r_06[1],
     io_r_06[0]}), .bot_op(net_6463[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_5237), .purst(purst), .slf_op(net_6603[0:7]),
     .pgate(pgate[287:272]), .bnr_op({io_r_05[3], io_r_05[2],
     io_r_05[1], io_r_05[0], io_r_05[3], io_r_05[2], io_r_05[1],
     io_r_05[0]}), .bnl_op(net_6519[0:7]), .tnr_op({io_r_07[3],
     io_r_07[2], io_r_07[1], io_r_07[0], io_r_07[3], io_r_07[2],
     io_r_07[1], io_r_07[0]}), .tnl_op(net_5903[0:7]));
ltile4rev I_23_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6581), .lft_op(net_6407[0:7]),
     .sp12_h_l(net_6531[0:23]), .sp4_h_l(net_6532[0:47]),
     .sp4_v_b(net_6535[0:47]), .sp12_v_b(net_6449[0:23]),
     .sp12_h_r(net_6587[0:23]), .sp4_h_r(net_6588[0:47]),
     .sp12_v_t(net_6589[0:23]), .sp4_v_t(net_5891[0:47]),
     .sp4_r_v_b(net_6591[0:47]), .wl(wl[303:288]),
     .top_op(net_5931[0:7]), .rgt_op(net_5847[0:7]),
     .bot_op(net_6547[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_6441), .purst(purst), .slf_op(net_5903[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6603[0:7]),
     .bnl_op(net_5177[0:7]), .tnr_op(net_5987[0:7]),
     .tnl_op(net_6409[0:7]));
ltile4rev I_23_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_6609), .lft_op(slf_op_22_11[7:0]),
     .sp12_h_l(net_6671[0:23]), .sp4_h_l(net_6672[0:47]),
     .sp4_v_b(sp4_v_b_23_11[47:0]), .sp12_v_b(sp12_v_b_23_11[23:0]),
     .sp12_h_r(net_6615[0:23]), .sp4_h_r(net_6616[0:47]),
     .sp12_v_t(net_6617[0:23]), .sp4_v_t(net_6703[0:47]),
     .sp4_r_v_b(sp4_v_b_24_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7303[0:7]), .rgt_op(slf_op_24_11[7:0]),
     .bot_op(bot_op_23_11[7:0]), .bl(bl[1239:1186]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(carry_in_23_11), .purst(purst),
     .slf_op(slf_op_23_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_23_11[7:0]), .bnl_op(bnl_op_23_11[7:0]),
     .tnr_op(net_7247[0:7]), .tnl_op(net_7219[0:7]));
ltile4rev I_24_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_6637), .lft_op(net_7303[0:7]),
     .sp12_h_l(net_6755[0:23]), .sp4_h_l(net_6756[0:47]),
     .sp4_v_b(net_6759[0:47]), .sp12_v_b(net_6729[0:23]),
     .sp12_h_r(net_6643[0:23]), .sp4_h_r(net_6644[0:47]),
     .sp12_v_t(net_6645[0:23]), .sp4_v_t(net_7235[0:47]),
     .sp4_r_v_b(net_6647[0:47]), .wl(wl[207:192]),
     .top_op(net_7387[0:7]), .rgt_op({io_r_01[3], io_r_01[2],
     io_r_01[1], io_r_01[0], io_r_01[3], io_r_01[2], io_r_01[1],
     io_r_01[0]}), .bot_op(slf_op_24_11[7:0]), .bl(bl[1293:1240]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_6721), .purst(purst), .slf_op(net_7247[0:7]),
     .pgate(pgate[207:192]), .bnr_op({io_r_00_24_11[3],
     io_r_00_24_11[2], io_r_00_24_11[1], io_r_00_24_11[0],
     io_r_00_24_11[3], io_r_00_24_11[2], io_r_00_24_11[1],
     io_r_00_24_11[0]}), .bnl_op(slf_op_23_11[7:0]),
     .tnr_op({io_r_02[3], io_r_02[2], io_r_02[1], io_r_02[0],
     io_r_02[3], io_r_02[2], io_r_02[1], io_r_02[0]}),
     .tnl_op(net_7331[0:7]));
ltile4rev I_22_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_6665), .lft_op(slf_op_21_11[7:0]),
     .sp12_h_l(net_4739[0:23]), .sp4_h_l(net_4740[0:47]),
     .sp4_v_b(sp4_v_b_22_11[47:0]), .sp12_v_b(sp12_v_b_22_11[23:0]),
     .sp12_h_r(net_6671[0:23]), .sp4_h_r(net_6672[0:47]),
     .sp12_v_t(net_6673[0:23]), .sp4_v_t(net_4715[0:47]),
     .sp4_r_v_b(sp4_v_b_23_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7219[0:7]), .rgt_op(slf_op_23_11[7:0]),
     .bot_op(bot_op_22_11[7:0]), .bl(bl[1185:1132]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(carry_in_22_11), .purst(purst),
     .slf_op(slf_op_22_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_22_11[7:0]), .bnl_op(bnl_op_22_11[7:0]),
     .tnr_op(net_7303[0:7]), .tnl_op(net_7135[0:7]));
ltile4rev I_22_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_6693), .lft_op(net_7135[0:7]),
     .sp12_h_l(net_4711[0:23]), .sp4_h_l(net_4712[0:47]),
     .sp4_v_b(net_4715[0:47]), .sp12_v_b(net_6673[0:23]),
     .sp12_h_r(net_6699[0:23]), .sp4_h_r(net_6700[0:47]),
     .sp12_v_t(net_6701[0:23]), .sp4_v_t(net_7207[0:47]),
     .sp4_r_v_b(net_6703[0:47]), .wl(wl[207:192]),
     .top_op(net_4729[0:7]), .rgt_op(net_7303[0:7]),
     .bot_op(slf_op_22_11[7:0]), .bl(bl[1185:1132]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_6665), .purst(purst), .slf_op(net_7219[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_23_11[7:0]),
     .bnl_op(slf_op_21_11[7:0]), .tnr_op(net_7331[0:7]),
     .tnl_op(net_7163[0:7]));
ltile4rev I_24_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_6721), .lft_op(slf_op_23_11[7:0]),
     .sp12_h_l(net_6615[0:23]), .sp4_h_l(net_6616[0:47]),
     .sp4_v_b(sp4_v_b_24_11[47:0]), .sp12_v_b(sp12_v_b_24_11[23:0]),
     .sp12_h_r(net_6727[0:23]), .sp4_h_r(net_6728[0:47]),
     .sp12_v_t(net_6729[0:23]), .sp4_v_t(net_6759[0:47]),
     .sp4_r_v_b(net_6731[0:47]), .wl(wl[191:176]),
     .top_op(net_7247[0:7]), .rgt_op({io_r_00_24_11[3],
     io_r_00_24_11[2], io_r_00_24_11[1], io_r_00_24_11[0],
     io_r_00_24_11[3], io_r_00_24_11[2], io_r_00_24_11[1],
     io_r_00_24_11[0]}), .bot_op(bot_op_24_11[7:0]),
     .bl(bl[1293:1240]), .reset_b(reset_b[191:176]),
     .glb_netwk(glb_netwk_24[7:0]), .carry_in(carry_in_24_11),
     .purst(purst), .slf_op(slf_op_24_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_24_11[7:0]), .bnl_op(bnl_op_24_11[7:0]),
     .tnr_op({io_r_01[3], io_r_01[2], io_r_01[1], io_r_01[0],
     io_r_01[3], io_r_01[2], io_r_01[1], io_r_01[0]}),
     .tnl_op(net_7303[0:7]));
ltile4rev I_23_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_6749), .lft_op(net_7219[0:7]),
     .sp12_h_l(net_6699[0:23]), .sp4_h_l(net_6700[0:47]),
     .sp4_v_b(net_6703[0:47]), .sp12_v_b(net_6617[0:23]),
     .sp12_h_r(net_6755[0:23]), .sp4_h_r(net_6756[0:47]),
     .sp12_v_t(net_6757[0:23]), .sp4_v_t(net_7291[0:47]),
     .sp4_r_v_b(net_6759[0:47]), .wl(wl[207:192]),
     .top_op(net_7331[0:7]), .rgt_op(net_7247[0:7]),
     .bot_op(slf_op_23_11[7:0]), .bl(bl[1239:1186]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_6609), .purst(purst), .slf_op(net_7303[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_24_11[7:0]),
     .bnl_op(slf_op_22_11[7:0]), .tnr_op(net_7387[0:7]),
     .tnl_op(net_4729[0:7]));
ltile4rev I_13_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_6777), .lft_op(lft_op_13_03[7:0]),
     .sp12_h_l(sp12_h_l_13_03[23:0]), .sp4_h_l(sp4_h_l_13_03[47:0]),
     .sp4_v_b(sp4_v_b_13_03[47:0]), .sp12_v_b(net_4573[0:23]),
     .sp12_h_r(net_6783[0:23]), .sp4_h_r(net_6784[0:47]),
     .sp12_v_t(net_6785[0:23]), .sp4_v_t(sp4_v_b_13_04[47:0]),
     .sp4_r_v_b(net_6787[0:47]), .wl(wl[223:208]),
     .top_op(slf_op_13_04[7:0]), .rgt_op(net_6827[0:7]),
     .bot_op(slf_op_13_02[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_4565), .purst(purst), .slf_op(slf_op_13_03[7:0]),
     .pgate(pgate[223:208]), .bnr_op(net_6799[0:7]),
     .bnl_op(lft_op_13_02[7:0]), .tnr_op(net_5063[0:7]),
     .tnl_op(lft_op_13_04[7:0]));
ltile4rev I_13_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_6805), .lft_op(lft_op_13_04[7:0]),
     .sp12_h_l(sp12_h_l_13_04[23:0]), .sp4_h_l(sp4_h_l_13_04[47:0]),
     .sp4_v_b(sp4_v_b_13_04[47:0]), .sp12_v_b(net_6785[0:23]),
     .sp12_h_r(net_6811[0:23]), .sp4_h_r(net_6812[0:47]),
     .sp12_v_t(net_6813[0:23]), .sp4_v_t(sp4_v_b_13_05[47:0]),
     .sp4_r_v_b(net_6815[0:47]), .wl(wl[239:224]),
     .top_op(slf_op_13_05[7:0]), .rgt_op(net_5063[0:7]),
     .bot_op(slf_op_13_03[7:0]), .bl(bl[711:658]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_13[7:0]),
     .carry_in(net_6777), .purst(purst), .slf_op(slf_op_13_04[7:0]),
     .pgate(pgate[239:224]), .bnr_op(net_6827[0:7]),
     .bnl_op(lft_op_13_03[7:0]), .tnr_op(net_5035[0:7]),
     .tnl_op(lft_op_13_05[7:0]));
ltile4rev I_14_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_6833), .lft_op(slf_op_13_04[7:0]),
     .sp12_h_l(net_6811[0:23]), .sp4_h_l(net_6812[0:47]),
     .sp4_v_b(net_6815[0:47]), .sp12_v_b(net_6869[0:23]),
     .sp12_h_r(net_6839[0:23]), .sp4_h_r(net_6840[0:47]),
     .sp12_v_t(net_6841[0:23]), .sp4_v_t(net_5051[0:47]),
     .sp4_r_v_b(net_6843[0:47]), .wl(wl[239:224]),
     .top_op(net_5035[0:7]), .rgt_op(net_4979[0:7]),
     .bot_op(net_6827[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_6861), .purst(purst), .slf_op(net_5063[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_6855[0:7]),
     .bnl_op(slf_op_13_03[7:0]), .tnr_op(net_5007[0:7]),
     .tnl_op(slf_op_13_05[7:0]));
ltile4rev I_14_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_6861), .lft_op(slf_op_13_03[7:0]),
     .sp12_h_l(net_6783[0:23]), .sp4_h_l(net_6784[0:47]),
     .sp4_v_b(net_6787[0:47]), .sp12_v_b(net_4545[0:23]),
     .sp12_h_r(net_6867[0:23]), .sp4_h_r(net_6868[0:47]),
     .sp12_v_t(net_6869[0:23]), .sp4_v_t(net_6815[0:47]),
     .sp4_r_v_b(net_6871[0:47]), .wl(wl[223:208]),
     .top_op(net_5063[0:7]), .rgt_op(net_6855[0:7]),
     .bot_op(net_6799[0:7]), .bl(bl[765:712]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_14[7:0]),
     .carry_in(net_4537), .purst(purst), .slf_op(net_6827[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_6883[0:7]),
     .bnl_op(slf_op_13_02[7:0]), .tnr_op(net_4979[0:7]),
     .tnl_op(slf_op_13_04[7:0]));
ltile4rev I_17_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_6889), .lft_op(net_6995[0:7]),
     .sp12_h_l(net_7035[0:23]), .sp4_h_l(net_7036[0:47]),
     .sp4_v_b(net_7039[0:47]), .sp12_v_b(net_4349[0:23]),
     .sp12_h_r(net_6895[0:23]), .sp4_h_r(net_6896[0:47]),
     .sp12_v_t(net_6897[0:23]), .sp4_v_t(net_7011[0:47]),
     .sp4_r_v_b(net_6899[0:47]), .wl(wl[223:208]),
     .top_op(net_4923[0:7]), .rgt_op(net_6939[0:7]),
     .bot_op(net_7051[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_4341), .purst(purst), .slf_op(net_7023[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_6911[0:7]),
     .bnl_op(net_6967[0:7]), .tnr_op(net_4783[0:7]),
     .tnl_op(net_4839[0:7]));
ltile4rev I_17_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_6917), .lft_op(net_4839[0:7]),
     .sp12_h_l(net_7007[0:23]), .sp4_h_l(net_7008[0:47]),
     .sp4_v_b(net_7011[0:47]), .sp12_v_b(net_6897[0:23]),
     .sp12_h_r(net_6923[0:23]), .sp4_h_r(net_6924[0:47]),
     .sp12_v_t(net_6925[0:23]), .sp4_v_t(net_4911[0:47]),
     .sp4_r_v_b(net_6927[0:47]), .wl(wl[239:224]),
     .top_op(net_4895[0:7]), .rgt_op(net_4783[0:7]),
     .bot_op(net_7023[0:7]), .bl(bl[927:874]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_17[7:0]),
     .carry_in(net_6889), .purst(purst), .slf_op(net_4923[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_6939[0:7]),
     .bnl_op(net_6995[0:7]), .tnr_op(net_4811[0:7]),
     .tnl_op(net_4867[0:7]));
ltile4rev I_15_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_6945), .lft_op(net_6827[0:7]),
     .sp12_h_l(net_6867[0:23]), .sp4_h_l(net_6868[0:47]),
     .sp4_v_b(net_6871[0:47]), .sp12_v_b(net_4405[0:23]),
     .sp12_h_r(net_6951[0:23]), .sp4_h_r(net_6952[0:47]),
     .sp12_v_t(net_6953[0:23]), .sp4_v_t(net_6843[0:47]),
     .sp4_r_v_b(net_6955[0:47]), .wl(wl[223:208]),
     .top_op(net_4979[0:7]), .rgt_op(net_6995[0:7]),
     .bot_op(net_6883[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_4397), .purst(purst), .slf_op(net_6855[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_6967[0:7]),
     .bnl_op(net_6799[0:7]), .tnr_op(net_4839[0:7]),
     .tnl_op(net_5063[0:7]));
ltile4rev I_15_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_6973), .lft_op(net_5063[0:7]),
     .sp12_h_l(net_6839[0:23]), .sp4_h_l(net_6840[0:47]),
     .sp4_v_b(net_6843[0:47]), .sp12_v_b(net_6953[0:23]),
     .sp12_h_r(net_6979[0:23]), .sp4_h_r(net_6980[0:47]),
     .sp12_v_t(net_6981[0:23]), .sp4_v_t(net_4967[0:47]),
     .sp4_r_v_b(net_6983[0:47]), .wl(wl[239:224]),
     .top_op(net_5007[0:7]), .rgt_op(net_4839[0:7]),
     .bot_op(net_6855[0:7]), .bl(bl[819:766]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_15[7:0]),
     .carry_in(net_6945), .purst(purst), .slf_op(net_4979[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_6995[0:7]),
     .bnl_op(net_6827[0:7]), .tnr_op(net_4867[0:7]),
     .tnl_op(net_5035[0:7]));
ltile4rev I_16_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7001), .lft_op(net_4979[0:7]),
     .sp12_h_l(net_6979[0:23]), .sp4_h_l(net_6980[0:47]),
     .sp4_v_b(net_6983[0:47]), .sp12_v_b(net_7037[0:23]),
     .sp12_h_r(net_7007[0:23]), .sp4_h_r(net_7008[0:47]),
     .sp12_v_t(net_7009[0:23]), .sp4_v_t(net_4827[0:47]),
     .sp4_r_v_b(net_7011[0:47]), .wl(wl[239:224]),
     .top_op(net_4867[0:7]), .rgt_op(net_4923[0:7]),
     .bot_op(net_6995[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_7029), .purst(purst), .slf_op(net_4839[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7023[0:7]),
     .bnl_op(net_6855[0:7]), .tnr_op(net_4895[0:7]),
     .tnl_op(net_5007[0:7]));
ltile4rev I_16_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7029), .lft_op(net_6855[0:7]),
     .sp12_h_l(net_6951[0:23]), .sp4_h_l(net_6952[0:47]),
     .sp4_v_b(net_6955[0:47]), .sp12_v_b(net_4433[0:23]),
     .sp12_h_r(net_7035[0:23]), .sp4_h_r(net_7036[0:47]),
     .sp12_v_t(net_7037[0:23]), .sp4_v_t(net_6983[0:47]),
     .sp4_r_v_b(net_7039[0:47]), .wl(wl[223:208]),
     .top_op(net_4839[0:7]), .rgt_op(net_7023[0:7]),
     .bot_op(net_6967[0:7]), .bl(bl[873:820]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_16[7:0]),
     .carry_in(net_4425), .purst(purst), .slf_op(net_6995[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7051[0:7]),
     .bnl_op(net_6883[0:7]), .tnr_op(net_4923[0:7]),
     .tnl_op(net_4979[0:7]));
ltile4rev I_18_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7057), .lft_op(net_4923[0:7]),
     .sp12_h_l(net_6923[0:23]), .sp4_h_l(net_6924[0:47]),
     .sp4_v_b(net_6927[0:47]), .sp12_v_b(net_7093[0:23]),
     .sp12_h_r(net_7063[0:23]), .sp4_h_r(net_7064[0:47]),
     .sp12_v_t(net_7065[0:23]), .sp4_v_t(net_4771[0:47]),
     .sp4_r_v_b(net_7067[0:47]), .wl(wl[239:224]),
     .top_op(net_4811[0:7]), .rgt_op(net_5091[0:7]),
     .bot_op(net_6939[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_7085), .purst(purst), .slf_op(net_4783[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_4262[0:7]),
     .bnl_op(net_7023[0:7]), .tnr_op(net_7081[0:7]),
     .tnl_op(net_4895[0:7]));
ltile4rev I_18_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7085), .lft_op(net_7023[0:7]),
     .sp12_h_l(net_6895[0:23]), .sp4_h_l(net_6896[0:47]),
     .sp4_v_b(net_6899[0:47]), .sp12_v_b(net_4489[0:23]),
     .sp12_h_r(net_7091[0:23]), .sp4_h_r(net_7092[0:47]),
     .sp12_v_t(net_7093[0:23]), .sp4_v_t(net_6927[0:47]),
     .sp4_r_v_b(net_7095[0:47]), .wl(wl[223:208]),
     .top_op(net_4783[0:7]), .rgt_op(net_4262[0:7]),
     .bot_op(net_6911[0:7]), .bl(bl[981:928]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_18[7:0]),
     .carry_in(net_4481), .purst(purst), .slf_op(net_6939[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_4645[0:7]),
     .bnl_op(net_7051[0:7]), .tnr_op(net_5091[0:7]),
     .tnl_op(net_4923[0:7]));
ltile4rev I_20_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7113), .lft_op(net_4262[0:7]),
     .sp12_h_l(net_4201[0:23]), .sp4_h_l(net_4202[0:47]),
     .sp4_v_b(net_4206[0:47]), .sp12_v_b(net_4685[0:23]),
     .sp12_h_r(net_7119[0:23]), .sp4_h_r(net_7120[0:47]),
     .sp12_v_t(net_7121[0:23]), .sp4_v_t(net_4205[0:47]),
     .sp4_r_v_b(net_7123[0:47]), .wl(wl[223:208]),
     .top_op(net_4155[0:7]), .rgt_op(net_7163[0:7]),
     .bot_op(net_4207[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_4677), .purst(purst), .slf_op(net_4689[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7135[0:7]),
     .bnl_op(net_4645[0:7]), .tnr_op(net_5119[0:7]),
     .tnl_op(net_5091[0:7]));
ltile4rev I_20_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7141), .lft_op(net_5091[0:7]),
     .sp12_h_l(net_4200[0:23]), .sp4_h_l(net_4203[0:47]),
     .sp4_v_b(net_4205[0:47]), .sp12_v_b(net_7121[0:23]),
     .sp12_h_r(net_7147[0:23]), .sp4_h_r(net_7148[0:47]),
     .sp12_v_t(net_7149[0:23]), .sp4_v_t(net_4169[0:47]),
     .sp4_r_v_b(net_7151[0:47]), .wl(wl[239:224]),
     .top_op(net_4198[0:7]), .rgt_op(net_5119[0:7]),
     .bot_op(net_4689[0:7]), .bl(bl[1077:1024]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_20[7:0]),
     .carry_in(net_7113), .purst(purst), .slf_op(net_4155[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7163[0:7]),
     .bnl_op(net_4262[0:7]), .tnr_op(net_5147[0:7]),
     .tnl_op(net_7081[0:7]));
ltile4rev I_21_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7169), .lft_op(net_4155[0:7]),
     .sp12_h_l(net_7147[0:23]), .sp4_h_l(net_7148[0:47]),
     .sp4_v_b(net_7151[0:47]), .sp12_v_b(net_7205[0:23]),
     .sp12_h_r(net_7175[0:23]), .sp4_h_r(net_7176[0:47]),
     .sp12_v_t(net_7177[0:23]), .sp4_v_t(net_5107[0:47]),
     .sp4_r_v_b(net_7179[0:47]), .wl(wl[239:224]),
     .top_op(net_5147[0:7]), .rgt_op(net_7191[0:7]),
     .bot_op(net_7163[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_7197), .purst(purst), .slf_op(net_5119[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_4729[0:7]),
     .bnl_op(net_4689[0:7]), .tnr_op(net_7193[0:7]),
     .tnl_op(net_4198[0:7]));
ltile4rev I_21_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7197), .lft_op(net_4689[0:7]),
     .sp12_h_l(net_7119[0:23]), .sp4_h_l(net_7120[0:47]),
     .sp4_v_b(net_7123[0:47]), .sp12_v_b(net_4713[0:23]),
     .sp12_h_r(net_7203[0:23]), .sp4_h_r(net_7204[0:47]),
     .sp12_v_t(net_7205[0:23]), .sp4_v_t(net_7151[0:47]),
     .sp4_r_v_b(net_7207[0:47]), .wl(wl[223:208]),
     .top_op(net_5119[0:7]), .rgt_op(net_4729[0:7]),
     .bot_op(net_7135[0:7]), .bl(bl[1131:1078]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_21[7:0]),
     .carry_in(net_4705), .purst(purst), .slf_op(net_7163[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7219[0:7]),
     .bnl_op(net_4207[0:7]), .tnr_op(net_7191[0:7]),
     .tnl_op(net_4155[0:7]));
ltile4rev I_23_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7225), .lft_op(net_4729[0:7]),
     .sp12_h_l(net_7287[0:23]), .sp4_h_l(net_7288[0:47]),
     .sp4_v_b(net_7291[0:47]), .sp12_v_b(net_6757[0:23]),
     .sp12_h_r(net_7231[0:23]), .sp4_h_r(net_7232[0:47]),
     .sp12_v_t(net_7233[0:23]), .sp4_v_t(net_7319[0:47]),
     .sp4_r_v_b(net_7235[0:47]), .wl(wl[223:208]),
     .top_op(net_5287[0:7]), .rgt_op(net_7387[0:7]),
     .bot_op(net_7303[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_6749), .purst(purst), .slf_op(net_7331[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7247[0:7]),
     .bnl_op(net_7219[0:7]), .tnr_op(net_5231[0:7]),
     .tnl_op(net_7191[0:7]));
ltile4rev I_24_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7253), .lft_op(net_5287[0:7]),
     .sp12_h_l(net_7371[0:23]), .sp4_h_l(net_7372[0:47]),
     .sp4_v_b(net_7375[0:47]), .sp12_v_b(net_7345[0:23]),
     .sp12_h_r(net_7259[0:23]), .sp4_h_r(net_7260[0:47]),
     .sp12_v_t(net_7261[0:23]), .sp4_v_t(net_5219[0:47]),
     .sp4_r_v_b(net_7263[0:47]), .wl(wl[239:224]),
     .top_op(net_5371[0:7]), .rgt_op({io_r_03[3], io_r_03[2],
     io_r_03[1], io_r_03[0], io_r_03[3], io_r_03[2], io_r_03[1],
     io_r_03[0]}), .bot_op(net_7387[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_7337), .purst(purst), .slf_op(net_5231[0:7]),
     .pgate(pgate[239:224]), .bnr_op({io_r_02[3], io_r_02[2],
     io_r_02[1], io_r_02[0], io_r_02[3], io_r_02[2], io_r_02[1],
     io_r_02[0]}), .bnl_op(net_7331[0:7]), .tnr_op({io_r_04[3],
     io_r_04[2], io_r_04[1], io_r_04[0], io_r_04[3], io_r_04[2],
     io_r_04[1], io_r_04[0]}), .tnl_op(net_5315[0:7]));
ltile4rev I_22_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7281), .lft_op(net_7163[0:7]),
     .sp12_h_l(net_7203[0:23]), .sp4_h_l(net_7204[0:47]),
     .sp4_v_b(net_7207[0:47]), .sp12_v_b(net_6701[0:23]),
     .sp12_h_r(net_7287[0:23]), .sp4_h_r(net_7288[0:47]),
     .sp12_v_t(net_7289[0:23]), .sp4_v_t(net_7179[0:47]),
     .sp4_r_v_b(net_7291[0:47]), .wl(wl[223:208]),
     .top_op(net_7191[0:7]), .rgt_op(net_7331[0:7]),
     .bot_op(net_7219[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_6693), .purst(purst), .slf_op(net_4729[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7303[0:7]),
     .bnl_op(net_7135[0:7]), .tnr_op(net_5287[0:7]),
     .tnl_op(net_5119[0:7]));
ltile4rev I_22_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7309), .lft_op(net_5119[0:7]),
     .sp12_h_l(net_7175[0:23]), .sp4_h_l(net_7176[0:47]),
     .sp4_v_b(net_7179[0:47]), .sp12_v_b(net_7289[0:23]),
     .sp12_h_r(net_7315[0:23]), .sp4_h_r(net_7316[0:47]),
     .sp12_v_t(net_7317[0:23]), .sp4_v_t(net_5191[0:47]),
     .sp4_r_v_b(net_7319[0:47]), .wl(wl[239:224]),
     .top_op(net_7193[0:7]), .rgt_op(net_5287[0:7]),
     .bot_op(net_4729[0:7]), .bl(bl[1185:1132]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_22[7:0]),
     .carry_in(net_7281), .purst(purst), .slf_op(net_7191[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7331[0:7]),
     .bnl_op(net_7163[0:7]), .tnr_op(net_5315[0:7]),
     .tnl_op(net_5147[0:7]));
ltile4rev I_24_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7337), .lft_op(net_7331[0:7]),
     .sp12_h_l(net_7231[0:23]), .sp4_h_l(net_7232[0:47]),
     .sp4_v_b(net_7235[0:47]), .sp12_v_b(net_6645[0:23]),
     .sp12_h_r(net_7343[0:23]), .sp4_h_r(net_7344[0:47]),
     .sp12_v_t(net_7345[0:23]), .sp4_v_t(net_7375[0:47]),
     .sp4_r_v_b(net_7347[0:47]), .wl(wl[223:208]),
     .top_op(net_5231[0:7]), .rgt_op({io_r_02[3], io_r_02[2],
     io_r_02[1], io_r_02[0], io_r_02[3], io_r_02[2], io_r_02[1],
     io_r_02[0]}), .bot_op(net_7247[0:7]), .bl(bl[1293:1240]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_24[7:0]),
     .carry_in(net_6637), .purst(purst), .slf_op(net_7387[0:7]),
     .pgate(pgate[223:208]), .bnr_op({io_r_01[3], io_r_01[2],
     io_r_01[1], io_r_01[0], io_r_01[3], io_r_01[2], io_r_01[1],
     io_r_01[0]}), .bnl_op(net_7303[0:7]), .tnr_op({io_r_03[3],
     io_r_03[2], io_r_03[1], io_r_03[0], io_r_03[3], io_r_03[2],
     io_r_03[1], io_r_03[0]}), .tnl_op(net_5287[0:7]));
ltile4rev I_23_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7365), .lft_op(net_7191[0:7]),
     .sp12_h_l(net_7315[0:23]), .sp4_h_l(net_7316[0:47]),
     .sp4_v_b(net_7319[0:47]), .sp12_v_b(net_7233[0:23]),
     .sp12_h_r(net_7371[0:23]), .sp4_h_r(net_7372[0:47]),
     .sp12_v_t(net_7373[0:23]), .sp4_v_t(net_5275[0:47]),
     .sp4_r_v_b(net_7375[0:47]), .wl(wl[239:224]),
     .top_op(net_5315[0:7]), .rgt_op(net_5231[0:7]),
     .bot_op(net_7331[0:7]), .bl(bl[1239:1186]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_23[7:0]),
     .carry_in(net_7225), .purst(purst), .slf_op(net_5287[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7387[0:7]),
     .bnl_op(net_4729[0:7]), .tnr_op(net_5371[0:7]),
     .tnl_op(net_7193[0:7]));
clk_colbufx8 I785 ( .clko(glb_netwk_13[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I786 ( .clko(glb_netwk_14[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I787 ( .clko(glb_netwk_16[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I788 ( .clko(glb_netwk_15[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I789 ( .clko(glb_netwk_19[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I790 ( .clko(glb_netwk_20[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I791 ( .clko(glb_netwk_18[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I792 ( .clko(glb_netwk_17[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I793 ( .clko(glb_netwk_io_r[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I797 ( .clko(glb_netwk_23[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I798 ( .clko(glb_netwk_24[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I799 ( .clko(glb_netwk_22[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I800 ( .clko(glb_netwk_21[7:0]),
     .clki(net2col_drivers[7:0]));
io_col4 I_14_21_iot27 ( .ceb(ceb_o), .cf(cf_t[335:312]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_8216), .sdo(net_8034), .sdi(net_7422),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[14]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[27:26]), .pado(pado_t[27:26]),
     .padeb(padeb_t[27:26]), .sp4_v_t(net_8058[0:15]),
     .sp4_h_l(net_7437[0:47]), .sp12_h_l(net_5609[0:23]), .prog(prog),
     .spi_ss_in_b(net_7440[0:1]), .tnl_op(slf_op_13_10[7:0]),
     .lft_op(net_8055[0:7]), .bnl_op(net_7443[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7446[0:15]), .wl(wl[351:336]), .bl({bl[713], bl[712],
     bl[751], bl[749], bl[740], bl[746], bl[745], bl[744], bl[743],
     bl[742], bl[723], bl[722], bl[721], bl[720], bl[719], bl[718],
     bl[753], bl[752]}), .slf_op(io_t_14[3:0]),
     .glb_netwk(glb_netwk_14[7:0]));
io_col4 I_15_21_iot29 ( .ceb(ceb_o), .cf(cf_t[359:336]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_8213), .sdo(net_7422), .sdi(net_7456),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[15]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[29:28]), .pado(pado_t[29:28]),
     .padeb(padeb_t[29:28]), .sp4_v_t(net_7446[0:15]),
     .sp4_h_l(net_7471[0:47]), .sp12_h_l(net_5469[0:23]), .prog(prog),
     .spi_ss_in_b(net_7474[0:1]), .tnl_op(net_8055[0:7]),
     .lft_op(net_7443[0:7]), .bnl_op(net_7477[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7480[0:15]), .wl(wl[351:336]), .bl({bl[767], bl[766],
     bl[805], bl[803], bl[794], bl[800], bl[799], bl[798], bl[797],
     bl[796], bl[777], bl[776], bl[775], bl[774], bl[773], bl[772],
     bl[807], bl[806]}), .slf_op(io_t_15[3:0]),
     .glb_netwk(glb_netwk_15[7:0]));
io_col4 I_16_21_iot31 ( .ceb(ceb_o), .cf(cf_t[383:360]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_8206), .sdo(net_7456), .sdi(net_7490),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[16]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[31:30]), .pado(pado_t[31:30]),
     .padeb(padeb_t[31:30]), .sp4_v_t(net_7480[0:15]),
     .sp4_h_l(net_7505[0:47]), .sp12_h_l(net_5497[0:23]), .prog(prog),
     .spi_ss_in_b(net_7508[0:1]), .tnl_op(net_7443[0:7]),
     .lft_op(net_7477[0:7]), .bnl_op(net_7511[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7514[0:15]), .wl(wl[351:336]), .bl({bl[821], bl[820],
     bl[859], bl[857], bl[848], bl[854], bl[853], bl[852], bl[851],
     bl[850], bl[831], bl[830], bl[829], bl[828], bl[827], bl[826],
     bl[861], bl[860]}), .slf_op(io_t_16[3:0]),
     .glb_netwk(glb_netwk_16[7:0]));
io_col4 I_17_21_iot33 ( .ceb(ceb_o), .cf(cf_t[407:384]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_7522), .sdo(net_7490), .sdi(net_7524),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[17]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[33:32]), .pado(pado_t[33:32]),
     .padeb(padeb_t[33:32]), .sp4_v_t(net_7514[0:15]),
     .sp4_h_l(net_7539[0:47]), .sp12_h_l(net_5413[0:23]), .prog(prog),
     .spi_ss_in_b(net_7542[0:1]), .tnl_op(net_7477[0:7]),
     .lft_op(net_7511[0:7]), .bnl_op(net_7545[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7548[0:15]), .wl(wl[351:336]), .bl({bl[875], bl[874],
     bl[913], bl[911], bl[902], bl[908], bl[907], bl[906], bl[905],
     bl[904], bl[885], bl[884], bl[883], bl[882], bl[881], bl[880],
     bl[915], bl[914]}), .slf_op(io_t_17[3:0]),
     .glb_netwk(glb_netwk_17[7:0]));
io_col4 I_19_21_iot37 ( .ceb(ceb_o), .cf(cf_t[455:432]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_8208), .sdo(net_8136), .sdi(net_7592),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[19]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[37:36]), .pado(pado_t[37:36]),
     .padeb(padeb_t[37:36]), .sp4_v_t(net_8160[0:15]),
     .sp4_h_l(net_7607[0:47]), .sp12_h_l(net_4034[0:23]), .prog(prog),
     .spi_ss_in_b(net_7610[0:1]), .tnl_op(net_7545[0:7]),
     .lft_op(net_8157[0:7]), .bnl_op(net_7613[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7616[0:15]), .wl(wl[351:336]), .bl({bl[983], bl[982],
     bl[1009], bl[1007], bl[998], bl[1004], bl[1003], bl[1002],
     bl[1001], bl[1000], bl[993], bl[992], bl[991], bl[990], bl[989],
     bl[988], bl[1011], bl[1010]}), .slf_op(io_t_19[3:0]),
     .glb_netwk(glb_netwk_19[7:0]));
io_col4 I_20_21_iot39 ( .ceb(ceb_o), .cf(cf_t[479:456]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_7658), .sdo(net_7592), .sdi(net_7660),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[20]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[39:38]), .pado(pado_t[39:38]),
     .padeb(padeb_t[39:38]), .sp4_v_t(net_7616[0:15]),
     .sp4_h_l(net_7675[0:47]), .sp12_h_l(net_5749[0:23]), .prog(prog),
     .spi_ss_in_b(net_7678[0:1]), .tnl_op(net_8157[0:7]),
     .lft_op(net_7613[0:7]), .bnl_op(net_7681[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7684[0:15]), .wl(wl[351:336]), .bl({bl[1025],
     bl[1024], bl[1063], bl[1061], bl[1052], bl[1058], bl[1057],
     bl[1056], bl[1055], bl[1054], bl[1035], bl[1034], bl[1033],
     bl[1032], bl[1031], bl[1030], bl[1065], bl[1064]}),
     .slf_op(io_t_20[3:0]), .glb_netwk(glb_netwk_20[7:0]));
io_col4 I_21_21_iot41 ( .ceb(ceb_o), .cf(cf_t[503:480]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_8190), .sdo(net_7660), .sdi(net_7694),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[21]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[41:40]), .pado(pado_t[41:40]),
     .padeb(padeb_t[41:40]), .sp4_v_t(net_7684[0:15]),
     .sp4_h_l(net_7709[0:47]), .sp12_h_l(net_5777[0:23]), .prog(prog),
     .spi_ss_in_b(net_7712[0:1]), .tnl_op(net_7613[0:7]),
     .lft_op(net_7681[0:7]), .bnl_op(net_7715[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7718[0:15]), .wl(wl[351:336]), .bl({bl[1079],
     bl[1078], bl[1117], bl[1115], bl[1106], bl[1112], bl[1111],
     bl[1110], bl[1109], bl[1108], bl[1089], bl[1088], bl[1087],
     bl[1086], bl[1085], bl[1084], bl[1119], bl[1118]}),
     .slf_op(io_t_21[3:0]), .glb_netwk(glb_netwk_21[7:0]));
io_col4 I_22_21_iot43 ( .ceb(ceb_o), .cf(cf_t[527:504]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_7726), .sdo(net_7694), .sdi(net_7728),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[22]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[43:42]), .pado(pado_t[43:42]),
     .padeb(padeb_t[43:42]), .sp4_v_t(net_7718[0:15]),
     .sp4_h_l(net_7743[0:47]), .sp12_h_l(net_5917[0:23]), .prog(prog),
     .spi_ss_in_b(net_7746[0:1]), .tnl_op(net_7681[0:7]),
     .lft_op(net_7715[0:7]), .bnl_op(net_7749[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7752[0:15]), .wl(wl[351:336]), .bl({bl[1133],
     bl[1132], bl[1171], bl[1169], bl[1160], bl[1166], bl[1165],
     bl[1164], bl[1163], bl[1162], bl[1143], bl[1142], bl[1141],
     bl[1140], bl[1139], bl[1138], bl[1173], bl[1172]}),
     .slf_op(io_t_22[3:0]), .glb_netwk(glb_netwk_22[7:0]));
io_col4 I_23_21_iot45 ( .ceb(ceb_o), .cf(cf_t[551:528]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_8211), .sdo(net_7728), .sdi(net_7762),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[23]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[45:44]), .pado(pado_t[45:44]),
     .padeb(padeb_t[45:44]), .sp4_v_t(net_7752[0:15]),
     .sp4_h_l(net_7777[0:47]), .sp12_h_l(net_5973[0:23]), .prog(prog),
     .spi_ss_in_b(net_7780[0:1]), .tnl_op(net_7715[0:7]),
     .lft_op(net_7749[0:7]), .bnl_op(net_7783[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7786[0:15]), .wl(wl[351:336]), .bl({bl[1187],
     bl[1186], bl[1225], bl[1223], bl[1214], bl[1220], bl[1219],
     bl[1218], bl[1217], bl[1216], bl[1197], bl[1196], bl[1195],
     bl[1194], bl[1193], bl[1192], bl[1227], bl[1226]}),
     .slf_op(io_t_23[3:0]), .glb_netwk(glb_netwk_23[7:0]));
io_col4 I_24_21_iot47 ( .ceb(ceb_o), .cf(cf_t[575:552]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_7794), .sdo(net_7762), .sdi(net_3950),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[24]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[47:46]), .pado(pado_t[47:46]),
     .padeb(padeb_t[47:46]), .sp4_v_t(net_7786[0:15]),
     .sp4_h_l(net_7811[0:47]), .sp12_h_l(net_5861[0:23]), .prog(prog),
     .spi_ss_in_b(net_7814[0:1]), .tnl_op(net_7749[0:7]),
     .lft_op(net_7783[0:7]), .bnl_op(net_8170[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7820[0:15]), .wl(wl[351:336]), .bl({bl[1241],
     bl[1240], bl[1279], bl[1277], bl[1268], bl[1274], bl[1273],
     bl[1272], bl[1271], bl[1270], bl[1251], bl[1250], bl[1249],
     bl[1248], bl[1247], bl[1246], bl[1281], bl[1280]}),
     .slf_op(io_t_24[3:0]), .glb_netwk(glb_netwk_24[7:0]));
io_col4 I_13_21_iot25 ( .ceb(ceb_o), .cf(cf_t[311:288]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_3997), .sdo(sdo), .sdi(net_8034), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_top_r[13]), .spioeb({tievdd,
     tievdd}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[25:24]), .pado(pado_t[25:24]),
     .padeb(padeb_t[25:24]), .sp4_v_t(sp4_h_l_13_21[15:0]),
     .sp4_h_l(net_8049[0:47]), .sp12_h_l(net_5637[0:23]), .prog(prog),
     .spi_ss_in_b(net_8052[0:1]), .tnl_op(lft_op_13_10[7:0]),
     .lft_op(slf_op_13_10[7:0]), .bnl_op(net_8055[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8058[0:15]), .wl(wl[351:336]), .bl({bl[659], bl[658],
     bl[697], bl[695], bl[686], bl[692], bl[691], bl[690], bl[689],
     bl[688], bl[669], bl[668], bl[667], bl[666], bl[665], bl[664],
     bl[699], bl[698]}), .slf_op(slf_op_13_21[3:0]),
     .glb_netwk(glb_netwk_13[7:0]));
io_col4 I_18_21_iob35 ( .ceb(ceb_o), .cf(cf_t[431:408]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_r),
     .fabric_out(net_8189), .sdo(net_7524), .sdi(net_8136),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_r[18]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_t[35:34]), .pado(pado_t[35:34]),
     .padeb(padeb_t[35:34]), .sp4_v_t(net_7548[0:15]),
     .sp4_h_l(net_5554[0:47]), .sp12_h_l(net_5553[0:23]), .prog(prog),
     .spi_ss_in_b(net_8154[0:1]), .tnl_op(net_7511[0:7]),
     .lft_op(net_7545[0:7]), .bnl_op(net_8157[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8160[0:15]), .wl(wl[351:336]), .bl({bl[929], bl[928],
     bl[967], bl[965], bl[956], bl[962], bl[961], bl[960], bl[959],
     bl[958], bl[939], bl[938], bl[937], bl[936], bl[935], bl[934],
     bl[969], bl[968]}), .slf_op(io_t_18[3:0]),
     .glb_netwk(glb_netwk_18[7:0]));

endmodule
// Library - io, Cell - io_col4_row, View - schematic
// LAST TIME SAVED: Feb  8 13:53:52 2008
// NETLIST TIME: Nov 14 16:12:04 2008
`timescale 1ns / 1ns 

module io_col4_row ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [1:0]  spi_ss_in_b;
output [1:0]  padeb;
output [3:0]  slf_op;
output [23:0]  cf;

inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;

input [1:0]  padin;
input [15:0]  vdd_cntl;
input [15:0]  reset;
input [15:0]  pgate;
input [15:0]  wl;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [1:0]  spiout;
input [7:0]  lft_op;
input [1:0]  spioeb;
input [7:0]  glb_netwk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



rm7  R14_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7  R14_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7  R14_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7  R14_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7  R14_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7  R14_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7  R14_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7  R14_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7  R14_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7  R14_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7  R14_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7  R14_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7  R14_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7  R14_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7  R14_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7  R14_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[17:14],
     sp4_h_l[47:0], sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1],
     slf_op[3]}, pgate[15:0], prog, reset[15:0], vdd_cntl[15:0],
     wl[15:0]);
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl(vdd_cntl[15:0]),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[13:8]), .wl(wl[15:0]),
     .reset(reset[15:0]), .pgate(pgate[15:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(prog),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl(vdd_cntl[15:0]), .outclk(outclk),
     .fabric_out(fabric_out), .min6({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .inclk_in({lc_trk_g1[3],
     lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0], glb_netwk[7:0]}),
     .ceb_in({lc_trk_g1[5], lc_trk_g1[2], lc_trk_g0[5], lc_trk_g0[2],
     glb_netwk[6], glb_netwk[4], glb_netwk[2], glb_netwk[0]}),
     .clk_in({lc_trk_g1[4], lc_trk_g1[1], lc_trk_g0[4], lc_trk_g0[1],
     glb_netwk[7:0]}), .update(update), .spiout(spiout[1:0]),
     .spioeb(spioeb[1:0]), .padin(padin[1:0]), .out(om[1:0]),
     .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[7:2]), .inclk(inclk), .wl(wl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]), .prog(prog));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl(vdd_cntl[15:0]),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl(wl[15:0]), .reset(reset[15:0]), .pgate(pgate[15:0]),
     .hiz_b(hiz_b), .update(enable_update), .ti(ti[5:0]), .tclk(tclk),
     .shift(shift), .sdi(sdi), .prog(prog), .padin(padin[1:0]),
     .mode(mode), .inclk(inclk), .bs_en(bs_en),
     .sp12_h_l(sp12_h_l[23:0]), .sdo(sdo), .pado(om[1:0]),
     .padeb(oenm[1:0]), .bl(bl[1:0]));

endmodule
// Library - leafcell, Cell - QUAD_BL, View - schematic
// LAST TIME SAVED: Sep 15 14:12:23 2008
// NETLIST TIME: Nov 14 16:12:04 2008
`timescale 1ns / 1ns 

module QUAD_BL ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_10, carry_out_02_10,
     carry_out_03_10, carry_out_04_10, carry_out_05_10,
     carry_out_07_10, carry_out_08_10, carry_out_09_10,
     carry_out_10_10, carry_out_11_10, carry_out_12_10, ceb_o, cf_b,
     cf_l, fabric_out_34, fabric_out_38, fabric_out_93, hiz_b_o,
     mode_o, padeb_b, padeb_l, padin_34, padin_93, pado_b, pado_l, r_o,
     sdo, shift_o, slf_op_00_10, slf_op_01_10, slf_op_02_10,
     slf_op_03_10, slf_op_04_10, slf_op_05_10, slf_op_06_10,
     slf_op_07_10, slf_op_08_10, slf_op_09_10, slf_op_10_10,
     slf_op_11_10, .cdsNet0(slf_op_12_00_clash[3]),
     .cdsNet0(slf_op_12_00_clash[2]), .cdsNet0(slf_op_12_00_clash[1]),
     .cdsNet0(slf_op_12_00_clash[0]), slf_op_12_01, slf_op_12_02,
     slf_op_12_03, slf_op_12_04, slf_op_12_05, slf_op_12_06,
     slf_op_12_07, slf_op_12_08, slf_op_12_09, slf_op_12_10,
     spi_ss_in_lft_b, tclk_o, update_o, bl, pgate, reset_b,
     sp4_h_l_12_00, sp4_h_r_12_01, sp4_h_r_12_02, sp4_h_r_12_03,
     sp4_h_r_12_04, sp4_h_r_12_05, sp4_h_r_12_06, sp4_h_r_12_07,
     sp4_h_r_12_08, sp4_h_r_12_09, sp4_h_r_12_10, sp4_r_v_b_12_01,
     sp4_r_v_b_12_02, sp4_r_v_b_12_03, sp4_r_v_b_12_04,
     sp4_r_v_b_12_05, sp4_r_v_b_12_06, sp4_r_v_b_12_07,
     sp4_r_v_b_12_08, sp4_r_v_b_12_09, sp4_r_v_b_12_10, sp4_v_t_00_10,
     sp4_v_t_01_10, sp4_v_t_02_10, sp4_v_t_03_10, sp4_v_t_04_10,
     sp4_v_t_05_10, sp4_v_t_06_10, sp4_v_t_07_10, sp4_v_t_08_10,
     sp4_v_t_09_10, sp4_v_t_10_10, sp4_v_t_11_10, sp4_v_t_12_10,
     sp12_h_r_12_01, sp12_h_r_12_02, sp12_h_r_12_03, sp12_h_r_12_04,
     sp12_h_r_12_05, sp12_h_r_12_06, sp12_h_r_12_07, sp12_h_r_12_08,
     sp12_h_r_12_09, sp12_h_r_12_10, sp12_v_t_01_10, sp12_v_t_02_10,
     sp12_v_t_03_10, sp12_v_t_04_10, sp12_v_t_05_10, sp12_v_t_06_10,
     sp12_v_t_07_10, sp12_v_t_08_10, sp12_v_t_09_10, sp12_v_t_10_10,
     sp12_v_t_11_10, sp12_v_t_12_10, vdd_cntl, wl, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnr_op_12_01,
     bs_en_i, ceb_i, end_of_startup_lft_b, glb_in, hiz_b_i, hold_b_l,
     hold_l_b, mode_i, padin_b, padin_l, prog, purst, r_i,
     rgt_op_12_01, rgt_op_12_02, rgt_op_12_03, rgt_op_12_04,
     rgt_op_12_05, rgt_op_12_06, rgt_op_12_07, rgt_op_12_08,
     rgt_op_12_09, rgt_op_12_10, sdi, shift_i, spioeb_lft_b,
     spiout_lft_b, tclk_i, tiegnd, tievdd, tnl_op_00_10, tnl_op_01_10,
     tnl_op_02_10, tnl_op_03_10, tnl_op_04_10, tnl_op_05_10,
     tnl_op_06_10, tnl_op_07_10, tnl_op_08_10, tnl_op_09_10,
     tnl_op_10_10, tnl_op_11_10, tnl_op_12_10, tnr_op_01_10,
     tnr_op_02_10, tnr_op_03_10, tnr_op_04_10, tnr_op_05_10,
     tnr_op_06_10, tnr_op_07_10, tnr_op_08_10, tnr_op_09_10,
     tnr_op_10_10, tnr_op_11_10, tnr_op_12_10, top_op_01_10,
     top_op_02_10, top_op_03_10, top_op_04_10, top_op_05_10,
     top_op_06_10, top_op_07_10, top_op_08_10, top_op_09_10,
     top_op_10_10, top_op_11_10, top_op_12_10, update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_10, carry_out_02_10,
     carry_out_03_10, carry_out_04_10, carry_out_05_10,
     carry_out_07_10, carry_out_08_10, carry_out_09_10,
     carry_out_10_10, carry_out_11_10, carry_out_12_10, ceb_o,
     fabric_out_34, fabric_out_38, fabric_out_93, hiz_b_o, mode_o,
     padin_34, padin_93, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, ceb_i, hiz_b_i, hold_b_l, hold_l_b,
     mode_i, prog, purst, r_i, sdi, shift_i, tclk_i, tiegnd, tievdd,
     update_i;

output [7:0]  slf_op_09_10;
output [7:0]  slf_op_12_01;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_03_10;
output [3:0]  slf_op_00_10;
output [7:0]  slf_op_04_10;
output [7:0]  slf_op_12_04;
output [7:0]  slf_op_12_06;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_12_09;
output [7:0]  slf_op_12_08;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_12_07;
output [7:0]  slf_op_12_05;
output [7:0]  slf_op_06_10;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_10_10;
output [7:0]  slf_op_07_10;
output [7:0]  slf_op_12_03;
output [7:0]  slf_op_05_10;
output [19:0]  padeb_l;
output [7:0]  slf_op_11_10;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_02_10;
output [7:0]  slf_op_12_10;
output [7:0]  slf_op_08_10;
output [23:0]  pado_b;
output [7:0]  slf_op_01_10;
output [19:0]  spi_ss_in_lft_b;
output [19:0]  pado_l;
output [287:0]  cf_b;
output [239:0]  cf_l;
output [3:0]  slf_op_12_00_clash;
output [7:0]  slf_op_12_02;
output [23:0]  padeb_b;

inout [47:0]  sp4_v_t_12_10;
inout [23:0]  sp12_h_r_12_01;
inout [23:0]  sp12_h_r_12_06;
inout [47:0]  sp4_h_r_12_01;
inout [23:0]  sp12_h_r_12_04;
inout [23:0]  sp12_h_r_12_09;
inout [23:0]  sp12_h_r_12_07;
inout [23:0]  sp12_v_t_05_10;
inout [47:0]  sp4_r_v_b_12_05;
inout [47:0]  sp4_r_v_b_12_02;
inout [23:0]  sp12_v_t_09_10;
inout [47:0]  sp4_r_v_b_12_04;
inout [23:0]  sp12_h_r_12_08;
inout [47:0]  sp4_v_t_11_10;
inout [47:0]  sp4_h_r_12_03;
inout [23:0]  sp12_v_t_04_10;
inout [47:0]  sp4_h_r_12_08;
inout [23:0]  sp12_v_t_02_10;
inout [23:0]  sp12_v_t_08_10;
inout [47:0]  sp4_v_t_02_10;
inout [23:0]  sp12_v_t_11_10;
inout [23:0]  sp12_v_t_12_10;
inout [47:0]  sp4_v_t_06_10;
inout [47:0]  sp4_v_t_09_10;
inout [47:0]  sp4_v_t_03_10;
inout [47:0]  sp4_h_r_12_06;
inout [47:0]  sp4_h_r_12_10;
inout [47:0]  sp4_r_v_b_12_06;
inout [23:0]  sp12_h_r_12_02;
inout [23:0]  sp12_h_r_12_03;
inout [47:0]  sp4_h_r_12_07;
inout [23:0]  sp12_v_t_07_10;
inout [47:0]  sp4_r_v_b_12_01;
inout [23:0]  sp12_v_t_06_10;
inout [47:0]  sp4_r_v_b_12_08;
inout [47:0]  sp4_h_r_12_04;
inout [47:0]  sp4_v_t_01_10;
inout [23:0]  sp12_h_r_12_05;
inout [47:0]  sp4_v_t_05_10;
inout [47:0]  sp4_v_t_08_10;
inout [47:0]  sp4_h_r_12_05;
inout [47:0]  sp4_r_v_b_12_07;
inout [47:0]  sp4_h_r_12_09;
inout [47:0]  sp4_r_v_b_12_09;
inout [47:0]  sp4_h_r_12_02;
inout [47:0]  sp4_r_v_b_12_03;
inout [15:0]  sp4_v_t_00_10;
inout [15:0]  sp4_h_l_12_00;
inout [175:0]  pgate;
inout [47:0]  sp4_r_v_b_12_10;
inout [47:0]  sp4_v_t_04_10;
inout [175:0]  vdd_cntl;
inout [23:0]  sp12_v_t_01_10;
inout [47:0]  sp4_v_t_07_10;
inout [23:0]  sp12_h_r_12_10;
inout [175:0]  wl;
inout [23:0]  sp12_v_t_10_10;
inout [47:0]  sp4_v_t_10_10;
inout [175:0]  reset_b;
inout [653:0]  bl;
inout [23:0]  sp12_v_t_03_10;

input [7:0]  top_op_06_10;
input [7:0]  rgt_op_12_08;
input [7:0]  tnr_op_01_10;
input [7:0]  top_op_02_10;
input [1:0]  bm_sdo_i;
input [7:0]  tnl_op_07_10;
input [7:0]  tnr_op_09_10;
input [1:0]  bm_sweb_i;
input [7:0]  tnl_op_01_10;
input [7:0]  top_op_03_10;
input [7:0]  tnr_op_02_10;
input [7:0]  top_op_08_10;
input [7:0]  tnl_op_12_10;
input [7:0]  tnl_op_00_10;
input [7:0]  tnl_op_10_10;
input [7:0]  rgt_op_12_06;
input [7:0]  tnl_op_09_10;
input [7:0]  tnr_op_05_10;
input [7:0]  top_op_01_10;
input [7:0]  top_op_11_10;
input [7:0]  tnl_op_11_10;
input [7:0]  tnr_op_03_10;
input [1:0]  bm_sclkrw_i;
input [7:0]  tnr_op_08_10;
input [7:0]  tnl_op_08_10;
input [7:0]  tnl_op_04_10;
input [7:0]  rgt_op_12_01;
input [7:0]  tnr_op_04_10;
input [7:0]  rgt_op_12_04;
input [7:0]  bm_sa_i;
input [7:0]  tnr_op_06_10;
input [7:0]  top_op_04_10;
input [7:0]  tnl_op_02_10;
input [7:0]  top_op_05_10;
input [7:0]  rgt_op_12_02;
input [7:0]  rgt_op_12_09;
input [7:0]  rgt_op_12_10;
input [7:0]  tnr_op_10_10;
input [7:0]  rgt_op_12_05;
input [1:0]  bm_sdi_i;
input [7:0]  top_op_07_10;
input [3:0]  bnr_op_12_01;
input [7:0]  tnr_op_07_10;
input [7:0]  tnl_op_05_10;
input [7:0]  top_op_09_10;
input [7:0]  rgt_op_12_03;
input [7:0]  top_op_10_10;
input [7:0]  tnr_op_11_10;
input [7:0]  rgt_op_12_07;
input [7:0]  tnl_op_03_10;
input [7:0]  tnl_op_06_10;
input [7:0]  tnr_op_12_10;
input [19:0]  padin_l;
input [7:0]  glb_in;
input [23:0]  padin_b;
input [19:0]  spioeb_lft_b;
input [10:1]  end_of_startup_lft_b;
input [19:0]  spiout_lft_b;
input [7:0]  top_op_12_10;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net4502;

wire  [0:23]  net7544;

wire  [0:7]  net6188;

wire  [0:47]  net5559;

wire  [7:0]  glb_netwk_05;

wire  [0:15]  net4607;

wire  [0:47]  net5053;

wire  [3:0]  io_l_28;

wire  [0:47]  net8079;

wire  [0:47]  net7520;

wire  [0:23]  net4942;

wire  [0:23]  net6622;

wire  [0:47]  net5840;

wire  [0:47]  net5140;

wire  [0:47]  net7324;

wire  [0:47]  net7573;

wire  [0:47]  net7237;

wire  [0:47]  net8202;

wire  [0:23]  net7042;

wire  [0:47]  net5000;

wire  [0:1]  net8145;

wire  [0:47]  net6565;

wire  [0:47]  net5700;

wire  [0:7]  net8121;

wire  [0:47]  net7769;

wire  [0:7]  net5236;

wire  [0:47]  net6453;

wire  [0:47]  net6596;

wire  [0:1]  net8026;

wire  [0:23]  net7404;

wire  [0:23]  net5948;

wire  [0:7]  net6748;

wire  [0:23]  net5808;

wire  [0:23]  net5334;

wire  [0:47]  net6537;

wire  [0:7]  net5096;

wire  [0:23]  net6284;

wire  [0:47]  net6341;

wire  [0:47]  net4156;

wire  [0:23]  net4886;

wire  [0:7]  net7985;

wire  [0:1]  net8159;

wire  [0:23]  net5446;

wire  [0:47]  net5252;

wire  [0:7]  net4740;

wire  [0:47]  net7629;

wire  [0:23]  net6172;

wire  [0:47]  net5392;

wire  [0:47]  net6540;

wire  [0:47]  net6148;

wire  [0:47]  net4054;

wire  [0:23]  net5670;

wire  [0:47]  net7657;

wire  [0:47]  net5672;

wire  [0:23]  net5668;

wire  [0:23]  net6984;

wire  [0:23]  net7154;

wire  [0:47]  net5277;

wire  [0:7]  net6664;

wire  [0:15]  net4573;

wire  [0:7]  net5488;

wire  [0:23]  net7768;

wire  [0:47]  net7797;

wire  [0:23]  net5696;

wire  [0:47]  net6509;

wire  [3:0]  io_l_24;

wire  [0:23]  net7628;

wire  [0:7]  net7084;

wire  [0:1]  net8010;

wire  [0:23]  net4735;

wire  [0:47]  net4913;

wire  [0:23]  net7910;

wire  [0:47]  net7377;

wire  [0:47]  net5756;

wire  [0:23]  net5724;

wire  [0:47]  net4258;

wire  [0:23]  net5026;

wire  [0:47]  net4969;

wire  [7:0]  glb_netwk_06;

wire  [0:23]  net7070;

wire  [0:47]  net8035;

wire  [0:47]  net6512;

wire  [0:47]  net5644;

wire  [0:23]  net4055;

wire  [0:1]  net8252;

wire  [0:23]  net6676;

wire  [0:23]  net6872;

wire  [0:23]  net8070;

wire  [0:7]  net6878;

wire  [0:47]  net6145;

wire  [0:47]  net4360;

wire  [0:7]  net6542;

wire  [0:47]  net5165;

wire  [0:7]  net4671;

wire  [0:47]  net6092;

wire  [0:47]  net5501;

wire  [0:47]  net5109;

wire  [0:47]  net8037;

wire  [0:23]  net5500;

wire  [0:47]  net5081;

wire  [0:7]  net6552;

wire  [0:47]  net8080;

wire  [0:23]  net5920;

wire  [0:23]  net4667;

wire  [0:15]  net4325;

wire  [0:47]  net4088;

wire  [3:0]  io_b_09;

wire  [0:47]  net6008;

wire  [0:47]  net7380;

wire  [0:23]  net7630;

wire  [0:47]  net5084;

wire  [0:7]  net5656;

wire  [0:23]  net4968;

wire  [0:47]  net6089;

wire  [0:47]  net7240;

wire  [0:23]  net7714;

wire  [0:7]  net5674;

wire  [0:47]  net8201;

wire  [0:47]  net7517;

wire  [0:23]  net7770;

wire  [0:1]  net8299;

wire  [0:47]  net6204;

wire  [0:23]  net6594;

wire  [0:47]  net6176;

wire  [0:7]  net5592;

wire  [0:23]  net4463;

wire  [0:23]  net7854;

wire  [0:7]  net5432;

wire  [0:23]  net7658;

wire  [0:23]  net7236;

wire  [0:47]  net5476;

wire  [0:47]  net6985;

wire  [0:47]  net4944;

wire  [0:47]  net7716;

wire  [0:23]  net8033;

wire  [0:47]  net6033;

wire  [0:47]  net5529;

wire  [0:23]  net6144;

wire  [0:47]  net5137;

wire  [0:47]  net6428;

wire  [0:23]  net5754;

wire  [0:7]  net6048;

wire  [0:23]  net5362;

wire  [0:7]  net5264;

wire  [0:47]  net5361;

wire  [7:0]  glb_netwk_07;

wire  [0:47]  net5305;

wire  [3:0]  io_l_30;

wire  [0:47]  net6201;

wire  [0:47]  net8078;

wire  [0:23]  net4812;

wire  [0:23]  net8195;

wire  [0:47]  net6789;

wire  [0:23]  net7124;

wire  [0:47]  net7212;

wire  [0:1]  net8291;

wire  [0:7]  net7420;

wire  [0:23]  net5836;

wire  [0:47]  net6621;

wire  [0:47]  net6229;

wire  [0:7]  net7784;

wire  [0:7]  net5600;

wire  [0:23]  net6340;

wire  [0:47]  net5221;

wire  [0:7]  net5012;

wire  [0:47]  net5445;

wire  [0:7]  net6804;

wire  [0:7]  net7662;

wire  [0:47]  net5420;

wire  [3:0]  io_b_08;

wire  [0:23]  net5418;

wire  [0:23]  net4123;

wire  [0:7]  net5544;

wire  [0:47]  net4820;

wire  [0:7]  net6160;

wire  [0:47]  net5753;

wire  [0:7]  net6822;

wire  [0:47]  net5056;

wire  [0:7]  net6776;

wire  [0:23]  net7742;

wire  [0:47]  net6369;

wire  [0:23]  net4912;

wire  [0:23]  net5556;

wire  [0:47]  net6285;

wire  [0:47]  net6960;

wire  [0:47]  net7352;

wire  [0:1]  net8207;

wire  [0:47]  net5111;

wire  [0:7]  net6906;

wire  [0:15]  net4155;

wire  [0:23]  net6424;

wire  [0:7]  net5684;

wire  [7:0]  glb_netwk_10;

wire  [0:47]  net4888;

wire  [0:47]  net7492;

wire  [0:23]  net7406;

wire  [0:47]  net6257;

wire  [0:7]  net7252;

wire  [0:23]  net5726;

wire  [0:23]  net7348;

wire  [0:23]  net4701;

wire  [0:47]  net6203;

wire  [0:23]  net7999;

wire  [0:23]  net6564;

wire  [0:23]  net5220;

wire  [0:23]  net8032;

wire  [0:47]  net4326;

wire  [0:23]  net7266;

wire  [0:23]  net5922;

wire  [0:23]  net5304;

wire  [0:23]  net5080;

wire  [0:47]  net7072;

wire  [0:23]  net7684;

wire  [0:47]  net7744;

wire  [0:47]  net5389;

wire  [0:7]  net6972;

wire  [0:7]  net8218;

wire  [0:23]  net5528;

wire  [0:47]  net6792;

wire  [0:7]  net6720;

wire  [0:23]  net5444;

wire  [0:23]  net4565;

wire  [0:23]  net7574;

wire  [0:23]  net5530;

wire  [0:23]  net6760;

wire  [0:15]  net4709;

wire  [0:47]  net6761;

wire  [0:23]  net5306;

wire  [0:23]  net6818;

wire  [0:23]  net7068;

wire  [0:47]  net5333;

wire  [0:23]  net5360;

wire  [0:7]  net8171;

wire  [0:23]  net6230;

wire  [0:7]  net7532;

wire  [0:23]  net5614;

wire  [7:0]  glb_netwk_01;

wire  [0:23]  net5642;

wire  [0:15]  net4233;

wire  [0:1]  net8288;

wire  [0:23]  net6060;

wire  [0:23]  net5640;

wire  [0:47]  net5669;

wire  [0:47]  net5924;

wire  [0:23]  net5082;

wire  [0:1]  net8083;

wire  [0:47]  net7713;

wire  [0:47]  net5896;

wire  [0:47]  net8112;

wire  [0:47]  net6680;

wire  [0:23]  net5052;

wire  [0:7]  net4984;

wire  [0:47]  net5025;

wire  [0:47]  net4972;

wire  [0:23]  net5136;

wire  [0:47]  net7128;

wire  [0:47]  net7464;

wire  [0:47]  net6736;

wire  [0:47]  net4916;

wire  [0:7]  net6440;

wire  [7:0]  glb_netwk_09;

wire  [0:23]  net4429;

wire  [0:15]  net4359;

wire  [0:23]  net6592;

wire  [0:7]  net5404;

wire  [0:7]  net6888;

wire  [0:7]  net5460;

wire  [0:1]  net8162;

wire  [0:23]  net4327;

wire  [0:23]  net6342;

wire  [0:47]  net5837;

wire  [0:7]  net7616;

wire  [0:1]  net8097;

wire  [0:47]  net5585;

wire  [0:47]  net7296;

wire  [0:47]  net6845;

wire  [0:1]  net8256;

wire  [0:1]  net8281;

wire  [0:47]  net5139;

wire  [0:23]  net6062;

wire  [0:23]  net7938;

wire  [0:23]  net5250;

wire  [0:23]  net4633;

wire  [0:47]  net7156;

wire  [0:23]  net7546;

wire  [0:23]  net4970;

wire  [3:0]  io_b_11;

wire  [3:0]  io_b_05;

wire  [0:47]  net5417;

wire  [0:23]  net7126;

wire  [0:47]  net7379;

wire  [0:7]  net6608;

wire  [7:0]  glb_netwk_08;

wire  [0:1]  net8273;

wire  [0:23]  net7656;

wire  [0:23]  net6538;

wire  [0:47]  net7545;

wire  [0:7]  net7560;

wire  [0:23]  net5222;

wire  [0:47]  net5224;

wire  [0:47]  net5473;

wire  [0:7]  net5992;

wire  [0:47]  net5588;

wire  [0:23]  net4293;

wire  [0:47]  net5028;

wire  [0:47]  net6817;

wire  [0:23]  net5388;

wire  [0:23]  net6426;

wire  [0:47]  net4941;

wire  [0:47]  net7685;

wire  [0:7]  net7392;

wire  [0:47]  net5280;

wire  [0:23]  net6620;

wire  [0:1]  net8146;

wire  [0:7]  net8094;

wire  [0:7]  net5572;

wire  [0:47]  net8111;

wire  [0:23]  net5752;

wire  [0:23]  net6228;

wire  [0:23]  net5472;

wire  [0:47]  net6456;

wire  [0:23]  net4191;

wire  [0:1]  net8009;

wire  [0:7]  net7056;

wire  [0:23]  net8135;

wire  [0:1]  net8208;

wire  [0:23]  net8067;

wire  [0:47]  net5728;

wire  [0:7]  net5226;

wire  [0:23]  net5698;

wire  [0:23]  net7880;

wire  [0:7]  net5646;

wire  [0:47]  net6820;

wire  [0:47]  net6904;

wire  [0:47]  net6957;

wire  [0:47]  net6372;

wire  [0:7]  net4536;

wire  [0:23]  net7376;

wire  [0:47]  net7548;

wire  [0:23]  net7098;

wire  [0:47]  net5949;

wire  [0:23]  net6790;

wire  [0:47]  net7433;

wire  [0:7]  net6944;

wire  [0:47]  net6652;

wire  [0:47]  net5725;

wire  [0:23]  net7040;

wire  [0:23]  net7208;

wire  [0:47]  net4122;

wire  [0:23]  net6648;

wire  [0:47]  net7688;

wire  [7:0]  glb_netwk_02;

wire  [0:23]  net6004;

wire  [0:23]  net6116;

wire  [0:1]  net8298;

wire  [0:23]  net5584;

wire  [0:23]  net4531;

wire  [0:23]  net5976;

wire  [0:23]  net7378;

wire  [0:23]  net5194;

wire  [0:47]  net7940;

wire  [0:7]  net7976;

wire  [0:47]  net5616;

wire  [0:7]  net6636;

wire  [0:23]  net6844;

wire  [0:23]  net7322;

wire  [0:7]  net7868;

wire  [0:23]  net6762;

wire  [0:47]  net7321;

wire  [0:7]  net6850;

wire  [0:7]  net5058;

wire  [0:7]  net5170;

wire  [0:7]  net6570;

wire  [0:23]  net6704;

wire  [0:23]  net4089;

wire  [0:47]  net8077;

wire  [0:47]  net7604;

wire  [7:0]  glb_netwk_04;

wire  [0:7]  net5852;

wire  [0:47]  net4292;

wire  [7:0]  glb_netwk_03;

wire  [0:47]  net7461;

wire  [0:47]  net7660;

wire  [0:23]  net5332;

wire  [0:7]  net6328;

wire  [0:1]  net8084;

wire  [0:7]  net6132;

wire  [0:47]  net6901;

wire  [0:7]  net5376;

wire  [0:23]  net6900;

wire  [0:47]  net5809;

wire  [0:47]  net5196;

wire  [0:47]  net7576;

wire  [0:15]  net4471;

wire  [0:47]  net5557;

wire  [0:23]  net5110;

wire  [0:23]  net6368;

wire  [0:23]  net5054;

wire  [0:7]  net5124;

wire  [0:47]  net7489;

wire  [0:7]  net5618;

wire  [0:7]  net6468;

wire  [0:47]  net5504;

wire  [0:7]  net6076;

wire  [0:47]  net5812;

wire  [0:7]  net7588;

wire  [3:0]  io_b_01;

wire  [0:47]  net5952;

wire  [0:23]  net4813;

wire  [0:47]  net7800;

wire  [0:47]  net6733;

wire  [0:7]  net8047;

wire  [0:1]  net8023;

wire  [0:1]  net8221;

wire  [0:23]  net5502;

wire  [0:7]  net5198;

wire  [0:47]  net4885;

wire  [0:23]  net7460;

wire  [3:0]  io_b_07;

wire  [0:23]  net5866;

wire  [0:47]  net6232;

wire  [0:47]  net5980;

wire  [0:47]  net5134;

wire  [0:23]  net4497;

wire  [0:23]  net6788;

wire  [0:15]  net4539;

wire  [0:23]  net6032;

wire  [0:23]  net7490;

wire  [0:23]  net6566;

wire  [0:47]  net6764;

wire  [0:23]  net6930;

wire  [0:23]  net7826;

wire  [0:47]  net4822;

wire  [0:47]  net5560;

wire  [0:47]  net7293;

wire  [0:23]  net7516;

wire  [0:7]  net5648;

wire  [0:23]  net5838;

wire  [0:23]  net6678;

wire  [0:23]  net6312;

wire  [0:23]  net7210;

wire  [0:7]  net7700;

wire  [0:23]  net5276;

wire  [0:23]  net7238;

wire  [0:47]  net8034;

wire  [0:47]  net5193;

wire  [0:47]  net6120;

wire  [0:23]  net5810;

wire  [0:23]  net5390;

wire  [0:15]  net4743;

wire  [0:23]  net6846;

wire  [0:23]  net8110;

wire  [0:7]  net5712;

wire  [0:23]  net5978;

wire  [0:23]  net7462;

wire  [0:23]  net7852;

wire  [0:23]  net6452;

wire  [0:47]  net5613;

wire  [0:23]  net6200;

wire  [0:47]  net7209;

wire  [0:7]  net5740;

wire  [0:47]  net4821;

wire  [0:23]  net6650;

wire  [0:23]  net4361;

wire  [0:1]  net8100;

wire  [0:23]  net5108;

wire  [0:7]  net7364;

wire  [0:47]  net8204;

wire  [0:1]  net8224;

wire  [0:23]  net7712;

wire  [0:7]  net5516;

wire  [0:15]  net4291;

wire  [0:47]  net6705;

wire  [0:47]  net7069;

wire  [0:23]  net6536;

wire  [0:23]  net8109;

wire  [0:47]  net6848;

wire  [0:47]  net8114;

wire  [0:23]  net6088;

wire  [0:23]  net6202;

wire  [0:23]  net5782;

wire  [0:7]  net7448;

wire  [3:0]  io_b_06;

wire  [3:0]  io_b_04;

wire  [0:47]  net6173;

wire  [0:23]  net5248;

wire  [0:7]  net6580;

wire  [0:47]  net7632;

wire  [0:47]  net7772;

wire  [0:23]  net7882;

wire  [0:47]  net5977;

wire  [0:23]  net4996;

wire  [0:47]  net6567;

wire  [0:47]  net7853;

wire  [0:23]  net6816;

wire  [0:7]  net5824;

wire  [0:23]  net5892;

wire  [3:0]  io_b_03;

wire  [0:23]  net6734;

wire  [0:23]  net7798;

wire  [0:47]  net5921;

wire  [0:23]  net4767;

wire  [0:7]  net7728;

wire  [0:47]  net6568;

wire  [0:23]  net7014;

wire  [0:7]  net7896;

wire  [0:47]  net5112;

wire  [0:7]  net4161;

wire  [0:23]  net8071;

wire  [0:23]  net5474;

wire  [0:1]  net8253;

wire  [0:47]  net7436;

wire  [0:47]  net6316;

wire  [0:23]  net8191;

wire  [3:0]  io_l_22;

wire  [0:23]  net6732;

wire  [0:7]  net6216;

wire  [3:0]  slf_op_00_11;

wire  [0:23]  net7572;

wire  [0:47]  net7153;

wire  [0:47]  net6260;

wire  [0:47]  net6313;

wire  [0:23]  net7434;

wire  [0:23]  net6258;

wire  [0:47]  net7741;

wire  [0:47]  net8038;

wire  [0:47]  net6624;

wire  [0:47]  net6425;

wire  [0:15]  net4121;

wire  [0:47]  net5308;

wire  [0:7]  net7478;

wire  [0:47]  net8115;

wire  [0:47]  net5168;

wire  [0:23]  net5166;

wire  [0:7]  net6272;

wire  [0:47]  net7856;

wire  [0:23]  net6902;

wire  [0:23]  net4225;

wire  [0:23]  net4157;

wire  [0:23]  net5192;

wire  [0:23]  net7796;

wire  [0:47]  net6876;

wire  [0:23]  net4599;

wire  [0:23]  net7320;

wire  [0:7]  net6300;

wire  [0:47]  net6061;

wire  [0:47]  net6873;

wire  [0:23]  net5164;

wire  [0:47]  net6988;

wire  [0:23]  net6986;

wire  [0:47]  net5336;

wire  [0:1]  net8279;

wire  [0:7]  net5478;

wire  [0:47]  net7408;

wire  [0:7]  net6666;

wire  [3:0]  io_l_14;

wire  [3:0]  io_l_16;

wire  [0:23]  net6958;

wire  [0:47]  net5249;

wire  [0:23]  net7294;

wire  [0:23]  net4884;

wire  [7:0]  glb_netwk_11;

wire  [0:23]  net5586;

wire  [0:23]  net7600;

wire  [0:7]  net8020;

wire  [0:23]  net5138;

wire  [0:7]  net5114;

wire  [0:23]  net7432;

wire  [0:47]  net7601;

wire  [0:23]  net4940;

wire  [0:23]  net8194;

wire  [0:47]  net6677;

wire  [0:15]  net4675;

wire  [0:23]  net7292;

wire  [7:0]  glb_netwk_12;

wire  [0:7]  net7756;

wire  [0:15]  net4257;

wire  [0:15]  net4189;

wire  [0:23]  net5416;

wire  [0:7]  net6020;

wire  [0:47]  net6932;

wire  [0:47]  net7349;

wire  [0:15]  net4437;

wire  [0:47]  net5641;

wire  [0:23]  net5612;

wire  [0:23]  net5024;

wire  [0:23]  net7686;

wire  [0:23]  net6508;

wire  [0:23]  net5558;

wire  [0:47]  net6036;

wire  [0:47]  net6593;

wire  [0:47]  net5587;

wire  [0:23]  net6256;

wire  [0:23]  net4998;

wire  [0:47]  net6539;

wire  [0:15]  net4641;

wire  [0:23]  net7518;

wire  [0:47]  net6344;

wire  [3:0]  io_b_02;

wire  [0:7]  net8156;

wire  [0:23]  net6874;

wire  [0:47]  net4819;

wire  [0:47]  net7937;

wire  [3:0]  io_b_10;

wire  [0:23]  net7740;

wire  [0:23]  net6956;

wire  [0:23]  net4395;

wire  [0:7]  net4902;

wire  [0:23]  net6370;

wire  [0:15]  net4087;

wire  [0:7]  net7634;

wire  [0:47]  net6288;

wire  [0:47]  net7351;

wire  [0:47]  net4997;

wire  [0:23]  net4259;

wire  [0:47]  net6064;

wire  [0:23]  net6706;

wire  [0:23]  net6482;

wire  [0:47]  net5532;

wire  [0:23]  net7488;

wire  [0:47]  net4190;

wire  [0:47]  net5893;

wire  [0:47]  net7884;

wire  [0:47]  net6708;

wire  [0:23]  net5278;

wire  [0:47]  net6649;

wire  [0:23]  net7350;

wire  [3:0]  io_l_26;

wire  [3:0]  io_l_32;

wire  [0:47]  net7405;

wire  [0:23]  net7602;

wire  [0:47]  net7044;

wire  [0:23]  net6928;

wire  [0:47]  net4224;

wire  [0:23]  net6118;

wire  [0:47]  net6929;

wire  [0:47]  net6005;

wire  [0:47]  net5448;

wire  [0:47]  net8203;

wire  [0:15]  net4223;

wire  [0:23]  net5894;

wire  [0:23]  net7182;

wire  [0:7]  net6916;

wire  [0:15]  net4505;

wire  [0:7]  net5590;

wire  [0:47]  net6117;

wire  [0:7]  net5142;

wire  [0:7]  net5562;

wire  [0:47]  net7041;

wire  [0:23]  net7152;

wire  [7:0]  glb_netwk_io_l;

wire  [0:47]  net5697;

wire  [0:1]  net8264;

wire  [0:23]  net7936;

wire  [0:47]  net7881;

wire  [0:7]  net6356;

wire  [0:1]  net8284;

wire  [0:47]  net7125;

wire  [0:15]  net4403;

wire  [0:47]  net5364;

wire  [0:23]  net4914;



bram_bufferx4x6 I1091 ( .in(sdi), .out(net04069));
bram_bufferx4x6 I1092 ( .in(net4208), .out(net04068));
lowla_modified I1087 ( .clk(tclk_i), .min(net04069), .lao(net4039));
lowla_modified I1089 ( .clk(net4860), .min(net04068), .lao(net4845));
io_col4_row I_00_10_iol19 ( .ceb(net04144), .cf(cf_l[239:216]),
     .vdd_cntl(vdd_cntl[175:160]), .hold(hold_l_b),
     .fabric_out(net7974), .sdo(net4073), .sdi(net4039),
     .spiout(spiout_lft_b[19:18]), .cdone_in(end_of_startup_lft_b[10]),
     .spioeb(spioeb_lft_b[19:18]), .mode(net4213), .shift(net4214),
     .hiz_b(net4215), .r(net4216), .bs_en(net4217), .tclk(net4860),
     .update(net4219), .padin(padin_l[19:18]), .pado(pado_l[19:18]),
     .padeb(padeb_l[19:18]), .sp4_v_t(sp4_v_t_00_10[15:0]),
     .sp4_h_l(net4054[0:47]), .sp12_h_l(net4055[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[19:18]), .tnl_op(tnl_op_00_10[7:0]),
     .lft_op(slf_op_01_10[7:0]), .bnl_op(net6570[0:7]),
     .pgate(pgate[175:160]), .reset(reset_b[175:160]),
     .sp4_v_b(net4087[0:15]), .wl(wl[175:160]), .bl(bl[17:0]),
     .slf_op(slf_op_00_10[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_09_iol17 ( .ceb(net04144), .cf(cf_l[215:192]),
     .vdd_cntl(vdd_cntl[159:144]), .hold(hold_l_b),
     .fabric_out(net7960), .sdo(net4311), .sdi(net4073),
     .spiout(spiout_lft_b[17:16]), .cdone_in(end_of_startup_lft_b[9]),
     .spioeb(spioeb_lft_b[17:16]), .mode(net4213), .shift(net4214),
     .hiz_b(net4215), .r(net4216), .bs_en(net4217), .tclk(net4860),
     .update(net4219), .padin(padin_l[17:16]), .pado(pado_l[17:16]),
     .padeb(padeb_l[17:16]), .sp4_v_t(net4087[0:15]),
     .sp4_h_l(net4088[0:47]), .sp12_h_l(net4089[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[17:16]), .tnl_op(slf_op_01_10[7:0]),
     .lft_op(net6570[0:7]), .bnl_op(net6542[0:7]),
     .pgate(pgate[159:144]), .reset(reset_b[159:144]),
     .sp4_v_b(net4325[0:15]), .wl(wl[159:144]), .bl(bl[17:0]),
     .slf_op(io_l_16[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_06_iol11 ( .ceb(net04144), .cf(cf_l[143:120]),
     .vdd_cntl(vdd_cntl[111:96]), .hold(hold_l_b),
     .fabric_out(net8258), .sdo(net4141), .sdi(net4107),
     .spiout(spiout_lft_b[11:10]), .cdone_in(end_of_startup_lft_b[6]),
     .spioeb(spioeb_lft_b[11:10]), .mode(net4213), .shift(net4214),
     .hiz_b(net4215), .r(net4216), .bs_en(net4217), .tclk(net4860),
     .update(net4219), .padin(padin_l[11:10]), .pado(pado_l[11:10]),
     .padeb(padeb_l[11:10]), .sp4_v_t(net4121[0:15]),
     .sp4_h_l(net4122[0:47]), .sp12_h_l(net4123[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[11:10]), .tnl_op(net5562[0:7]),
     .lft_op(net5590[0:7]), .bnl_op(net4161[0:7]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net4155[0:15]), .wl(wl[111:96]), .bl(bl[17:0]),
     .slf_op(io_l_30[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_05_iol09 ( .ceb(net04144), .cf(cf_l[119:96]),
     .vdd_cntl(vdd_cntl[95:80]), .hold(hold_l_b), .fabric_out(net8275),
     .sdo(net4140), .sdi(net4141), .spiout(spiout_lft_b[9:8]),
     .cdone_in(end_of_startup_lft_b[5]), .spioeb(spioeb_lft_b[9:8]),
     .mode(net4213), .shift(net4214), .hiz_b(net4215), .r(net4216),
     .bs_en(net4217), .tclk(net4860), .update(net4219),
     .padin(padin_l[9:8]), .pado(pado_l[9:8]), .padeb(padeb_l[9:8]),
     .sp4_v_t(net4155[0:15]), .sp4_h_l(net4156[0:47]),
     .sp12_h_l(net4157[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[9:8]), .tnl_op(net5590[0:7]),
     .lft_op(net4161[0:7]), .bnl_op(net5592[0:7]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net4257[0:15]), .wl(wl[95:80]), .bl(bl[17:0]),
     .slf_op(io_l_28[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_02_iol03 ( .ceb(net04144), .cf(cf_l[47:24]),
     .vdd_cntl(vdd_cntl[47:32]), .hold(hold_l_b), .fabric_out(net8301),
     .sdo(net4174), .sdi(net4175), .spiout(spiout_lft_b[3:2]),
     .cdone_in(end_of_startup_lft_b[2]), .spioeb(spioeb_lft_b[3:2]),
     .mode(net4213), .shift(net4214), .hiz_b(net4215), .r(net4216),
     .bs_en(net4217), .tclk(net4860), .update(net4219),
     .padin(padin_l[3:2]), .pado(pado_l[3:2]), .padeb(padeb_l[3:2]),
     .sp4_v_t(net4189[0:15]), .sp4_h_l(net4190[0:47]),
     .sp12_h_l(net4191[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[3:2]), .tnl_op(net5114[0:7]),
     .lft_op(net5142[0:7]), .bnl_op(net4671[0:7]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net4223[0:15]), .wl(wl[47:32]), .bl(bl[17:0]),
     .slf_op(io_l_22[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_01iol01 ( .ceb(net04144), .cf(cf_l[23:0]),
     .vdd_cntl(vdd_cntl[31:16]), .hold(hold_l_b), .fabric_out(net8274),
     .sdo(net4208), .sdi(net4174), .spiout(spiout_lft_b[1:0]),
     .cdone_in(end_of_startup_lft_b[1]), .spioeb(spioeb_lft_b[1:0]),
     .mode(net4213), .shift(net4214), .hiz_b(net4215), .r(net4216),
     .bs_en(net4217), .tclk(net4860), .update(net4219),
     .padin(padin_l[1:0]), .pado(pado_l[1:0]), .padeb(padeb_l[1:0]),
     .sp4_v_t(net4223[0:15]), .sp4_h_l(net4224[0:47]),
     .sp12_h_l(net4225[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[1:0]), .tnl_op(net5142[0:7]),
     .lft_op(net4671[0:7]), .bnl_op({io_b_01[3], io_b_01[2],
     io_b_01[1], io_b_01[0], io_b_01[3], io_b_01[2], io_b_01[1],
     io_b_01[0]}), .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(net4233[0:15]), .wl(wl[31:16]), .bl(bl[17:0]),
     .slf_op(slf_op_00_11[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_04_iol07 ( .ceb(net04144), .cf(cf_l[95:72]),
     .vdd_cntl(vdd_cntl[79:64]), .hold(hold_l_b), .fabric_out(net8289),
     .sdo(net4242), .sdi(net4140), .spiout(spiout_lft_b[7:6]),
     .cdone_in(end_of_startup_lft_b[4]), .spioeb(spioeb_lft_b[7:6]),
     .mode(net4213), .shift(net4214), .hiz_b(net4215), .r(net4216),
     .bs_en(net4217), .tclk(net4860), .update(net4219),
     .padin(padin_l[7:6]), .pado(pado_l[7:6]), .padeb(padeb_l[7:6]),
     .sp4_v_t(net4257[0:15]), .sp4_h_l(net4258[0:47]),
     .sp12_h_l(net4259[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[7:6]), .tnl_op(net4161[0:7]),
     .lft_op(net5592[0:7]), .bnl_op(net5114[0:7]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net4291[0:15]), .wl(wl[79:64]), .bl(bl[17:0]),
     .slf_op(io_l_26[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_03_iol05 ( .ceb(net04144), .cf(cf_l[71:48]),
     .vdd_cntl(vdd_cntl[63:48]), .hold(hold_l_b), .fabric_out(net8294),
     .sdo(net4175), .sdi(net4242), .spiout(spiout_lft_b[5:4]),
     .cdone_in(end_of_startup_lft_b[3]), .spioeb(spioeb_lft_b[5:4]),
     .mode(net4213), .shift(net4214), .hiz_b(net4215), .r(net4216),
     .bs_en(net4217), .tclk(net4860), .update(net4219),
     .padin(padin_l[5:4]), .pado(pado_l[5:4]), .padeb(padeb_l[5:4]),
     .sp4_v_t(net4291[0:15]), .sp4_h_l(net4292[0:47]),
     .sp12_h_l(net4293[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[5:4]), .tnl_op(net5592[0:7]),
     .lft_op(net5114[0:7]), .bnl_op(net5142[0:7]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net4189[0:15]), .wl(wl[63:48]), .bl(bl[17:0]),
     .slf_op(io_l_24[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_08_iol15 ( .ceb(net04144), .cf(cf_l[191:168]),
     .vdd_cntl(vdd_cntl[143:128]), .hold(hold_l_b),
     .fabric_out(net8303), .sdo(net4345), .sdi(net4311),
     .spiout(spiout_lft_b[15:14]), .cdone_in(end_of_startup_lft_b[8]),
     .spioeb(spioeb_lft_b[15:14]), .mode(net4213), .shift(net4214),
     .hiz_b(net4215), .r(net4216), .bs_en(net4217), .tclk(net4860),
     .update(net4219), .padin(padin_l[15:14]), .pado(pado_l[15:14]),
     .padeb(padeb_l[15:14]), .sp4_v_t(net4325[0:15]),
     .sp4_h_l(net4326[0:47]), .sp12_h_l(net4327[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[15:14]), .tnl_op(net6570[0:7]),
     .lft_op(net6542[0:7]), .bnl_op(net5562[0:7]),
     .pgate(pgate[143:128]), .reset(reset_b[143:128]),
     .sp4_v_b(net4359[0:15]), .wl(wl[143:128]), .bl(bl[17:0]),
     .slf_op(io_l_14[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_07_iol13 ( .ceb(net04144), .cf(cf_l[167:144]),
     .vdd_cntl(vdd_cntl[127:112]), .hold(hold_l_b),
     .fabric_out(net8254), .sdo(net4107), .sdi(net4345),
     .spiout(spiout_lft_b[13:12]), .cdone_in(end_of_startup_lft_b[7]),
     .spioeb(spioeb_lft_b[13:12]), .mode(net4213), .shift(net4214),
     .hiz_b(net4215), .r(net4216), .bs_en(net4217), .tclk(net4860),
     .update(net4219), .padin(padin_l[13:12]), .pado(pado_l[13:12]),
     .padeb(padeb_l[13:12]), .sp4_v_t(net4359[0:15]),
     .sp4_h_l(net4360[0:47]), .sp12_h_l(net4361[0:23]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_lft_b[13:12]), .tnl_op(net6542[0:7]),
     .lft_op(net5562[0:7]), .bnl_op(net5590[0:7]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net4121[0:15]), .wl(wl[127:112]), .bl(bl[17:0]),
     .slf_op(io_l_32[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_lb I_10_00_iob19 ( .ceb(ceb_o), .cf(cf_b[239:216]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8260),
     .sdo(net4378), .sdi(net4446), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[19:18]),
     .pado(pado_b[19:18]), .padeb(padeb_b[19:18]),
     .sp4_v_t(net4471[0:15]), .sp4_h_l(net5280[0:47]),
     .sp12_h_l(net4395[0:23]), .prog(prog), .spi_ss_in_b(net8273[0:1]),
     .tnl_op(net5236[0:7]), .lft_op(net5264[0:7]),
     .bnl_op(net7252[0:7]), .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net4403[0:15]), .wl(wl[15:0]), .bl({bl[493], bl[492],
     bl[531], bl[529], bl[520], bl[526], bl[525], bl[524], bl[523],
     bl[522], bl[503], bl[502], bl[501], bl[500], bl[499], bl[498],
     bl[533], bl[532]}), .slf_op(io_b_10[3:0]),
     .glb_netwk(glb_netwk_10[7:0]));
io_col4_lb I_11_00_iob21 ( .ceb(ceb_o), .cf(cf_b[263:240]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8285),
     .sdo(net4412), .sdi(net4378), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[21:20]),
     .pado(pado_b[21:20]), .padeb(padeb_b[21:20]),
     .sp4_v_t(net4403[0:15]), .sp4_h_l(net7212[0:47]),
     .sp12_h_l(net4429[0:23]), .prog(prog), .spi_ss_in_b(net8281[0:1]),
     .tnl_op(net5264[0:7]), .lft_op(net7252[0:7]),
     .bnl_op(slf_op_12_01[7:0]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(net4437[0:15]), .wl(wl[15:0]),
     .bl({bl[547], bl[546], bl[585], bl[583], bl[574], bl[580],
     bl[579], bl[578], bl[577], bl[576], bl[557], bl[556], bl[555],
     bl[554], bl[553], bl[552], bl[587], bl[586]}),
     .slf_op(io_b_11[3:0]), .glb_netwk(glb_netwk_11[7:0]));
io_col4_lb I_09_00_iob17 ( .ceb(ceb_o), .cf(cf_b[215:192]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8280),
     .sdo(net4446), .sdi(net4684), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[17:16]),
     .pado(pado_b[17:16]), .padeb(padeb_b[17:16]),
     .sp4_v_t(net4709[0:15]), .sp4_h_l(net5196[0:47]),
     .sp12_h_l(net4463[0:23]), .prog(prog), .spi_ss_in_b(net8291[0:1]),
     .tnl_op(net4740[0:7]), .lft_op(net5236[0:7]),
     .bnl_op(net5264[0:7]), .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net4471[0:15]), .wl(wl[15:0]), .bl({bl[439], bl[438],
     bl[477], bl[475], bl[466], bl[472], bl[471], bl[470], bl[469],
     bl[468], bl[449], bl[448], bl[447], bl[446], bl[445], bl[444],
     bl[479], bl[478]}), .slf_op(io_b_09[3:0]),
     .glb_netwk(glb_netwk_09[7:0]));
io_col4_lb I_06_00_iob11 ( .ceb(ceb_o), .cf(cf_b[143:120]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8300),
     .sdo(net4480), .sdi(net4514), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[11:10]),
     .pado(pado_b[11:10]), .padeb(padeb_b[11:10]),
     .sp4_v_t(net4539[0:15]), .sp4_h_l(net4888[0:47]),
     .sp12_h_l(net4497[0:23]), .prog(prog), .spi_ss_in_b(net8253[0:1]),
     .tnl_op(net5012[0:7]), .lft_op(net4536[0:7]),
     .bnl_op(net4502[0:7]), .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net4505[0:15]), .wl(wl[15:0]), .bl({bl[289], bl[288],
     bl[315], bl[313], bl[304], bl[310], bl[309], bl[308], bl[307],
     bl[306], bl[299], bl[298], bl[297], bl[296], bl[295], bl[294],
     bl[317], bl[316]}), .slf_op(io_b_06[3:0]),
     .glb_netwk(glb_netwk_06[7:0]));
io_col4_lb I_05_00_iob09 ( .ceb(ceb_o), .cf(cf_b[119:96]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8277),
     .sdo(net4514), .sdi(net4548), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[9:8]),
     .pado(pado_b[9:8]), .padeb(padeb_b[9:8]), .sp4_v_t(net4573[0:15]),
     .sp4_h_l(net5028[0:47]), .sp12_h_l(net4531[0:23]), .prog(prog),
     .spi_ss_in_b(net8284[0:1]), .tnl_op(net4984[0:7]),
     .lft_op(net5012[0:7]), .bnl_op(net4536[0:7]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(net4539[0:15]), .wl(wl[15:0]),
     .bl({bl[235], bl[234], bl[273], bl[271], bl[262], bl[268],
     bl[267], bl[266], bl[265], bl[264], bl[245], bl[244], bl[243],
     bl[242], bl[241], bl[240], bl[275], bl[274]}),
     .slf_op(io_b_05[3:0]), .glb_netwk(glb_netwk_05[7:0]));
io_col4_lb I_04_00_iob_07 ( .ceb(ceb_o), .cf(cf_b[95:72]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8283),
     .sdo(net4548), .sdi(net4582), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[7:6]),
     .pado(pado_b[7:6]), .padeb(padeb_b[7:6]), .sp4_v_t(net4607[0:15]),
     .sp4_h_l(net4944[0:47]), .sp12_h_l(net4565[0:23]), .prog(prog),
     .spi_ss_in_b(net8256[0:1]), .tnl_op(net5096[0:7]),
     .lft_op(net4984[0:7]), .bnl_op(net5012[0:7]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(net4573[0:15]), .wl(wl[15:0]),
     .bl({bl[181], bl[180], bl[219], bl[217], bl[208], bl[214],
     bl[213], bl[212], bl[211], bl[210], bl[191], bl[190], bl[189],
     bl[188], bl[187], bl[186], bl[221], bl[220]}),
     .slf_op(io_b_04[3:0]), .glb_netwk(glb_netwk_04[7:0]));
io_col4_lb I_03_00_iob05 ( .ceb(ceb_o), .cf(cf_b[71:48]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8302),
     .sdo(net4582), .sdi(net4616), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[5:4]),
     .pado(pado_b[5:4]), .padeb(padeb_b[5:4]), .sp4_v_t(net4641[0:15]),
     .sp4_h_l(net7324[0:47]), .sp12_h_l(net4599[0:23]), .prog(prog),
     .spi_ss_in_b(net8264[0:1]), .tnl_op(net5124[0:7]),
     .lft_op(net5096[0:7]), .bnl_op(net4984[0:7]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(net4607[0:15]), .wl(wl[15:0]),
     .bl({bl[127], bl[126], bl[165], bl[163], bl[154], bl[160],
     bl[159], bl[158], bl[157], bl[156], bl[137], bl[136], bl[135],
     bl[134], bl[133], bl[132], bl[167], bl[166]}),
     .slf_op(io_b_03[3:0]), .glb_netwk(glb_netwk_03[7:0]));
io_col4_lb I_02_00_iob03 ( .ceb(ceb_o), .cf(cf_b[47:24]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8282),
     .sdo(net4616), .sdi(net4650), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[3:2]),
     .pado(pado_b[3:2]), .padeb(padeb_b[3:2]), .sp4_v_t(net4675[0:15]),
     .sp4_h_l(net5140[0:47]), .sp12_h_l(net4633[0:23]), .prog(prog),
     .spi_ss_in_b(net8252[0:1]), .tnl_op(net4671[0:7]),
     .lft_op(net5124[0:7]), .bnl_op(net5096[0:7]), .pgate(pgate[15:0]),
     .reset(reset_b[15:0]), .sp4_v_b(net4641[0:15]), .wl(wl[15:0]),
     .bl({bl[73], bl[72], bl[111], bl[109], bl[100], bl[106], bl[105],
     bl[104], bl[103], bl[102], bl[83], bl[82], bl[81], bl[80], bl[79],
     bl[78], bl[113], bl[112]}), .slf_op(io_b_02[3:0]),
     .glb_netwk(glb_netwk_02[7:0]));
io_col4_lb I_01_00_iob01 ( .ceb(ceb_o), .cf(cf_b[23:0]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8262),
     .sdo(net4650), .sdi(net4845), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[1:0]),
     .pado(pado_b[1:0]), .padeb(padeb_b[1:0]), .sp4_v_t(net4233[0:15]),
     .sp4_h_l(net5134[0:47]), .sp12_h_l(net4667[0:23]), .prog(prog),
     .spi_ss_in_b(net8288[0:1]), .tnl_op({slf_op_00_11[3],
     slf_op_00_11[2], slf_op_00_11[1], slf_op_00_11[0],
     slf_op_00_11[3], slf_op_00_11[2], slf_op_00_11[1],
     slf_op_00_11[0]}), .lft_op(net4671[0:7]), .bnl_op(net5124[0:7]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net4675[0:15]), .wl(wl[15:0]), .bl({bl[19], bl[18],
     bl[57], bl[55], bl[46], bl[52], bl[51], bl[50], bl[49], bl[48],
     bl[29], bl[28], bl[27], bl[26], bl[25], bl[24], bl[59], bl[58]}),
     .slf_op(io_b_01[3:0]), .glb_netwk(glb_netwk_01[7:0]));
io_col4_lb I_08_00_iob15 ( .ceb(ceb_o), .cf(cf_b[191:168]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8266),
     .sdo(net4684), .sdi(net4718), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[15:14]),
     .pado(pado_b[15:14]), .padeb(padeb_b[15:14]),
     .sp4_v_t(net4743[0:15]), .sp4_h_l(net5168[0:47]),
     .sp12_h_l(net4701[0:23]), .prog(prog), .spi_ss_in_b(net8298[0:1]),
     .tnl_op(net4502[0:7]), .lft_op(net4740[0:7]),
     .bnl_op(net5236[0:7]), .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net4709[0:15]), .wl(wl[15:0]), .bl({bl[385], bl[384],
     bl[423], bl[421], bl[412], bl[418], bl[417], bl[416], bl[415],
     bl[414], bl[395], bl[394], bl[393], bl[392], bl[391], bl[390],
     bl[425], bl[424]}), .slf_op(io_b_08[3:0]),
     .glb_netwk(glb_netwk_08[7:0]));
io_col4_lb I_07_00_iob13 ( .ceb(ceb_o), .cf(cf_b[167:144]),
     .vdd_cntl(vdd_cntl[15:0]), .hold(hold_b_l), .fabric_out(net8278),
     .sdo(net4718), .sdi(net4480), .spiout({tiegnd, tiegnd}),
     .cdone_in(tievdd), .spioeb({tievdd, tievdd}), .mode(mode_o),
     .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o),
     .tclk(tclk_o), .update(update_o), .padin(padin_b[13:12]),
     .pado(pado_b[13:12]), .padeb(padeb_b[13:12]),
     .sp4_v_t(net4505[0:15]), .sp4_h_l(net8202[0:47]),
     .sp12_h_l(net4735[0:23]), .prog(prog), .spi_ss_in_b(net8279[0:1]),
     .tnl_op(net4536[0:7]), .lft_op(net4502[0:7]),
     .bnl_op(net4740[0:7]), .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(net4743[0:15]), .wl(wl[15:0]), .bl({bl[331], bl[330],
     bl[369], bl[367], bl[358], bl[364], bl[363], bl[362], bl[361],
     bl[360], bl[341], bl[340], bl[339], bl[338], bl[337], bl[336],
     bl[371], bl[370]}), .slf_op(io_b_07[3:0]),
     .glb_netwk(glb_netwk_07[7:0]));
io_col4_lb I_12_00_iob23 ( .ceb(ceb_o), .cf(cf_b[287:264]),
     .vdd_cntl(vdd_cntl[15:0]), .sdo(sdo), .sdi(net4412),
     .spiout({tiegnd, tiegnd}), .cdone_in(tievdd), .spioeb({tievdd,
     tievdd}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_b[23:22]), .pado(pado_b[23:22]),
     .padeb(padeb_b[23:22]), .sp4_v_t(net4437[0:15]),
     .sp4_h_l(net7156[0:47]), .sp12_h_l(net4767[0:23]), .prog(prog),
     .spi_ss_in_b(net8299[0:1]), .tnl_op(net7252[0:7]),
     .lft_op(slf_op_12_01[7:0]), .bnl_op(rgt_op_12_01[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_h_l_12_00[15:0]), .wl(wl[15:0]), .bl({bl[601],
     bl[600], bl[639], bl[637], bl[628], bl[634], bl[633], bl[632],
     bl[631], bl[630], bl[611], bl[610], bl[609], bl[608], bl[607],
     bl[606], bl[641], bl[640]}), .slf_op(slf_op_12_00_clash[3:0]),
     .glb_netwk(glb_netwk_12[7:0]), .hold(hold_b_l),
     .fabric_out(net4781));
bram_4kprouting_bbankin I_bram_0609 ( .glb_netwk(glb_netwk_06[7:0]),
     .vdd_cntl_bot(vdd_cntl[159:144]),
     .vdd_cntl_top(vdd_cntl[175:160]), .slf_op_top(slf_op_06_10[7:0]),
     .slf_op_bot(net7985[0:7]), .wl_top(wl[175:160]),
     .wl_bot(wl[159:144]), .top_op_top(top_op_06_10[7:0]),
     .tnr_op_top(tnr_op_06_10[7:0]), .tnr_op_bot(slf_op_07_10[7:0]),
     .tnl_op_top(tnl_op_06_10[7:0]), .tnl_op_bot(slf_op_05_10[7:0]),
     .rgt_op_top(slf_op_07_10[7:0]), .rgt_op_bot(net6822[0:7]),
     .reset_b_top(reset_b[175:160]), .reset_b_bot(reset_b[159:144]),
     .prog(prog), .pgate_top(pgate[175:160]),
     .pgate_bot(pgate[159:144]), .lft_op_top(slf_op_05_10[7:0]),
     .lft_op_bot(net6048[0:7]), .bm_wdummymux_en_i(net8024),
     .bot_op_bot(net6666[0:7]), .bnr_op_top(net6822[0:7]),
     .bnr_op_bot(net6850[0:7]), .bnl_op_top(net6048[0:7]),
     .bnl_op_bot(net6076[0:7]), .sp12_v_t_top(sp12_v_t_06_10[23:0]),
     .sp12_v_b_bot(net7999[0:23]), .bm_init_i(net8019),
     .sp12_h_r_top(net4812[0:23]), .sp12_h_r_bot(net4813[0:23]),
     .sp12_h_l_top(net5948[0:23]), .sp12_h_l_bot(net5920[0:23]),
     .sp4_v_t_top(sp4_v_t_06_10[47:0]), .sp4_v_b_top(net5952[0:47]),
     .sp4_v_b_bot(net5924[0:47]), .sp4_r_v_b_top(net4819[0:47]),
     .sp4_r_v_b_bot(net4820[0:47]), .sp4_h_r_top(net4821[0:47]),
     .sp4_h_r_bot(net4822[0:47]), .sp4_h_l_top(net5949[0:47]),
     .sp4_h_l_bot(net5921[0:47]), .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(net8018), .bm_sa_i(net8020[0:7]),
     .bm_sclk_i(net8021), .bm_sclkrw_i(net8010[0:1]),
     .bm_sreb_i(net8022), .bm_sweb_i(net8023[0:1]),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sdi_i(net8009[0:1]),
     .bm_sdo_i(bm_sdo_i[1:0]), .bm_sdo_o(net8026[0:1]));
bram_bufferx4 I1069 ( .in(net4214), .out(shift_o));
bram_bufferx4 I1070 ( .in(net4213), .out(mode_o));
bram_bufferx4 I1071 ( .in(net4215), .out(hiz_b_o));
bram_bufferx4 I1072 ( .in(net4219), .out(update_o));
bram_bufferx4 I1073 ( .in(net4216), .out(r_o));
bram_bufferx4 I1074 ( .in(net4217), .out(bs_en_o));
bram_bufferx4 I885 ( .in(net4860), .out(tclk_o));
bram_bufferx4 I1088 ( .in(ceb_i), .out(net04144));
bram_bufferx4 I1076 ( .in(mode_i), .out(net4213));
bram_bufferx4 I1078 ( .in(shift_i), .out(net4214));
bram_bufferx4 I1080 ( .in(r_i), .out(net4216));
bram_bufferx4 I1081 ( .in(hiz_b_i), .out(net4215));
bram_bufferx4 I1090 ( .in(net04144), .out(ceb_o));
bram_bufferx4 I1082 ( .in(update_i), .out(net4219));
bram_bufferx4 I1077 ( .in(tclk_i), .out(net4860));
bram_bufferx4 I1079 ( .in(bs_en_i), .out(net4217));
ltile4rev I_05_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net4878), .lft_op(net4984[0:7]),
     .sp12_h_l(net5024[0:23]), .sp4_h_l(net5025[0:47]),
     .sp4_v_b(net5028[0:47]), .sp12_v_b(net4531[0:23]),
     .sp12_h_r(net4884[0:23]), .sp4_h_r(net4885[0:47]),
     .sp12_v_t(net4886[0:23]), .sp4_v_t(net5000[0:47]),
     .sp4_r_v_b(net4888[0:47]), .wl(wl[31:16]), .top_op(net7616[0:7]),
     .rgt_op(net4536[0:7]), .bot_op({io_b_05[3], io_b_05[2],
     io_b_05[1], io_b_05[0], io_b_05[3], io_b_05[2], io_b_05[1],
     io_b_05[0]}), .bl(bl[287:234]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_05[7:0]), .carry_in(net8295), .purst(purst),
     .slf_op(net5012[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_06[3],
     io_b_06[2], io_b_06[1], io_b_06[0], io_b_06[3], io_b_06[2],
     io_b_06[1], io_b_06[0]}), .bnl_op({io_b_04[3], io_b_04[2],
     io_b_04[1], io_b_04[0], io_b_04[3], io_b_04[2], io_b_04[1],
     io_b_04[0]}), .tnr_op(net4902[0:7]), .tnl_op(net7532[0:7]));
ltile4rev I_05_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net4906), .lft_op(net7532[0:7]),
     .sp12_h_l(net4996[0:23]), .sp4_h_l(net4997[0:47]),
     .sp4_v_b(net5000[0:47]), .sp12_v_b(net4886[0:23]),
     .sp12_h_r(net4912[0:23]), .sp4_h_r(net4913[0:47]),
     .sp12_v_t(net4914[0:23]), .sp4_v_t(net7604[0:47]),
     .sp4_r_v_b(net4916[0:47]), .wl(wl[47:32]), .top_op(net7588[0:7]),
     .rgt_op(net4902[0:7]), .bot_op(net5012[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net4878), .purst(purst), .slf_op(net7616[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net4536[0:7]),
     .bnl_op(net4984[0:7]), .tnr_op(net8171[0:7]),
     .tnl_op(net7560[0:7]));
ltile4rev I_03_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net4934), .lft_op(net5124[0:7]),
     .sp12_h_l(net7320[0:23]), .sp4_h_l(net7321[0:47]),
     .sp4_v_b(net7324[0:47]), .sp12_v_b(net4599[0:23]),
     .sp12_h_r(net4940[0:23]), .sp4_h_r(net4941[0:47]),
     .sp12_v_t(net4942[0:23]), .sp4_v_t(net5084[0:47]),
     .sp4_r_v_b(net4944[0:47]), .wl(wl[31:16]), .top_op(net7448[0:7]),
     .rgt_op(net4984[0:7]), .bot_op({io_b_03[3], io_b_03[2],
     io_b_03[1], io_b_03[0], io_b_03[3], io_b_03[2], io_b_03[1],
     io_b_03[0]}), .bl(bl[179:126]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_03[7:0]), .carry_in(net8269), .purst(purst),
     .slf_op(net5096[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_04[3],
     io_b_04[2], io_b_04[1], io_b_04[0], io_b_04[3], io_b_04[2],
     io_b_04[1], io_b_04[0]}), .bnl_op({io_b_02[3], io_b_02[2],
     io_b_02[1], io_b_02[0], io_b_02[3], io_b_02[2], io_b_02[1],
     io_b_02[0]}), .tnr_op(net7532[0:7]), .tnl_op(net7364[0:7]));
ltile4rev I_03_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net4962), .lft_op(net7364[0:7]),
     .sp12_h_l(net5080[0:23]), .sp4_h_l(net5081[0:47]),
     .sp4_v_b(net5084[0:47]), .sp12_v_b(net4942[0:23]),
     .sp12_h_r(net4968[0:23]), .sp4_h_r(net4969[0:47]),
     .sp12_v_t(net4970[0:23]), .sp4_v_t(net7436[0:47]),
     .sp4_r_v_b(net4972[0:47]), .wl(wl[47:32]), .top_op(net7420[0:7]),
     .rgt_op(net7532[0:7]), .bot_op(net5096[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net4934), .purst(purst), .slf_op(net7448[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net4984[0:7]),
     .bnl_op(net5124[0:7]), .tnr_op(net7560[0:7]),
     .tnl_op(net7392[0:7]));
ltile4rev I_04_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net4990), .lft_op(net7448[0:7]),
     .sp12_h_l(net4968[0:23]), .sp4_h_l(net4969[0:47]),
     .sp4_v_b(net4972[0:47]), .sp12_v_b(net5026[0:23]),
     .sp12_h_r(net4996[0:23]), .sp4_h_r(net4997[0:47]),
     .sp12_v_t(net4998[0:23]), .sp4_v_t(net7520[0:47]),
     .sp4_r_v_b(net5000[0:47]), .wl(wl[47:32]), .top_op(net7560[0:7]),
     .rgt_op(net7616[0:7]), .bot_op(net4984[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net5018), .purst(purst), .slf_op(net7532[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net5012[0:7]),
     .bnl_op(net5096[0:7]), .tnr_op(net7588[0:7]),
     .tnl_op(net7420[0:7]));
ltile4rev I_04_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net5018), .lft_op(net5096[0:7]),
     .sp12_h_l(net4940[0:23]), .sp4_h_l(net4941[0:47]),
     .sp4_v_b(net4944[0:47]), .sp12_v_b(net4565[0:23]),
     .sp12_h_r(net5024[0:23]), .sp4_h_r(net5025[0:47]),
     .sp12_v_t(net5026[0:23]), .sp4_v_t(net4972[0:47]),
     .sp4_r_v_b(net5028[0:47]), .wl(wl[31:16]), .top_op(net7532[0:7]),
     .rgt_op(net5012[0:7]), .bot_op({io_b_04[3], io_b_04[2],
     io_b_04[1], io_b_04[0], io_b_04[3], io_b_04[2], io_b_04[1],
     io_b_04[0]}), .bl(bl[233:180]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_04[7:0]), .carry_in(net8293), .purst(purst),
     .slf_op(net4984[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_05[3],
     io_b_05[2], io_b_05[1], io_b_05[0], io_b_05[3], io_b_05[2],
     io_b_05[1], io_b_05[0]}), .bnl_op({io_b_03[3], io_b_03[2],
     io_b_03[1], io_b_03[0], io_b_03[3], io_b_03[2], io_b_03[1],
     io_b_03[0]}), .tnr_op(net7616[0:7]), .tnl_op(net7448[0:7]));
ltile4rev I_07_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net5046), .lft_op(net4902[0:7]),
     .sp12_h_l(net8194[0:23]), .sp4_h_l(net8203[0:47]),
     .sp4_v_b(net8201[0:47]), .sp12_v_b(net5166[0:23]),
     .sp12_h_r(net5052[0:23]), .sp4_h_r(net5053[0:47]),
     .sp12_v_t(net5054[0:23]), .sp4_v_t(net8115[0:47]),
     .sp4_r_v_b(net5056[0:47]), .wl(wl[47:32]), .top_op(net5058[0:7]),
     .rgt_op(net5198[0:7]), .bot_op(net4502[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net5158), .purst(purst), .slf_op(net5170[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net4740[0:7]),
     .bnl_op(net4536[0:7]), .tnr_op(net5226[0:7]),
     .tnl_op(net8171[0:7]));
ltile4rev I_02_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net5074), .lft_op(net5142[0:7]),
     .sp12_h_l(net5108[0:23]), .sp4_h_l(net5109[0:47]),
     .sp4_v_b(net5112[0:47]), .sp12_v_b(net7322[0:23]),
     .sp12_h_r(net5080[0:23]), .sp4_h_r(net5081[0:47]),
     .sp12_v_t(net5082[0:23]), .sp4_v_t(net7352[0:47]),
     .sp4_r_v_b(net5084[0:47]), .wl(wl[47:32]), .top_op(net7392[0:7]),
     .rgt_op(net7448[0:7]), .bot_op(net5124[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net7314), .purst(purst), .slf_op(net7364[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net5096[0:7]),
     .bnl_op(net4671[0:7]), .tnr_op(net7420[0:7]),
     .tnl_op(net5114[0:7]));
ltile4rev I_01_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net5102), .lft_op({io_l_22[3], io_l_22[2], io_l_22[1],
     io_l_22[0], io_l_22[3], io_l_22[2], io_l_22[1], io_l_22[0]}),
     .sp12_h_l(net4191[0:23]), .sp4_h_l(net4190[0:47]),
     .sp4_v_b(net5139[0:47]), .sp12_v_b(net5138[0:23]),
     .sp12_h_r(net5108[0:23]), .sp4_h_r(net5109[0:47]),
     .sp12_v_t(net5110[0:23]), .sp4_v_t(net5111[0:47]),
     .sp4_r_v_b(net5112[0:47]), .wl(wl[47:32]), .top_op(net5114[0:7]),
     .rgt_op(net7364[0:7]), .bot_op(net4671[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net5130), .purst(purst), .slf_op(net5142[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net5124[0:7]),
     .bnl_op({slf_op_00_11[3], slf_op_00_11[2], slf_op_00_11[1],
     slf_op_00_11[0], slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0]}), .tnr_op(net7392[0:7]),
     .tnl_op({io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0],
     io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0]}));
ltile4rev I_01_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net5130), .lft_op({slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0], slf_op_00_11[3],
     slf_op_00_11[2], slf_op_00_11[1], slf_op_00_11[0]}),
     .sp12_h_l(net4225[0:23]), .sp4_h_l(net4224[0:47]),
     .sp4_v_b(net5134[0:47]), .sp12_v_b(net4667[0:23]),
     .sp12_h_r(net5136[0:23]), .sp4_h_r(net5137[0:47]),
     .sp12_v_t(net5138[0:23]), .sp4_v_t(net5139[0:47]),
     .sp4_r_v_b(net5140[0:47]), .wl(wl[31:16]), .top_op(net5142[0:7]),
     .rgt_op(net5124[0:7]), .bot_op({io_b_01[3], io_b_01[2],
     io_b_01[1], io_b_01[0], io_b_01[3], io_b_01[2], io_b_01[1],
     io_b_01[0]}), .bl(bl[71:18]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_01[7:0]), .carry_in(net8272), .purst(purst),
     .slf_op(net4671[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_02[3],
     io_b_02[2], io_b_02[1], io_b_02[0], io_b_02[3], io_b_02[2],
     io_b_02[1], io_b_02[0]}), .bnl_op({tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd}), .tnr_op(net7364[0:7]),
     .tnl_op({io_l_22[3], io_l_22[2], io_l_22[1], io_l_22[0],
     io_l_22[3], io_l_22[2], io_l_22[1], io_l_22[0]}));
ltile4rev I_07_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net5158), .lft_op(net4536[0:7]),
     .sp12_h_l(net8195[0:23]), .sp4_h_l(net8204[0:47]),
     .sp4_v_b(net8202[0:47]), .sp12_v_b(net4735[0:23]),
     .sp12_h_r(net5164[0:23]), .sp4_h_r(net5165[0:47]),
     .sp12_v_t(net5166[0:23]), .sp4_v_t(net8201[0:47]),
     .sp4_r_v_b(net5168[0:47]), .wl(wl[31:16]), .top_op(net5170[0:7]),
     .rgt_op(net4740[0:7]), .bot_op({io_b_07[3], io_b_07[2],
     io_b_07[1], io_b_07[0], io_b_07[3], io_b_07[2], io_b_07[1],
     io_b_07[0]}), .bl(bl[383:330]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_07[7:0]), .carry_in(net8271), .purst(purst),
     .slf_op(net4502[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_08[3],
     io_b_08[2], io_b_08[1], io_b_08[0], io_b_08[3], io_b_08[2],
     io_b_08[1], io_b_08[0]}), .bnl_op({io_b_06[3], io_b_06[2],
     io_b_06[1], io_b_06[0], io_b_06[3], io_b_06[2], io_b_06[1],
     io_b_06[0]}), .tnr_op(net5198[0:7]), .tnl_op(net4902[0:7]));
ltile4rev I_08_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net5186), .lft_op(net4502[0:7]),
     .sp12_h_l(net5164[0:23]), .sp4_h_l(net5165[0:47]),
     .sp4_v_b(net5168[0:47]), .sp12_v_b(net4701[0:23]),
     .sp12_h_r(net5192[0:23]), .sp4_h_r(net5193[0:47]),
     .sp12_v_t(net5194[0:23]), .sp4_v_t(net5056[0:47]),
     .sp4_r_v_b(net5196[0:47]), .wl(wl[31:16]), .top_op(net5198[0:7]),
     .rgt_op(net5236[0:7]), .bot_op({io_b_08[3], io_b_08[2],
     io_b_08[1], io_b_08[0], io_b_08[3], io_b_08[2], io_b_08[1],
     io_b_08[0]}), .bl(bl[437:384]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_08[7:0]), .carry_in(net8276), .purst(purst),
     .slf_op(net4740[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_09[3],
     io_b_09[2], io_b_09[1], io_b_09[0], io_b_09[3], io_b_09[2],
     io_b_09[1], io_b_09[0]}), .bnl_op({io_b_07[3], io_b_07[2],
     io_b_07[1], io_b_07[0], io_b_07[3], io_b_07[2], io_b_07[1],
     io_b_07[0]}), .tnr_op(net7700[0:7]), .tnl_op(net5170[0:7]));
ltile4rev I_08_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net5214), .lft_op(net5170[0:7]),
     .sp12_h_l(net5052[0:23]), .sp4_h_l(net5053[0:47]),
     .sp4_v_b(net5056[0:47]), .sp12_v_b(net5194[0:23]),
     .sp12_h_r(net5220[0:23]), .sp4_h_r(net5221[0:47]),
     .sp12_v_t(net5222[0:23]), .sp4_v_t(net7660[0:47]),
     .sp4_r_v_b(net5224[0:47]), .wl(wl[47:32]), .top_op(net5226[0:7]),
     .rgt_op(net7700[0:7]), .bot_op(net4740[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net5186), .purst(purst), .slf_op(net5198[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net5236[0:7]),
     .bnl_op(net4502[0:7]), .tnr_op(net7728[0:7]),
     .tnl_op(net5058[0:7]));
ltile4rev I_09_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net5242), .lft_op(net5198[0:7]),
     .sp12_h_l(net5220[0:23]), .sp4_h_l(net5221[0:47]),
     .sp4_v_b(net5224[0:47]), .sp12_v_b(net5278[0:23]),
     .sp12_h_r(net5248[0:23]), .sp4_h_r(net5249[0:47]),
     .sp12_v_t(net5250[0:23]), .sp4_v_t(net7688[0:47]),
     .sp4_r_v_b(net5252[0:47]), .wl(wl[47:32]), .top_op(net7728[0:7]),
     .rgt_op(net7784[0:7]), .bot_op(net5236[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net5270), .purst(purst), .slf_op(net7700[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net5264[0:7]),
     .bnl_op(net4740[0:7]), .tnr_op(net7756[0:7]),
     .tnl_op(net5226[0:7]));
ltile4rev I_09_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net5270), .lft_op(net4740[0:7]),
     .sp12_h_l(net5192[0:23]), .sp4_h_l(net5193[0:47]),
     .sp4_v_b(net5196[0:47]), .sp12_v_b(net4463[0:23]),
     .sp12_h_r(net5276[0:23]), .sp4_h_r(net5277[0:47]),
     .sp12_v_t(net5278[0:23]), .sp4_v_t(net5224[0:47]),
     .sp4_r_v_b(net5280[0:47]), .wl(wl[31:16]), .top_op(net7700[0:7]),
     .rgt_op(net5264[0:7]), .bot_op({io_b_09[3], io_b_09[2],
     io_b_09[1], io_b_09[0], io_b_09[3], io_b_09[2], io_b_09[1],
     io_b_09[0]}), .bl(bl[491:438]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_09[7:0]), .carry_in(net8286), .purst(purst),
     .slf_op(net5236[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_10[3],
     io_b_10[2], io_b_10[1], io_b_10[0], io_b_10[3], io_b_10[2],
     io_b_10[1], io_b_10[0]}), .bnl_op({io_b_08[3], io_b_08[2],
     io_b_08[1], io_b_08[0], io_b_08[3], io_b_08[2], io_b_08[1],
     io_b_08[0]}), .tnr_op(net7784[0:7]), .tnl_op(net5198[0:7]));
ltile4rev I_05_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5298), .lft_op(net5404[0:7]),
     .sp12_h_l(net5444[0:23]), .sp4_h_l(net5445[0:47]),
     .sp4_v_b(net5448[0:47]), .sp12_v_b(net7490[0:23]),
     .sp12_h_r(net5304[0:23]), .sp4_h_r(net5305[0:47]),
     .sp12_v_t(net5306[0:23]), .sp4_v_t(net5420[0:47]),
     .sp4_r_v_b(net5308[0:47]), .wl(wl[95:80]), .top_op(net6804[0:7]),
     .rgt_op(net8121[0:7]), .bot_op(net5460[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net7482), .purst(purst), .slf_op(net5432[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net7478[0:7]),
     .bnl_op(net5376[0:7]), .tnr_op(net6664[0:7]),
     .tnl_op(net6720[0:7]));
ltile4rev I_05_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5326), .lft_op(net6720[0:7]),
     .sp12_h_l(net5416[0:23]), .sp4_h_l(net5417[0:47]),
     .sp4_v_b(net5420[0:47]), .sp12_v_b(net5306[0:23]),
     .sp12_h_r(net5332[0:23]), .sp4_h_r(net5333[0:47]),
     .sp12_v_t(net5334[0:23]), .sp4_v_t(net6792[0:47]),
     .sp4_r_v_b(net5336[0:47]), .wl(wl[111:96]), .top_op(net6776[0:7]),
     .rgt_op(net6664[0:7]), .bot_op(net5432[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net5298), .purst(purst), .slf_op(net6804[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net8121[0:7]),
     .bnl_op(net5404[0:7]), .tnr_op(net8047[0:7]),
     .tnl_op(net6748[0:7]));
ltile4rev I_03_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5354), .lft_op(net5572[0:7]),
     .sp12_h_l(net5500[0:23]), .sp4_h_l(net5501[0:47]),
     .sp4_v_b(net5504[0:47]), .sp12_v_b(net7546[0:23]),
     .sp12_h_r(net5360[0:23]), .sp4_h_r(net5361[0:47]),
     .sp12_v_t(net5362[0:23]), .sp4_v_t(net5532[0:47]),
     .sp4_r_v_b(net5364[0:47]), .wl(wl[95:80]), .top_op(net6636[0:7]),
     .rgt_op(net5404[0:7]), .bot_op(net5516[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net7538), .purst(purst), .slf_op(net5544[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5376[0:7]),
     .bnl_op(net5600[0:7]), .tnr_op(net6720[0:7]),
     .tnl_op(net6552[0:7]));
ltile4rev I_03_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5382), .lft_op(net6552[0:7]),
     .sp12_h_l(net5528[0:23]), .sp4_h_l(net5529[0:47]),
     .sp4_v_b(net5532[0:47]), .sp12_v_b(net5362[0:23]),
     .sp12_h_r(net5388[0:23]), .sp4_h_r(net5389[0:47]),
     .sp12_v_t(net5390[0:23]), .sp4_v_t(net6624[0:47]),
     .sp4_r_v_b(net5392[0:47]), .wl(wl[111:96]), .top_op(net6608[0:7]),
     .rgt_op(net6720[0:7]), .bot_op(net5544[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net5354), .purst(purst), .slf_op(net6636[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5404[0:7]),
     .bnl_op(net5572[0:7]), .tnr_op(net6748[0:7]),
     .tnl_op(net6580[0:7]));
ltile4rev I_04_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5410), .lft_op(net6636[0:7]),
     .sp12_h_l(net5388[0:23]), .sp4_h_l(net5389[0:47]),
     .sp4_v_b(net5392[0:47]), .sp12_v_b(net5446[0:23]),
     .sp12_h_r(net5416[0:23]), .sp4_h_r(net5417[0:47]),
     .sp12_v_t(net5418[0:23]), .sp4_v_t(net6708[0:47]),
     .sp4_r_v_b(net5420[0:47]), .wl(wl[111:96]), .top_op(net6748[0:7]),
     .rgt_op(net6804[0:7]), .bot_op(net5404[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net5438), .purst(purst), .slf_op(net6720[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5432[0:7]),
     .bnl_op(net5544[0:7]), .tnr_op(net6776[0:7]),
     .tnl_op(net6608[0:7]));
ltile4rev I_04_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5438), .lft_op(net5544[0:7]),
     .sp12_h_l(net5360[0:23]), .sp4_h_l(net5361[0:47]),
     .sp4_v_b(net5364[0:47]), .sp12_v_b(net7574[0:23]),
     .sp12_h_r(net5444[0:23]), .sp4_h_r(net5445[0:47]),
     .sp12_v_t(net5446[0:23]), .sp4_v_t(net5392[0:47]),
     .sp4_r_v_b(net5448[0:47]), .wl(wl[95:80]), .top_op(net6720[0:7]),
     .rgt_op(net5432[0:7]), .bot_op(net5376[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net7566), .purst(purst), .slf_op(net5404[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5460[0:7]),
     .bnl_op(net5516[0:7]), .tnr_op(net6804[0:7]),
     .tnl_op(net6636[0:7]));
ltile4rev I_07_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5466), .lft_op(net6664[0:7]),
     .sp12_h_l(net8070[0:23]), .sp4_h_l(net8079[0:47]),
     .sp4_v_b(net8077[0:47]), .sp12_v_b(net5614[0:23]),
     .sp12_h_r(net5472[0:23]), .sp4_h_r(net5473[0:47]),
     .sp12_v_t(net5474[0:23]), .sp4_v_t(net8038[0:47]),
     .sp4_r_v_b(net5476[0:47]), .wl(wl[111:96]), .top_op(net5478[0:7]),
     .rgt_op(net5646[0:7]), .bot_op(net7634[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net5606), .purst(purst), .slf_op(net5618[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5488[0:7]),
     .bnl_op(net8121[0:7]), .tnr_op(net5674[0:7]),
     .tnl_op(net8047[0:7]));
ltile4rev I_02_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5494), .lft_op(net4161[0:7]),
     .sp12_h_l(net5584[0:23]), .sp4_h_l(net5585[0:47]),
     .sp4_v_b(net5588[0:47]), .sp12_v_b(net7406[0:23]),
     .sp12_h_r(net5500[0:23]), .sp4_h_r(net5501[0:47]),
     .sp12_v_t(net5502[0:23]), .sp4_v_t(net5560[0:47]),
     .sp4_r_v_b(net5504[0:47]), .wl(wl[95:80]), .top_op(net6552[0:7]),
     .rgt_op(net5544[0:7]), .bot_op(net5600[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net7398), .purst(purst), .slf_op(net5572[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5516[0:7]),
     .bnl_op(net5592[0:7]), .tnr_op(net6636[0:7]),
     .tnl_op(net5590[0:7]));
ltile4rev I_02_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5522), .lft_op(net5590[0:7]),
     .sp12_h_l(net5556[0:23]), .sp4_h_l(net5557[0:47]),
     .sp4_v_b(net5560[0:47]), .sp12_v_b(net5502[0:23]),
     .sp12_h_r(net5528[0:23]), .sp4_h_r(net5529[0:47]),
     .sp12_v_t(net5530[0:23]), .sp4_v_t(net6540[0:47]),
     .sp4_r_v_b(net5532[0:47]), .wl(wl[111:96]), .top_op(net6580[0:7]),
     .rgt_op(net6636[0:7]), .bot_op(net5572[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net5494), .purst(purst), .slf_op(net6552[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5544[0:7]),
     .bnl_op(net4161[0:7]), .tnr_op(net6608[0:7]),
     .tnl_op(net5562[0:7]));
ltile4rev I_01_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5550), .lft_op({io_l_30[3], io_l_30[2], io_l_30[1],
     io_l_30[0], io_l_30[3], io_l_30[2], io_l_30[1], io_l_30[0]}),
     .sp12_h_l(net4123[0:23]), .sp4_h_l(net4122[0:47]),
     .sp4_v_b(net5587[0:47]), .sp12_v_b(net5586[0:23]),
     .sp12_h_r(net5556[0:23]), .sp4_h_r(net5557[0:47]),
     .sp12_v_t(net5558[0:23]), .sp4_v_t(net5559[0:47]),
     .sp4_r_v_b(net5560[0:47]), .wl(wl[111:96]), .top_op(net5562[0:7]),
     .rgt_op(net6552[0:7]), .bot_op(net4161[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net5578), .purst(purst), .slf_op(net5590[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5572[0:7]), .bnl_op({io_l_28[3],
     io_l_28[2], io_l_28[1], io_l_28[0], io_l_28[3], io_l_28[2],
     io_l_28[1], io_l_28[0]}), .tnr_op(net6580[0:7]),
     .tnl_op({io_l_32[3], io_l_32[2], io_l_32[1], io_l_32[0],
     io_l_32[3], io_l_32[2], io_l_32[1], io_l_32[0]}));
ltile4rev I_01_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5578), .lft_op({io_l_28[3], io_l_28[2], io_l_28[1],
     io_l_28[0], io_l_28[3], io_l_28[2], io_l_28[1], io_l_28[0]}),
     .sp12_h_l(net4157[0:23]), .sp4_h_l(net4156[0:47]),
     .sp4_v_b(net7379[0:47]), .sp12_v_b(net7378[0:23]),
     .sp12_h_r(net5584[0:23]), .sp4_h_r(net5585[0:47]),
     .sp12_v_t(net5586[0:23]), .sp4_v_t(net5587[0:47]),
     .sp4_r_v_b(net5588[0:47]), .wl(wl[95:80]), .top_op(net5590[0:7]),
     .rgt_op(net5572[0:7]), .bot_op(net5592[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net7370), .purst(purst), .slf_op(net4161[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5600[0:7]), .bnl_op({io_l_26[3],
     io_l_26[2], io_l_26[1], io_l_26[0], io_l_26[3], io_l_26[2],
     io_l_26[1], io_l_26[0]}), .tnr_op(net6552[0:7]),
     .tnl_op({io_l_30[3], io_l_30[2], io_l_30[1], io_l_30[0],
     io_l_30[3], io_l_30[2], io_l_30[1], io_l_30[0]}));
ltile4rev I_07_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5606), .lft_op(net8121[0:7]),
     .sp12_h_l(net8071[0:23]), .sp4_h_l(net8080[0:47]),
     .sp4_v_b(net8078[0:47]), .sp12_v_b(net7630[0:23]),
     .sp12_h_r(net5612[0:23]), .sp4_h_r(net5613[0:47]),
     .sp12_v_t(net5614[0:23]), .sp4_v_t(net8077[0:47]),
     .sp4_r_v_b(net5616[0:47]), .wl(wl[95:80]), .top_op(net5618[0:7]),
     .rgt_op(net5488[0:7]), .bot_op(net7662[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net7622), .purst(purst), .slf_op(net7634[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5648[0:7]),
     .bnl_op(net7478[0:7]), .tnr_op(net5646[0:7]),
     .tnl_op(net6664[0:7]));
ltile4rev I_08_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5634), .lft_op(net7634[0:7]),
     .sp12_h_l(net5612[0:23]), .sp4_h_l(net5613[0:47]),
     .sp4_v_b(net5616[0:47]), .sp12_v_b(net7714[0:23]),
     .sp12_h_r(net5640[0:23]), .sp4_h_r(net5641[0:47]),
     .sp12_v_t(net5642[0:23]), .sp4_v_t(net5476[0:47]),
     .sp4_r_v_b(net5644[0:47]), .wl(wl[95:80]), .top_op(net5646[0:7]),
     .rgt_op(net5684[0:7]), .bot_op(net5648[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net7706), .purst(purst), .slf_op(net5488[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5656[0:7]),
     .bnl_op(net7662[0:7]), .tnr_op(net6888[0:7]),
     .tnl_op(net5618[0:7]));
ltile4rev I_08_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5662), .lft_op(net5618[0:7]),
     .sp12_h_l(net5472[0:23]), .sp4_h_l(net5473[0:47]),
     .sp4_v_b(net5476[0:47]), .sp12_v_b(net5642[0:23]),
     .sp12_h_r(net5668[0:23]), .sp4_h_r(net5669[0:47]),
     .sp12_v_t(net5670[0:23]), .sp4_v_t(net6848[0:47]),
     .sp4_r_v_b(net5672[0:47]), .wl(wl[111:96]), .top_op(net5674[0:7]),
     .rgt_op(net6888[0:7]), .bot_op(net5488[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net5634), .purst(purst), .slf_op(net5646[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5684[0:7]),
     .bnl_op(net7634[0:7]), .tnr_op(net6916[0:7]),
     .tnl_op(net5478[0:7]));
ltile4rev I_09_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5690), .lft_op(net5646[0:7]),
     .sp12_h_l(net5668[0:23]), .sp4_h_l(net5669[0:47]),
     .sp4_v_b(net5672[0:47]), .sp12_v_b(net5726[0:23]),
     .sp12_h_r(net5696[0:23]), .sp4_h_r(net5697[0:47]),
     .sp12_v_t(net5698[0:23]), .sp4_v_t(net6876[0:47]),
     .sp4_r_v_b(net5700[0:47]), .wl(wl[111:96]), .top_op(net6916[0:7]),
     .rgt_op(net6972[0:7]), .bot_op(net5684[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net5718), .purst(purst), .slf_op(net6888[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5712[0:7]),
     .bnl_op(net5488[0:7]), .tnr_op(net6944[0:7]),
     .tnl_op(net5674[0:7]));
ltile4rev I_09_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5718), .lft_op(net5488[0:7]),
     .sp12_h_l(net5640[0:23]), .sp4_h_l(net5641[0:47]),
     .sp4_v_b(net5644[0:47]), .sp12_v_b(net7742[0:23]),
     .sp12_h_r(net5724[0:23]), .sp4_h_r(net5725[0:47]),
     .sp12_v_t(net5726[0:23]), .sp4_v_t(net5672[0:47]),
     .sp4_r_v_b(net5728[0:47]), .wl(wl[95:80]), .top_op(net6888[0:7]),
     .rgt_op(net5712[0:7]), .bot_op(net5656[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net7734), .purst(purst), .slf_op(net5684[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5740[0:7]),
     .bnl_op(net5648[0:7]), .tnr_op(net6972[0:7]),
     .tnl_op(net5646[0:7]));
ltile4rev I_11_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5746), .lft_op(net5712[0:7]),
     .sp12_h_l(net5808[0:23]), .sp4_h_l(net5809[0:47]),
     .sp4_v_b(net5812[0:47]), .sp12_v_b(net7938[0:23]),
     .sp12_h_r(net5752[0:23]), .sp4_h_r(net5753[0:47]),
     .sp12_v_t(net5754[0:23]), .sp4_v_t(net5840[0:47]),
     .sp4_r_v_b(net5756[0:47]), .wl(wl[95:80]), .top_op(net7056[0:7]),
     .rgt_op(slf_op_12_05[7:0]), .bot_op(net5824[0:7]),
     .bl(bl[599:546]), .reset_b(reset_b[95:80]),
     .glb_netwk(glb_netwk_11[7:0]), .carry_in(net7930), .purst(purst),
     .slf_op(net5852[0:7]), .pgate(pgate[95:80]),
     .bnr_op(slf_op_12_04[7:0]), .bnl_op(net5740[0:7]),
     .tnr_op(slf_op_12_06[7:0]), .tnl_op(net6972[0:7]));
ltile4rev I_12_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net7108), .lft_op(net7056[0:7]),
     .sp12_h_l(net5892[0:23]), .sp4_h_l(net5893[0:47]),
     .sp4_v_b(net5896[0:47]), .sp12_v_b(net5866[0:23]),
     .sp12_h_r(sp12_h_r_12_06[23:0]), .sp4_h_r(sp4_h_r_12_06[47:0]),
     .sp12_v_t(net5782[0:23]), .sp4_v_t(net6988[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_06[47:0]), .wl(wl[111:96]),
     .top_op(slf_op_12_07[7:0]), .rgt_op(rgt_op_12_06[7:0]),
     .bot_op(slf_op_12_05[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net5858), .purst(purst), .slf_op(slf_op_12_06[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_12_05[7:0]),
     .bnl_op(net5852[0:7]), .tnr_op(rgt_op_12_07[7:0]),
     .tnl_op(net7084[0:7]));
ltile4rev I_10_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5802), .lft_op(net5684[0:7]),
     .sp12_h_l(net5724[0:23]), .sp4_h_l(net5725[0:47]),
     .sp4_v_b(net5728[0:47]), .sp12_v_b(net7882[0:23]),
     .sp12_h_r(net5808[0:23]), .sp4_h_r(net5809[0:47]),
     .sp12_v_t(net5810[0:23]), .sp4_v_t(net5700[0:47]),
     .sp4_r_v_b(net5812[0:47]), .wl(wl[95:80]), .top_op(net6972[0:7]),
     .rgt_op(net5852[0:7]), .bot_op(net5740[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net7874), .purst(purst), .slf_op(net5712[0:7]),
     .pgate(pgate[95:80]), .bnr_op(net5824[0:7]),
     .bnl_op(net5656[0:7]), .tnr_op(net7056[0:7]),
     .tnl_op(net6888[0:7]));
ltile4rev I_10_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5830), .lft_op(net6888[0:7]),
     .sp12_h_l(net5696[0:23]), .sp4_h_l(net5697[0:47]),
     .sp4_v_b(net5700[0:47]), .sp12_v_b(net5810[0:23]),
     .sp12_h_r(net5836[0:23]), .sp4_h_r(net5837[0:47]),
     .sp12_v_t(net5838[0:23]), .sp4_v_t(net6960[0:47]),
     .sp4_r_v_b(net5840[0:47]), .wl(wl[111:96]), .top_op(net6944[0:7]),
     .rgt_op(net7056[0:7]), .bot_op(net5712[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[111:96]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net5802), .purst(purst), .slf_op(net6972[0:7]),
     .pgate(pgate[111:96]), .bnr_op(net5852[0:7]),
     .bnl_op(net5684[0:7]), .tnr_op(net7084[0:7]),
     .tnl_op(net6916[0:7]));
ltile4rev I_12_05 ( .vdd_cntl(vdd_cntl[95:80]), .prog(prog),
     .carry_out(net5858), .lft_op(net5852[0:7]),
     .sp12_h_l(net5752[0:23]), .sp4_h_l(net5753[0:47]),
     .sp4_v_b(net5756[0:47]), .sp12_v_b(net7826[0:23]),
     .sp12_h_r(sp12_h_r_12_05[23:0]), .sp4_h_r(sp4_h_r_12_05[47:0]),
     .sp12_v_t(net5866[0:23]), .sp4_v_t(net5896[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_05[47:0]), .wl(wl[95:80]),
     .top_op(slf_op_12_06[7:0]), .rgt_op(rgt_op_12_05[7:0]),
     .bot_op(slf_op_12_04[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[95:80]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net7818), .purst(purst), .slf_op(slf_op_12_05[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_12_04[7:0]),
     .bnl_op(net5824[0:7]), .tnr_op(rgt_op_12_06[7:0]),
     .tnl_op(net7056[0:7]));
ltile4rev I_11_06 ( .vdd_cntl(vdd_cntl[111:96]), .prog(prog),
     .carry_out(net5886), .lft_op(net6972[0:7]),
     .sp12_h_l(net5836[0:23]), .sp4_h_l(net5837[0:47]),
     .sp4_v_b(net5840[0:47]), .sp12_v_b(net5754[0:23]),
     .sp12_h_r(net5892[0:23]), .sp4_h_r(net5893[0:47]),
     .sp12_v_t(net5894[0:23]), .sp4_v_t(net7044[0:47]),
     .sp4_r_v_b(net5896[0:47]), .wl(wl[111:96]), .top_op(net7084[0:7]),
     .rgt_op(slf_op_12_06[7:0]), .bot_op(net5852[0:7]),
     .bl(bl[599:546]), .reset_b(reset_b[111:96]),
     .glb_netwk(glb_netwk_11[7:0]), .carry_in(net5746), .purst(purst),
     .slf_op(net7056[0:7]), .pgate(pgate[111:96]),
     .bnr_op(slf_op_12_05[7:0]), .bnl_op(net5712[0:7]),
     .tnr_op(slf_op_12_07[7:0]), .tnl_op(net6944[0:7]));
ltile4rev I_05_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net5914), .lft_op(net6020[0:7]),
     .sp12_h_l(net6060[0:23]), .sp4_h_l(net6061[0:47]),
     .sp4_v_b(net6064[0:47]), .sp12_v_b(net6678[0:23]),
     .sp12_h_r(net5920[0:23]), .sp4_h_r(net5921[0:47]),
     .sp12_v_t(net5922[0:23]), .sp4_v_t(net6036[0:47]),
     .sp4_r_v_b(net5924[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_05_10[7:0]), .rgt_op(net7985[0:7]),
     .bot_op(net6076[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net6670), .purst(purst), .slf_op(net6048[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net6666[0:7]),
     .bnl_op(net5992[0:7]), .tnr_op(slf_op_06_10[7:0]),
     .tnl_op(slf_op_04_10[7:0]));
ltile4rev I_05_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_05_10), .lft_op(slf_op_04_10[7:0]),
     .sp12_h_l(net6032[0:23]), .sp4_h_l(net6033[0:47]),
     .sp4_v_b(net6036[0:47]), .sp12_v_b(net5922[0:23]),
     .sp12_h_r(net5948[0:23]), .sp4_h_r(net5949[0:47]),
     .sp12_v_t(sp12_v_t_05_10[23:0]), .sp4_v_t(sp4_v_t_05_10[47:0]),
     .sp4_r_v_b(net5952[0:47]), .wl(wl[175:160]),
     .top_op(top_op_05_10[7:0]), .rgt_op(slf_op_06_10[7:0]),
     .bot_op(net6048[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net5914), .purst(purst), .slf_op(slf_op_05_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net7985[0:7]),
     .bnl_op(net6020[0:7]), .tnr_op(tnr_op_05_10[7:0]),
     .tnl_op(tnl_op_05_10[7:0]));
ltile4rev I_03_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net5970), .lft_op(net6188[0:7]),
     .sp12_h_l(net6116[0:23]), .sp4_h_l(net6117[0:47]),
     .sp4_v_b(net6120[0:47]), .sp12_v_b(net6734[0:23]),
     .sp12_h_r(net5976[0:23]), .sp4_h_r(net5977[0:47]),
     .sp12_v_t(net5978[0:23]), .sp4_v_t(net6148[0:47]),
     .sp4_r_v_b(net5980[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_03_10[7:0]), .rgt_op(net6020[0:7]),
     .bot_op(net6132[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net6726), .purst(purst), .slf_op(net6160[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net5992[0:7]),
     .bnl_op(net6216[0:7]), .tnr_op(slf_op_04_10[7:0]),
     .tnl_op(slf_op_02_10[7:0]));
ltile4rev I_03_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_03_10), .lft_op(slf_op_02_10[7:0]),
     .sp12_h_l(net6144[0:23]), .sp4_h_l(net6145[0:47]),
     .sp4_v_b(net6148[0:47]), .sp12_v_b(net5978[0:23]),
     .sp12_h_r(net6004[0:23]), .sp4_h_r(net6005[0:47]),
     .sp12_v_t(sp12_v_t_03_10[23:0]), .sp4_v_t(sp4_v_t_03_10[47:0]),
     .sp4_r_v_b(net6008[0:47]), .wl(wl[175:160]),
     .top_op(top_op_03_10[7:0]), .rgt_op(slf_op_04_10[7:0]),
     .bot_op(net6160[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net5970), .purst(purst), .slf_op(slf_op_03_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6020[0:7]),
     .bnl_op(net6188[0:7]), .tnr_op(tnr_op_03_10[7:0]),
     .tnl_op(tnl_op_03_10[7:0]));
ltile4rev I_04_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_04_10), .lft_op(slf_op_03_10[7:0]),
     .sp12_h_l(net6004[0:23]), .sp4_h_l(net6005[0:47]),
     .sp4_v_b(net6008[0:47]), .sp12_v_b(net6062[0:23]),
     .sp12_h_r(net6032[0:23]), .sp4_h_r(net6033[0:47]),
     .sp12_v_t(sp12_v_t_04_10[23:0]), .sp4_v_t(sp4_v_t_04_10[47:0]),
     .sp4_r_v_b(net6036[0:47]), .wl(wl[175:160]),
     .top_op(top_op_04_10[7:0]), .rgt_op(slf_op_05_10[7:0]),
     .bot_op(net6020[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net6054), .purst(purst), .slf_op(slf_op_04_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6048[0:7]),
     .bnl_op(net6160[0:7]), .tnr_op(tnr_op_04_10[7:0]),
     .tnl_op(tnl_op_04_10[7:0]));
ltile4rev I_04_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6054), .lft_op(net6160[0:7]),
     .sp12_h_l(net5976[0:23]), .sp4_h_l(net5977[0:47]),
     .sp4_v_b(net5980[0:47]), .sp12_v_b(net6762[0:23]),
     .sp12_h_r(net6060[0:23]), .sp4_h_r(net6061[0:47]),
     .sp12_v_t(net6062[0:23]), .sp4_v_t(net6008[0:47]),
     .sp4_r_v_b(net6064[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_04_10[7:0]), .rgt_op(net6048[0:7]),
     .bot_op(net5992[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net6754), .purst(purst), .slf_op(net6020[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net6076[0:7]),
     .bnl_op(net6132[0:7]), .tnr_op(slf_op_05_10[7:0]),
     .tnl_op(slf_op_03_10[7:0]));
ltile4rev I_07_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_07_10), .lft_op(slf_op_06_10[7:0]),
     .sp12_h_l(net4812[0:23]), .sp4_h_l(net4821[0:47]),
     .sp4_v_b(net4819[0:47]), .sp12_v_b(net6230[0:23]),
     .sp12_h_r(net6088[0:23]), .sp4_h_r(net6089[0:47]),
     .sp12_v_t(sp12_v_t_07_10[23:0]), .sp4_v_t(sp4_v_t_07_10[47:0]),
     .sp4_r_v_b(net6092[0:47]), .wl(wl[175:160]),
     .top_op(top_op_07_10[7:0]), .rgt_op(slf_op_08_10[7:0]),
     .bot_op(net6822[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net6222), .purst(purst), .slf_op(slf_op_07_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6906[0:7]),
     .bnl_op(net7985[0:7]), .tnr_op(tnr_op_07_10[7:0]),
     .tnl_op(tnl_op_07_10[7:0]));
ltile4rev I_02_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6110), .lft_op(net6570[0:7]),
     .sp12_h_l(net6200[0:23]), .sp4_h_l(net6201[0:47]),
     .sp4_v_b(net6204[0:47]), .sp12_v_b(net6594[0:23]),
     .sp12_h_r(net6116[0:23]), .sp4_h_r(net6117[0:47]),
     .sp12_v_t(net6118[0:23]), .sp4_v_t(net6176[0:47]),
     .sp4_r_v_b(net6120[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_02_10[7:0]), .rgt_op(net6160[0:7]),
     .bot_op(net6216[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net6586), .purst(purst), .slf_op(net6188[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net6132[0:7]),
     .bnl_op(net6542[0:7]), .tnr_op(slf_op_03_10[7:0]),
     .tnl_op(slf_op_01_10[7:0]));
ltile4rev I_02_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_02_10), .lft_op(slf_op_01_10[7:0]),
     .sp12_h_l(net6172[0:23]), .sp4_h_l(net6173[0:47]),
     .sp4_v_b(net6176[0:47]), .sp12_v_b(net6118[0:23]),
     .sp12_h_r(net6144[0:23]), .sp4_h_r(net6145[0:47]),
     .sp12_v_t(sp12_v_t_02_10[23:0]), .sp4_v_t(sp4_v_t_02_10[47:0]),
     .sp4_r_v_b(net6148[0:47]), .wl(wl[175:160]),
     .top_op(top_op_02_10[7:0]), .rgt_op(slf_op_03_10[7:0]),
     .bot_op(net6188[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net6110), .purst(purst), .slf_op(slf_op_02_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6160[0:7]),
     .bnl_op(net6570[0:7]), .tnr_op(tnr_op_02_10[7:0]),
     .tnl_op(tnl_op_02_10[7:0]));
ltile4rev I_01_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_01_10), .lft_op({slf_op_00_10[3],
     slf_op_00_10[2], slf_op_00_10[1], slf_op_00_10[0],
     slf_op_00_10[3], slf_op_00_10[2], slf_op_00_10[1],
     slf_op_00_10[0]}), .sp12_h_l(net4055[0:23]),
     .sp4_h_l(net4054[0:47]), .sp4_v_b(net6203[0:47]),
     .sp12_v_b(net6202[0:23]), .sp12_h_r(net6172[0:23]),
     .sp4_h_r(net6173[0:47]), .sp12_v_t(sp12_v_t_01_10[23:0]),
     .sp4_v_t(sp4_v_t_01_10[47:0]), .sp4_r_v_b(net6176[0:47]),
     .wl(wl[175:160]), .top_op(top_op_01_10[7:0]),
     .rgt_op(slf_op_02_10[7:0]), .bot_op(net6570[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net6194), .purst(purst), .slf_op(slf_op_01_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6188[0:7]),
     .bnl_op({io_l_16[3], io_l_16[2], io_l_16[1], io_l_16[0],
     io_l_16[3], io_l_16[2], io_l_16[1], io_l_16[0]}),
     .tnr_op(tnr_op_01_10[7:0]), .tnl_op(tnl_op_01_10[7:0]));
ltile4rev I_01_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6194), .lft_op({io_l_16[3], io_l_16[2], io_l_16[1],
     io_l_16[0], io_l_16[3], io_l_16[2], io_l_16[1], io_l_16[0]}),
     .sp12_h_l(net4089[0:23]), .sp4_h_l(net4088[0:47]),
     .sp4_v_b(net6567[0:47]), .sp12_v_b(net6566[0:23]),
     .sp12_h_r(net6200[0:23]), .sp4_h_r(net6201[0:47]),
     .sp12_v_t(net6202[0:23]), .sp4_v_t(net6203[0:47]),
     .sp4_r_v_b(net6204[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_01_10[7:0]), .rgt_op(net6188[0:7]),
     .bot_op(net6542[0:7]), .bl(bl[71:18]), .reset_b(reset_b[159:144]),
     .glb_netwk(glb_netwk_01[7:0]), .carry_in(net6558), .purst(purst),
     .slf_op(net6570[0:7]), .pgate(pgate[159:144]),
     .bnr_op(net6216[0:7]), .bnl_op({io_l_14[3], io_l_14[2],
     io_l_14[1], io_l_14[0], io_l_14[3], io_l_14[2], io_l_14[1],
     io_l_14[0]}), .tnr_op(slf_op_02_10[7:0]),
     .tnl_op({slf_op_00_10[3], slf_op_00_10[2], slf_op_00_10[1],
     slf_op_00_10[0], slf_op_00_10[3], slf_op_00_10[2],
     slf_op_00_10[1], slf_op_00_10[0]}));
ltile4rev I_07_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6222), .lft_op(net7985[0:7]),
     .sp12_h_l(net4813[0:23]), .sp4_h_l(net4822[0:47]),
     .sp4_v_b(net4820[0:47]), .sp12_v_b(net6818[0:23]),
     .sp12_h_r(net6228[0:23]), .sp4_h_r(net6229[0:47]),
     .sp12_v_t(net6230[0:23]), .sp4_v_t(net4819[0:47]),
     .sp4_r_v_b(net6232[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_07_10[7:0]), .rgt_op(net6906[0:7]),
     .bot_op(net6850[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net6810), .purst(purst), .slf_op(net6822[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net6878[0:7]),
     .bnl_op(net6666[0:7]), .tnr_op(slf_op_08_10[7:0]),
     .tnl_op(slf_op_06_10[7:0]));
ltile4rev I_08_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6250), .lft_op(net6822[0:7]),
     .sp12_h_l(net6228[0:23]), .sp4_h_l(net6229[0:47]),
     .sp4_v_b(net6232[0:47]), .sp12_v_b(net6902[0:23]),
     .sp12_h_r(net6256[0:23]), .sp4_h_r(net6257[0:47]),
     .sp12_v_t(net6258[0:23]), .sp4_v_t(net6092[0:47]),
     .sp4_r_v_b(net6260[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_08_10[7:0]), .rgt_op(net6300[0:7]),
     .bot_op(net6878[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net6894), .purst(purst), .slf_op(net6906[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net6272[0:7]),
     .bnl_op(net6850[0:7]), .tnr_op(slf_op_09_10[7:0]),
     .tnl_op(slf_op_07_10[7:0]));
ltile4rev I_08_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_08_10), .lft_op(slf_op_07_10[7:0]),
     .sp12_h_l(net6088[0:23]), .sp4_h_l(net6089[0:47]),
     .sp4_v_b(net6092[0:47]), .sp12_v_b(net6258[0:23]),
     .sp12_h_r(net6284[0:23]), .sp4_h_r(net6285[0:47]),
     .sp12_v_t(sp12_v_t_08_10[23:0]), .sp4_v_t(sp4_v_t_08_10[47:0]),
     .sp4_r_v_b(net6288[0:47]), .wl(wl[175:160]),
     .top_op(top_op_08_10[7:0]), .rgt_op(slf_op_09_10[7:0]),
     .bot_op(net6906[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net6250), .purst(purst), .slf_op(slf_op_08_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6300[0:7]),
     .bnl_op(net6822[0:7]), .tnr_op(tnr_op_08_10[7:0]),
     .tnl_op(tnl_op_08_10[7:0]));
ltile4rev I_09_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_09_10), .lft_op(slf_op_08_10[7:0]),
     .sp12_h_l(net6284[0:23]), .sp4_h_l(net6285[0:47]),
     .sp4_v_b(net6288[0:47]), .sp12_v_b(net6342[0:23]),
     .sp12_h_r(net6312[0:23]), .sp4_h_r(net6313[0:47]),
     .sp12_v_t(sp12_v_t_09_10[23:0]), .sp4_v_t(sp4_v_t_09_10[47:0]),
     .sp4_r_v_b(net6316[0:47]), .wl(wl[175:160]),
     .top_op(top_op_09_10[7:0]), .rgt_op(slf_op_10_10[7:0]),
     .bot_op(net6300[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net6334), .purst(purst), .slf_op(slf_op_09_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6328[0:7]),
     .bnl_op(net6906[0:7]), .tnr_op(tnr_op_09_10[7:0]),
     .tnl_op(tnl_op_09_10[7:0]));
ltile4rev I_09_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6334), .lft_op(net6906[0:7]),
     .sp12_h_l(net6256[0:23]), .sp4_h_l(net6257[0:47]),
     .sp4_v_b(net6260[0:47]), .sp12_v_b(net6930[0:23]),
     .sp12_h_r(net6340[0:23]), .sp4_h_r(net6341[0:47]),
     .sp12_v_t(net6342[0:23]), .sp4_v_t(net6288[0:47]),
     .sp4_r_v_b(net6344[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_09_10[7:0]), .rgt_op(net6328[0:7]),
     .bot_op(net6272[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net6922), .purst(purst), .slf_op(net6300[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net6356[0:7]),
     .bnl_op(net6878[0:7]), .tnr_op(slf_op_10_10[7:0]),
     .tnl_op(slf_op_08_10[7:0]));
ltile4rev I_11_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6362), .lft_op(net6328[0:7]),
     .sp12_h_l(net6424[0:23]), .sp4_h_l(net6425[0:47]),
     .sp4_v_b(net6428[0:47]), .sp12_v_b(net7126[0:23]),
     .sp12_h_r(net6368[0:23]), .sp4_h_r(net6369[0:47]),
     .sp12_v_t(net6370[0:23]), .sp4_v_t(net6456[0:47]),
     .sp4_r_v_b(net6372[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_11_10[7:0]), .rgt_op(slf_op_12_09[7:0]),
     .bot_op(net6440[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net7118), .purst(purst), .slf_op(net6468[0:7]),
     .pgate(pgate[159:144]), .bnr_op(slf_op_12_08[7:0]),
     .bnl_op(net6356[0:7]), .tnr_op(slf_op_12_10[7:0]),
     .tnl_op(slf_op_10_10[7:0]));
ltile4rev I_12_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_12_10), .lft_op(slf_op_11_10[7:0]),
     .sp12_h_l(net6508[0:23]), .sp4_h_l(net6509[0:47]),
     .sp4_v_b(net6512[0:47]), .sp12_v_b(net6482[0:23]),
     .sp12_h_r(sp12_h_r_12_10[23:0]), .sp4_h_r(sp4_h_r_12_10[47:0]),
     .sp12_v_t(sp12_v_t_12_10[23:0]), .sp4_v_t(sp4_v_t_12_10[47:0]),
     .sp4_r_v_b(sp4_r_v_b_12_10[47:0]), .wl(wl[175:160]),
     .top_op(top_op_12_10[7:0]), .rgt_op(rgt_op_12_10[7:0]),
     .bot_op(slf_op_12_09[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net6474), .purst(purst), .slf_op(slf_op_12_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(rgt_op_12_09[7:0]),
     .bnl_op(net6468[0:7]), .tnr_op(tnr_op_12_10[7:0]),
     .tnl_op(tnl_op_12_10[7:0]));
ltile4rev I_10_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6418), .lft_op(net6300[0:7]),
     .sp12_h_l(net6340[0:23]), .sp4_h_l(net6341[0:47]),
     .sp4_v_b(net6344[0:47]), .sp12_v_b(net7070[0:23]),
     .sp12_h_r(net6424[0:23]), .sp4_h_r(net6425[0:47]),
     .sp12_v_t(net6426[0:23]), .sp4_v_t(net6316[0:47]),
     .sp4_r_v_b(net6428[0:47]), .wl(wl[159:144]),
     .top_op(slf_op_10_10[7:0]), .rgt_op(net6468[0:7]),
     .bot_op(net6356[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net7062), .purst(purst), .slf_op(net6328[0:7]),
     .pgate(pgate[159:144]), .bnr_op(net6440[0:7]),
     .bnl_op(net6272[0:7]), .tnr_op(slf_op_11_10[7:0]),
     .tnl_op(slf_op_09_10[7:0]));
ltile4rev I_10_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_10_10), .lft_op(slf_op_09_10[7:0]),
     .sp12_h_l(net6312[0:23]), .sp4_h_l(net6313[0:47]),
     .sp4_v_b(net6316[0:47]), .sp12_v_b(net6426[0:23]),
     .sp12_h_r(net6452[0:23]), .sp4_h_r(net6453[0:47]),
     .sp12_v_t(sp12_v_t_10_10[23:0]), .sp4_v_t(sp4_v_t_10_10[47:0]),
     .sp4_r_v_b(net6456[0:47]), .wl(wl[175:160]),
     .top_op(top_op_10_10[7:0]), .rgt_op(slf_op_11_10[7:0]),
     .bot_op(net6328[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net6418), .purst(purst), .slf_op(slf_op_10_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(net6468[0:7]),
     .bnl_op(net6300[0:7]), .tnr_op(tnr_op_10_10[7:0]),
     .tnl_op(tnl_op_10_10[7:0]));
ltile4rev I_12_09 ( .vdd_cntl(vdd_cntl[159:144]), .prog(prog),
     .carry_out(net6474), .lft_op(net6468[0:7]),
     .sp12_h_l(net6368[0:23]), .sp4_h_l(net6369[0:47]),
     .sp4_v_b(net6372[0:47]), .sp12_v_b(net7014[0:23]),
     .sp12_h_r(sp12_h_r_12_09[23:0]), .sp4_h_r(sp4_h_r_12_09[47:0]),
     .sp12_v_t(net6482[0:23]), .sp4_v_t(net6512[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_09[47:0]), .wl(wl[159:144]),
     .top_op(slf_op_12_10[7:0]), .rgt_op(rgt_op_12_09[7:0]),
     .bot_op(slf_op_12_08[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[159:144]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net7006), .purst(purst), .slf_op(slf_op_12_09[7:0]),
     .pgate(pgate[159:144]), .bnr_op(rgt_op_12_08[7:0]),
     .bnl_op(net6440[0:7]), .tnr_op(rgt_op_12_10[7:0]),
     .tnl_op(slf_op_11_10[7:0]));
ltile4rev I_11_10 ( .vdd_cntl(vdd_cntl[175:160]), .prog(prog),
     .carry_out(carry_out_11_10), .lft_op(slf_op_10_10[7:0]),
     .sp12_h_l(net6452[0:23]), .sp4_h_l(net6453[0:47]),
     .sp4_v_b(net6456[0:47]), .sp12_v_b(net6370[0:23]),
     .sp12_h_r(net6508[0:23]), .sp4_h_r(net6509[0:47]),
     .sp12_v_t(sp12_v_t_11_10[23:0]), .sp4_v_t(sp4_v_t_11_10[47:0]),
     .sp4_r_v_b(net6512[0:47]), .wl(wl[175:160]),
     .top_op(top_op_11_10[7:0]), .rgt_op(slf_op_12_10[7:0]),
     .bot_op(net6468[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[175:160]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net6362), .purst(purst), .slf_op(slf_op_11_10[7:0]),
     .pgate(pgate[175:160]), .bnr_op(slf_op_12_09[7:0]),
     .bnl_op(net6328[0:7]), .tnr_op(tnr_op_11_10[7:0]),
     .tnl_op(tnl_op_11_10[7:0]));
ltile4rev I_01_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6530), .lft_op({io_l_32[3], io_l_32[2], io_l_32[1],
     io_l_32[0], io_l_32[3], io_l_32[2], io_l_32[1], io_l_32[0]}),
     .sp12_h_l(net4361[0:23]), .sp4_h_l(net4360[0:47]),
     .sp4_v_b(net5559[0:47]), .sp12_v_b(net5558[0:23]),
     .sp12_h_r(net6536[0:23]), .sp4_h_r(net6537[0:47]),
     .sp12_v_t(net6538[0:23]), .sp4_v_t(net6539[0:47]),
     .sp4_r_v_b(net6540[0:47]), .wl(wl[127:112]),
     .top_op(net6542[0:7]), .rgt_op(net6580[0:7]),
     .bot_op(net5590[0:7]), .bl(bl[71:18]), .reset_b(reset_b[127:112]),
     .glb_netwk(glb_netwk_01[7:0]), .carry_in(net5550), .purst(purst),
     .slf_op(net5562[0:7]), .pgate(pgate[127:112]),
     .bnr_op(net6552[0:7]), .bnl_op({io_l_30[3], io_l_30[2],
     io_l_30[1], io_l_30[0], io_l_30[3], io_l_30[2], io_l_30[1],
     io_l_30[0]}), .tnr_op(net6216[0:7]), .tnl_op({io_l_14[3],
     io_l_14[2], io_l_14[1], io_l_14[0], io_l_14[3], io_l_14[2],
     io_l_14[1], io_l_14[0]}));
ltile4rev I_01_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6558), .lft_op({io_l_14[3], io_l_14[2], io_l_14[1],
     io_l_14[0], io_l_14[3], io_l_14[2], io_l_14[1], io_l_14[0]}),
     .sp12_h_l(net4327[0:23]), .sp4_h_l(net4326[0:47]),
     .sp4_v_b(net6539[0:47]), .sp12_v_b(net6538[0:23]),
     .sp12_h_r(net6564[0:23]), .sp4_h_r(net6565[0:47]),
     .sp12_v_t(net6566[0:23]), .sp4_v_t(net6567[0:47]),
     .sp4_r_v_b(net6568[0:47]), .wl(wl[143:128]),
     .top_op(net6570[0:7]), .rgt_op(net6216[0:7]),
     .bot_op(net5562[0:7]), .bl(bl[71:18]), .reset_b(reset_b[143:128]),
     .glb_netwk(glb_netwk_01[7:0]), .carry_in(net6530), .purst(purst),
     .slf_op(net6542[0:7]), .pgate(pgate[143:128]),
     .bnr_op(net6580[0:7]), .bnl_op({io_l_32[3], io_l_32[2],
     io_l_32[1], io_l_32[0], io_l_32[3], io_l_32[2], io_l_32[1],
     io_l_32[0]}), .tnr_op(net6188[0:7]), .tnl_op({io_l_16[3],
     io_l_16[2], io_l_16[1], io_l_16[0], io_l_16[3], io_l_16[2],
     io_l_16[1], io_l_16[0]}));
ltile4rev I_02_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6586), .lft_op(net6542[0:7]),
     .sp12_h_l(net6564[0:23]), .sp4_h_l(net6565[0:47]),
     .sp4_v_b(net6568[0:47]), .sp12_v_b(net6622[0:23]),
     .sp12_h_r(net6592[0:23]), .sp4_h_r(net6593[0:47]),
     .sp12_v_t(net6594[0:23]), .sp4_v_t(net6204[0:47]),
     .sp4_r_v_b(net6596[0:47]), .wl(wl[143:128]),
     .top_op(net6188[0:7]), .rgt_op(net6132[0:7]),
     .bot_op(net6580[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net6614), .purst(purst), .slf_op(net6216[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net6608[0:7]),
     .bnl_op(net5562[0:7]), .tnr_op(net6160[0:7]),
     .tnl_op(net6570[0:7]));
ltile4rev I_02_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6614), .lft_op(net5562[0:7]),
     .sp12_h_l(net6536[0:23]), .sp4_h_l(net6537[0:47]),
     .sp4_v_b(net6540[0:47]), .sp12_v_b(net5530[0:23]),
     .sp12_h_r(net6620[0:23]), .sp4_h_r(net6621[0:47]),
     .sp12_v_t(net6622[0:23]), .sp4_v_t(net6568[0:47]),
     .sp4_r_v_b(net6624[0:47]), .wl(wl[127:112]),
     .top_op(net6216[0:7]), .rgt_op(net6608[0:7]),
     .bot_op(net6552[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net5522), .purst(purst), .slf_op(net6580[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net6636[0:7]),
     .bnl_op(net5590[0:7]), .tnr_op(net6132[0:7]),
     .tnl_op(net6542[0:7]));
ltile4rev I_05_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6642), .lft_op(net6748[0:7]),
     .sp12_h_l(net6788[0:23]), .sp4_h_l(net6789[0:47]),
     .sp4_v_b(net6792[0:47]), .sp12_v_b(net5334[0:23]),
     .sp12_h_r(net6648[0:23]), .sp4_h_r(net6649[0:47]),
     .sp12_v_t(net6650[0:23]), .sp4_v_t(net6764[0:47]),
     .sp4_r_v_b(net6652[0:47]), .wl(wl[127:112]),
     .top_op(net6076[0:7]), .rgt_op(net8047[0:7]),
     .bot_op(net6804[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net5326), .purst(purst), .slf_op(net6776[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net6664[0:7]),
     .bnl_op(net6720[0:7]), .tnr_op(net6666[0:7]),
     .tnl_op(net5992[0:7]));
ltile4rev I_05_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6670), .lft_op(net5992[0:7]),
     .sp12_h_l(net6760[0:23]), .sp4_h_l(net6761[0:47]),
     .sp4_v_b(net6764[0:47]), .sp12_v_b(net6650[0:23]),
     .sp12_h_r(net6676[0:23]), .sp4_h_r(net6677[0:47]),
     .sp12_v_t(net6678[0:23]), .sp4_v_t(net6064[0:47]),
     .sp4_r_v_b(net6680[0:47]), .wl(wl[143:128]),
     .top_op(net6048[0:7]), .rgt_op(net6666[0:7]),
     .bot_op(net6776[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net6642), .purst(purst), .slf_op(net6076[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net8047[0:7]),
     .bnl_op(net6748[0:7]), .tnr_op(net7985[0:7]),
     .tnl_op(net6020[0:7]));
ltile4rev I_03_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6698), .lft_op(net6580[0:7]),
     .sp12_h_l(net6620[0:23]), .sp4_h_l(net6621[0:47]),
     .sp4_v_b(net6624[0:47]), .sp12_v_b(net5390[0:23]),
     .sp12_h_r(net6704[0:23]), .sp4_h_r(net6705[0:47]),
     .sp12_v_t(net6706[0:23]), .sp4_v_t(net6596[0:47]),
     .sp4_r_v_b(net6708[0:47]), .wl(wl[127:112]),
     .top_op(net6132[0:7]), .rgt_op(net6748[0:7]),
     .bot_op(net6636[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net5382), .purst(purst), .slf_op(net6608[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net6720[0:7]),
     .bnl_op(net6552[0:7]), .tnr_op(net5992[0:7]),
     .tnl_op(net6216[0:7]));
ltile4rev I_03_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6726), .lft_op(net6216[0:7]),
     .sp12_h_l(net6592[0:23]), .sp4_h_l(net6593[0:47]),
     .sp4_v_b(net6596[0:47]), .sp12_v_b(net6706[0:23]),
     .sp12_h_r(net6732[0:23]), .sp4_h_r(net6733[0:47]),
     .sp12_v_t(net6734[0:23]), .sp4_v_t(net6120[0:47]),
     .sp4_r_v_b(net6736[0:47]), .wl(wl[143:128]),
     .top_op(net6160[0:7]), .rgt_op(net5992[0:7]),
     .bot_op(net6608[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net6698), .purst(purst), .slf_op(net6132[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net6748[0:7]),
     .bnl_op(net6580[0:7]), .tnr_op(net6020[0:7]),
     .tnl_op(net6188[0:7]));
ltile4rev I_04_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6754), .lft_op(net6132[0:7]),
     .sp12_h_l(net6732[0:23]), .sp4_h_l(net6733[0:47]),
     .sp4_v_b(net6736[0:47]), .sp12_v_b(net6790[0:23]),
     .sp12_h_r(net6760[0:23]), .sp4_h_r(net6761[0:47]),
     .sp12_v_t(net6762[0:23]), .sp4_v_t(net5980[0:47]),
     .sp4_r_v_b(net6764[0:47]), .wl(wl[143:128]),
     .top_op(net6020[0:7]), .rgt_op(net6076[0:7]),
     .bot_op(net6748[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net6782), .purst(purst), .slf_op(net5992[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net6776[0:7]),
     .bnl_op(net6608[0:7]), .tnr_op(net6048[0:7]),
     .tnl_op(net6160[0:7]));
ltile4rev I_04_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6782), .lft_op(net6608[0:7]),
     .sp12_h_l(net6704[0:23]), .sp4_h_l(net6705[0:47]),
     .sp4_v_b(net6708[0:47]), .sp12_v_b(net5418[0:23]),
     .sp12_h_r(net6788[0:23]), .sp4_h_r(net6789[0:47]),
     .sp12_v_t(net6790[0:23]), .sp4_v_t(net6736[0:47]),
     .sp4_r_v_b(net6792[0:47]), .wl(wl[127:112]),
     .top_op(net5992[0:7]), .rgt_op(net6776[0:7]),
     .bot_op(net6720[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net5410), .purst(purst), .slf_op(net6748[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net6804[0:7]),
     .bnl_op(net6636[0:7]), .tnr_op(net6076[0:7]),
     .tnl_op(net6132[0:7]));
ltile4rev I_07_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6810), .lft_op(net6666[0:7]),
     .sp12_h_l(net8032[0:23]), .sp4_h_l(net8035[0:47]),
     .sp4_v_b(net8037[0:47]), .sp12_v_b(net6846[0:23]),
     .sp12_h_r(net6816[0:23]), .sp4_h_r(net6817[0:47]),
     .sp12_v_t(net6818[0:23]), .sp4_v_t(net4820[0:47]),
     .sp4_r_v_b(net6820[0:47]), .wl(wl[143:128]),
     .top_op(net6822[0:7]), .rgt_op(net6878[0:7]),
     .bot_op(net5478[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net6838), .purst(purst), .slf_op(net6850[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net5674[0:7]),
     .bnl_op(net8047[0:7]), .tnr_op(net6906[0:7]),
     .tnl_op(net7985[0:7]));
ltile4rev I_07_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6838), .lft_op(net8047[0:7]),
     .sp12_h_l(net8033[0:23]), .sp4_h_l(net8034[0:47]),
     .sp4_v_b(net8038[0:47]), .sp12_v_b(net5474[0:23]),
     .sp12_h_r(net6844[0:23]), .sp4_h_r(net6845[0:47]),
     .sp12_v_t(net6846[0:23]), .sp4_v_t(net8037[0:47]),
     .sp4_r_v_b(net6848[0:47]), .wl(wl[127:112]),
     .top_op(net6850[0:7]), .rgt_op(net5674[0:7]),
     .bot_op(net5618[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net5466), .purst(purst), .slf_op(net5478[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net5646[0:7]),
     .bnl_op(net6664[0:7]), .tnr_op(net6878[0:7]),
     .tnl_op(net6666[0:7]));
ltile4rev I_08_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6866), .lft_op(net5478[0:7]),
     .sp12_h_l(net6844[0:23]), .sp4_h_l(net6845[0:47]),
     .sp4_v_b(net6848[0:47]), .sp12_v_b(net5670[0:23]),
     .sp12_h_r(net6872[0:23]), .sp4_h_r(net6873[0:47]),
     .sp12_v_t(net6874[0:23]), .sp4_v_t(net6820[0:47]),
     .sp4_r_v_b(net6876[0:47]), .wl(wl[127:112]),
     .top_op(net6878[0:7]), .rgt_op(net6916[0:7]),
     .bot_op(net5646[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net5662), .purst(purst), .slf_op(net5674[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net6888[0:7]),
     .bnl_op(net5618[0:7]), .tnr_op(net6272[0:7]),
     .tnl_op(net6850[0:7]));
ltile4rev I_08_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6894), .lft_op(net6850[0:7]),
     .sp12_h_l(net6816[0:23]), .sp4_h_l(net6817[0:47]),
     .sp4_v_b(net6820[0:47]), .sp12_v_b(net6874[0:23]),
     .sp12_h_r(net6900[0:23]), .sp4_h_r(net6901[0:47]),
     .sp12_v_t(net6902[0:23]), .sp4_v_t(net6232[0:47]),
     .sp4_r_v_b(net6904[0:47]), .wl(wl[143:128]),
     .top_op(net6906[0:7]), .rgt_op(net6272[0:7]),
     .bot_op(net5674[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net6866), .purst(purst), .slf_op(net6878[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net6916[0:7]),
     .bnl_op(net5478[0:7]), .tnr_op(net6300[0:7]),
     .tnl_op(net6822[0:7]));
ltile4rev I_09_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net6922), .lft_op(net6878[0:7]),
     .sp12_h_l(net6900[0:23]), .sp4_h_l(net6901[0:47]),
     .sp4_v_b(net6904[0:47]), .sp12_v_b(net6958[0:23]),
     .sp12_h_r(net6928[0:23]), .sp4_h_r(net6929[0:47]),
     .sp12_v_t(net6930[0:23]), .sp4_v_t(net6260[0:47]),
     .sp4_r_v_b(net6932[0:47]), .wl(wl[143:128]),
     .top_op(net6300[0:7]), .rgt_op(net6356[0:7]),
     .bot_op(net6916[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net6950), .purst(purst), .slf_op(net6272[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net6944[0:7]),
     .bnl_op(net5674[0:7]), .tnr_op(net6328[0:7]),
     .tnl_op(net6906[0:7]));
ltile4rev I_09_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6950), .lft_op(net5674[0:7]),
     .sp12_h_l(net6872[0:23]), .sp4_h_l(net6873[0:47]),
     .sp4_v_b(net6876[0:47]), .sp12_v_b(net5698[0:23]),
     .sp12_h_r(net6956[0:23]), .sp4_h_r(net6957[0:47]),
     .sp12_v_t(net6958[0:23]), .sp4_v_t(net6904[0:47]),
     .sp4_r_v_b(net6960[0:47]), .wl(wl[127:112]),
     .top_op(net6272[0:7]), .rgt_op(net6944[0:7]),
     .bot_op(net6888[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net5690), .purst(purst), .slf_op(net6916[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net6972[0:7]),
     .bnl_op(net5646[0:7]), .tnr_op(net6356[0:7]),
     .tnl_op(net6878[0:7]));
ltile4rev I_11_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net6978), .lft_op(net6944[0:7]),
     .sp12_h_l(net7040[0:23]), .sp4_h_l(net7041[0:47]),
     .sp4_v_b(net7044[0:47]), .sp12_v_b(net5894[0:23]),
     .sp12_h_r(net6984[0:23]), .sp4_h_r(net6985[0:47]),
     .sp12_v_t(net6986[0:23]), .sp4_v_t(net7072[0:47]),
     .sp4_r_v_b(net6988[0:47]), .wl(wl[127:112]),
     .top_op(net6440[0:7]), .rgt_op(slf_op_12_07[7:0]),
     .bot_op(net7056[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net5886), .purst(purst), .slf_op(net7084[0:7]),
     .pgate(pgate[127:112]), .bnr_op(slf_op_12_06[7:0]),
     .bnl_op(net6972[0:7]), .tnr_op(slf_op_12_08[7:0]),
     .tnl_op(net6356[0:7]));
ltile4rev I_12_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net7006), .lft_op(net6440[0:7]),
     .sp12_h_l(net7124[0:23]), .sp4_h_l(net7125[0:47]),
     .sp4_v_b(net7128[0:47]), .sp12_v_b(net7098[0:23]),
     .sp12_h_r(sp12_h_r_12_08[23:0]), .sp4_h_r(sp4_h_r_12_08[47:0]),
     .sp12_v_t(net7014[0:23]), .sp4_v_t(net6372[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_08[47:0]), .wl(wl[143:128]),
     .top_op(slf_op_12_09[7:0]), .rgt_op(rgt_op_12_08[7:0]),
     .bot_op(slf_op_12_07[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net7090), .purst(purst), .slf_op(slf_op_12_08[7:0]),
     .pgate(pgate[143:128]), .bnr_op(rgt_op_12_07[7:0]),
     .bnl_op(net7084[0:7]), .tnr_op(rgt_op_12_09[7:0]),
     .tnl_op(net6468[0:7]));
ltile4rev I_10_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net7034), .lft_op(net6916[0:7]),
     .sp12_h_l(net6956[0:23]), .sp4_h_l(net6957[0:47]),
     .sp4_v_b(net6960[0:47]), .sp12_v_b(net5838[0:23]),
     .sp12_h_r(net7040[0:23]), .sp4_h_r(net7041[0:47]),
     .sp12_v_t(net7042[0:23]), .sp4_v_t(net6932[0:47]),
     .sp4_r_v_b(net7044[0:47]), .wl(wl[127:112]),
     .top_op(net6356[0:7]), .rgt_op(net7084[0:7]),
     .bot_op(net6972[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net5830), .purst(purst), .slf_op(net6944[0:7]),
     .pgate(pgate[127:112]), .bnr_op(net7056[0:7]),
     .bnl_op(net6888[0:7]), .tnr_op(net6440[0:7]),
     .tnl_op(net6272[0:7]));
ltile4rev I_10_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net7062), .lft_op(net6272[0:7]),
     .sp12_h_l(net6928[0:23]), .sp4_h_l(net6929[0:47]),
     .sp4_v_b(net6932[0:47]), .sp12_v_b(net7042[0:23]),
     .sp12_h_r(net7068[0:23]), .sp4_h_r(net7069[0:47]),
     .sp12_v_t(net7070[0:23]), .sp4_v_t(net6344[0:47]),
     .sp4_r_v_b(net7072[0:47]), .wl(wl[143:128]),
     .top_op(net6328[0:7]), .rgt_op(net6440[0:7]),
     .bot_op(net6944[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net7034), .purst(purst), .slf_op(net6356[0:7]),
     .pgate(pgate[143:128]), .bnr_op(net7084[0:7]),
     .bnl_op(net6916[0:7]), .tnr_op(net6468[0:7]),
     .tnl_op(net6300[0:7]));
ltile4rev I_12_07 ( .vdd_cntl(vdd_cntl[127:112]), .prog(prog),
     .carry_out(net7090), .lft_op(net7084[0:7]),
     .sp12_h_l(net6984[0:23]), .sp4_h_l(net6985[0:47]),
     .sp4_v_b(net6988[0:47]), .sp12_v_b(net5782[0:23]),
     .sp12_h_r(sp12_h_r_12_07[23:0]), .sp4_h_r(sp4_h_r_12_07[47:0]),
     .sp12_v_t(net7098[0:23]), .sp4_v_t(net7128[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_07[47:0]), .wl(wl[127:112]),
     .top_op(slf_op_12_08[7:0]), .rgt_op(rgt_op_12_07[7:0]),
     .bot_op(slf_op_12_06[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[127:112]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net7108), .purst(purst), .slf_op(slf_op_12_07[7:0]),
     .pgate(pgate[127:112]), .bnr_op(rgt_op_12_06[7:0]),
     .bnl_op(net7056[0:7]), .tnr_op(rgt_op_12_08[7:0]),
     .tnl_op(net6440[0:7]));
ltile4rev I_11_08 ( .vdd_cntl(vdd_cntl[143:128]), .prog(prog),
     .carry_out(net7118), .lft_op(net6356[0:7]),
     .sp12_h_l(net7068[0:23]), .sp4_h_l(net7069[0:47]),
     .sp4_v_b(net7072[0:47]), .sp12_v_b(net6986[0:23]),
     .sp12_h_r(net7124[0:23]), .sp4_h_r(net7125[0:47]),
     .sp12_v_t(net7126[0:23]), .sp4_v_t(net6428[0:47]),
     .sp4_r_v_b(net7128[0:47]), .wl(wl[143:128]),
     .top_op(net6468[0:7]), .rgt_op(slf_op_12_08[7:0]),
     .bot_op(net7084[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[143:128]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net6978), .purst(purst), .slf_op(net6440[0:7]),
     .pgate(pgate[143:128]), .bnr_op(slf_op_12_07[7:0]),
     .bnl_op(net6944[0:7]), .tnr_op(slf_op_12_09[7:0]),
     .tnl_op(net6328[0:7]));
ltile4rev I_11_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net7146), .lft_op(net5264[0:7]),
     .sp12_h_l(net7208[0:23]), .sp4_h_l(net7209[0:47]),
     .sp4_v_b(net7212[0:47]), .sp12_v_b(net4429[0:23]),
     .sp12_h_r(net7152[0:23]), .sp4_h_r(net7153[0:47]),
     .sp12_v_t(net7154[0:23]), .sp4_v_t(net7240[0:47]),
     .sp4_r_v_b(net7156[0:47]), .wl(wl[31:16]), .top_op(net7868[0:7]),
     .rgt_op(slf_op_12_01[7:0]), .bot_op({io_b_11[3], io_b_11[2],
     io_b_11[1], io_b_11[0], io_b_11[3], io_b_11[2], io_b_11[1],
     io_b_11[0]}), .bl(bl[599:546]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_11[7:0]), .carry_in(net8296), .purst(purst),
     .slf_op(net7252[0:7]), .pgate(pgate[31:16]),
     .bnr_op({slf_op_12_00_clash[3], slf_op_12_00_clash[2],
     slf_op_12_00_clash[1], slf_op_12_00_clash[0],
     slf_op_12_00_clash[3], slf_op_12_00_clash[2],
     slf_op_12_00_clash[1], slf_op_12_00_clash[0]}),
     .bnl_op({io_b_10[3], io_b_10[2], io_b_10[1], io_b_10[0],
     io_b_10[3], io_b_10[2], io_b_10[1], io_b_10[0]}),
     .tnr_op(slf_op_12_02[7:0]), .tnl_op(net7784[0:7]));
ltile4rev I_12_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net7920), .lft_op(net7868[0:7]),
     .sp12_h_l(net7292[0:23]), .sp4_h_l(net7293[0:47]),
     .sp4_v_b(net7296[0:47]), .sp12_v_b(net7266[0:23]),
     .sp12_h_r(sp12_h_r_12_02[23:0]), .sp4_h_r(sp4_h_r_12_02[47:0]),
     .sp12_v_t(net7182[0:23]), .sp4_v_t(net7800[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_02[47:0]), .wl(wl[47:32]),
     .top_op(slf_op_12_03[7:0]), .rgt_op(rgt_op_12_02[7:0]),
     .bot_op(slf_op_12_01[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net7258), .purst(purst), .slf_op(slf_op_12_02[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_12_01[7:0]),
     .bnl_op(net7252[0:7]), .tnr_op(rgt_op_12_03[7:0]),
     .tnl_op(net7896[0:7]));
ltile4rev I_10_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net7202), .lft_op(net5236[0:7]),
     .sp12_h_l(net5276[0:23]), .sp4_h_l(net5277[0:47]),
     .sp4_v_b(net5280[0:47]), .sp12_v_b(net4395[0:23]),
     .sp12_h_r(net7208[0:23]), .sp4_h_r(net7209[0:47]),
     .sp12_v_t(net7210[0:23]), .sp4_v_t(net5252[0:47]),
     .sp4_r_v_b(net7212[0:47]), .wl(wl[31:16]), .top_op(net7784[0:7]),
     .rgt_op(net7252[0:7]), .bot_op({io_b_10[3], io_b_10[2],
     io_b_10[1], io_b_10[0], io_b_10[3], io_b_10[2], io_b_10[1],
     io_b_10[0]}), .bl(bl[545:492]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_10[7:0]), .carry_in(net8297), .purst(purst),
     .slf_op(net5264[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_11[3],
     io_b_11[2], io_b_11[1], io_b_11[0], io_b_11[3], io_b_11[2],
     io_b_11[1], io_b_11[0]}), .bnl_op({io_b_09[3], io_b_09[2],
     io_b_09[1], io_b_09[0], io_b_09[3], io_b_09[2], io_b_09[1],
     io_b_09[0]}), .tnr_op(net7868[0:7]), .tnl_op(net7700[0:7]));
ltile4rev I_10_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net7230), .lft_op(net7700[0:7]),
     .sp12_h_l(net5248[0:23]), .sp4_h_l(net5249[0:47]),
     .sp4_v_b(net5252[0:47]), .sp12_v_b(net7210[0:23]),
     .sp12_h_r(net7236[0:23]), .sp4_h_r(net7237[0:47]),
     .sp12_v_t(net7238[0:23]), .sp4_v_t(net7772[0:47]),
     .sp4_r_v_b(net7240[0:47]), .wl(wl[47:32]), .top_op(net7756[0:7]),
     .rgt_op(net7868[0:7]), .bot_op(net5264[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[47:32]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net7202), .purst(purst), .slf_op(net7784[0:7]),
     .pgate(pgate[47:32]), .bnr_op(net7252[0:7]),
     .bnl_op(net5236[0:7]), .tnr_op(net7896[0:7]),
     .tnl_op(net7728[0:7]));
ltile4rev I_12_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net7258), .lft_op(net7252[0:7]),
     .sp12_h_l(net7152[0:23]), .sp4_h_l(net7153[0:47]),
     .sp4_v_b(net7156[0:47]), .sp12_v_b(net4767[0:23]),
     .sp12_h_r(sp12_h_r_12_01[23:0]), .sp4_h_r(sp4_h_r_12_01[47:0]),
     .sp12_v_t(net7266[0:23]), .sp4_v_t(net7296[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_01[47:0]), .wl(wl[31:16]),
     .top_op(slf_op_12_02[7:0]), .rgt_op(rgt_op_12_01[7:0]),
     .bot_op({slf_op_12_00_clash[3], slf_op_12_00_clash[2],
     slf_op_12_00_clash[1], slf_op_12_00_clash[0],
     slf_op_12_00_clash[3], slf_op_12_00_clash[2],
     slf_op_12_00_clash[1], slf_op_12_00_clash[0]}), .bl(bl[653:600]),
     .reset_b(reset_b[31:16]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net8261), .purst(purst), .slf_op(slf_op_12_01[7:0]),
     .pgate(pgate[31:16]), .bnr_op({bnr_op_12_01[3], bnr_op_12_01[2],
     bnr_op_12_01[1], bnr_op_12_01[0], bnr_op_12_01[3],
     bnr_op_12_01[2], bnr_op_12_01[1], bnr_op_12_01[0]}),
     .bnl_op({io_b_11[3], io_b_11[2], io_b_11[1], io_b_11[0],
     io_b_11[3], io_b_11[2], io_b_11[1], io_b_11[0]}),
     .tnr_op(rgt_op_12_02[7:0]), .tnl_op(net7868[0:7]));
ltile4rev I_11_02 ( .vdd_cntl(vdd_cntl[47:32]), .prog(prog),
     .carry_out(net7286), .lft_op(net7784[0:7]),
     .sp12_h_l(net7236[0:23]), .sp4_h_l(net7237[0:47]),
     .sp4_v_b(net7240[0:47]), .sp12_v_b(net7154[0:23]),
     .sp12_h_r(net7292[0:23]), .sp4_h_r(net7293[0:47]),
     .sp12_v_t(net7294[0:23]), .sp4_v_t(net7856[0:47]),
     .sp4_r_v_b(net7296[0:47]), .wl(wl[47:32]), .top_op(net7896[0:7]),
     .rgt_op(slf_op_12_02[7:0]), .bot_op(net7252[0:7]),
     .bl(bl[599:546]), .reset_b(reset_b[47:32]),
     .glb_netwk(glb_netwk_11[7:0]), .carry_in(net7146), .purst(purst),
     .slf_op(net7868[0:7]), .pgate(pgate[47:32]),
     .bnr_op(slf_op_12_01[7:0]), .bnl_op(net5264[0:7]),
     .tnr_op(slf_op_12_03[7:0]), .tnl_op(net7756[0:7]));
ltile4rev I_02_01 ( .vdd_cntl(vdd_cntl[31:16]), .prog(prog),
     .carry_out(net7314), .lft_op(net4671[0:7]),
     .sp12_h_l(net5136[0:23]), .sp4_h_l(net5137[0:47]),
     .sp4_v_b(net5140[0:47]), .sp12_v_b(net4633[0:23]),
     .sp12_h_r(net7320[0:23]), .sp4_h_r(net7321[0:47]),
     .sp12_v_t(net7322[0:23]), .sp4_v_t(net5112[0:47]),
     .sp4_r_v_b(net7324[0:47]), .wl(wl[31:16]), .top_op(net7364[0:7]),
     .rgt_op(net5096[0:7]), .bot_op({io_b_02[3], io_b_02[2],
     io_b_02[1], io_b_02[0], io_b_02[3], io_b_02[2], io_b_02[1],
     io_b_02[0]}), .bl(bl[125:72]), .reset_b(reset_b[31:16]),
     .glb_netwk(glb_netwk_02[7:0]), .carry_in(net8287), .purst(purst),
     .slf_op(net5124[0:7]), .pgate(pgate[31:16]), .bnr_op({io_b_03[3],
     io_b_03[2], io_b_03[1], io_b_03[0], io_b_03[3], io_b_03[2],
     io_b_03[1], io_b_03[0]}), .bnl_op({io_b_01[3], io_b_01[2],
     io_b_01[1], io_b_01[0], io_b_01[3], io_b_01[2], io_b_01[1],
     io_b_01[0]}), .tnr_op(net7448[0:7]), .tnl_op(net5142[0:7]));
ltile4rev I_01_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7342), .lft_op({io_l_24[3], io_l_24[2], io_l_24[1],
     io_l_24[0], io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0]}),
     .sp12_h_l(net4293[0:23]), .sp4_h_l(net4292[0:47]),
     .sp4_v_b(net5111[0:47]), .sp12_v_b(net5110[0:23]),
     .sp12_h_r(net7348[0:23]), .sp4_h_r(net7349[0:47]),
     .sp12_v_t(net7350[0:23]), .sp4_v_t(net7351[0:47]),
     .sp4_r_v_b(net7352[0:47]), .wl(wl[63:48]), .top_op(net5592[0:7]),
     .rgt_op(net7392[0:7]), .bot_op(net5142[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net5102), .purst(purst), .slf_op(net5114[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net7364[0:7]), .bnl_op({io_l_22[3],
     io_l_22[2], io_l_22[1], io_l_22[0], io_l_22[3], io_l_22[2],
     io_l_22[1], io_l_22[0]}), .tnr_op(net5600[0:7]),
     .tnl_op({io_l_26[3], io_l_26[2], io_l_26[1], io_l_26[0],
     io_l_26[3], io_l_26[2], io_l_26[1], io_l_26[0]}));
ltile4rev I_01_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7370), .lft_op({io_l_26[3], io_l_26[2], io_l_26[1],
     io_l_26[0], io_l_26[3], io_l_26[2], io_l_26[1], io_l_26[0]}),
     .sp12_h_l(net4259[0:23]), .sp4_h_l(net4258[0:47]),
     .sp4_v_b(net7351[0:47]), .sp12_v_b(net7350[0:23]),
     .sp12_h_r(net7376[0:23]), .sp4_h_r(net7377[0:47]),
     .sp12_v_t(net7378[0:23]), .sp4_v_t(net7379[0:47]),
     .sp4_r_v_b(net7380[0:47]), .wl(wl[79:64]), .top_op(net4161[0:7]),
     .rgt_op(net5600[0:7]), .bot_op(net5114[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net7342), .purst(purst), .slf_op(net5592[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net7392[0:7]), .bnl_op({io_l_24[3],
     io_l_24[2], io_l_24[1], io_l_24[0], io_l_24[3], io_l_24[2],
     io_l_24[1], io_l_24[0]}), .tnr_op(net5572[0:7]),
     .tnl_op({io_l_28[3], io_l_28[2], io_l_28[1], io_l_28[0],
     io_l_28[3], io_l_28[2], io_l_28[1], io_l_28[0]}));
ltile4rev I_02_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7398), .lft_op(net5592[0:7]),
     .sp12_h_l(net7376[0:23]), .sp4_h_l(net7377[0:47]),
     .sp4_v_b(net7380[0:47]), .sp12_v_b(net7434[0:23]),
     .sp12_h_r(net7404[0:23]), .sp4_h_r(net7405[0:47]),
     .sp12_v_t(net7406[0:23]), .sp4_v_t(net5588[0:47]),
     .sp4_r_v_b(net7408[0:47]), .wl(wl[79:64]), .top_op(net5572[0:7]),
     .rgt_op(net5516[0:7]), .bot_op(net7392[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net7426), .purst(purst), .slf_op(net5600[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net7420[0:7]),
     .bnl_op(net5114[0:7]), .tnr_op(net5544[0:7]),
     .tnl_op(net4161[0:7]));
ltile4rev I_02_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7426), .lft_op(net5114[0:7]),
     .sp12_h_l(net7348[0:23]), .sp4_h_l(net7349[0:47]),
     .sp4_v_b(net7352[0:47]), .sp12_v_b(net5082[0:23]),
     .sp12_h_r(net7432[0:23]), .sp4_h_r(net7433[0:47]),
     .sp12_v_t(net7434[0:23]), .sp4_v_t(net7380[0:47]),
     .sp4_r_v_b(net7436[0:47]), .wl(wl[63:48]), .top_op(net5600[0:7]),
     .rgt_op(net7420[0:7]), .bot_op(net7364[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net5074), .purst(purst), .slf_op(net7392[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net7448[0:7]),
     .bnl_op(net5142[0:7]), .tnr_op(net5516[0:7]),
     .tnl_op(net5592[0:7]));
ltile4rev I_05_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7454), .lft_op(net7560[0:7]),
     .sp12_h_l(net7600[0:23]), .sp4_h_l(net7601[0:47]),
     .sp4_v_b(net7604[0:47]), .sp12_v_b(net4914[0:23]),
     .sp12_h_r(net7460[0:23]), .sp4_h_r(net7461[0:47]),
     .sp12_v_t(net7462[0:23]), .sp4_v_t(net7576[0:47]),
     .sp4_r_v_b(net7464[0:47]), .wl(wl[63:48]), .top_op(net5460[0:7]),
     .rgt_op(net8171[0:7]), .bot_op(net7616[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net4906), .purst(purst), .slf_op(net7588[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net4902[0:7]),
     .bnl_op(net7532[0:7]), .tnr_op(net7478[0:7]),
     .tnl_op(net5376[0:7]));
ltile4rev I_05_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7482), .lft_op(net5376[0:7]),
     .sp12_h_l(net7572[0:23]), .sp4_h_l(net7573[0:47]),
     .sp4_v_b(net7576[0:47]), .sp12_v_b(net7462[0:23]),
     .sp12_h_r(net7488[0:23]), .sp4_h_r(net7489[0:47]),
     .sp12_v_t(net7490[0:23]), .sp4_v_t(net5448[0:47]),
     .sp4_r_v_b(net7492[0:47]), .wl(wl[79:64]), .top_op(net5432[0:7]),
     .rgt_op(net7478[0:7]), .bot_op(net7588[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_05[7:0]),
     .carry_in(net7454), .purst(purst), .slf_op(net5460[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net8171[0:7]),
     .bnl_op(net7560[0:7]), .tnr_op(net8121[0:7]),
     .tnl_op(net5404[0:7]));
ltile4rev I_03_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7510), .lft_op(net7392[0:7]),
     .sp12_h_l(net7432[0:23]), .sp4_h_l(net7433[0:47]),
     .sp4_v_b(net7436[0:47]), .sp12_v_b(net4970[0:23]),
     .sp12_h_r(net7516[0:23]), .sp4_h_r(net7517[0:47]),
     .sp12_v_t(net7518[0:23]), .sp4_v_t(net7408[0:47]),
     .sp4_r_v_b(net7520[0:47]), .wl(wl[63:48]), .top_op(net5516[0:7]),
     .rgt_op(net7560[0:7]), .bot_op(net7448[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net4962), .purst(purst), .slf_op(net7420[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net7532[0:7]),
     .bnl_op(net7364[0:7]), .tnr_op(net5376[0:7]),
     .tnl_op(net5600[0:7]));
ltile4rev I_03_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7538), .lft_op(net5600[0:7]),
     .sp12_h_l(net7404[0:23]), .sp4_h_l(net7405[0:47]),
     .sp4_v_b(net7408[0:47]), .sp12_v_b(net7518[0:23]),
     .sp12_h_r(net7544[0:23]), .sp4_h_r(net7545[0:47]),
     .sp12_v_t(net7546[0:23]), .sp4_v_t(net5504[0:47]),
     .sp4_r_v_b(net7548[0:47]), .wl(wl[79:64]), .top_op(net5544[0:7]),
     .rgt_op(net5376[0:7]), .bot_op(net7420[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net7510), .purst(purst), .slf_op(net5516[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net7560[0:7]),
     .bnl_op(net7392[0:7]), .tnr_op(net5404[0:7]),
     .tnl_op(net5572[0:7]));
ltile4rev I_04_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7566), .lft_op(net5516[0:7]),
     .sp12_h_l(net7544[0:23]), .sp4_h_l(net7545[0:47]),
     .sp4_v_b(net7548[0:47]), .sp12_v_b(net7602[0:23]),
     .sp12_h_r(net7572[0:23]), .sp4_h_r(net7573[0:47]),
     .sp12_v_t(net7574[0:23]), .sp4_v_t(net5364[0:47]),
     .sp4_r_v_b(net7576[0:47]), .wl(wl[79:64]), .top_op(net5404[0:7]),
     .rgt_op(net5460[0:7]), .bot_op(net7560[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net7594), .purst(purst), .slf_op(net5376[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net7588[0:7]),
     .bnl_op(net7420[0:7]), .tnr_op(net5432[0:7]),
     .tnl_op(net5544[0:7]));
ltile4rev I_04_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7594), .lft_op(net7420[0:7]),
     .sp12_h_l(net7516[0:23]), .sp4_h_l(net7517[0:47]),
     .sp4_v_b(net7520[0:47]), .sp12_v_b(net4998[0:23]),
     .sp12_h_r(net7600[0:23]), .sp4_h_r(net7601[0:47]),
     .sp12_v_t(net7602[0:23]), .sp4_v_t(net7548[0:47]),
     .sp4_r_v_b(net7604[0:47]), .wl(wl[63:48]), .top_op(net5376[0:7]),
     .rgt_op(net7588[0:7]), .bot_op(net7532[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net4990), .purst(purst), .slf_op(net7560[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net7616[0:7]),
     .bnl_op(net7448[0:7]), .tnr_op(net5460[0:7]),
     .tnl_op(net5516[0:7]));
ltile4rev I_07_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7622), .lft_op(net7478[0:7]),
     .sp12_h_l(net8109[0:23]), .sp4_h_l(net8112[0:47]),
     .sp4_v_b(net8114[0:47]), .sp12_v_b(net7658[0:23]),
     .sp12_h_r(net7628[0:23]), .sp4_h_r(net7629[0:47]),
     .sp12_v_t(net7630[0:23]), .sp4_v_t(net8078[0:47]),
     .sp4_r_v_b(net7632[0:47]), .wl(wl[79:64]), .top_op(net7634[0:7]),
     .rgt_op(net5648[0:7]), .bot_op(net5058[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net7650), .purst(purst), .slf_op(net7662[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net5226[0:7]),
     .bnl_op(net8171[0:7]), .tnr_op(net5488[0:7]),
     .tnl_op(net8121[0:7]));
ltile4rev I_07_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7650), .lft_op(net8171[0:7]),
     .sp12_h_l(net8110[0:23]), .sp4_h_l(net8111[0:47]),
     .sp4_v_b(net8115[0:47]), .sp12_v_b(net5054[0:23]),
     .sp12_h_r(net7656[0:23]), .sp4_h_r(net7657[0:47]),
     .sp12_v_t(net7658[0:23]), .sp4_v_t(net8114[0:47]),
     .sp4_r_v_b(net7660[0:47]), .wl(wl[63:48]), .top_op(net7662[0:7]),
     .rgt_op(net5226[0:7]), .bot_op(net5170[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net5046), .purst(purst), .slf_op(net5058[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net5198[0:7]),
     .bnl_op(net4902[0:7]), .tnr_op(net5648[0:7]),
     .tnl_op(net7478[0:7]));
ltile4rev I_08_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7678), .lft_op(net5058[0:7]),
     .sp12_h_l(net7656[0:23]), .sp4_h_l(net7657[0:47]),
     .sp4_v_b(net7660[0:47]), .sp12_v_b(net5222[0:23]),
     .sp12_h_r(net7684[0:23]), .sp4_h_r(net7685[0:47]),
     .sp12_v_t(net7686[0:23]), .sp4_v_t(net7632[0:47]),
     .sp4_r_v_b(net7688[0:47]), .wl(wl[63:48]), .top_op(net5648[0:7]),
     .rgt_op(net7728[0:7]), .bot_op(net5198[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net5214), .purst(purst), .slf_op(net5226[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net7700[0:7]),
     .bnl_op(net5170[0:7]), .tnr_op(net5656[0:7]),
     .tnl_op(net7662[0:7]));
ltile4rev I_08_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7706), .lft_op(net7662[0:7]),
     .sp12_h_l(net7628[0:23]), .sp4_h_l(net7629[0:47]),
     .sp4_v_b(net7632[0:47]), .sp12_v_b(net7686[0:23]),
     .sp12_h_r(net7712[0:23]), .sp4_h_r(net7713[0:47]),
     .sp12_v_t(net7714[0:23]), .sp4_v_t(net5616[0:47]),
     .sp4_r_v_b(net7716[0:47]), .wl(wl[79:64]), .top_op(net5488[0:7]),
     .rgt_op(net5656[0:7]), .bot_op(net5226[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net7678), .purst(purst), .slf_op(net5648[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net7728[0:7]),
     .bnl_op(net5058[0:7]), .tnr_op(net5684[0:7]),
     .tnl_op(net7634[0:7]));
ltile4rev I_09_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7734), .lft_op(net5648[0:7]),
     .sp12_h_l(net7712[0:23]), .sp4_h_l(net7713[0:47]),
     .sp4_v_b(net7716[0:47]), .sp12_v_b(net7770[0:23]),
     .sp12_h_r(net7740[0:23]), .sp4_h_r(net7741[0:47]),
     .sp12_v_t(net7742[0:23]), .sp4_v_t(net5644[0:47]),
     .sp4_r_v_b(net7744[0:47]), .wl(wl[79:64]), .top_op(net5684[0:7]),
     .rgt_op(net5740[0:7]), .bot_op(net7728[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net7762), .purst(purst), .slf_op(net5656[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net7756[0:7]),
     .bnl_op(net5226[0:7]), .tnr_op(net5712[0:7]),
     .tnl_op(net5488[0:7]));
ltile4rev I_09_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7762), .lft_op(net5226[0:7]),
     .sp12_h_l(net7684[0:23]), .sp4_h_l(net7685[0:47]),
     .sp4_v_b(net7688[0:47]), .sp12_v_b(net5250[0:23]),
     .sp12_h_r(net7768[0:23]), .sp4_h_r(net7769[0:47]),
     .sp12_v_t(net7770[0:23]), .sp4_v_t(net7716[0:47]),
     .sp4_r_v_b(net7772[0:47]), .wl(wl[63:48]), .top_op(net5656[0:7]),
     .rgt_op(net7756[0:7]), .bot_op(net7700[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net5242), .purst(purst), .slf_op(net7728[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net7784[0:7]),
     .bnl_op(net5198[0:7]), .tnr_op(net5740[0:7]),
     .tnl_op(net5648[0:7]));
ltile4rev I_11_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7790), .lft_op(net7756[0:7]),
     .sp12_h_l(net7852[0:23]), .sp4_h_l(net7853[0:47]),
     .sp4_v_b(net7856[0:47]), .sp12_v_b(net7294[0:23]),
     .sp12_h_r(net7796[0:23]), .sp4_h_r(net7797[0:47]),
     .sp12_v_t(net7798[0:23]), .sp4_v_t(net7884[0:47]),
     .sp4_r_v_b(net7800[0:47]), .wl(wl[63:48]), .top_op(net5824[0:7]),
     .rgt_op(slf_op_12_03[7:0]), .bot_op(net7868[0:7]),
     .bl(bl[599:546]), .reset_b(reset_b[63:48]),
     .glb_netwk(glb_netwk_11[7:0]), .carry_in(net7286), .purst(purst),
     .slf_op(net7896[0:7]), .pgate(pgate[63:48]),
     .bnr_op(slf_op_12_02[7:0]), .bnl_op(net7784[0:7]),
     .tnr_op(slf_op_12_04[7:0]), .tnl_op(net5740[0:7]));
ltile4rev I_12_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7818), .lft_op(net5824[0:7]),
     .sp12_h_l(net7936[0:23]), .sp4_h_l(net7937[0:47]),
     .sp4_v_b(net7940[0:47]), .sp12_v_b(net7910[0:23]),
     .sp12_h_r(sp12_h_r_12_04[23:0]), .sp4_h_r(sp4_h_r_12_04[47:0]),
     .sp12_v_t(net7826[0:23]), .sp4_v_t(net5756[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_04[47:0]), .wl(wl[79:64]),
     .top_op(slf_op_12_05[7:0]), .rgt_op(rgt_op_12_04[7:0]),
     .bot_op(slf_op_12_03[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net7902), .purst(purst), .slf_op(slf_op_12_04[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_12_03[7:0]),
     .bnl_op(net7896[0:7]), .tnr_op(rgt_op_12_05[7:0]),
     .tnl_op(net5852[0:7]));
ltile4rev I_10_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7846), .lft_op(net7728[0:7]),
     .sp12_h_l(net7768[0:23]), .sp4_h_l(net7769[0:47]),
     .sp4_v_b(net7772[0:47]), .sp12_v_b(net7238[0:23]),
     .sp12_h_r(net7852[0:23]), .sp4_h_r(net7853[0:47]),
     .sp12_v_t(net7854[0:23]), .sp4_v_t(net7744[0:47]),
     .sp4_r_v_b(net7856[0:47]), .wl(wl[63:48]), .top_op(net5740[0:7]),
     .rgt_op(net7896[0:7]), .bot_op(net7784[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net7230), .purst(purst), .slf_op(net7756[0:7]),
     .pgate(pgate[63:48]), .bnr_op(net7868[0:7]),
     .bnl_op(net7700[0:7]), .tnr_op(net5824[0:7]),
     .tnl_op(net5656[0:7]));
ltile4rev I_10_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7874), .lft_op(net5656[0:7]),
     .sp12_h_l(net7740[0:23]), .sp4_h_l(net7741[0:47]),
     .sp4_v_b(net7744[0:47]), .sp12_v_b(net7854[0:23]),
     .sp12_h_r(net7880[0:23]), .sp4_h_r(net7881[0:47]),
     .sp12_v_t(net7882[0:23]), .sp4_v_t(net5728[0:47]),
     .sp4_r_v_b(net7884[0:47]), .wl(wl[79:64]), .top_op(net5712[0:7]),
     .rgt_op(net5824[0:7]), .bot_op(net7756[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[79:64]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net7846), .purst(purst), .slf_op(net5740[0:7]),
     .pgate(pgate[79:64]), .bnr_op(net7896[0:7]),
     .bnl_op(net7728[0:7]), .tnr_op(net5852[0:7]),
     .tnl_op(net5684[0:7]));
ltile4rev I_12_03 ( .vdd_cntl(vdd_cntl[63:48]), .prog(prog),
     .carry_out(net7902), .lft_op(net7896[0:7]),
     .sp12_h_l(net7796[0:23]), .sp4_h_l(net7797[0:47]),
     .sp4_v_b(net7800[0:47]), .sp12_v_b(net7182[0:23]),
     .sp12_h_r(sp12_h_r_12_03[23:0]), .sp4_h_r(sp4_h_r_12_03[47:0]),
     .sp12_v_t(net7910[0:23]), .sp4_v_t(net7940[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_03[47:0]), .wl(wl[63:48]),
     .top_op(slf_op_12_04[7:0]), .rgt_op(rgt_op_12_03[7:0]),
     .bot_op(slf_op_12_02[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[63:48]), .glb_netwk(glb_netwk_12[7:0]),
     .carry_in(net7920), .purst(purst), .slf_op(slf_op_12_03[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_12_02[7:0]),
     .bnl_op(net7868[0:7]), .tnr_op(rgt_op_12_04[7:0]),
     .tnl_op(net5824[0:7]));
ltile4rev I_11_04 ( .vdd_cntl(vdd_cntl[79:64]), .prog(prog),
     .carry_out(net7930), .lft_op(net5740[0:7]),
     .sp12_h_l(net7880[0:23]), .sp4_h_l(net7881[0:47]),
     .sp4_v_b(net7884[0:47]), .sp12_v_b(net7798[0:23]),
     .sp12_h_r(net7936[0:23]), .sp4_h_r(net7937[0:47]),
     .sp12_v_t(net7938[0:23]), .sp4_v_t(net5812[0:47]),
     .sp4_r_v_b(net7940[0:47]), .wl(wl[79:64]), .top_op(net5852[0:7]),
     .rgt_op(slf_op_12_04[7:0]), .bot_op(net7896[0:7]),
     .bl(bl[599:546]), .reset_b(reset_b[79:64]),
     .glb_netwk(glb_netwk_11[7:0]), .carry_in(net7790), .purst(purst),
     .slf_op(net5824[0:7]), .pgate(pgate[79:64]),
     .bnr_op(slf_op_12_03[7:0]), .bnl_op(net7756[0:7]),
     .tnr_op(slf_op_12_05[7:0]), .tnl_op(net5712[0:7]));
inv_hvt I1017 ( .A(net7959), .Y(padin_93));
inv_hvt I1018 ( .A(padin_b[23]), .Y(net7959));
inv_hvt I1015 ( .A(net7960), .Y(net7966));
inv_hvt I1014 ( .A(net7962), .Y(fabric_out_34));
inv_hvt I1021 ( .A(net7971), .Y(fabric_out_93));
inv_hvt I1016 ( .A(net7966), .Y(fabric_out_38));
inv_hvt I1019 ( .A(net7968), .Y(padin_34));
inv_hvt I1022 ( .A(net4781), .Y(net7971));
inv_hvt I1020 ( .A(padin_l[19]), .Y(net7968));
inv_hvt I1013 ( .A(net7974), .Y(net7962));
clk_quad_bufx8 I_quad_driver ( .clko(net7976[0:7]),
     .clki(glb_in[7:0]));
bram_4kprouting_bbank I_bram0607 ( .glb_netwk(glb_netwk_06[7:0]),
     .vdd_cntl_top(vdd_cntl[143:128]),
     .vdd_cntl_bot(vdd_cntl[127:112]), .slf_op_top(net6666[0:7]),
     .slf_op_bot(net8047[0:7]), .wl_top(wl[143:128]),
     .wl_bot(wl[127:112]), .top_op_top(net7985[0:7]),
     .tnl_op_top(net6048[0:7]), .tnl_op_bot(net6076[0:7]),
     .reset_b_top(reset_b[143:128]), .reset_b_bot(reset_b[127:112]),
     .prog(prog), .pgate_top(pgate[143:128]),
     .pgate_bot(pgate[127:112]), .lft_op_top(net6076[0:7]),
     .lft_op_bot(net6776[0:7]), .bm_wdummymux_en_i(net8098),
     .bot_op_bot(net6664[0:7]), .bnl_op_top(net6776[0:7]),
     .bnl_op_bot(net6804[0:7]), .sp12_v_t_top(net7999[0:23]),
     .sp12_v_b_bot(net8067[0:23]), .bm_init_i(net8093),
     .sp12_h_l_top(net6676[0:23]), .sp12_h_l_bot(net6648[0:23]),
     .sp4_v_t_top(net5924[0:47]), .sp4_v_b_top(net6680[0:47]),
     .sp4_v_b_bot(net6652[0:47]), .sp4_h_l_top(net6677[0:47]),
     .sp4_h_l_bot(net6649[0:47]), .bm_sdi_o(net8009[0:1]),
     .bm_sclkrw_o(net8010[0:1]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(net8092), .bm_sa_i(net8094[0:7]),
     .bm_sclk_i(net8095), .bm_sclkrw_i(net8084[0:1]),
     .bm_sreb_i(net8096), .bm_sweb_i(net8097[0:1]),
     .bm_rcapmux_en_o(net8018), .bm_init_o(net8019),
     .bm_sa_o(net8020[0:7]), .bm_sclk_o(net8021), .bm_sreb_o(net8022),
     .bm_sweb_o(net8023[0:1]), .bm_wdummymux_en_o(net8024),
     .bm_sdi_i(net8083[0:1]), .bm_sdo_i(net8026[0:1]),
     .bm_sdo_o(net8100[0:1]), .bnr_op_top(net5478[0:7]),
     .rgt_op_top(net6850[0:7]), .tnr_op_top(net6822[0:7]),
     .tnr_op_bot(net6850[0:7]), .sp12_h_r_top(net8032[0:23]),
     .sp12_h_r_bot(net8033[0:23]), .sp4_h_r_bot(net8034[0:47]),
     .sp4_h_r_top(net8035[0:47]), .rgt_op_bot(net5478[0:7]),
     .sp4_r_v_b_top(net8037[0:47]), .sp4_r_v_b_bot(net8038[0:47]),
     .bnr_op_bot(net5618[0:7]));
bram_4kprouting_bbank I_bram_0605 ( .glb_netwk(glb_netwk_06[7:0]),
     .vdd_cntl_bot(vdd_cntl[95:80]), .vdd_cntl_top(vdd_cntl[111:96]),
     .slf_op_top(net6664[0:7]), .slf_op_bot(net8121[0:7]),
     .wl_top(wl[111:96]), .wl_bot(wl[95:80]),
     .top_op_top(net8047[0:7]), .tnr_op_top(net5478[0:7]),
     .tnr_op_bot(net5618[0:7]), .tnl_op_top(net6776[0:7]),
     .tnl_op_bot(net6804[0:7]), .rgt_op_top(net5618[0:7]),
     .rgt_op_bot(net7634[0:7]), .reset_b_top(reset_b[111:96]),
     .reset_b_bot(reset_b[95:80]), .prog(prog),
     .pgate_top(pgate[111:96]), .pgate_bot(pgate[95:80]),
     .lft_op_top(net6804[0:7]), .lft_op_bot(net5432[0:7]),
     .bm_wdummymux_en_i(net8160), .bot_op_bot(net7478[0:7]),
     .bnr_op_top(net7634[0:7]), .bnr_op_bot(net7662[0:7]),
     .bnl_op_top(net5432[0:7]), .bnl_op_bot(net5460[0:7]),
     .sp12_v_t_top(net8067[0:23]), .sp12_v_b_bot(net8135[0:23]),
     .bm_init_i(net8155), .sp12_h_r_top(net8070[0:23]),
     .sp12_h_r_bot(net8071[0:23]), .sp12_h_l_top(net5332[0:23]),
     .sp12_h_l_bot(net5304[0:23]), .sp4_v_t_top(net6652[0:47]),
     .sp4_v_b_top(net5336[0:47]), .sp4_v_b_bot(net5308[0:47]),
     .sp4_r_v_b_top(net8077[0:47]), .sp4_r_v_b_bot(net8078[0:47]),
     .sp4_h_r_top(net8079[0:47]), .sp4_h_r_bot(net8080[0:47]),
     .sp4_h_l_top(net5333[0:47]), .sp4_h_l_bot(net5305[0:47]),
     .bm_sdi_o(net8083[0:1]), .bm_sclkrw_o(net8084[0:1]),
     .bl(bl[329:288]), .bm_rcapmux_en_i(net8154),
     .bm_sa_i(net8156[0:7]), .bm_sclk_i(net8157),
     .bm_sclkrw_i(net8146[0:1]), .bm_sreb_i(net8158),
     .bm_sweb_i(net8159[0:1]), .bm_rcapmux_en_o(net8092),
     .bm_init_o(net8093), .bm_sa_o(net8094[0:7]), .bm_sclk_o(net8095),
     .bm_sreb_o(net8096), .bm_sweb_o(net8097[0:1]),
     .bm_wdummymux_en_o(net8098), .bm_sdi_i(net8145[0:1]),
     .bm_sdo_i(net8100[0:1]), .bm_sdo_o(net8162[0:1]));
bram_4kprouting_bbank I_bram0603 ( .glb_netwk(glb_netwk_06[7:0]),
     .vdd_cntl_top(vdd_cntl[79:64]), .vdd_cntl_bot(vdd_cntl[63:48]),
     .bnr_op_top(net5058[0:7]), .rgt_op_top(net7662[0:7]),
     .tnr_op_top(net7634[0:7]), .tnr_op_bot(net7662[0:7]),
     .sp12_h_r_top(net8109[0:23]), .sp12_h_r_bot(net8110[0:23]),
     .sp4_h_r_bot(net8111[0:47]), .sp4_h_r_top(net8112[0:47]),
     .rgt_op_bot(net5058[0:7]), .sp4_r_v_b_top(net8114[0:47]),
     .sp4_r_v_b_bot(net8115[0:47]), .bnr_op_bot(net5170[0:7]),
     .slf_op_top(net7478[0:7]), .slf_op_bot(net8171[0:7]),
     .wl_top(wl[79:64]), .wl_bot(wl[63:48]), .top_op_top(net8121[0:7]),
     .tnl_op_top(net5432[0:7]), .tnl_op_bot(net5460[0:7]),
     .reset_b_top(reset_b[79:64]), .reset_b_bot(reset_b[63:48]),
     .prog(prog), .pgate_top(pgate[79:64]), .pgate_bot(pgate[63:48]),
     .lft_op_top(net5460[0:7]), .lft_op_bot(net7588[0:7]),
     .bm_wdummymux_en_i(net8222), .bot_op_bot(net4902[0:7]),
     .bnl_op_top(net7588[0:7]), .bnl_op_bot(net7616[0:7]),
     .sp12_v_t_top(net8135[0:23]), .sp12_v_b_bot(net8191[0:23]),
     .bm_init_i(net8217), .sp12_h_l_top(net7488[0:23]),
     .sp12_h_l_bot(net7460[0:23]), .sp4_v_t_top(net5308[0:47]),
     .sp4_v_b_top(net7492[0:47]), .sp4_v_b_bot(net7464[0:47]),
     .sp4_h_l_top(net7489[0:47]), .sp4_h_l_bot(net7461[0:47]),
     .bm_sdi_o(net8145[0:1]), .bm_sclkrw_o(net8146[0:1]),
     .bl(bl[329:288]), .bm_rcapmux_en_i(net8216),
     .bm_sa_i(net8218[0:7]), .bm_sclk_i(net8219),
     .bm_sclkrw_i(net8208[0:1]), .bm_sreb_i(net8220),
     .bm_sweb_i(net8221[0:1]), .bm_rcapmux_en_o(net8154),
     .bm_init_o(net8155), .bm_sa_o(net8156[0:7]), .bm_sclk_o(net8157),
     .bm_sreb_o(net8158), .bm_sweb_o(net8159[0:1]),
     .bm_wdummymux_en_o(net8160), .bm_sdi_i(net8207[0:1]),
     .bm_sdo_i(net8162[0:1]), .bm_sdo_o(net8224[0:1]));
bram_4kprouting_bbankout I_bram0601 ( .glb_netwk(glb_netwk_06[7:0]),
     .vdd_cntl_bot(vdd_cntl[31:16]), .vdd_cntl_top(vdd_cntl[47:32]),
     .slf_op_top(net4902[0:7]), .slf_op_bot(net4536[0:7]),
     .wl_top(wl[47:32]), .wl_bot(wl[31:16]), .top_op_top(net8171[0:7]),
     .tnr_op_top(net5058[0:7]), .tnr_op_bot(net5170[0:7]),
     .tnl_op_top(net7588[0:7]), .tnl_op_bot(net7616[0:7]),
     .rgt_op_top(net5170[0:7]), .rgt_op_bot(net4502[0:7]),
     .reset_b_top(reset_b[47:32]), .reset_b_bot(reset_b[31:16]),
     .prog(prog), .pgate_top(pgate[47:32]), .pgate_bot(pgate[31:16]),
     .lft_op_top(net7616[0:7]), .lft_op_bot(net5012[0:7]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bot_op_bot({io_b_06[3],
     io_b_06[2], io_b_06[1], io_b_06[0], io_b_06[3], io_b_06[2],
     io_b_06[1], io_b_06[0]}), .bnr_op_top(net4502[0:7]),
     .bnr_op_bot({io_b_07[3], io_b_07[2], io_b_07[1], io_b_07[0],
     io_b_07[3], io_b_07[2], io_b_07[1], io_b_07[0]}),
     .bnl_op_top(net5012[0:7]), .bnl_op_bot({io_b_05[3], io_b_05[2],
     io_b_05[1], io_b_05[0], io_b_05[3], io_b_05[2], io_b_05[1],
     io_b_05[0]}), .sp12_v_t_top(net8191[0:23]),
     .sp12_v_b_bot(net4497[0:23]), .bm_init_i(bm_init_i),
     .sp12_h_r_top(net8194[0:23]), .sp12_h_r_bot(net8195[0:23]),
     .sp12_h_l_top(net4912[0:23]), .sp12_h_l_bot(net4884[0:23]),
     .sp4_v_t_top(net7464[0:47]), .sp4_v_b_top(net4916[0:47]),
     .sp4_v_b_bot(net4888[0:47]), .sp4_r_v_b_top(net8201[0:47]),
     .sp4_r_v_b_bot(net8202[0:47]), .sp4_h_r_top(net8203[0:47]),
     .sp4_h_r_bot(net8204[0:47]), .sp4_h_l_top(net4913[0:47]),
     .sp4_h_l_bot(net4885[0:47]), .bm_sdi_o(net8207[0:1]),
     .bm_sclkrw_o(net8208[0:1]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i[1:0]),
     .bm_rcapmux_en_o(net8216), .bm_init_o(net8217),
     .bm_sa_o(net8218[0:7]), .bm_sclk_o(net8219), .bm_sreb_o(net8220),
     .bm_sweb_o(net8221[0:1]), .bm_wdummymux_en_o(net8222),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sdo_i(net8224[0:1]),
     .bm_sdo_o(bm_sdo_o[1:0]));
clk_colbufx8 I790 ( .clko(glb_netwk_08[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I798 ( .clko(glb_netwk_12[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I787 ( .clko(glb_netwk_04[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I791 ( .clko(glb_netwk_06[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I788 ( .clko(glb_netwk_03[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I800 ( .clko(glb_netwk_09[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I786 ( .clko(glb_netwk_02[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I789 ( .clko(glb_netwk_07[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I799 ( .clko(glb_netwk_10[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I797 ( .clko(glb_netwk_11[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I793 ( .clko(glb_netwk_io_l[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I792 ( .clko(glb_netwk_05[7:0]), .clki(net7976[0:7]));
clk_colbufx8 I785 ( .clko(glb_netwk_01[7:0]), .clki(net7976[0:7]));

endmodule
// Library - leafcell, Cell - QUAD_TL, View - schematic
// LAST TIME SAVED: Sep 15 14:08:44 2008
// NETLIST TIME: Nov 14 16:12:04 2008
`timescale 1ns / 1ns 

module QUAD_TL ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, ceb_o, cf_l, cf_t, fabric_out_30,
     fabric_out_226, fabric_out_228, hiz_b_o, mode_o, padeb_l, padeb_t,
     padin_30, padin_226, pado_l, pado_t, r_o, sdo, shift_o,
     slf_op_00_11, slf_op_01_11, slf_op_02_11, slf_op_03_11,
     slf_op_04_11, slf_op_05_11, slf_op_06_11, slf_op_07_11,
     slf_op_08_11, slf_op_09_11, slf_op_10_11, slf_op_11_11,
     slf_op_12_11, slf_op_12_12, slf_op_12_13, slf_op_12_14,
     slf_op_12_15, slf_op_12_16, slf_op_12_17, slf_op_12_18,
     slf_op_12_19, slf_op_12_20, slf_op_12_21, tclk_o, update_o, bl,
     pgate, reset_b, sp4_h_r_12_11, sp4_h_r_12_12, sp4_h_r_12_13,
     sp4_h_r_12_14, sp4_h_r_12_15, sp4_h_r_12_16, sp4_h_r_12_17,
     sp4_h_r_12_18, sp4_h_r_12_19, sp4_h_r_12_20, sp4_h_r_12_21,
     sp4_r_v_b_12_11, sp4_r_v_b_12_12, sp4_r_v_b_12_13,
     sp4_r_v_b_12_14, sp4_r_v_b_12_15, sp4_r_v_b_12_16,
     sp4_r_v_b_12_17, sp4_r_v_b_12_18, sp4_r_v_b_12_19,
     sp4_r_v_b_12_20, sp4_v_b_00_11, sp4_v_b_01_11, sp4_v_b_02_11,
     sp4_v_b_03_11, sp4_v_b_04_11, sp4_v_b_05_11, sp4_v_b_06_11,
     sp4_v_b_07_11, sp4_v_b_08_11, sp4_v_b_09_11, sp4_v_b_10_11,
     sp4_v_b_11_11, sp4_v_b_12_11, sp12_h_r_12_11, sp12_h_r_12_12,
     sp12_h_r_12_13, sp12_h_r_12_14, sp12_h_r_12_15, sp12_h_r_12_16,
     sp12_h_r_12_17, sp12_h_r_12_18, sp12_h_r_12_19, sp12_h_r_12_20,
     sp12_v_b_01_11, sp12_v_b_02_11, sp12_v_b_03_11, sp12_v_b_04_11,
     sp12_v_b_05_11, sp12_v_b_06_11, sp12_v_b_07_11, sp12_v_b_08_11,
     sp12_v_b_09_11, sp12_v_b_10_11, sp12_v_b_11_11, sp12_v_b_12_11,
     vdd_cntl, wl, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_01_11, bnl_op_02_11, bnl_op_03_11,
     bnl_op_04_11, bnl_op_05_11, bnl_op_06_11, bnl_op_07_11,
     bnl_op_08_11, bnl_op_09_11, bnl_op_10_11, bnl_op_11_11,
     bnl_op_12_11, bnr_op_00_11, bnr_op_01_11, bnr_op_02_11,
     bnr_op_03_11, bnr_op_04_11, bnr_op_05_11, bnr_op_06_11,
     bnr_op_07_11, bnr_op_08_11, bnr_op_09_11, bnr_op_10_11,
     bnr_op_11_11, bnr_op_12_11, bot_op_01_11, bot_op_02_11,
     bot_op_03_11, bot_op_04_11, bot_op_05_11, bot_op_06_11,
     bot_op_07_11, bot_op_08_11, bot_op_09_11, bot_op_10_11,
     bot_op_11_11, bot_op_12_11, bs_en_i, carry_in_01_11,
     carry_in_02_11, carry_in_03_11, carry_in_04_11, carry_in_05_11,
     carry_in_07_11, carry_in_08_11, carry_in_09_11, carry_in_10_11,
     carry_in_11_11, carry_in_12_11, ceb_i, end_of_startup_lft_t,
     end_of_startup_top_l, glb_in, hiz_b_i, hold_l_t, hold_t_l, mode_i,
     padin_l, padin_t, prog, purst, r_i, rgt_op_12_11, rgt_op_12_12,
     rgt_op_12_13, rgt_op_12_14, rgt_op_12_15, rgt_op_12_16,
     rgt_op_12_17, rgt_op_12_18, rgt_op_12_19, rgt_op_12_20, sdi,
     shift_i, tclk_i, tiegnd, tievdd, tnr_op_12_20, update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bs_en_o, ceb_o,
     fabric_out_30, fabric_out_226, fabric_out_228, hiz_b_o, mode_o,
     padin_30, padin_226, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en_i,
     carry_in_01_11, carry_in_02_11, carry_in_03_11, carry_in_04_11,
     carry_in_05_11, carry_in_07_11, carry_in_08_11, carry_in_09_11,
     carry_in_10_11, carry_in_11_11, carry_in_12_11, ceb_i, hiz_b_i,
     hold_l_t, hold_t_l, mode_i, prog, purst, r_i, sdi, shift_i,
     tclk_i, tiegnd, tievdd, update_i;

output [7:0]  slf_op_04_11;
output [7:0]  slf_op_05_11;
output [7:0]  slf_op_02_11;
output [7:0]  slf_op_12_13;
output [7:0]  slf_op_12_19;
output [7:0]  slf_op_12_12;
output [7:0]  slf_op_10_11;
output [7:0]  slf_op_12_16;
output [7:0]  slf_op_12_20;
output [7:0]  slf_op_12_15;
output [7:0]  slf_op_11_11;
output [3:0]  slf_op_00_11;
output [7:0]  slf_op_06_11;
output [7:0]  slf_op_01_11;
output [7:0]  slf_op_07_11;
output [7:0]  slf_op_09_11;
output [7:0]  slf_op_08_11;
output [7:0]  slf_op_12_14;
output [39:20]  pado_l;
output [7:0]  slf_op_12_17;
output [287:0]  cf_t;
output [7:0]  slf_op_12_18;
output [23:0]  padeb_t;
output [39:20]  padeb_l;
output [479:240]  cf_l;
output [7:0]  bm_sa_o;
output [23:0]  pado_t;
output [3:0]  slf_op_12_21;
output [7:0]  slf_op_12_11;
output [7:0]  slf_op_03_11;

inout [47:0]  sp4_h_r_12_19;
inout [47:0]  sp4_r_v_b_12_18;
inout [23:0]  sp12_h_r_12_20;
inout [47:0]  sp4_r_v_b_12_19;
inout [47:0]  sp4_v_b_08_11;
inout [47:0]  sp4_v_b_05_11;
inout [23:0]  sp12_h_r_12_19;
inout [47:0]  sp4_h_r_12_16;
inout [23:0]  sp12_h_r_12_12;
inout [23:0]  sp12_v_b_11_11;
inout [23:0]  sp12_h_r_12_16;
inout [47:0]  sp4_h_r_12_18;
inout [23:0]  sp12_h_r_12_18;
inout [23:0]  sp12_h_r_12_14;
inout [23:0]  sp12_h_r_12_15;
inout [47:0]  sp4_v_b_04_11;
inout [47:0]  sp4_h_r_12_20;
inout [23:0]  sp12_v_b_06_11;
inout [47:0]  sp4_r_v_b_12_16;
inout [47:0]  sp4_h_r_12_17;
inout [23:0]  sp12_v_b_04_11;
inout [23:0]  sp12_v_b_12_11;
inout [23:0]  sp12_v_b_05_11;
inout [47:0]  sp4_r_v_b_12_15;
inout [47:0]  sp4_r_v_b_12_17;
inout [23:0]  sp12_v_b_10_11;
inout [47:0]  sp4_r_v_b_12_12;
inout [47:0]  sp4_h_r_12_11;
inout [47:0]  sp4_h_r_12_12;
inout [47:0]  sp4_v_b_02_11;
inout [47:0]  sp4_r_v_b_12_14;
inout [47:0]  sp4_v_b_10_11;
inout [47:0]  sp4_r_v_b_12_20;
inout [23:0]  sp12_v_b_03_11;
inout [23:0]  sp12_v_b_08_11;
inout [23:0]  sp12_v_b_07_11;
inout [351:176]  vdd_cntl;
inout [47:0]  sp4_v_b_06_11;
inout [47:0]  sp4_h_r_12_14;
inout [47:0]  sp4_v_b_03_11;
inout [23:0]  sp12_v_b_01_11;
inout [47:0]  sp4_v_b_12_11;
inout [47:0]  sp4_r_v_b_12_13;
inout [351:176]  wl;
inout [23:0]  sp12_v_b_09_11;
inout [23:0]  sp12_v_b_02_11;
inout [47:0]  sp4_v_b_01_11;
inout [23:0]  sp12_h_r_12_13;
inout [23:0]  sp12_h_r_12_11;
inout [47:0]  sp4_v_b_07_11;
inout [351:176]  pgate;
inout [653:0]  bl;
inout [351:176]  reset_b;
inout [47:0]  sp4_h_r_12_15;
inout [47:0]  sp4_h_r_12_13;
inout [47:0]  sp4_r_v_b_12_11;
inout [15:0]  sp4_h_r_12_21;
inout [47:0]  sp4_v_b_11_11;
inout [15:0]  sp4_v_b_00_11;
inout [23:0]  sp12_h_r_12_17;
inout [47:0]  sp4_v_b_09_11;

input [7:0]  bnr_op_11_11;
input [7:0]  bot_op_10_11;
input [7:0]  bot_op_03_11;
input [7:0]  bot_op_07_11;
input [7:0]  bnl_op_03_11;
input [7:0]  rgt_op_12_13;
input [7:0]  bot_op_09_11;
input [7:0]  bm_sa_i;
input [7:0]  bnr_op_12_11;
input [7:0]  bnl_op_08_11;
input [7:0]  bnr_op_07_11;
input [7:0]  bnr_op_05_11;
input [7:0]  bnl_op_02_11;
input [7:0]  bnl_op_12_11;
input [7:0]  bot_op_11_11;
input [7:0]  bnl_op_09_11;
input [7:0]  bot_op_05_11;
input [7:0]  rgt_op_12_19;
input [7:0]  bnr_op_02_11;
input [7:0]  bnr_op_04_11;
input [7:0]  rgt_op_12_11;
input [7:0]  bnr_op_03_11;
input [7:0]  bnl_op_01_11;
input [7:0]  bnl_op_04_11;
input [7:0]  glb_in;
input [7:0]  rgt_op_12_14;
input [7:0]  bnl_op_06_11;
input [7:0]  bnr_op_01_11;
input [7:0]  bnl_op_07_11;
input [7:0]  bnl_op_10_11;
input [7:0]  bot_op_08_11;
input [7:0]  bnr_op_10_11;
input [7:0]  rgt_op_12_18;
input [7:0]  rgt_op_12_20;
input [7:0]  bot_op_02_11;
input [7:0]  rgt_op_12_12;
input [7:0]  bnr_op_08_11;
input [7:0]  bot_op_04_11;
input [7:0]  rgt_op_12_15;
input [39:20]  padin_l;
input [7:0]  bot_op_01_11;
input [23:0]  padin_t;
input [7:0]  bnr_op_09_11;
input [3:0]  tnr_op_12_20;
input [11:0]  end_of_startup_top_l;
input [9:0]  end_of_startup_lft_t;
input [7:0]  bnl_op_11_11;
input [7:0]  bot_op_06_11;
input [7:0]  bot_op_12_11;
input [7:0]  bnr_op_00_11;
input [7:0]  rgt_op_12_17;
input [7:0]  rgt_op_12_16;
input [7:0]  bnr_op_06_11;
input [7:0]  bnl_op_05_11;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:23]  net_7758;

wire  [0:47]  net_8171;

wire  [0:23]  net_4807;

wire  [0:23]  net_5227;

wire  [0:23]  net_4723;

wire  [0:7]  net_7147;

wire  [0:47]  net_6967;

wire  [0:23]  net_5593;

wire  [0:7]  net_5551;

wire  [0:23]  net_6685;

wire  [0:23]  net_6349;

wire  [0:23]  net_6993;

wire  [0:47]  net_4892;

wire  [0:47]  net_5315;

wire  [0:7]  net_6979;

wire  [0:23]  net_5255;

wire  [0:47]  net_5147;

wire  [0:23]  net_5845;

wire  [0:23]  net_7105;

wire  [0:1]  net_8272;

wire  [0:23]  net_4022;

wire  [0:23]  net_5257;

wire  [0:23]  net_7327;

wire  [0:23]  net_5285;

wire  [0:23]  net_6683;

wire  [0:23]  net_5369;

wire  [0:23]  net_5451;

wire  [0:15]  net_7874;

wire  [0:47]  net_4531;

wire  [0:47]  net_5928;

wire  [0:47]  net_7594;

wire  [0:47]  net_4867;

wire  [0:23]  net_4613;

wire  [0:1]  net_7902;

wire  [0:23]  net_4226;

wire  [0:47]  net_5200;

wire  [0:47]  net_8035;

wire  [0:47]  net_4500;

wire  [0:7]  net_6409;

wire  [0:7]  net_5915;

wire  [0:47]  net_5483;

wire  [0:47]  net_5203;

wire  [0:23]  net_4445;

wire  [0:47]  net_4021;

wire  [0:47]  net_7415;

wire  [0:47]  net_4225;

wire  [0:23]  net_4192;

wire  [0:47]  net_6519;

wire  [0:15]  net_4258;

wire  [0:47]  net_7933;

wire  [0:23]  net_6545;

wire  [0:7]  net_5149;

wire  [0:7]  net_5103;

wire  [0:7]  net_7175;

wire  [0:23]  net_5283;

wire  [0:7]  net_7315;

wire  [0:7]  net_6027;

wire  [0:47]  net_6911;

wire  [0:7]  net_6531;

wire  [0:23]  net_4641;

wire  [0:23]  net_7591;

wire  [0:47]  net_6992;

wire  [0:47]  net_7644;

wire  [0:47]  net_6155;

wire  [0:47]  net_7107;

wire  [0:47]  net_6407;

wire  [0:47]  net_6938;

wire  [0:47]  net_5592;

wire  [0:47]  net_7247;

wire  [0:23]  net_4557;

wire  [0:7]  net_7427;

wire  [0:47]  net_7593;

wire  [0:15]  net_7908;

wire  [0:47]  net_6015;

wire  [0:23]  net_4667;

wire  [0:47]  net_6323;

wire  [0:47]  net_5480;

wire  [0:47]  net_6320;

wire  [0:47]  net_4920;

wire  [0:15]  net_4326;

wire  [0:47]  net_6351;

wire  [0:23]  net_6237;

wire  [0:23]  net_5087;

wire  [0:23]  net_5817;

wire  [0:23]  net_7385;

wire  [0:23]  net_5927;

wire  [0:23]  net_4583;

wire  [0:47]  net_6936;

wire  [0:7]  net_6951;

wire  [0:23]  net_6907;

wire  [0:47]  net_5844;

wire  [0:23]  net_4753;

wire  [0:23]  net_5229;

wire  [0:47]  net_6908;

wire  [7:0]  net2col_drivers;

wire  [7:0]  glb_netwk_02;

wire  [7:0]  glb_netwk_00;

wire  [7:0]  glb_netwk_08;

wire  [7:0]  glb_netwk_07;

wire  [7:0]  glb_netwk_05;

wire  [0:23]  net_6179;

wire  [7:0]  glb_netwk_01;

wire  [3:0]  io_t_6;

wire  [3:0]  io_t_8;

wire  [0:23]  net_6347;

wire  [7:0]  glb_netwk_09;

wire  [7:0]  glb_netwk_06;

wire  [7:0]  glb_netwk_io_l;

wire  [3:0]  io_t_4;

wire  [0:23]  net_7329;

wire  [0:7]  net_5159;

wire  [7:0]  glb_netwk_10;

wire  [0:23]  net_6797;

wire  [0:7]  net_6223;

wire  [0:7]  net_5607;

wire  [0:47]  net_7244;

wire  [0:23]  net_7355;

wire  [7:0]  glb_netwk_04;

wire  [0:23]  net_6543;

wire  [0:7]  net_4461;

wire  [0:47]  net_6488;

wire  [0:7]  net_7688;

wire  [0:47]  net_5648;

wire  [0:47]  net_4979;

wire  [0:47]  net_5118;

wire  [0:23]  net_7495;

wire  [0:23]  net_5677;

wire  [0:47]  net_4387;

wire  [0:47]  net_4123;

wire  [0:23]  net_5761;

wire  [0:15]  net_4122;

wire  [0:23]  net_7469;

wire  [0:23]  net_6853;

wire  [0:1]  net_8238;

wire  [0:47]  net_4559;

wire  [0:7]  net_7973;

wire  [0:23]  net_4501;

wire  [0:47]  net_6491;

wire  [0:7]  net_5887;

wire  [0:47]  net_7771;

wire  [0:23]  net_6067;

wire  [0:23]  net_5983;

wire  [0:23]  net_7299;

wire  [0:47]  net_6600;

wire  [0:47]  net_6124;

wire  [0:47]  net_7135;

wire  [0:23]  net_5509;

wire  [0:47]  net_7300;

wire  [0:47]  net_6099;

wire  [0:23]  net_4124;

wire  [0:47]  net_4615;

wire  [0:23]  net_6123;

wire  [0:47]  net_5900;

wire  [0:23]  net_5535;

wire  [0:47]  net_6404;

wire  [0:47]  net_6267;

wire  [0:47]  net_7132;

wire  [0:23]  net_7566;

wire  [0:47]  net_7020;

wire  [0:47]  net_5256;

wire  [0:23]  net_6405;

wire  [0:7]  net_4935;

wire  [0:1]  net_8275;

wire  [0:23]  net_5537;

wire  [3:0]  io_l_34;

wire  [0:7]  net_7871;

wire  [7:0]  glb_netwk_03;

wire  [0:47]  net_5536;

wire  [3:0]  io_t_2;

wire  [0:23]  net_5061;

wire  [0:15]  net_8044;

wire  [0:47]  net_7328;

wire  [0:7]  net_6129;

wire  [0:47]  net_4670;

wire  [0:23]  net_6599;

wire  [0:47]  net_4698;

wire  [0:23]  net_7131;

wire  [0:7]  net_5121;

wire  [0:47]  net_7597;

wire  [0:47]  net_5119;

wire  [0:47]  net_4327;

wire  [0:7]  net_7552;

wire  [0:23]  net_6769;

wire  [0:47]  net_5259;

wire  [0:47]  net_7272;

wire  [0:47]  net_5620;

wire  [0:23]  net_7077;

wire  [0:47]  net_7496;

wire  [0:23]  net_5621;

wire  [0:47]  net_5032;

wire  [0:47]  net_4389;

wire  [0:15]  net_4224;

wire  [0:1]  net_8174;

wire  [0:7]  net_6111;

wire  [0:15]  net_8010;

wire  [0:23]  net_5929;

wire  [0:23]  net_6573;

wire  [0:47]  net_5396;

wire  [0:23]  net_6487;

wire  [0:47]  net_5312;

wire  [0:47]  net_5567;

wire  [0:47]  net_7048;

wire  [0:23]  net_4893;

wire  [0:1]  net_7936;

wire  [0:47]  net_5676;

wire  [0:23]  net_4977;

wire  [0:23]  net_4090;

wire  [0:7]  net_6363;

wire  [0:23]  net_6767;

wire  [0:47]  net_7865;

wire  [0:47]  net_4584;

wire  [0:23]  net_5871;

wire  [0:47]  net_5060;

wire  [0:47]  net_4923;

wire  [0:47]  net_5762;

wire  [0:7]  net_7455;

wire  [0:23]  net_5649;

wire  [0:47]  net_7359;

wire  [0:47]  net_4388;

wire  [0:23]  net_6879;

wire  [0:7]  net_6615;

wire  [0:23]  net_6461;

wire  [0:23]  net_5563;

wire  [0:23]  net_6151;

wire  [0:7]  net_6101;

wire  [0:47]  net_6880;

wire  [0:23]  net_4809;

wire  [0:23]  net_5089;

wire  [0:47]  net_7647;

wire  [0:47]  net_4864;

wire  [0:23]  net_6963;

wire  [0:47]  net_6348;

wire  [0:23]  net_5481;

wire  [0:23]  net_7049;

wire  [0:7]  net_5299;

wire  [0:1]  net_8267;

wire  [0:23]  net_4529;

wire  [0:47]  net_5847;

wire  [0:7]  net_7277;

wire  [0:47]  net_7216;

wire  [0:47]  net_5284;

wire  [0:23]  net_6125;

wire  [0:23]  net_5899;

wire  [0:23]  net_4585;

wire  [0:7]  net_6913;

wire  [0:23]  net_7676;

wire  [0:23]  net_5901;

wire  [0:15]  net_7840;

wire  [0:23]  net_6403;

wire  [0:47]  net_6432;

wire  [0:47]  net_6127;

wire  [0:47]  net_5984;

wire  [0:7]  net_7091;

wire  [0:23]  net_6713;

wire  [0:47]  net_7104;

wire  [0:7]  net_4785;

wire  [0:7]  net_7719;

wire  [0:23]  net_6627;

wire  [0:47]  net_4668;

wire  [0:23]  net_5395;

wire  [0:23]  net_6235;

wire  [0:15]  net_4190;

wire  [0:47]  net_7596;

wire  [0:47]  net_5875;

wire  [0:47]  net_4808;

wire  [0:47]  net_6603;

wire  [0:7]  net_5205;

wire  [0:7]  net_5999;

wire  [0:23]  net_6097;

wire  [0:23]  net_6657;

wire  [0:1]  net_7970;

wire  [0:23]  net_6095;

wire  [0:7]  net_7614;

wire  [0:7]  net_7287;

wire  [0:47]  net_6684;

wire  [0:23]  net_5171;

wire  [0:23]  net_7677;

wire  [0:23]  net_6209;

wire  [0:23]  net_5565;

wire  [0:23]  net_6041;

wire  [0:47]  net_4612;

wire  [0:23]  net_5201;

wire  [0:1]  net_8230;

wire  [0:23]  net_4725;

wire  [0:7]  net_5579;

wire  [0:7]  net_7119;

wire  [0:23]  net_7634;

wire  [0:23]  net_4695;

wire  [0:47]  net_7023;

wire  [0:23]  net_7217;

wire  [0:23]  net_5479;

wire  [0:23]  net_6825;

wire  [0:15]  net_8180;

wire  [0:47]  net_5595;

wire  [0:47]  net_4191;

wire  [0:23]  net_5787;

wire  [0:47]  net_5763;

wire  [0:23]  net_4751;

wire  [0:47]  net_6435;

wire  [0:47]  net_4472;

wire  [0:7]  net_5037;

wire  [0:47]  net_7443;

wire  [0:23]  net_5733;

wire  [0:7]  net_5691;

wire  [0:47]  net_5732;

wire  [0:23]  net_6741;

wire  [0:23]  net_7133;

wire  [0:23]  net_6517;

wire  [0:47]  net_4836;

wire  [0:7]  net_4617;

wire  [0:7]  net_5131;

wire  [0:23]  net_6433;

wire  [3:0]  io_l_22;

wire  [0:7]  net_6503;

wire  [3:0]  io_l_38;

wire  [0:47]  net_6239;

wire  [0:47]  net_4780;

wire  [0:47]  net_6068;

wire  [0:47]  net_4556;

wire  [0:47]  net_4783;

wire  [0:23]  net_5619;

wire  [0:47]  net_5228;

wire  [0:47]  net_4528;

wire  [3:0]  io_l_32;

wire  [0:23]  net_6459;

wire  [0:23]  net_4697;

wire  [0:23]  net_5031;

wire  [0:23]  net_5703;

wire  [0:47]  net_7160;

wire  [0:47]  net_4259;

wire  [0:7]  net_7905;

wire  [0:7]  net_6381;

wire  [3:0]  io_l_28;

wire  [0:23]  net_5005;

wire  [0:1]  net_8261;

wire  [0:47]  net_7051;

wire  [0:47]  net_7967;

wire  [0:47]  net_7499;

wire  [0:47]  net_6152;

wire  [0:47]  net_6463;

wire  [0:47]  net_6855;

wire  [0:23]  net_5705;

wire  [0:47]  net_4383;

wire  [0:47]  net_6295;

wire  [0:47]  net_7076;

wire  [3:0]  io_l_36;

wire  [0:47]  net_7678;

wire  [0:1]  net_8004;

wire  [0:23]  net_4919;

wire  [0:7]  net_6643;

wire  [0:47]  net_5903;

wire  [0:23]  net_5985;

wire  [0:7]  net_7037;

wire  [0:7]  net_7249;

wire  [0:47]  net_4643;

wire  [0:47]  net_8137;

wire  [0:7]  net_6167;

wire  [0:47]  net_6208;

wire  [0:23]  net_5425;

wire  [0:7]  net_5383;

wire  [0:23]  net_6991;

wire  [0:7]  net_7837;

wire  [0:47]  net_6547;

wire  [0:7]  net_7343;

wire  [0:47]  net_5508;

wire  [0:23]  net_5173;

wire  [0:23]  net_4376;

wire  [0:7]  net_7193;

wire  [0:47]  net_5679;

wire  [0:47]  net_4444;

wire  [3:0]  io_t_20;

wire  [0:47]  net_5399;

wire  [0:7]  net_5075;

wire  [0:47]  net_4811;

wire  [0:47]  net_6852;

wire  [0:23]  net_6909;

wire  [0:47]  net_7188;

wire  [0:47]  net_5091;

wire  [0:15]  net_4292;

wire  [0:23]  net_5789;

wire  [0:23]  net_5003;

wire  [0:23]  net_6851;

wire  [3:0]  io_l_24;

wire  [3:0]  io_l_30;

wire  [0:47]  net_6126;

wire  [0:23]  net_6321;

wire  [7:0]  glb_netwk_11;

wire  [3:0]  io_t_16;

wire  [0:1]  net_8245;

wire  [0:23]  net_6711;

wire  [0:1]  net_8072;

wire  [0:23]  net_4158;

wire  [0:47]  net_5707;

wire  [0:1]  net_8234;

wire  [0:47]  net_5819;

wire  [0:7]  net_4673;

wire  [0:23]  net_7637;

wire  [0:23]  net_6013;

wire  [0:47]  net_6712;

wire  [0:47]  net_4475;

wire  [0:47]  net_4055;

wire  [0:23]  net_5313;

wire  [0:47]  net_7163;

wire  [0:23]  net_4863;

wire  [0:15]  net_4020;

wire  [0:23]  net_5843;

wire  [0:47]  net_5371;

wire  [0:23]  net_6881;

wire  [0:23]  net_6601;

wire  [0:23]  net_7357;

wire  [0:23]  net_6181;

wire  [0:47]  net_4640;

wire  [0:23]  net_5199;

wire  [0:23]  net_6965;

wire  [0:23]  net_7271;

wire  [0:47]  net_6460;

wire  [0:23]  net_5591;

wire  [0:7]  net_7781;

wire  [0:23]  net_4527;

wire  [0:47]  net_7681;

wire  [0:47]  net_8069;

wire  [0:15]  net_4054;

wire  [0:47]  net_5791;

wire  [0:7]  net_5019;

wire  [0:23]  net_5675;

wire  [0:23]  net_4779;

wire  [0:7]  net_6335;

wire  [0:23]  net_7413;

wire  [0:7]  net_5215;

wire  [0:47]  net_4293;

wire  [0:47]  net_6799;

wire  [0:47]  net_5623;

wire  [0:47]  net_6964;

wire  [0:23]  net_4380;

wire  [0:7]  net_6307;

wire  [0:47]  net_5564;

wire  [0:47]  net_7831;

wire  [0:23]  net_4056;

wire  [0:23]  net_7047;

wire  [0:23]  net_6069;

wire  [0:7]  net_6195;

wire  [0:23]  net_4443;

wire  [0:47]  net_4895;

wire  [0:47]  net_4157;

wire  [0:23]  net_7761;

wire  [0:47]  net_5231;

wire  [0:23]  net_7019;

wire  [0:23]  net_5311;

wire  [0:47]  net_6631;

wire  [0:23]  net_7592;

wire  [0:23]  net_7187;

wire  [0:7]  net_4991;

wire  [0:23]  net_7075;

wire  [0:47]  net_5816;

wire  [0:47]  net_6995;

wire  [0:47]  net_4948;

wire  [0:47]  net_5872;

wire  [0:7]  net_6447;

wire  [0:47]  net_7899;

wire  [0:47]  net_4976;

wire  [0:23]  net_4781;

wire  [0:23]  net_5341;

wire  [0:47]  net_7191;

wire  [0:23]  net_6153;

wire  [0:23]  net_5367;

wire  [0:23]  net_7441;

wire  [0:47]  net_6796;

wire  [0:47]  net_7646;

wire  [0:47]  net_6376;

wire  [0:47]  net_5063;

wire  [0:23]  net_4379;

wire  [0:23]  net_7702;

wire  [0:23]  net_6265;

wire  [0:23]  net_7273;

wire  [0:23]  net_4975;

wire  [0:23]  net_7301;

wire  [0:47]  net_5172;

wire  [0:47]  net_6379;

wire  [0:7]  net_4963;

wire  [0:47]  net_5651;

wire  [0:23]  net_4865;

wire  [0:47]  net_5007;

wire  [0:47]  net_7440;

wire  [0:23]  net_6795;

wire  [0:7]  net_6923;

wire  [0:23]  net_4949;

wire  [0:47]  net_5175;

wire  [0:7]  net_8177;

wire  [0:47]  net_4696;

wire  [3:0]  io_l_26;

wire  [0:7]  net_7583;

wire  [0:23]  net_6629;

wire  [0:47]  net_5455;

wire  [0:7]  net_5411;

wire  [0:47]  net_6098;

wire  [0:47]  net_5144;

wire  [0:23]  net_6431;

wire  [0:23]  net_6011;

wire  [0:47]  net_5368;

wire  [0:15]  net_8078;

wire  [0:47]  net_7219;

wire  [0:23]  net_6319;

wire  [0:23]  net_7411;

wire  [0:47]  net_5035;

wire  [0:23]  net_4471;

wire  [0:47]  net_4386;

wire  [0:47]  net_6096;

wire  [0:47]  net_7770;

wire  [0:23]  net_7439;

wire  [0:47]  net_6516;

wire  [0:7]  net_7221;

wire  [0:23]  net_4499;

wire  [0:47]  net_5146;

wire  [0:23]  net_5759;

wire  [0:47]  net_6939;

wire  [0:23]  net_7497;

wire  [0:23]  net_7021;

wire  [0:1]  net_8106;

wire  [0:47]  net_5931;

wire  [0:47]  net_5760;

wire  [0:23]  net_6377;

wire  [0:1]  net_8266;

wire  [0:23]  net_7189;

wire  [0:47]  net_6292;

wire  [0:47]  net_5116;

wire  [0:23]  net_6515;

wire  [0:23]  net_5059;

wire  [0:7]  net_7738;

wire  [0:7]  net_5775;

wire  [0:23]  net_5115;

wire  [0:1]  net_7868;

wire  [0:23]  net_4947;

wire  [0:47]  net_6071;

wire  [0:23]  net_5731;

wire  [0:23]  net_7161;

wire  [0:47]  net_8103;

wire  [0:47]  net_5539;

wire  [0:47]  net_6236;

wire  [0:1]  net_8250;

wire  [0:47]  net_7356;

wire  [0:7]  net_6475;

wire  [0:23]  net_6291;

wire  [0:23]  net_4473;

wire  [0:1]  net_8208;

wire  [0:47]  net_6768;

wire  [0:23]  net_5957;

wire  [0:7]  net_5747;

wire  [0:23]  net_7638;

wire  [0:23]  net_5815;

wire  [0:23]  net_7103;

wire  [0:47]  net_7412;

wire  [0:23]  net_4611;

wire  [0:47]  net_8001;

wire  [0:23]  net_5873;

wire  [0:23]  net_4921;

wire  [0:23]  net_4837;

wire  [0:23]  net_5647;

wire  [0:7]  net_5831;

wire  [0:47]  net_5788;

wire  [0:47]  net_7768;

wire  [0:47]  net_7331;

wire  [0:47]  net_6910;

wire  [0:7]  net_6279;

wire  [0:23]  net_6263;

wire  [0:47]  net_6628;

wire  [0:15]  net_7942;

wire  [0:7]  net_6225;

wire  [0:7]  net_5859;

wire  [0:7]  net_8143;

wire  [0:7]  net_4701;

wire  [0:47]  net_5452;

wire  [0:7]  net_7259;

wire  [0:7]  net_5765;

wire  [0:23]  net_4328;

wire  [0:23]  net_4891;

wire  [0:7]  net_5635;

wire  [0:7]  net_6465;

wire  [3:0]  io_t_0;

wire  [0:23]  net_4260;

wire  [3:0]  io_t_10;

wire  [0:23]  net_4555;

wire  [0:7]  net_6941;

wire  [0:47]  net_6183;

wire  [0:7]  net_8211;

wire  [0:7]  net_7939;

wire  [0:23]  net_5117;

wire  [0:47]  net_7275;

wire  [0:47]  net_6264;

wire  [0:7]  net_4729;

wire  [0:7]  net_5271;

wire  [0:23]  net_5145;

wire  [0:15]  net_4156;

wire  [0:47]  net_5987;

wire  [0:23]  net_4639;

wire  [0:47]  net_4089;

wire  [0:47]  net_6687;

wire  [0:7]  net_7007;

wire  [0:7]  net_5719;

wire  [0:47]  net_7303;

wire  [0:47]  net_7682;

wire  [0:23]  net_5397;

wire  [0:23]  net_7243;

wire  [0:23]  net_6207;

wire  [0:1]  net_7834;

wire  [0:7]  net_5233;

wire  [0:47]  net_6180;

wire  [0:7]  net_4757;

wire  [0:47]  net_5511;

wire  [0:7]  net_5177;

wire  [0:23]  net_7159;

wire  [0:23]  net_6935;

wire  [0:1]  net_8140;

wire  [0:47]  net_4752;

wire  [0:15]  net_8146;

wire  [0:23]  net_5143;

wire  [0:7]  net_5243;

wire  [0:23]  net_6293;

wire  [0:23]  net_7762;

wire  [0:7]  net_6139;

wire  [0:23]  net_5453;

wire  [0:47]  net_7679;

wire  [0:47]  net_4724;

wire  [0:15]  net_8214;

wire  [0:47]  net_5735;

wire  [3:0]  io_t_14;

wire  [0:47]  net_6544;

wire  [0:47]  net_5704;

wire  [0:23]  net_4835;

wire  [0:47]  net_7645;

wire  [0:47]  net_5287;

wire  [0:23]  net_5507;

wire  [0:23]  net_6489;

wire  [0:47]  net_7079;

wire  [0:47]  net_5004;

wire  [0:23]  net_7215;

wire  [0:7]  net_8007;

wire  [0:15]  net_7976;

wire  [0:23]  net_7245;

wire  [0:47]  net_5088;

wire  [0:15]  net_4088;

wire  [0:23]  net_5033;

wire  [3:0]  io_t_18;

wire  [0:1]  net_8038;

wire  [3:0]  io_t_12;

wire  [0:23]  net_6937;

wire  [0:7]  net_8041;

wire  [0:47]  net_6211;

wire  [0:23]  net_4294;

wire  [0:7]  net_6437;

wire  [0:47]  net_6012;

wire  [0:23]  net_4669;

wire  [0:23]  net_6375;

wire  [0:47]  net_4951;

wire  [0:47]  net_4671;

wire  [0:7]  net_7657;



bram_bufferx4x6 I1070 ( .in(sdi), .out(net_04041));
bram_bufferx4x6 I1071 ( .in(net_4405), .out(net_04038));
lowla_modified I1068 ( .clk(net_4407), .min(net_04038),
     .lao(net_4006));
lowla_modified I1066 ( .clk(tclk_i), .min(net_04041), .lao(net_8088));
io_col4_row I_00_20_iol39 ( .ceb(ceb_o), .cf(cf_l[263:240]),
     .vdd_cntl(vdd_cntl[335:320]), .hold(hold_l_t),
     .fabric_out(net_8252), .sdo(net_4040), .sdi(net_4006),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[9]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[39:38]), .pado(pado_l[39:38]),
     .padeb(padeb_l[39:38]), .sp4_v_t(net_4020[0:15]),
     .sp4_h_l(net_4021[0:47]), .sp12_h_l(net_4022[0:23]), .prog(prog),
     .spi_ss_in_b(net_8275[0:1]), .tnl_op({io_t_0[3], io_t_0[2],
     io_t_0[1], io_t_0[0], io_t_0[3], io_t_0[2], io_t_0[1],
     io_t_0[0]}), .lft_op(net_5765[0:7]), .bnl_op(net_6129[0:7]),
     .pgate(pgate[335:320]), .reset(reset_b[335:320]),
     .sp4_v_b(net_4054[0:15]), .wl(wl[335:320]), .bl(bl[17:0]),
     .slf_op(io_l_38[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_19_iol37 ( .ceb(ceb_o), .cf(cf_l[287:264]),
     .vdd_cntl(vdd_cntl[319:304]), .hold(hold_l_t),
     .fabric_out(net_8264), .sdo(net_4278), .sdi(net_4040),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[8]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[37:36]), .pado(pado_l[37:36]),
     .padeb(padeb_l[37:36]), .sp4_v_t(net_4054[0:15]),
     .sp4_h_l(net_4055[0:47]), .sp12_h_l(net_4056[0:23]), .prog(prog),
     .spi_ss_in_b(net_8238[0:1]), .tnl_op(net_5765[0:7]),
     .lft_op(net_6129[0:7]), .bnl_op(net_6101[0:7]),
     .pgate(pgate[319:304]), .reset(reset_b[319:304]),
     .sp4_v_b(net_4292[0:15]), .wl(wl[319:304]), .bl(bl[17:0]),
     .slf_op(io_l_36[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_16_iol31 ( .ceb(ceb_o), .cf(cf_l[359:336]),
     .vdd_cntl(vdd_cntl[271:256]), .hold(hold_l_t),
     .fabric_out(net_8228), .sdo(net_4108), .sdi(net_4074),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[5]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[31:30]), .pado(pado_l[31:30]),
     .padeb(padeb_l[31:30]), .sp4_v_t(net_4088[0:15]),
     .sp4_h_l(net_4089[0:47]), .sp12_h_l(net_4090[0:23]), .prog(prog),
     .spi_ss_in_b(net_8261[0:1]), .tnl_op(net_5121[0:7]),
     .lft_op(net_5149[0:7]), .bnl_op(net_6941[0:7]),
     .pgate(pgate[271:256]), .reset(reset_b[271:256]),
     .sp4_v_b(net_4122[0:15]), .wl(wl[271:256]), .bl(bl[17:0]),
     .slf_op(io_l_30[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_15_iol29 ( .ceb(ceb_o), .cf(cf_l[383:360]),
     .vdd_cntl(vdd_cntl[255:240]), .hold(hold_l_t),
     .fabric_out(net_8255), .sdo(net_4107), .sdi(net_4108),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[4]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[29:28]), .pado(pado_l[29:28]),
     .padeb(padeb_l[29:28]), .sp4_v_t(net_4122[0:15]),
     .sp4_h_l(net_4123[0:47]), .sp12_h_l(net_4124[0:23]), .prog(prog),
     .spi_ss_in_b(net_8250[0:1]), .tnl_op(net_5149[0:7]),
     .lft_op(net_6941[0:7]), .bnl_op(net_6913[0:7]),
     .pgate(pgate[255:240]), .reset(reset_b[255:240]),
     .sp4_v_b(net_4224[0:15]), .wl(wl[255:240]), .bl(bl[17:0]),
     .slf_op(io_l_28[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_12_iol23 ( .ceb(ceb_o), .cf(cf_l[455:432]),
     .vdd_cntl(vdd_cntl[207:192]), .hold(hold_l_t),
     .fabric_out(net_8278), .sdo(net_4141), .sdi(net_4142),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[1]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[23:22]), .pado(pado_l[23:22]),
     .padeb(padeb_l[23:22]), .sp4_v_t(net_4156[0:15]),
     .sp4_h_l(net_4157[0:47]), .sp12_h_l(net_4158[0:23]), .prog(prog),
     .spi_ss_in_b(net_8267[0:1]), .tnl_op(net_4673[0:7]),
     .lft_op(net_4701[0:7]), .bnl_op(slf_op_01_11[7:0]),
     .pgate(pgate[207:192]), .reset(reset_b[207:192]),
     .sp4_v_b(net_4190[0:15]), .wl(wl[207:192]), .bl(bl[17:0]),
     .slf_op(io_l_22[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_11_iol21 ( .ceb(ceb_o), .cf(cf_l[479:456]),
     .vdd_cntl(vdd_cntl[191:176]), .hold(hold_l_t),
     .fabric_out(net_7531), .sdo(sdo), .sdi(net_4141), .spiout({tiegnd,
     tiegnd}), .cdone_in(end_of_startup_lft_t[0]), .spioeb({tievdd,
     tievdd}), .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o),
     .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_l[21:20]), .pado(pado_l[21:20]),
     .padeb(padeb_l[21:20]), .sp4_v_t(net_4190[0:15]),
     .sp4_h_l(net_4191[0:47]), .sp12_h_l(net_4192[0:23]), .prog(prog),
     .spi_ss_in_b(net_8234[0:1]), .tnl_op(net_4701[0:7]),
     .lft_op(slf_op_01_11[7:0]), .bnl_op(bnr_op_00_11[7:0]),
     .pgate(pgate[191:176]), .reset(reset_b[191:176]),
     .sp4_v_b(sp4_v_b_00_11[15:0]), .wl(wl[191:176]), .bl(bl[17:0]),
     .slf_op(slf_op_00_11[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_14_iol27 ( .ceb(ceb_o), .cf(cf_l[407:384]),
     .vdd_cntl(vdd_cntl[239:224]), .hold(hold_l_t),
     .fabric_out(net_8270), .sdo(net_4209), .sdi(net_4107),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[3]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[27:26]), .pado(pado_l[27:26]),
     .padeb(padeb_l[27:26]), .sp4_v_t(net_4224[0:15]),
     .sp4_h_l(net_4225[0:47]), .sp12_h_l(net_4226[0:23]), .prog(prog),
     .spi_ss_in_b(net_8230[0:1]), .tnl_op(net_6941[0:7]),
     .lft_op(net_6913[0:7]), .bnl_op(net_4673[0:7]),
     .pgate(pgate[239:224]), .reset(reset_b[239:224]),
     .sp4_v_b(net_4258[0:15]), .wl(wl[239:224]), .bl(bl[17:0]),
     .slf_op(io_l_26[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_13_iol25 ( .ceb(ceb_o), .cf(cf_l[431:408]),
     .vdd_cntl(vdd_cntl[223:208]), .hold(hold_l_t),
     .fabric_out(net_8274), .sdo(net_4142), .sdi(net_4209),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[2]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[25:24]), .pado(pado_l[25:24]),
     .padeb(padeb_l[25:24]), .sp4_v_t(net_4258[0:15]),
     .sp4_h_l(net_4259[0:47]), .sp12_h_l(net_4260[0:23]), .prog(prog),
     .spi_ss_in_b(net_8245[0:1]), .tnl_op(net_6913[0:7]),
     .lft_op(net_4673[0:7]), .bnl_op(net_4701[0:7]),
     .pgate(pgate[223:208]), .reset(reset_b[223:208]),
     .sp4_v_b(net_4156[0:15]), .wl(wl[223:208]), .bl(bl[17:0]),
     .slf_op(io_l_24[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_18_iol35 ( .ceb(ceb_o), .cf(cf_l[311:288]),
     .vdd_cntl(vdd_cntl[303:288]), .hold(hold_l_t),
     .fabric_out(net_8280), .sdo(net_4312), .sdi(net_4278),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[7]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[35:34]), .pado(pado_l[35:34]),
     .padeb(padeb_l[35:34]), .sp4_v_t(net_4292[0:15]),
     .sp4_h_l(net_4293[0:47]), .sp12_h_l(net_4294[0:23]), .prog(prog),
     .spi_ss_in_b(net_8266[0:1]), .tnl_op(net_6129[0:7]),
     .lft_op(net_6101[0:7]), .bnl_op(net_5121[0:7]),
     .pgate(pgate[303:288]), .reset(reset_b[303:288]),
     .sp4_v_b(net_4326[0:15]), .wl(wl[303:288]), .bl(bl[17:0]),
     .slf_op(io_l_34[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
io_col4_row I_00_17_iol33 ( .ceb(ceb_o), .cf(cf_l[335:312]),
     .vdd_cntl(vdd_cntl[287:272]), .hold(hold_l_t),
     .fabric_out(net_8224), .sdo(net_4074), .sdi(net_4312),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_lft_t[6]),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_l[33:32]), .pado(pado_l[33:32]),
     .padeb(padeb_l[33:32]), .sp4_v_t(net_4326[0:15]),
     .sp4_h_l(net_4327[0:47]), .sp12_h_l(net_4328[0:23]), .prog(prog),
     .spi_ss_in_b(net_8272[0:1]), .tnl_op(net_6101[0:7]),
     .lft_op(net_5121[0:7]), .bnl_op(net_5149[0:7]),
     .pgate(pgate[287:272]), .reset(reset_b[287:272]),
     .sp4_v_b(net_4088[0:15]), .wl(wl[287:272]), .bl(bl[17:0]),
     .slf_op(io_l_32[3:0]), .glb_netwk(glb_netwk_io_l[7:0]));
bram_4kprouting_tbankin I_bram0619 ( .glb_netwk(glb_netwk_05[7:0]),
     .vdd_cntl_bot(vdd_cntl[319:304]),
     .vdd_cntl_top(vdd_cntl[335:320]), .bm_sdo_o(net_7543),
     .bm_sdi_i(net_7545), .bm_sclkrw_i(net_7546), .bm_sdo_i(bm_sdo_i),
     .bm_sweb_i(net_7547), .bm_sdi_o(bm_sdi_o),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_sweb_o(bm_sweb_o),
     .slf_op_top(net_8177[0:7]), .slf_op_bot(net_7552[0:7]),
     .wl_top(wl[335:320]), .wl_bot(wl[319:304]),
     .top_op_top({io_t_10[3], io_t_10[2], io_t_10[1], io_t_10[0],
     io_t_10[3], io_t_10[2], io_t_10[1], io_t_10[0]}),
     .tnr_op_top({io_t_12[3], io_t_12[2], io_t_12[1], io_t_12[0],
     io_t_12[3], io_t_12[2], io_t_12[1], io_t_12[0]}),
     .tnr_op_bot(net_8211[0:7]), .tnl_op_top({io_t_8[3], io_t_8[2],
     io_t_8[1], io_t_8[0], io_t_8[3], io_t_8[2], io_t_8[1],
     io_t_8[0]}), .tnl_op_bot(net_7905[0:7]),
     .rgt_op_top(net_8211[0:7]), .rgt_op_bot(net_6381[0:7]),
     .reset_b_top(reset_b[335:320]), .reset_b_bot(reset_b[319:304]),
     .prog(prog), .pgate_top(pgate[335:320]),
     .pgate_bot(pgate[319:304]), .lft_op_top(net_7905[0:7]),
     .lft_op_bot(net_5607[0:7]), .bm_wdummymux_en_i(net_7586),
     .bot_op_bot(net_6225[0:7]), .bnr_op_top(net_6381[0:7]),
     .bnr_op_bot(net_6409[0:7]), .bnl_op_top(net_5607[0:7]),
     .bnl_op_bot(net_5635[0:7]), .sp12_v_t_top(net_4376[0:23]),
     .sp12_v_b_bot(net_7566[0:23]), .bm_init_i(net_7582),
     .sp12_h_r_top(net_4379[0:23]), .sp12_h_r_bot(net_4380[0:23]),
     .sp12_h_l_top(net_5507[0:23]), .sp12_h_l_bot(net_5479[0:23]),
     .sp4_v_t_top(net_4383[0:47]), .sp4_v_b_top(net_5511[0:47]),
     .sp4_v_b_bot(net_5483[0:47]), .sp4_r_v_b_top(net_4386[0:47]),
     .sp4_r_v_b_bot(net_4387[0:47]), .sp4_h_r_top(net_4388[0:47]),
     .sp4_h_r_bot(net_4389[0:47]), .sp4_h_l_top(net_5508[0:47]),
     .sp4_h_l_bot(net_5480[0:47]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(net_7581), .bm_sa_i(net_7583[0:7]),
     .bm_sclk_i(net_7584), .bm_sreb_i(net_7585),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_bufferx4 I1067 ( .in(ceb_i), .out(net_04420));
bram_bufferx4 I1069 ( .in(net_04420), .out(ceb_o));
bram_bufferx4 I1057 ( .in(net_4407), .out(tclk_o));
bram_bufferx4 I1080 ( .in(r_i), .out(net_4419));
bram_bufferx4 I1077 ( .in(tclk_i), .out(net_4407));
bram_bufferx4 I1078 ( .in(shift_i), .out(net_4429));
bram_bufferx4 I1056 ( .in(net_4415), .out(mode_o));
bram_bufferx4 I1079 ( .in(bs_en_i), .out(net_4427));
bram_bufferx4 I1054 ( .in(net_4419), .out(r_o));
bram_bufferx4 I1082 ( .in(update_i), .out(net_4431));
bram_bufferx4 I1076 ( .in(mode_i), .out(net_4415));
bram_bufferx4 I1081 ( .in(hiz_b_i), .out(net_4433));
bram_bufferx4 I1051 ( .in(net_4427), .out(bs_en_o));
bram_bufferx4 I1055 ( .in(net_4429), .out(shift_o));
bram_bufferx4 I1052 ( .in(net_4431), .out(update_o));
bram_bufferx4 I1053 ( .in(net_4433), .out(hiz_b_o));
ltile4rev I_05_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4437), .lft_op(slf_op_04_11[7:0]),
     .sp12_h_l(net_4583[0:23]), .sp4_h_l(net_4584[0:47]),
     .sp4_v_b(sp4_v_b_05_11[47:0]), .sp12_v_b(sp12_v_b_05_11[23:0]),
     .sp12_h_r(net_4443[0:23]), .sp4_h_r(net_4444[0:47]),
     .sp12_v_t(net_4445[0:23]), .sp4_v_t(net_4559[0:47]),
     .sp4_r_v_b(sp4_v_b_06_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7175[0:7]), .rgt_op(slf_op_06_11[7:0]),
     .bot_op(bot_op_05_11[7:0]), .bl(bl[287:234]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(carry_in_05_11), .purst(purst),
     .slf_op(slf_op_05_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_05_11[7:0]), .bnl_op(bnl_op_05_11[7:0]),
     .tnr_op(net_4461[0:7]), .tnl_op(net_7091[0:7]));
ltile4rev I_05_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4465), .lft_op(net_7091[0:7]),
     .sp12_h_l(net_4555[0:23]), .sp4_h_l(net_4556[0:47]),
     .sp4_v_b(net_4559[0:47]), .sp12_v_b(net_4445[0:23]),
     .sp12_h_r(net_4471[0:23]), .sp4_h_r(net_4472[0:47]),
     .sp12_v_t(net_4473[0:23]), .sp4_v_t(net_7163[0:47]),
     .sp4_r_v_b(net_4475[0:47]), .wl(wl[207:192]),
     .top_op(net_7147[0:7]), .rgt_op(net_4461[0:7]),
     .bot_op(slf_op_05_11[7:0]), .bl(bl[287:234]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_4437), .purst(purst), .slf_op(net_7175[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_06_11[7:0]),
     .bnl_op(slf_op_04_11[7:0]), .tnr_op(net_7738[0:7]),
     .tnl_op(net_7119[0:7]));
ltile4rev I_03_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4493), .lft_op(slf_op_02_11[7:0]),
     .sp12_h_l(net_6879[0:23]), .sp4_h_l(net_6880[0:47]),
     .sp4_v_b(sp4_v_b_03_11[47:0]), .sp12_v_b(sp12_v_b_03_11[23:0]),
     .sp12_h_r(net_4499[0:23]), .sp4_h_r(net_4500[0:47]),
     .sp12_v_t(net_4501[0:23]), .sp4_v_t(net_4643[0:47]),
     .sp4_r_v_b(sp4_v_b_04_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7007[0:7]), .rgt_op(slf_op_04_11[7:0]),
     .bot_op(bot_op_03_11[7:0]), .bl(bl[179:126]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(carry_in_03_11), .purst(purst),
     .slf_op(slf_op_03_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_03_11[7:0]), .bnl_op(bnl_op_03_11[7:0]),
     .tnr_op(net_7091[0:7]), .tnl_op(net_6923[0:7]));
ltile4rev I_03_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4521), .lft_op(net_6923[0:7]),
     .sp12_h_l(net_4639[0:23]), .sp4_h_l(net_4640[0:47]),
     .sp4_v_b(net_4643[0:47]), .sp12_v_b(net_4501[0:23]),
     .sp12_h_r(net_4527[0:23]), .sp4_h_r(net_4528[0:47]),
     .sp12_v_t(net_4529[0:23]), .sp4_v_t(net_6995[0:47]),
     .sp4_r_v_b(net_4531[0:47]), .wl(wl[207:192]),
     .top_op(net_6979[0:7]), .rgt_op(net_7091[0:7]),
     .bot_op(slf_op_03_11[7:0]), .bl(bl[179:126]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_4493), .purst(purst), .slf_op(net_7007[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_04_11[7:0]),
     .bnl_op(slf_op_02_11[7:0]), .tnr_op(net_7119[0:7]),
     .tnl_op(net_6951[0:7]));
ltile4rev I_04_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4549), .lft_op(net_7007[0:7]),
     .sp12_h_l(net_4527[0:23]), .sp4_h_l(net_4528[0:47]),
     .sp4_v_b(net_4531[0:47]), .sp12_v_b(net_4585[0:23]),
     .sp12_h_r(net_4555[0:23]), .sp4_h_r(net_4556[0:47]),
     .sp12_v_t(net_4557[0:23]), .sp4_v_t(net_7079[0:47]),
     .sp4_r_v_b(net_4559[0:47]), .wl(wl[207:192]),
     .top_op(net_7119[0:7]), .rgt_op(net_7175[0:7]),
     .bot_op(slf_op_04_11[7:0]), .bl(bl[233:180]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_4577), .purst(purst), .slf_op(net_7091[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_05_11[7:0]),
     .bnl_op(slf_op_03_11[7:0]), .tnr_op(net_7147[0:7]),
     .tnl_op(net_6979[0:7]));
ltile4rev I_04_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4577), .lft_op(slf_op_03_11[7:0]),
     .sp12_h_l(net_4499[0:23]), .sp4_h_l(net_4500[0:47]),
     .sp4_v_b(sp4_v_b_04_11[47:0]), .sp12_v_b(sp12_v_b_04_11[23:0]),
     .sp12_h_r(net_4583[0:23]), .sp4_h_r(net_4584[0:47]),
     .sp12_v_t(net_4585[0:23]), .sp4_v_t(net_4531[0:47]),
     .sp4_r_v_b(sp4_v_b_05_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7091[0:7]), .rgt_op(slf_op_05_11[7:0]),
     .bot_op(bot_op_04_11[7:0]), .bl(bl[233:180]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(carry_in_04_11), .purst(purst),
     .slf_op(slf_op_04_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_04_11[7:0]), .bnl_op(bnl_op_04_11[7:0]),
     .tnr_op(net_7175[0:7]), .tnl_op(net_7007[0:7]));
ltile4rev I_07_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4605), .lft_op(net_4461[0:7]),
     .sp12_h_l(net_7761[0:23]), .sp4_h_l(net_7770[0:47]),
     .sp4_v_b(net_7768[0:47]), .sp12_v_b(net_4725[0:23]),
     .sp12_h_r(net_4611[0:23]), .sp4_h_r(net_4612[0:47]),
     .sp12_v_t(net_4613[0:23]), .sp4_v_t(net_7682[0:47]),
     .sp4_r_v_b(net_4615[0:47]), .wl(wl[207:192]),
     .top_op(net_4617[0:7]), .rgt_op(net_4757[0:7]),
     .bot_op(slf_op_07_11[7:0]), .bl(bl[383:330]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_4717), .purst(purst), .slf_op(net_4729[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_08_11[7:0]),
     .bnl_op(slf_op_06_11[7:0]), .tnr_op(net_4785[0:7]),
     .tnl_op(net_7738[0:7]));
ltile4rev I_02_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4633), .lft_op(net_4701[0:7]),
     .sp12_h_l(net_4667[0:23]), .sp4_h_l(net_4668[0:47]),
     .sp4_v_b(net_4671[0:47]), .sp12_v_b(net_6881[0:23]),
     .sp12_h_r(net_4639[0:23]), .sp4_h_r(net_4640[0:47]),
     .sp12_v_t(net_4641[0:23]), .sp4_v_t(net_6911[0:47]),
     .sp4_r_v_b(net_4643[0:47]), .wl(wl[207:192]),
     .top_op(net_6951[0:7]), .rgt_op(net_7007[0:7]),
     .bot_op(slf_op_02_11[7:0]), .bl(bl[125:72]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_6873), .purst(purst), .slf_op(net_6923[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_03_11[7:0]),
     .bnl_op(slf_op_01_11[7:0]), .tnr_op(net_6979[0:7]),
     .tnl_op(net_4673[0:7]));
ltile4rev I_01_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4661), .lft_op({io_l_22[3], io_l_22[2], io_l_22[1],
     io_l_22[0], io_l_22[3], io_l_22[2], io_l_22[1], io_l_22[0]}),
     .sp12_h_l(net_4158[0:23]), .sp4_h_l(net_4157[0:47]),
     .sp4_v_b(net_4698[0:47]), .sp12_v_b(net_4697[0:23]),
     .sp12_h_r(net_4667[0:23]), .sp4_h_r(net_4668[0:47]),
     .sp12_v_t(net_4669[0:23]), .sp4_v_t(net_4670[0:47]),
     .sp4_r_v_b(net_4671[0:47]), .wl(wl[207:192]),
     .top_op(net_4673[0:7]), .rgt_op(net_6923[0:7]),
     .bot_op(slf_op_01_11[7:0]), .bl(bl[71:18]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_4689), .purst(purst), .slf_op(net_4701[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_02_11[7:0]),
     .bnl_op({slf_op_00_11[3], slf_op_00_11[2], slf_op_00_11[1],
     slf_op_00_11[0], slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0]}), .tnr_op(net_6951[0:7]),
     .tnl_op({io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0],
     io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0]}));
ltile4rev I_01_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4689), .lft_op({slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0], slf_op_00_11[3],
     slf_op_00_11[2], slf_op_00_11[1], slf_op_00_11[0]}),
     .sp12_h_l(net_4192[0:23]), .sp4_h_l(net_4191[0:47]),
     .sp4_v_b(sp4_v_b_01_11[47:0]), .sp12_v_b(sp12_v_b_01_11[23:0]),
     .sp12_h_r(net_4695[0:23]), .sp4_h_r(net_4696[0:47]),
     .sp12_v_t(net_4697[0:23]), .sp4_v_t(net_4698[0:47]),
     .sp4_r_v_b(sp4_v_b_02_11[47:0]), .wl(wl[191:176]),
     .top_op(net_4701[0:7]), .rgt_op(slf_op_02_11[7:0]),
     .bot_op(bot_op_01_11[7:0]), .bl(bl[71:18]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(carry_in_01_11), .purst(purst),
     .slf_op(slf_op_01_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_01_11[7:0]), .bnl_op(bnl_op_01_11[7:0]),
     .tnr_op(net_6923[0:7]), .tnl_op({io_l_22[3], io_l_22[2],
     io_l_22[1], io_l_22[0], io_l_22[3], io_l_22[2], io_l_22[1],
     io_l_22[0]}));
ltile4rev I_07_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4717), .lft_op(slf_op_06_11[7:0]),
     .sp12_h_l(net_7762[0:23]), .sp4_h_l(net_7771[0:47]),
     .sp4_v_b(sp4_v_b_07_11[47:0]), .sp12_v_b(sp12_v_b_07_11[23:0]),
     .sp12_h_r(net_4723[0:23]), .sp4_h_r(net_4724[0:47]),
     .sp12_v_t(net_4725[0:23]), .sp4_v_t(net_7768[0:47]),
     .sp4_r_v_b(sp4_v_b_08_11[47:0]), .wl(wl[191:176]),
     .top_op(net_4729[0:7]), .rgt_op(slf_op_08_11[7:0]),
     .bot_op(bot_op_07_11[7:0]), .bl(bl[383:330]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(carry_in_07_11), .purst(purst),
     .slf_op(slf_op_07_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_07_11[7:0]), .bnl_op(bnl_op_07_11[7:0]),
     .tnr_op(net_4757[0:7]), .tnl_op(net_4461[0:7]));
ltile4rev I_08_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4745), .lft_op(slf_op_07_11[7:0]),
     .sp12_h_l(net_4723[0:23]), .sp4_h_l(net_4724[0:47]),
     .sp4_v_b(sp4_v_b_08_11[47:0]), .sp12_v_b(sp12_v_b_08_11[23:0]),
     .sp12_h_r(net_4751[0:23]), .sp4_h_r(net_4752[0:47]),
     .sp12_v_t(net_4753[0:23]), .sp4_v_t(net_4615[0:47]),
     .sp4_r_v_b(sp4_v_b_09_11[47:0]), .wl(wl[191:176]),
     .top_op(net_4757[0:7]), .rgt_op(slf_op_09_11[7:0]),
     .bot_op(bot_op_08_11[7:0]), .bl(bl[437:384]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(carry_in_08_11), .purst(purst),
     .slf_op(slf_op_08_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_08_11[7:0]), .bnl_op(bnl_op_08_11[7:0]),
     .tnr_op(net_7259[0:7]), .tnl_op(net_4729[0:7]));
ltile4rev I_08_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4773), .lft_op(net_4729[0:7]),
     .sp12_h_l(net_4611[0:23]), .sp4_h_l(net_4612[0:47]),
     .sp4_v_b(net_4615[0:47]), .sp12_v_b(net_4753[0:23]),
     .sp12_h_r(net_4779[0:23]), .sp4_h_r(net_4780[0:47]),
     .sp12_v_t(net_4781[0:23]), .sp4_v_t(net_7219[0:47]),
     .sp4_r_v_b(net_4783[0:47]), .wl(wl[207:192]),
     .top_op(net_4785[0:7]), .rgt_op(net_7259[0:7]),
     .bot_op(slf_op_08_11[7:0]), .bl(bl[437:384]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_4745), .purst(purst), .slf_op(net_4757[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_09_11[7:0]),
     .bnl_op(slf_op_07_11[7:0]), .tnr_op(net_7287[0:7]),
     .tnl_op(net_4617[0:7]));
ltile4rev I_09_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_4801), .lft_op(net_4757[0:7]),
     .sp12_h_l(net_4779[0:23]), .sp4_h_l(net_4780[0:47]),
     .sp4_v_b(net_4783[0:47]), .sp12_v_b(net_4837[0:23]),
     .sp12_h_r(net_4807[0:23]), .sp4_h_r(net_4808[0:47]),
     .sp12_v_t(net_4809[0:23]), .sp4_v_t(net_7247[0:47]),
     .sp4_r_v_b(net_4811[0:47]), .wl(wl[207:192]),
     .top_op(net_7287[0:7]), .rgt_op(net_7343[0:7]),
     .bot_op(slf_op_09_11[7:0]), .bl(bl[491:438]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_4829), .purst(purst), .slf_op(net_7259[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_10_11[7:0]),
     .bnl_op(slf_op_08_11[7:0]), .tnr_op(net_7315[0:7]),
     .tnl_op(net_4785[0:7]));
ltile4rev I_09_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_4829), .lft_op(slf_op_08_11[7:0]),
     .sp12_h_l(net_4751[0:23]), .sp4_h_l(net_4752[0:47]),
     .sp4_v_b(sp4_v_b_09_11[47:0]), .sp12_v_b(sp12_v_b_09_11[23:0]),
     .sp12_h_r(net_4835[0:23]), .sp4_h_r(net_4836[0:47]),
     .sp12_v_t(net_4837[0:23]), .sp4_v_t(net_4783[0:47]),
     .sp4_r_v_b(sp4_v_b_10_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7259[0:7]), .rgt_op(slf_op_10_11[7:0]),
     .bot_op(bot_op_09_11[7:0]), .bl(bl[491:438]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(carry_in_09_11), .purst(purst),
     .slf_op(slf_op_09_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_09_11[7:0]), .bnl_op(bnl_op_09_11[7:0]),
     .tnr_op(net_7343[0:7]), .tnl_op(net_4757[0:7]));
ltile4rev I_05_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_4857), .lft_op(net_4963[0:7]),
     .sp12_h_l(net_5003[0:23]), .sp4_h_l(net_5004[0:47]),
     .sp4_v_b(net_5007[0:47]), .sp12_v_b(net_7049[0:23]),
     .sp12_h_r(net_4863[0:23]), .sp4_h_r(net_4864[0:47]),
     .sp12_v_t(net_4865[0:23]), .sp4_v_t(net_4979[0:47]),
     .sp4_r_v_b(net_4867[0:47]), .wl(wl[255:240]),
     .top_op(net_6363[0:7]), .rgt_op(net_7688[0:7]),
     .bot_op(net_5019[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_7041), .purst(purst), .slf_op(net_4991[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_7037[0:7]),
     .bnl_op(net_4935[0:7]), .tnr_op(net_6223[0:7]),
     .tnl_op(net_6279[0:7]));
ltile4rev I_05_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4885), .lft_op(net_6279[0:7]),
     .sp12_h_l(net_4975[0:23]), .sp4_h_l(net_4976[0:47]),
     .sp4_v_b(net_4979[0:47]), .sp12_v_b(net_4865[0:23]),
     .sp12_h_r(net_4891[0:23]), .sp4_h_r(net_4892[0:47]),
     .sp12_v_t(net_4893[0:23]), .sp4_v_t(net_6351[0:47]),
     .sp4_r_v_b(net_4895[0:47]), .wl(wl[271:256]),
     .top_op(net_6335[0:7]), .rgt_op(net_6223[0:7]),
     .bot_op(net_4991[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_4857), .purst(purst), .slf_op(net_6363[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_7688[0:7]),
     .bnl_op(net_4963[0:7]), .tnr_op(net_7614[0:7]),
     .tnl_op(net_6307[0:7]));
ltile4rev I_03_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_4913), .lft_op(net_5131[0:7]),
     .sp12_h_l(net_5059[0:23]), .sp4_h_l(net_5060[0:47]),
     .sp4_v_b(net_5063[0:47]), .sp12_v_b(net_7105[0:23]),
     .sp12_h_r(net_4919[0:23]), .sp4_h_r(net_4920[0:47]),
     .sp12_v_t(net_4921[0:23]), .sp4_v_t(net_5091[0:47]),
     .sp4_r_v_b(net_4923[0:47]), .wl(wl[255:240]),
     .top_op(net_6195[0:7]), .rgt_op(net_4963[0:7]),
     .bot_op(net_5075[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_7097), .purst(purst), .slf_op(net_5103[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_4935[0:7]),
     .bnl_op(net_5159[0:7]), .tnr_op(net_6279[0:7]),
     .tnl_op(net_6111[0:7]));
ltile4rev I_03_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4941), .lft_op(net_6111[0:7]),
     .sp12_h_l(net_5087[0:23]), .sp4_h_l(net_5088[0:47]),
     .sp4_v_b(net_5091[0:47]), .sp12_v_b(net_4921[0:23]),
     .sp12_h_r(net_4947[0:23]), .sp4_h_r(net_4948[0:47]),
     .sp12_v_t(net_4949[0:23]), .sp4_v_t(net_6183[0:47]),
     .sp4_r_v_b(net_4951[0:47]), .wl(wl[271:256]),
     .top_op(net_6167[0:7]), .rgt_op(net_6279[0:7]),
     .bot_op(net_5103[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_4913), .purst(purst), .slf_op(net_6195[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_4963[0:7]),
     .bnl_op(net_5131[0:7]), .tnr_op(net_6307[0:7]),
     .tnl_op(net_6139[0:7]));
ltile4rev I_04_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_4969), .lft_op(net_6195[0:7]),
     .sp12_h_l(net_4947[0:23]), .sp4_h_l(net_4948[0:47]),
     .sp4_v_b(net_4951[0:47]), .sp12_v_b(net_5005[0:23]),
     .sp12_h_r(net_4975[0:23]), .sp4_h_r(net_4976[0:47]),
     .sp12_v_t(net_4977[0:23]), .sp4_v_t(net_6267[0:47]),
     .sp4_r_v_b(net_4979[0:47]), .wl(wl[271:256]),
     .top_op(net_6307[0:7]), .rgt_op(net_6363[0:7]),
     .bot_op(net_4963[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_4997), .purst(purst), .slf_op(net_6279[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_4991[0:7]),
     .bnl_op(net_5103[0:7]), .tnr_op(net_6335[0:7]),
     .tnl_op(net_6167[0:7]));
ltile4rev I_04_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_4997), .lft_op(net_5103[0:7]),
     .sp12_h_l(net_4919[0:23]), .sp4_h_l(net_4920[0:47]),
     .sp4_v_b(net_4923[0:47]), .sp12_v_b(net_7133[0:23]),
     .sp12_h_r(net_5003[0:23]), .sp4_h_r(net_5004[0:47]),
     .sp12_v_t(net_5005[0:23]), .sp4_v_t(net_4951[0:47]),
     .sp4_r_v_b(net_5007[0:47]), .wl(wl[255:240]),
     .top_op(net_6279[0:7]), .rgt_op(net_4991[0:7]),
     .bot_op(net_4935[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_7125), .purst(purst), .slf_op(net_4963[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5019[0:7]),
     .bnl_op(net_5075[0:7]), .tnr_op(net_6363[0:7]),
     .tnl_op(net_6195[0:7]));
ltile4rev I_07_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5025), .lft_op(net_6223[0:7]),
     .sp12_h_l(net_7637[0:23]), .sp4_h_l(net_7646[0:47]),
     .sp4_v_b(net_7644[0:47]), .sp12_v_b(net_5173[0:23]),
     .sp12_h_r(net_5031[0:23]), .sp4_h_r(net_5032[0:47]),
     .sp12_v_t(net_5033[0:23]), .sp4_v_t(net_7597[0:47]),
     .sp4_r_v_b(net_5035[0:47]), .wl(wl[271:256]),
     .top_op(net_5037[0:7]), .rgt_op(net_5205[0:7]),
     .bot_op(net_7193[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_5165), .purst(purst), .slf_op(net_5177[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_7277[0:7]),
     .bnl_op(net_7688[0:7]), .tnr_op(net_5233[0:7]),
     .tnl_op(net_7614[0:7]));
ltile4rev I_02_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5053), .lft_op(net_6941[0:7]),
     .sp12_h_l(net_5143[0:23]), .sp4_h_l(net_5144[0:47]),
     .sp4_v_b(net_5147[0:47]), .sp12_v_b(net_6965[0:23]),
     .sp12_h_r(net_5059[0:23]), .sp4_h_r(net_5060[0:47]),
     .sp12_v_t(net_5061[0:23]), .sp4_v_t(net_5119[0:47]),
     .sp4_r_v_b(net_5063[0:47]), .wl(wl[255:240]),
     .top_op(net_6111[0:7]), .rgt_op(net_5103[0:7]),
     .bot_op(net_5159[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_6957), .purst(purst), .slf_op(net_5131[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5075[0:7]),
     .bnl_op(net_6913[0:7]), .tnr_op(net_6195[0:7]),
     .tnl_op(net_5149[0:7]));
ltile4rev I_02_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5081), .lft_op(net_5149[0:7]),
     .sp12_h_l(net_5115[0:23]), .sp4_h_l(net_5116[0:47]),
     .sp4_v_b(net_5119[0:47]), .sp12_v_b(net_5061[0:23]),
     .sp12_h_r(net_5087[0:23]), .sp4_h_r(net_5088[0:47]),
     .sp12_v_t(net_5089[0:23]), .sp4_v_t(net_6099[0:47]),
     .sp4_r_v_b(net_5091[0:47]), .wl(wl[271:256]),
     .top_op(net_6139[0:7]), .rgt_op(net_6195[0:7]),
     .bot_op(net_5131[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_5053), .purst(purst), .slf_op(net_6111[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5103[0:7]),
     .bnl_op(net_6941[0:7]), .tnr_op(net_6167[0:7]),
     .tnl_op(net_5121[0:7]));
ltile4rev I_01_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5109), .lft_op({io_l_30[3], io_l_30[2], io_l_30[1],
     io_l_30[0], io_l_30[3], io_l_30[2], io_l_30[1], io_l_30[0]}),
     .sp12_h_l(net_4090[0:23]), .sp4_h_l(net_4089[0:47]),
     .sp4_v_b(net_5146[0:47]), .sp12_v_b(net_5145[0:23]),
     .sp12_h_r(net_5115[0:23]), .sp4_h_r(net_5116[0:47]),
     .sp12_v_t(net_5117[0:23]), .sp4_v_t(net_5118[0:47]),
     .sp4_r_v_b(net_5119[0:47]), .wl(wl[271:256]),
     .top_op(net_5121[0:7]), .rgt_op(net_6111[0:7]),
     .bot_op(net_6941[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_5137), .purst(purst), .slf_op(net_5149[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5131[0:7]),
     .bnl_op({io_l_28[3], io_l_28[2], io_l_28[1], io_l_28[0],
     io_l_28[3], io_l_28[2], io_l_28[1], io_l_28[0]}),
     .tnr_op(net_6139[0:7]), .tnl_op({io_l_32[3], io_l_32[2],
     io_l_32[1], io_l_32[0], io_l_32[3], io_l_32[2], io_l_32[1],
     io_l_32[0]}));
ltile4rev I_01_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5137), .lft_op({io_l_28[3], io_l_28[2], io_l_28[1],
     io_l_28[0], io_l_28[3], io_l_28[2], io_l_28[1], io_l_28[0]}),
     .sp12_h_l(net_4124[0:23]), .sp4_h_l(net_4123[0:47]),
     .sp4_v_b(net_6938[0:47]), .sp12_v_b(net_6937[0:23]),
     .sp12_h_r(net_5143[0:23]), .sp4_h_r(net_5144[0:47]),
     .sp12_v_t(net_5145[0:23]), .sp4_v_t(net_5146[0:47]),
     .sp4_r_v_b(net_5147[0:47]), .wl(wl[255:240]),
     .top_op(net_5149[0:7]), .rgt_op(net_5131[0:7]),
     .bot_op(net_6913[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_6929), .purst(purst), .slf_op(net_6941[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5159[0:7]),
     .bnl_op({io_l_26[3], io_l_26[2], io_l_26[1], io_l_26[0],
     io_l_26[3], io_l_26[2], io_l_26[1], io_l_26[0]}),
     .tnr_op(net_6111[0:7]), .tnl_op({io_l_30[3], io_l_30[2],
     io_l_30[1], io_l_30[0], io_l_30[3], io_l_30[2], io_l_30[1],
     io_l_30[0]}));
ltile4rev I_07_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5165), .lft_op(net_7688[0:7]),
     .sp12_h_l(net_7638[0:23]), .sp4_h_l(net_7647[0:47]),
     .sp4_v_b(net_7645[0:47]), .sp12_v_b(net_7189[0:23]),
     .sp12_h_r(net_5171[0:23]), .sp4_h_r(net_5172[0:47]),
     .sp12_v_t(net_5173[0:23]), .sp4_v_t(net_7644[0:47]),
     .sp4_r_v_b(net_5175[0:47]), .wl(wl[255:240]),
     .top_op(net_5177[0:7]), .rgt_op(net_7277[0:7]),
     .bot_op(net_7221[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_7181), .purst(purst), .slf_op(net_7193[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_7249[0:7]),
     .bnl_op(net_7037[0:7]), .tnr_op(net_5205[0:7]),
     .tnl_op(net_6223[0:7]));
ltile4rev I_08_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5193), .lft_op(net_7193[0:7]),
     .sp12_h_l(net_5171[0:23]), .sp4_h_l(net_5172[0:47]),
     .sp4_v_b(net_5175[0:47]), .sp12_v_b(net_7273[0:23]),
     .sp12_h_r(net_5199[0:23]), .sp4_h_r(net_5200[0:47]),
     .sp12_v_t(net_5201[0:23]), .sp4_v_t(net_5035[0:47]),
     .sp4_r_v_b(net_5203[0:47]), .wl(wl[255:240]),
     .top_op(net_5205[0:7]), .rgt_op(net_5243[0:7]),
     .bot_op(net_7249[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_7265), .purst(purst), .slf_op(net_7277[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5215[0:7]),
     .bnl_op(net_7221[0:7]), .tnr_op(net_6447[0:7]),
     .tnl_op(net_5177[0:7]));
ltile4rev I_08_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5221), .lft_op(net_5177[0:7]),
     .sp12_h_l(net_5031[0:23]), .sp4_h_l(net_5032[0:47]),
     .sp4_v_b(net_5035[0:47]), .sp12_v_b(net_5201[0:23]),
     .sp12_h_r(net_5227[0:23]), .sp4_h_r(net_5228[0:47]),
     .sp12_v_t(net_5229[0:23]), .sp4_v_t(net_6407[0:47]),
     .sp4_r_v_b(net_5231[0:47]), .wl(wl[271:256]),
     .top_op(net_5233[0:7]), .rgt_op(net_6447[0:7]),
     .bot_op(net_7277[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_5193), .purst(purst), .slf_op(net_5205[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5243[0:7]),
     .bnl_op(net_7193[0:7]), .tnr_op(net_6475[0:7]),
     .tnl_op(net_5037[0:7]));
ltile4rev I_09_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5249), .lft_op(net_5205[0:7]),
     .sp12_h_l(net_5227[0:23]), .sp4_h_l(net_5228[0:47]),
     .sp4_v_b(net_5231[0:47]), .sp12_v_b(net_5285[0:23]),
     .sp12_h_r(net_5255[0:23]), .sp4_h_r(net_5256[0:47]),
     .sp12_v_t(net_5257[0:23]), .sp4_v_t(net_6435[0:47]),
     .sp4_r_v_b(net_5259[0:47]), .wl(wl[271:256]),
     .top_op(net_6475[0:7]), .rgt_op(net_6531[0:7]),
     .bot_op(net_5243[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_5277), .purst(purst), .slf_op(net_6447[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5271[0:7]),
     .bnl_op(net_7277[0:7]), .tnr_op(net_6503[0:7]),
     .tnl_op(net_5233[0:7]));
ltile4rev I_09_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5277), .lft_op(net_7277[0:7]),
     .sp12_h_l(net_5199[0:23]), .sp4_h_l(net_5200[0:47]),
     .sp4_v_b(net_5203[0:47]), .sp12_v_b(net_7301[0:23]),
     .sp12_h_r(net_5283[0:23]), .sp4_h_r(net_5284[0:47]),
     .sp12_v_t(net_5285[0:23]), .sp4_v_t(net_5231[0:47]),
     .sp4_r_v_b(net_5287[0:47]), .wl(wl[255:240]),
     .top_op(net_6447[0:7]), .rgt_op(net_5271[0:7]),
     .bot_op(net_5215[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_7293), .purst(purst), .slf_op(net_5243[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5299[0:7]),
     .bnl_op(net_7249[0:7]), .tnr_op(net_6531[0:7]),
     .tnl_op(net_5205[0:7]));
ltile4rev I_11_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5305), .lft_op(net_5271[0:7]),
     .sp12_h_l(net_5367[0:23]), .sp4_h_l(net_5368[0:47]),
     .sp4_v_b(net_5371[0:47]), .sp12_v_b(net_7497[0:23]),
     .sp12_h_r(net_5311[0:23]), .sp4_h_r(net_5312[0:47]),
     .sp12_v_t(net_5313[0:23]), .sp4_v_t(net_5399[0:47]),
     .sp4_r_v_b(net_5315[0:47]), .wl(wl[255:240]),
     .top_op(net_6615[0:7]), .rgt_op(slf_op_12_15[7:0]),
     .bot_op(net_5383[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_7489), .purst(purst), .slf_op(net_5411[0:7]),
     .pgate(pgate[255:240]), .bnr_op(slf_op_12_14[7:0]),
     .bnl_op(net_5299[0:7]), .tnr_op(slf_op_12_16[7:0]),
     .tnl_op(net_6531[0:7]));
ltile4rev I_12_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_6667), .lft_op(net_6615[0:7]),
     .sp12_h_l(net_5451[0:23]), .sp4_h_l(net_5452[0:47]),
     .sp4_v_b(net_5455[0:47]), .sp12_v_b(net_5425[0:23]),
     .sp12_h_r(sp12_h_r_12_16[23:0]), .sp4_h_r(sp4_h_r_12_16[47:0]),
     .sp12_v_t(net_5341[0:23]), .sp4_v_t(net_6547[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_16[47:0]), .wl(wl[271:256]),
     .top_op(slf_op_12_17[7:0]), .rgt_op(rgt_op_12_16[7:0]),
     .bot_op(slf_op_12_15[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_5417), .purst(purst), .slf_op(slf_op_12_16[7:0]),
     .pgate(pgate[271:256]), .bnr_op(rgt_op_12_15[7:0]),
     .bnl_op(net_5411[0:7]), .tnr_op(rgt_op_12_17[7:0]),
     .tnl_op(net_6643[0:7]));
ltile4rev I_10_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5361), .lft_op(net_5243[0:7]),
     .sp12_h_l(net_5283[0:23]), .sp4_h_l(net_5284[0:47]),
     .sp4_v_b(net_5287[0:47]), .sp12_v_b(net_7441[0:23]),
     .sp12_h_r(net_5367[0:23]), .sp4_h_r(net_5368[0:47]),
     .sp12_v_t(net_5369[0:23]), .sp4_v_t(net_5259[0:47]),
     .sp4_r_v_b(net_5371[0:47]), .wl(wl[255:240]),
     .top_op(net_6531[0:7]), .rgt_op(net_5411[0:7]),
     .bot_op(net_5299[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_7433), .purst(purst), .slf_op(net_5271[0:7]),
     .pgate(pgate[255:240]), .bnr_op(net_5383[0:7]),
     .bnl_op(net_5215[0:7]), .tnr_op(net_6615[0:7]),
     .tnl_op(net_6447[0:7]));
ltile4rev I_10_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5389), .lft_op(net_6447[0:7]),
     .sp12_h_l(net_5255[0:23]), .sp4_h_l(net_5256[0:47]),
     .sp4_v_b(net_5259[0:47]), .sp12_v_b(net_5369[0:23]),
     .sp12_h_r(net_5395[0:23]), .sp4_h_r(net_5396[0:47]),
     .sp12_v_t(net_5397[0:23]), .sp4_v_t(net_6519[0:47]),
     .sp4_r_v_b(net_5399[0:47]), .wl(wl[271:256]),
     .top_op(net_6503[0:7]), .rgt_op(net_6615[0:7]),
     .bot_op(net_5271[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_5361), .purst(purst), .slf_op(net_6531[0:7]),
     .pgate(pgate[271:256]), .bnr_op(net_5411[0:7]),
     .bnl_op(net_5243[0:7]), .tnr_op(net_6643[0:7]),
     .tnl_op(net_6475[0:7]));
ltile4rev I_12_15 ( .vdd_cntl(vdd_cntl[255:240]), .prog(prog),
     .carry_out(net_5417), .lft_op(net_5411[0:7]),
     .sp12_h_l(net_5311[0:23]), .sp4_h_l(net_5312[0:47]),
     .sp4_v_b(net_5315[0:47]), .sp12_v_b(net_7385[0:23]),
     .sp12_h_r(sp12_h_r_12_15[23:0]), .sp4_h_r(sp4_h_r_12_15[47:0]),
     .sp12_v_t(net_5425[0:23]), .sp4_v_t(net_5455[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_15[47:0]), .wl(wl[255:240]),
     .top_op(slf_op_12_16[7:0]), .rgt_op(rgt_op_12_15[7:0]),
     .bot_op(slf_op_12_14[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[255:240]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_7377), .purst(purst), .slf_op(slf_op_12_15[7:0]),
     .pgate(pgate[255:240]), .bnr_op(rgt_op_12_14[7:0]),
     .bnl_op(net_5383[0:7]), .tnr_op(rgt_op_12_16[7:0]),
     .tnl_op(net_6615[0:7]));
ltile4rev I_11_16 ( .vdd_cntl(vdd_cntl[271:256]), .prog(prog),
     .carry_out(net_5445), .lft_op(net_6531[0:7]),
     .sp12_h_l(net_5395[0:23]), .sp4_h_l(net_5396[0:47]),
     .sp4_v_b(net_5399[0:47]), .sp12_v_b(net_5313[0:23]),
     .sp12_h_r(net_5451[0:23]), .sp4_h_r(net_5452[0:47]),
     .sp12_v_t(net_5453[0:23]), .sp4_v_t(net_6603[0:47]),
     .sp4_r_v_b(net_5455[0:47]), .wl(wl[271:256]),
     .top_op(net_6643[0:7]), .rgt_op(slf_op_12_16[7:0]),
     .bot_op(net_5411[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[271:256]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_5305), .purst(purst), .slf_op(net_6615[0:7]),
     .pgate(pgate[271:256]), .bnr_op(slf_op_12_15[7:0]),
     .bnl_op(net_5271[0:7]), .tnr_op(slf_op_12_17[7:0]),
     .tnl_op(net_6503[0:7]));
ltile4rev I_05_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5473), .lft_op(net_5579[0:7]),
     .sp12_h_l(net_5619[0:23]), .sp4_h_l(net_5620[0:47]),
     .sp4_v_b(net_5623[0:47]), .sp12_v_b(net_6237[0:23]),
     .sp12_h_r(net_5479[0:23]), .sp4_h_r(net_5480[0:47]),
     .sp12_v_t(net_5481[0:23]), .sp4_v_t(net_5595[0:47]),
     .sp4_r_v_b(net_5483[0:47]), .wl(wl[319:304]),
     .top_op(net_7905[0:7]), .rgt_op(net_7552[0:7]),
     .bot_op(net_5635[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_6229), .purst(purst), .slf_op(net_5607[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_6225[0:7]),
     .bnl_op(net_5551[0:7]), .tnr_op(net_8177[0:7]),
     .tnl_op(net_7837[0:7]));
ltile4rev I_05_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_5501), .lft_op(net_7837[0:7]),
     .sp12_h_l(net_5591[0:23]), .sp4_h_l(net_5592[0:47]),
     .sp4_v_b(net_5595[0:47]), .sp12_v_b(net_5481[0:23]),
     .sp12_h_r(net_5507[0:23]), .sp4_h_r(net_5508[0:47]),
     .sp12_v_t(net_5509[0:23]), .sp4_v_t(net_8171[0:47]),
     .sp4_r_v_b(net_5511[0:47]), .wl(wl[335:320]), .top_op({io_t_8[3],
     io_t_8[2], io_t_8[1], io_t_8[0], io_t_8[3], io_t_8[2], io_t_8[1],
     io_t_8[0]}), .rgt_op(net_8177[0:7]), .bot_op(net_5607[0:7]),
     .bl(bl[287:234]), .reset_b(reset_b[335:320]),
     .glb_netwk(glb_netwk_04[7:0]), .carry_in(net_5473), .purst(purst),
     .slf_op(net_7905[0:7]), .pgate(pgate[335:320]),
     .bnr_op(net_7552[0:7]), .bnl_op(net_5579[0:7]),
     .tnr_op({io_t_10[3], io_t_10[2], io_t_10[1], io_t_10[0],
     io_t_10[3], io_t_10[2], io_t_10[1], io_t_10[0]}),
     .tnl_op({io_t_6[3], io_t_6[2], io_t_6[1], io_t_6[0], io_t_6[3],
     io_t_6[2], io_t_6[1], io_t_6[0]}));
ltile4rev I_03_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5529), .lft_op(net_5747[0:7]),
     .sp12_h_l(net_5675[0:23]), .sp4_h_l(net_5676[0:47]),
     .sp4_v_b(net_5679[0:47]), .sp12_v_b(net_6293[0:23]),
     .sp12_h_r(net_5535[0:23]), .sp4_h_r(net_5536[0:47]),
     .sp12_v_t(net_5537[0:23]), .sp4_v_t(net_5707[0:47]),
     .sp4_r_v_b(net_5539[0:47]), .wl(wl[319:304]),
     .top_op(net_7871[0:7]), .rgt_op(net_5579[0:7]),
     .bot_op(net_5691[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_6285), .purst(purst), .slf_op(net_5719[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5551[0:7]),
     .bnl_op(net_5775[0:7]), .tnr_op(net_7837[0:7]),
     .tnl_op(net_8143[0:7]));
ltile4rev I_03_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8243), .lft_op(net_8143[0:7]),
     .sp12_h_l(net_5703[0:23]), .sp4_h_l(net_5704[0:47]),
     .sp4_v_b(net_5707[0:47]), .sp12_v_b(net_5537[0:23]),
     .sp12_h_r(net_5563[0:23]), .sp4_h_r(net_5564[0:47]),
     .sp12_v_t(net_5565[0:23]), .sp4_v_t(net_7831[0:47]),
     .sp4_r_v_b(net_5567[0:47]), .wl(wl[335:320]), .top_op({io_t_4[3],
     io_t_4[2], io_t_4[1], io_t_4[0], io_t_4[3], io_t_4[2], io_t_4[1],
     io_t_4[0]}), .rgt_op(net_7837[0:7]), .bot_op(net_5719[0:7]),
     .bl(bl[179:126]), .reset_b(reset_b[335:320]),
     .glb_netwk(glb_netwk_02[7:0]), .carry_in(net_5529), .purst(purst),
     .slf_op(net_7871[0:7]), .pgate(pgate[335:320]),
     .bnr_op(net_5579[0:7]), .bnl_op(net_5747[0:7]),
     .tnr_op({io_t_6[3], io_t_6[2], io_t_6[1], io_t_6[0], io_t_6[3],
     io_t_6[2], io_t_6[1], io_t_6[0]}), .tnl_op({io_t_2[3], io_t_2[2],
     io_t_2[1], io_t_2[0], io_t_2[3], io_t_2[2], io_t_2[1],
     io_t_2[0]}));
ltile4rev I_04_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8254), .lft_op(net_7871[0:7]),
     .sp12_h_l(net_5563[0:23]), .sp4_h_l(net_5564[0:47]),
     .sp4_v_b(net_5567[0:47]), .sp12_v_b(net_5621[0:23]),
     .sp12_h_r(net_5591[0:23]), .sp4_h_r(net_5592[0:47]),
     .sp12_v_t(net_5593[0:23]), .sp4_v_t(net_7899[0:47]),
     .sp4_r_v_b(net_5595[0:47]), .wl(wl[335:320]), .top_op({io_t_6[3],
     io_t_6[2], io_t_6[1], io_t_6[0], io_t_6[3], io_t_6[2], io_t_6[1],
     io_t_6[0]}), .rgt_op(net_7905[0:7]), .bot_op(net_5579[0:7]),
     .bl(bl[233:180]), .reset_b(reset_b[335:320]),
     .glb_netwk(glb_netwk_03[7:0]), .carry_in(net_5613), .purst(purst),
     .slf_op(net_7837[0:7]), .pgate(pgate[335:320]),
     .bnr_op(net_5607[0:7]), .bnl_op(net_5719[0:7]),
     .tnr_op({io_t_8[3], io_t_8[2], io_t_8[1], io_t_8[0], io_t_8[3],
     io_t_8[2], io_t_8[1], io_t_8[0]}), .tnl_op({io_t_4[3], io_t_4[2],
     io_t_4[1], io_t_4[0], io_t_4[3], io_t_4[2], io_t_4[1],
     io_t_4[0]}));
ltile4rev I_04_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5613), .lft_op(net_5719[0:7]),
     .sp12_h_l(net_5535[0:23]), .sp4_h_l(net_5536[0:47]),
     .sp4_v_b(net_5539[0:47]), .sp12_v_b(net_6321[0:23]),
     .sp12_h_r(net_5619[0:23]), .sp4_h_r(net_5620[0:47]),
     .sp12_v_t(net_5621[0:23]), .sp4_v_t(net_5567[0:47]),
     .sp4_r_v_b(net_5623[0:47]), .wl(wl[319:304]),
     .top_op(net_7837[0:7]), .rgt_op(net_5607[0:7]),
     .bot_op(net_5551[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_6313), .purst(purst), .slf_op(net_5579[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5635[0:7]),
     .bnl_op(net_5691[0:7]), .tnr_op(net_7905[0:7]),
     .tnl_op(net_7871[0:7]));
ltile4rev I_07_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8246), .lft_op(net_8177[0:7]),
     .sp12_h_l(net_4379[0:23]), .sp4_h_l(net_4388[0:47]),
     .sp4_v_b(net_4386[0:47]), .sp12_v_b(net_5789[0:23]),
     .sp12_h_r(net_5647[0:23]), .sp4_h_r(net_5648[0:47]),
     .sp12_v_t(net_5649[0:23]), .sp4_v_t(net_7933[0:47]),
     .sp4_r_v_b(net_5651[0:47]), .wl(wl[335:320]), .top_op({io_t_12[3],
     io_t_12[2], io_t_12[1], io_t_12[0], io_t_12[3], io_t_12[2],
     io_t_12[1], io_t_12[0]}), .rgt_op(net_7939[0:7]),
     .bot_op(net_6381[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_5781), .purst(purst), .slf_op(net_8211[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_6465[0:7]),
     .bnl_op(net_7552[0:7]), .tnr_op({io_t_14[3], io_t_14[2],
     io_t_14[1], io_t_14[0], io_t_14[3], io_t_14[2], io_t_14[1],
     io_t_14[0]}), .tnl_op({io_t_10[3], io_t_10[2], io_t_10[1],
     io_t_10[0], io_t_10[3], io_t_10[2], io_t_10[1], io_t_10[0]}));
ltile4rev I_02_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5669), .lft_op(net_6129[0:7]),
     .sp12_h_l(net_5759[0:23]), .sp4_h_l(net_5760[0:47]),
     .sp4_v_b(net_5763[0:47]), .sp12_v_b(net_6153[0:23]),
     .sp12_h_r(net_5675[0:23]), .sp4_h_r(net_5676[0:47]),
     .sp12_v_t(net_5677[0:23]), .sp4_v_t(net_5735[0:47]),
     .sp4_r_v_b(net_5679[0:47]), .wl(wl[319:304]),
     .top_op(net_8143[0:7]), .rgt_op(net_5719[0:7]),
     .bot_op(net_5775[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_6145), .purst(purst), .slf_op(net_5747[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5691[0:7]),
     .bnl_op(net_6101[0:7]), .tnr_op(net_7871[0:7]),
     .tnl_op(net_5765[0:7]));
ltile4rev I_02_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_5697), .lft_op(net_5765[0:7]),
     .sp12_h_l(net_5731[0:23]), .sp4_h_l(net_5732[0:47]),
     .sp4_v_b(net_5735[0:47]), .sp12_v_b(net_5677[0:23]),
     .sp12_h_r(net_5703[0:23]), .sp4_h_r(net_5704[0:47]),
     .sp12_v_t(net_5705[0:23]), .sp4_v_t(net_7865[0:47]),
     .sp4_r_v_b(net_5707[0:47]), .wl(wl[335:320]), .top_op({io_t_2[3],
     io_t_2[2], io_t_2[1], io_t_2[0], io_t_2[3], io_t_2[2], io_t_2[1],
     io_t_2[0]}), .rgt_op(net_7871[0:7]), .bot_op(net_5747[0:7]),
     .bl(bl[125:72]), .reset_b(reset_b[335:320]),
     .glb_netwk(glb_netwk_01[7:0]), .carry_in(net_5669), .purst(purst),
     .slf_op(net_8143[0:7]), .pgate(pgate[335:320]),
     .bnr_op(net_5719[0:7]), .bnl_op(net_6129[0:7]),
     .tnr_op({io_t_4[3], io_t_4[2], io_t_4[1], io_t_4[0], io_t_4[3],
     io_t_4[2], io_t_4[1], io_t_4[0]}), .tnl_op({io_t_0[3], io_t_0[2],
     io_t_0[1], io_t_0[0], io_t_0[3], io_t_0[2], io_t_0[1],
     io_t_0[0]}));
ltile4rev I_01_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_5725), .lft_op({io_l_38[3], io_l_38[2], io_l_38[1],
     io_l_38[0], io_l_38[3], io_l_38[2], io_l_38[1], io_l_38[0]}),
     .sp12_h_l(net_4022[0:23]), .sp4_h_l(net_4021[0:47]),
     .sp4_v_b(net_5762[0:47]), .sp12_v_b(net_5761[0:23]),
     .sp12_h_r(net_5731[0:23]), .sp4_h_r(net_5732[0:47]),
     .sp12_v_t(net_5733[0:23]), .sp4_v_t(net_8137[0:47]),
     .sp4_r_v_b(net_5735[0:47]), .wl(wl[335:320]), .top_op({io_t_0[3],
     io_t_0[2], io_t_0[1], io_t_0[0], io_t_0[3], io_t_0[2], io_t_0[1],
     io_t_0[0]}), .rgt_op(net_8143[0:7]), .bot_op(net_6129[0:7]),
     .bl(bl[71:18]), .reset_b(reset_b[335:320]),
     .glb_netwk(glb_netwk_00[7:0]), .carry_in(net_5753), .purst(purst),
     .slf_op(net_5765[0:7]), .pgate(pgate[335:320]),
     .bnr_op(net_5747[0:7]), .bnl_op({io_l_36[3], io_l_36[2],
     io_l_36[1], io_l_36[0], io_l_36[3], io_l_36[2], io_l_36[1],
     io_l_36[0]}), .tnr_op({io_t_2[3], io_t_2[2], io_t_2[1], io_t_2[0],
     io_t_2[3], io_t_2[2], io_t_2[1], io_t_2[0]}), .tnl_op({tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}));
ltile4rev I_01_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5753), .lft_op({io_l_36[3], io_l_36[2], io_l_36[1],
     io_l_36[0], io_l_36[3], io_l_36[2], io_l_36[1], io_l_36[0]}),
     .sp12_h_l(net_4056[0:23]), .sp4_h_l(net_4055[0:47]),
     .sp4_v_b(net_6126[0:47]), .sp12_v_b(net_6125[0:23]),
     .sp12_h_r(net_5759[0:23]), .sp4_h_r(net_5760[0:47]),
     .sp12_v_t(net_5761[0:23]), .sp4_v_t(net_5762[0:47]),
     .sp4_r_v_b(net_5763[0:47]), .wl(wl[319:304]),
     .top_op(net_5765[0:7]), .rgt_op(net_5747[0:7]),
     .bot_op(net_6101[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_6117), .purst(purst), .slf_op(net_6129[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5775[0:7]),
     .bnl_op({io_l_34[3], io_l_34[2], io_l_34[1], io_l_34[0],
     io_l_34[3], io_l_34[2], io_l_34[1], io_l_34[0]}),
     .tnr_op(net_8143[0:7]), .tnl_op({io_l_38[3], io_l_38[2],
     io_l_38[1], io_l_38[0], io_l_38[3], io_l_38[2], io_l_38[1],
     io_l_38[0]}));
ltile4rev I_07_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5781), .lft_op(net_7552[0:7]),
     .sp12_h_l(net_4380[0:23]), .sp4_h_l(net_4389[0:47]),
     .sp4_v_b(net_4387[0:47]), .sp12_v_b(net_6377[0:23]),
     .sp12_h_r(net_5787[0:23]), .sp4_h_r(net_5788[0:47]),
     .sp12_v_t(net_5789[0:23]), .sp4_v_t(net_4386[0:47]),
     .sp4_r_v_b(net_5791[0:47]), .wl(wl[319:304]),
     .top_op(net_8211[0:7]), .rgt_op(net_6465[0:7]),
     .bot_op(net_6409[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_6369), .purst(purst), .slf_op(net_6381[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_6437[0:7]),
     .bnl_op(net_6225[0:7]), .tnr_op(net_7939[0:7]),
     .tnl_op(net_8177[0:7]));
ltile4rev I_08_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5809), .lft_op(net_6381[0:7]),
     .sp12_h_l(net_5787[0:23]), .sp4_h_l(net_5788[0:47]),
     .sp4_v_b(net_5791[0:47]), .sp12_v_b(net_6461[0:23]),
     .sp12_h_r(net_5815[0:23]), .sp4_h_r(net_5816[0:47]),
     .sp12_v_t(net_5817[0:23]), .sp4_v_t(net_5651[0:47]),
     .sp4_r_v_b(net_5819[0:47]), .wl(wl[319:304]),
     .top_op(net_7939[0:7]), .rgt_op(net_5859[0:7]),
     .bot_op(net_6437[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_6453), .purst(purst), .slf_op(net_6465[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5831[0:7]),
     .bnl_op(net_6409[0:7]), .tnr_op(net_7973[0:7]),
     .tnl_op(net_8211[0:7]));
ltile4rev I_08_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_5837), .lft_op(net_8211[0:7]),
     .sp12_h_l(net_5647[0:23]), .sp4_h_l(net_5648[0:47]),
     .sp4_v_b(net_5651[0:47]), .sp12_v_b(net_5817[0:23]),
     .sp12_h_r(net_5843[0:23]), .sp4_h_r(net_5844[0:47]),
     .sp12_v_t(net_5845[0:23]), .sp4_v_t(net_7967[0:47]),
     .sp4_r_v_b(net_5847[0:47]), .wl(wl[335:320]), .top_op({io_t_14[3],
     io_t_14[2], io_t_14[1], io_t_14[0], io_t_14[3], io_t_14[2],
     io_t_14[1], io_t_14[0]}), .rgt_op(net_7973[0:7]),
     .bot_op(net_6465[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_5809), .purst(purst), .slf_op(net_7939[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5859[0:7]),
     .bnl_op(net_6381[0:7]), .tnr_op({io_t_16[3], io_t_16[2],
     io_t_16[1], io_t_16[0], io_t_16[3], io_t_16[2], io_t_16[1],
     io_t_16[0]}), .tnl_op({io_t_12[3], io_t_12[2], io_t_12[1],
     io_t_12[0], io_t_12[3], io_t_12[2], io_t_12[1], io_t_12[0]}));
ltile4rev I_09_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_5865), .lft_op(net_7939[0:7]),
     .sp12_h_l(net_5843[0:23]), .sp4_h_l(net_5844[0:47]),
     .sp4_v_b(net_5847[0:47]), .sp12_v_b(net_5901[0:23]),
     .sp12_h_r(net_5871[0:23]), .sp4_h_r(net_5872[0:47]),
     .sp12_v_t(net_5873[0:23]), .sp4_v_t(net_8001[0:47]),
     .sp4_r_v_b(net_5875[0:47]), .wl(wl[335:320]), .top_op({io_t_16[3],
     io_t_16[2], io_t_16[1], io_t_16[0], io_t_16[3], io_t_16[2],
     io_t_16[1], io_t_16[0]}), .rgt_op(net_8007[0:7]),
     .bot_op(net_5859[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_5893), .purst(purst), .slf_op(net_7973[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_5887[0:7]),
     .bnl_op(net_6465[0:7]), .tnr_op({io_t_18[3], io_t_18[2],
     io_t_18[1], io_t_18[0], io_t_18[3], io_t_18[2], io_t_18[1],
     io_t_18[0]}), .tnl_op({io_t_14[3], io_t_14[2], io_t_14[1],
     io_t_14[0], io_t_14[3], io_t_14[2], io_t_14[1], io_t_14[0]}));
ltile4rev I_09_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5893), .lft_op(net_6465[0:7]),
     .sp12_h_l(net_5815[0:23]), .sp4_h_l(net_5816[0:47]),
     .sp4_v_b(net_5819[0:47]), .sp12_v_b(net_6489[0:23]),
     .sp12_h_r(net_5899[0:23]), .sp4_h_r(net_5900[0:47]),
     .sp12_v_t(net_5901[0:23]), .sp4_v_t(net_5847[0:47]),
     .sp4_r_v_b(net_5903[0:47]), .wl(wl[319:304]),
     .top_op(net_7973[0:7]), .rgt_op(net_5887[0:7]),
     .bot_op(net_5831[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_6481), .purst(purst), .slf_op(net_5859[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5915[0:7]),
     .bnl_op(net_6437[0:7]), .tnr_op(net_8007[0:7]),
     .tnl_op(net_7939[0:7]));
ltile4rev I_11_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5921), .lft_op(net_5887[0:7]),
     .sp12_h_l(net_5983[0:23]), .sp4_h_l(net_5984[0:47]),
     .sp4_v_b(net_5987[0:47]), .sp12_v_b(net_6685[0:23]),
     .sp12_h_r(net_5927[0:23]), .sp4_h_r(net_5928[0:47]),
     .sp12_v_t(net_5929[0:23]), .sp4_v_t(net_6015[0:47]),
     .sp4_r_v_b(net_5931[0:47]), .wl(wl[319:304]),
     .top_op(net_8041[0:7]), .rgt_op(slf_op_12_19[7:0]),
     .bot_op(net_5999[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_6677), .purst(purst), .slf_op(net_6027[0:7]),
     .pgate(pgate[319:304]), .bnr_op(slf_op_12_18[7:0]),
     .bnl_op(net_5915[0:7]), .tnr_op(slf_op_12_20[7:0]),
     .tnl_op(net_8007[0:7]));
ltile4rev I_12_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_8257), .lft_op(net_8041[0:7]),
     .sp12_h_l(net_6067[0:23]), .sp4_h_l(net_6068[0:47]),
     .sp4_v_b(net_6071[0:47]), .sp12_v_b(net_6041[0:23]),
     .sp12_h_r(sp12_h_r_12_20[23:0]), .sp4_h_r(sp4_h_r_12_20[47:0]),
     .sp12_v_t(net_5957[0:23]), .sp4_v_t(net_8103[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_20[47:0]), .wl(wl[335:320]),
     .top_op({slf_op_12_21[3], slf_op_12_21[2], slf_op_12_21[1],
     slf_op_12_21[0], slf_op_12_21[3], slf_op_12_21[2],
     slf_op_12_21[1], slf_op_12_21[0]}), .rgt_op(rgt_op_12_20[7:0]),
     .bot_op(slf_op_12_19[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_6033), .purst(purst), .slf_op(slf_op_12_20[7:0]),
     .pgate(pgate[335:320]), .bnr_op(rgt_op_12_19[7:0]),
     .bnl_op(net_6027[0:7]), .tnr_op({tnr_op_12_20[3], tnr_op_12_20[2],
     tnr_op_12_20[1], tnr_op_12_20[0], tnr_op_12_20[3],
     tnr_op_12_20[2], tnr_op_12_20[1], tnr_op_12_20[0]}),
     .tnl_op({io_t_20[3], io_t_20[2], io_t_20[1], io_t_20[0],
     io_t_20[3], io_t_20[2], io_t_20[1], io_t_20[0]}));
ltile4rev I_10_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_5977), .lft_op(net_5859[0:7]),
     .sp12_h_l(net_5899[0:23]), .sp4_h_l(net_5900[0:47]),
     .sp4_v_b(net_5903[0:47]), .sp12_v_b(net_6629[0:23]),
     .sp12_h_r(net_5983[0:23]), .sp4_h_r(net_5984[0:47]),
     .sp12_v_t(net_5985[0:23]), .sp4_v_t(net_5875[0:47]),
     .sp4_r_v_b(net_5987[0:47]), .wl(wl[319:304]),
     .top_op(net_8007[0:7]), .rgt_op(net_6027[0:7]),
     .bot_op(net_5915[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_6621), .purst(purst), .slf_op(net_5887[0:7]),
     .pgate(pgate[319:304]), .bnr_op(net_5999[0:7]),
     .bnl_op(net_5831[0:7]), .tnr_op(net_8041[0:7]),
     .tnl_op(net_7973[0:7]));
ltile4rev I_10_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_6005), .lft_op(net_7973[0:7]),
     .sp12_h_l(net_5871[0:23]), .sp4_h_l(net_5872[0:47]),
     .sp4_v_b(net_5875[0:47]), .sp12_v_b(net_5985[0:23]),
     .sp12_h_r(net_6011[0:23]), .sp4_h_r(net_6012[0:47]),
     .sp12_v_t(net_6013[0:23]), .sp4_v_t(net_8035[0:47]),
     .sp4_r_v_b(net_6015[0:47]), .wl(wl[335:320]), .top_op({io_t_18[3],
     io_t_18[2], io_t_18[1], io_t_18[0], io_t_18[3], io_t_18[2],
     io_t_18[1], io_t_18[0]}), .rgt_op(net_8041[0:7]),
     .bot_op(net_5887[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_5977), .purst(purst), .slf_op(net_8007[0:7]),
     .pgate(pgate[335:320]), .bnr_op(net_6027[0:7]),
     .bnl_op(net_5859[0:7]), .tnr_op({io_t_20[3], io_t_20[2],
     io_t_20[1], io_t_20[0], io_t_20[3], io_t_20[2], io_t_20[1],
     io_t_20[0]}), .tnl_op({io_t_16[3], io_t_16[2], io_t_16[1],
     io_t_16[0], io_t_16[3], io_t_16[2], io_t_16[1], io_t_16[0]}));
ltile4rev I_12_19 ( .vdd_cntl(vdd_cntl[319:304]), .prog(prog),
     .carry_out(net_6033), .lft_op(net_6027[0:7]),
     .sp12_h_l(net_5927[0:23]), .sp4_h_l(net_5928[0:47]),
     .sp4_v_b(net_5931[0:47]), .sp12_v_b(net_6573[0:23]),
     .sp12_h_r(sp12_h_r_12_19[23:0]), .sp4_h_r(sp4_h_r_12_19[47:0]),
     .sp12_v_t(net_6041[0:23]), .sp4_v_t(net_6071[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_19[47:0]), .wl(wl[319:304]),
     .top_op(slf_op_12_20[7:0]), .rgt_op(rgt_op_12_19[7:0]),
     .bot_op(slf_op_12_18[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[319:304]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_6565), .purst(purst), .slf_op(slf_op_12_19[7:0]),
     .pgate(pgate[319:304]), .bnr_op(rgt_op_12_18[7:0]),
     .bnl_op(net_5999[0:7]), .tnr_op(rgt_op_12_20[7:0]),
     .tnl_op(net_8041[0:7]));
ltile4rev I_11_20 ( .vdd_cntl(vdd_cntl[335:320]), .prog(prog),
     .carry_out(net_6061), .lft_op(net_8007[0:7]),
     .sp12_h_l(net_6011[0:23]), .sp4_h_l(net_6012[0:47]),
     .sp4_v_b(net_6015[0:47]), .sp12_v_b(net_5929[0:23]),
     .sp12_h_r(net_6067[0:23]), .sp4_h_r(net_6068[0:47]),
     .sp12_v_t(net_6069[0:23]), .sp4_v_t(net_8069[0:47]),
     .sp4_r_v_b(net_6071[0:47]), .wl(wl[335:320]), .top_op({io_t_20[3],
     io_t_20[2], io_t_20[1], io_t_20[0], io_t_20[3], io_t_20[2],
     io_t_20[1], io_t_20[0]}), .rgt_op(slf_op_12_20[7:0]),
     .bot_op(net_6027[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[335:320]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_5921), .purst(purst), .slf_op(net_8041[0:7]),
     .pgate(pgate[335:320]), .bnr_op(slf_op_12_19[7:0]),
     .bnl_op(net_5887[0:7]), .tnr_op({slf_op_12_21[3], slf_op_12_21[2],
     slf_op_12_21[1], slf_op_12_21[0], slf_op_12_21[3],
     slf_op_12_21[2], slf_op_12_21[1], slf_op_12_21[0]}),
     .tnl_op({io_t_18[3], io_t_18[2], io_t_18[1], io_t_18[0],
     io_t_18[3], io_t_18[2], io_t_18[1], io_t_18[0]}));
ltile4rev I_01_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6089), .lft_op({io_l_32[3], io_l_32[2], io_l_32[1],
     io_l_32[0], io_l_32[3], io_l_32[2], io_l_32[1], io_l_32[0]}),
     .sp12_h_l(net_4328[0:23]), .sp4_h_l(net_4327[0:47]),
     .sp4_v_b(net_5118[0:47]), .sp12_v_b(net_5117[0:23]),
     .sp12_h_r(net_6095[0:23]), .sp4_h_r(net_6096[0:47]),
     .sp12_v_t(net_6097[0:23]), .sp4_v_t(net_6098[0:47]),
     .sp4_r_v_b(net_6099[0:47]), .wl(wl[287:272]),
     .top_op(net_6101[0:7]), .rgt_op(net_6139[0:7]),
     .bot_op(net_5149[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_5109), .purst(purst), .slf_op(net_5121[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6111[0:7]),
     .bnl_op({io_l_30[3], io_l_30[2], io_l_30[1], io_l_30[0],
     io_l_30[3], io_l_30[2], io_l_30[1], io_l_30[0]}),
     .tnr_op(net_5775[0:7]), .tnl_op({io_l_34[3], io_l_34[2],
     io_l_34[1], io_l_34[0], io_l_34[3], io_l_34[2], io_l_34[1],
     io_l_34[0]}));
ltile4rev I_01_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6117), .lft_op({io_l_34[3], io_l_34[2], io_l_34[1],
     io_l_34[0], io_l_34[3], io_l_34[2], io_l_34[1], io_l_34[0]}),
     .sp12_h_l(net_4294[0:23]), .sp4_h_l(net_4293[0:47]),
     .sp4_v_b(net_6098[0:47]), .sp12_v_b(net_6097[0:23]),
     .sp12_h_r(net_6123[0:23]), .sp4_h_r(net_6124[0:47]),
     .sp12_v_t(net_6125[0:23]), .sp4_v_t(net_6126[0:47]),
     .sp4_r_v_b(net_6127[0:47]), .wl(wl[303:288]),
     .top_op(net_6129[0:7]), .rgt_op(net_5775[0:7]),
     .bot_op(net_5121[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_6089), .purst(purst), .slf_op(net_6101[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6139[0:7]),
     .bnl_op({io_l_32[3], io_l_32[2], io_l_32[1], io_l_32[0],
     io_l_32[3], io_l_32[2], io_l_32[1], io_l_32[0]}),
     .tnr_op(net_5747[0:7]), .tnl_op({io_l_36[3], io_l_36[2],
     io_l_36[1], io_l_36[0], io_l_36[3], io_l_36[2], io_l_36[1],
     io_l_36[0]}));
ltile4rev I_02_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6145), .lft_op(net_6101[0:7]),
     .sp12_h_l(net_6123[0:23]), .sp4_h_l(net_6124[0:47]),
     .sp4_v_b(net_6127[0:47]), .sp12_v_b(net_6181[0:23]),
     .sp12_h_r(net_6151[0:23]), .sp4_h_r(net_6152[0:47]),
     .sp12_v_t(net_6153[0:23]), .sp4_v_t(net_5763[0:47]),
     .sp4_r_v_b(net_6155[0:47]), .wl(wl[303:288]),
     .top_op(net_5747[0:7]), .rgt_op(net_5691[0:7]),
     .bot_op(net_6139[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_6173), .purst(purst), .slf_op(net_5775[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6167[0:7]),
     .bnl_op(net_5121[0:7]), .tnr_op(net_5719[0:7]),
     .tnl_op(net_6129[0:7]));
ltile4rev I_02_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6173), .lft_op(net_5121[0:7]),
     .sp12_h_l(net_6095[0:23]), .sp4_h_l(net_6096[0:47]),
     .sp4_v_b(net_6099[0:47]), .sp12_v_b(net_5089[0:23]),
     .sp12_h_r(net_6179[0:23]), .sp4_h_r(net_6180[0:47]),
     .sp12_v_t(net_6181[0:23]), .sp4_v_t(net_6127[0:47]),
     .sp4_r_v_b(net_6183[0:47]), .wl(wl[287:272]),
     .top_op(net_5775[0:7]), .rgt_op(net_6167[0:7]),
     .bot_op(net_6111[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_5081), .purst(purst), .slf_op(net_6139[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6195[0:7]),
     .bnl_op(net_5149[0:7]), .tnr_op(net_5691[0:7]),
     .tnl_op(net_6101[0:7]));
ltile4rev I_05_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6201), .lft_op(net_6307[0:7]),
     .sp12_h_l(net_6347[0:23]), .sp4_h_l(net_6348[0:47]),
     .sp4_v_b(net_6351[0:47]), .sp12_v_b(net_4893[0:23]),
     .sp12_h_r(net_6207[0:23]), .sp4_h_r(net_6208[0:47]),
     .sp12_v_t(net_6209[0:23]), .sp4_v_t(net_6323[0:47]),
     .sp4_r_v_b(net_6211[0:47]), .wl(wl[287:272]),
     .top_op(net_5635[0:7]), .rgt_op(net_7614[0:7]),
     .bot_op(net_6363[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_4885), .purst(purst), .slf_op(net_6335[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6223[0:7]),
     .bnl_op(net_6279[0:7]), .tnr_op(net_6225[0:7]),
     .tnl_op(net_5551[0:7]));
ltile4rev I_05_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6229), .lft_op(net_5551[0:7]),
     .sp12_h_l(net_6319[0:23]), .sp4_h_l(net_6320[0:47]),
     .sp4_v_b(net_6323[0:47]), .sp12_v_b(net_6209[0:23]),
     .sp12_h_r(net_6235[0:23]), .sp4_h_r(net_6236[0:47]),
     .sp12_v_t(net_6237[0:23]), .sp4_v_t(net_5623[0:47]),
     .sp4_r_v_b(net_6239[0:47]), .wl(wl[303:288]),
     .top_op(net_5607[0:7]), .rgt_op(net_6225[0:7]),
     .bot_op(net_6335[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_6201), .purst(purst), .slf_op(net_5635[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_7614[0:7]),
     .bnl_op(net_6307[0:7]), .tnr_op(net_7552[0:7]),
     .tnl_op(net_5579[0:7]));
ltile4rev I_03_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6257), .lft_op(net_6139[0:7]),
     .sp12_h_l(net_6179[0:23]), .sp4_h_l(net_6180[0:47]),
     .sp4_v_b(net_6183[0:47]), .sp12_v_b(net_4949[0:23]),
     .sp12_h_r(net_6263[0:23]), .sp4_h_r(net_6264[0:47]),
     .sp12_v_t(net_6265[0:23]), .sp4_v_t(net_6155[0:47]),
     .sp4_r_v_b(net_6267[0:47]), .wl(wl[287:272]),
     .top_op(net_5691[0:7]), .rgt_op(net_6307[0:7]),
     .bot_op(net_6195[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_4941), .purst(purst), .slf_op(net_6167[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6279[0:7]),
     .bnl_op(net_6111[0:7]), .tnr_op(net_5551[0:7]),
     .tnl_op(net_5775[0:7]));
ltile4rev I_03_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6285), .lft_op(net_5775[0:7]),
     .sp12_h_l(net_6151[0:23]), .sp4_h_l(net_6152[0:47]),
     .sp4_v_b(net_6155[0:47]), .sp12_v_b(net_6265[0:23]),
     .sp12_h_r(net_6291[0:23]), .sp4_h_r(net_6292[0:47]),
     .sp12_v_t(net_6293[0:23]), .sp4_v_t(net_5679[0:47]),
     .sp4_r_v_b(net_6295[0:47]), .wl(wl[303:288]),
     .top_op(net_5719[0:7]), .rgt_op(net_5551[0:7]),
     .bot_op(net_6167[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_6257), .purst(purst), .slf_op(net_5691[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6307[0:7]),
     .bnl_op(net_6139[0:7]), .tnr_op(net_5579[0:7]),
     .tnl_op(net_5747[0:7]));
ltile4rev I_04_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6313), .lft_op(net_5691[0:7]),
     .sp12_h_l(net_6291[0:23]), .sp4_h_l(net_6292[0:47]),
     .sp4_v_b(net_6295[0:47]), .sp12_v_b(net_6349[0:23]),
     .sp12_h_r(net_6319[0:23]), .sp4_h_r(net_6320[0:47]),
     .sp12_v_t(net_6321[0:23]), .sp4_v_t(net_5539[0:47]),
     .sp4_r_v_b(net_6323[0:47]), .wl(wl[303:288]),
     .top_op(net_5579[0:7]), .rgt_op(net_5635[0:7]),
     .bot_op(net_6307[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_6341), .purst(purst), .slf_op(net_5551[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6335[0:7]),
     .bnl_op(net_6167[0:7]), .tnr_op(net_5607[0:7]),
     .tnl_op(net_5719[0:7]));
ltile4rev I_04_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6341), .lft_op(net_6167[0:7]),
     .sp12_h_l(net_6263[0:23]), .sp4_h_l(net_6264[0:47]),
     .sp4_v_b(net_6267[0:47]), .sp12_v_b(net_4977[0:23]),
     .sp12_h_r(net_6347[0:23]), .sp4_h_r(net_6348[0:47]),
     .sp12_v_t(net_6349[0:23]), .sp4_v_t(net_6295[0:47]),
     .sp4_r_v_b(net_6351[0:47]), .wl(wl[287:272]),
     .top_op(net_5551[0:7]), .rgt_op(net_6335[0:7]),
     .bot_op(net_6279[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_4969), .purst(purst), .slf_op(net_6307[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6363[0:7]),
     .bnl_op(net_6195[0:7]), .tnr_op(net_5635[0:7]),
     .tnl_op(net_5691[0:7]));
ltile4rev I_07_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6369), .lft_op(net_6225[0:7]),
     .sp12_h_l(net_7591[0:23]), .sp4_h_l(net_7594[0:47]),
     .sp4_v_b(net_7596[0:47]), .sp12_v_b(net_6405[0:23]),
     .sp12_h_r(net_6375[0:23]), .sp4_h_r(net_6376[0:47]),
     .sp12_v_t(net_6377[0:23]), .sp4_v_t(net_4387[0:47]),
     .sp4_r_v_b(net_6379[0:47]), .wl(wl[303:288]),
     .top_op(net_6381[0:7]), .rgt_op(net_6437[0:7]),
     .bot_op(net_5037[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_6397), .purst(purst), .slf_op(net_6409[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_5233[0:7]),
     .bnl_op(net_7614[0:7]), .tnr_op(net_6465[0:7]),
     .tnl_op(net_7552[0:7]));
ltile4rev I_07_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6397), .lft_op(net_7614[0:7]),
     .sp12_h_l(net_7592[0:23]), .sp4_h_l(net_7593[0:47]),
     .sp4_v_b(net_7597[0:47]), .sp12_v_b(net_5033[0:23]),
     .sp12_h_r(net_6403[0:23]), .sp4_h_r(net_6404[0:47]),
     .sp12_v_t(net_6405[0:23]), .sp4_v_t(net_7596[0:47]),
     .sp4_r_v_b(net_6407[0:47]), .wl(wl[287:272]),
     .top_op(net_6409[0:7]), .rgt_op(net_5233[0:7]),
     .bot_op(net_5177[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_5025), .purst(purst), .slf_op(net_5037[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_5205[0:7]),
     .bnl_op(net_6223[0:7]), .tnr_op(net_6437[0:7]),
     .tnl_op(net_6225[0:7]));
ltile4rev I_08_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6425), .lft_op(net_5037[0:7]),
     .sp12_h_l(net_6403[0:23]), .sp4_h_l(net_6404[0:47]),
     .sp4_v_b(net_6407[0:47]), .sp12_v_b(net_5229[0:23]),
     .sp12_h_r(net_6431[0:23]), .sp4_h_r(net_6432[0:47]),
     .sp12_v_t(net_6433[0:23]), .sp4_v_t(net_6379[0:47]),
     .sp4_r_v_b(net_6435[0:47]), .wl(wl[287:272]),
     .top_op(net_6437[0:7]), .rgt_op(net_6475[0:7]),
     .bot_op(net_5205[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_5221), .purst(purst), .slf_op(net_5233[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6447[0:7]),
     .bnl_op(net_5177[0:7]), .tnr_op(net_5831[0:7]),
     .tnl_op(net_6409[0:7]));
ltile4rev I_08_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6453), .lft_op(net_6409[0:7]),
     .sp12_h_l(net_6375[0:23]), .sp4_h_l(net_6376[0:47]),
     .sp4_v_b(net_6379[0:47]), .sp12_v_b(net_6433[0:23]),
     .sp12_h_r(net_6459[0:23]), .sp4_h_r(net_6460[0:47]),
     .sp12_v_t(net_6461[0:23]), .sp4_v_t(net_5791[0:47]),
     .sp4_r_v_b(net_6463[0:47]), .wl(wl[303:288]),
     .top_op(net_6465[0:7]), .rgt_op(net_5831[0:7]),
     .bot_op(net_5233[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_6425), .purst(purst), .slf_op(net_6437[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6475[0:7]),
     .bnl_op(net_5037[0:7]), .tnr_op(net_5859[0:7]),
     .tnl_op(net_6381[0:7]));
ltile4rev I_09_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6481), .lft_op(net_6437[0:7]),
     .sp12_h_l(net_6459[0:23]), .sp4_h_l(net_6460[0:47]),
     .sp4_v_b(net_6463[0:47]), .sp12_v_b(net_6517[0:23]),
     .sp12_h_r(net_6487[0:23]), .sp4_h_r(net_6488[0:47]),
     .sp12_v_t(net_6489[0:23]), .sp4_v_t(net_5819[0:47]),
     .sp4_r_v_b(net_6491[0:47]), .wl(wl[303:288]),
     .top_op(net_5859[0:7]), .rgt_op(net_5915[0:7]),
     .bot_op(net_6475[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_6509), .purst(purst), .slf_op(net_5831[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6503[0:7]),
     .bnl_op(net_5233[0:7]), .tnr_op(net_5887[0:7]),
     .tnl_op(net_6465[0:7]));
ltile4rev I_09_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6509), .lft_op(net_5233[0:7]),
     .sp12_h_l(net_6431[0:23]), .sp4_h_l(net_6432[0:47]),
     .sp4_v_b(net_6435[0:47]), .sp12_v_b(net_5257[0:23]),
     .sp12_h_r(net_6515[0:23]), .sp4_h_r(net_6516[0:47]),
     .sp12_v_t(net_6517[0:23]), .sp4_v_t(net_6463[0:47]),
     .sp4_r_v_b(net_6519[0:47]), .wl(wl[287:272]),
     .top_op(net_5831[0:7]), .rgt_op(net_6503[0:7]),
     .bot_op(net_6447[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_5249), .purst(purst), .slf_op(net_6475[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6531[0:7]),
     .bnl_op(net_5205[0:7]), .tnr_op(net_5915[0:7]),
     .tnl_op(net_6437[0:7]));
ltile4rev I_11_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6537), .lft_op(net_6503[0:7]),
     .sp12_h_l(net_6599[0:23]), .sp4_h_l(net_6600[0:47]),
     .sp4_v_b(net_6603[0:47]), .sp12_v_b(net_5453[0:23]),
     .sp12_h_r(net_6543[0:23]), .sp4_h_r(net_6544[0:47]),
     .sp12_v_t(net_6545[0:23]), .sp4_v_t(net_6631[0:47]),
     .sp4_r_v_b(net_6547[0:47]), .wl(wl[287:272]),
     .top_op(net_5999[0:7]), .rgt_op(slf_op_12_17[7:0]),
     .bot_op(net_6615[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_5445), .purst(purst), .slf_op(net_6643[0:7]),
     .pgate(pgate[287:272]), .bnr_op(slf_op_12_16[7:0]),
     .bnl_op(net_6531[0:7]), .tnr_op(slf_op_12_18[7:0]),
     .tnl_op(net_5915[0:7]));
ltile4rev I_12_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6565), .lft_op(net_5999[0:7]),
     .sp12_h_l(net_6683[0:23]), .sp4_h_l(net_6684[0:47]),
     .sp4_v_b(net_6687[0:47]), .sp12_v_b(net_6657[0:23]),
     .sp12_h_r(sp12_h_r_12_18[23:0]), .sp4_h_r(sp4_h_r_12_18[47:0]),
     .sp12_v_t(net_6573[0:23]), .sp4_v_t(net_5931[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_18[47:0]), .wl(wl[303:288]),
     .top_op(slf_op_12_19[7:0]), .rgt_op(rgt_op_12_18[7:0]),
     .bot_op(slf_op_12_17[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_6649), .purst(purst), .slf_op(slf_op_12_18[7:0]),
     .pgate(pgate[303:288]), .bnr_op(rgt_op_12_17[7:0]),
     .bnl_op(net_6643[0:7]), .tnr_op(rgt_op_12_19[7:0]),
     .tnl_op(net_6027[0:7]));
ltile4rev I_10_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6593), .lft_op(net_6475[0:7]),
     .sp12_h_l(net_6515[0:23]), .sp4_h_l(net_6516[0:47]),
     .sp4_v_b(net_6519[0:47]), .sp12_v_b(net_5397[0:23]),
     .sp12_h_r(net_6599[0:23]), .sp4_h_r(net_6600[0:47]),
     .sp12_v_t(net_6601[0:23]), .sp4_v_t(net_6491[0:47]),
     .sp4_r_v_b(net_6603[0:47]), .wl(wl[287:272]),
     .top_op(net_5915[0:7]), .rgt_op(net_6643[0:7]),
     .bot_op(net_6531[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_5389), .purst(purst), .slf_op(net_6503[0:7]),
     .pgate(pgate[287:272]), .bnr_op(net_6615[0:7]),
     .bnl_op(net_6447[0:7]), .tnr_op(net_5999[0:7]),
     .tnl_op(net_5831[0:7]));
ltile4rev I_10_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6621), .lft_op(net_5831[0:7]),
     .sp12_h_l(net_6487[0:23]), .sp4_h_l(net_6488[0:47]),
     .sp4_v_b(net_6491[0:47]), .sp12_v_b(net_6601[0:23]),
     .sp12_h_r(net_6627[0:23]), .sp4_h_r(net_6628[0:47]),
     .sp12_v_t(net_6629[0:23]), .sp4_v_t(net_5903[0:47]),
     .sp4_r_v_b(net_6631[0:47]), .wl(wl[303:288]),
     .top_op(net_5887[0:7]), .rgt_op(net_5999[0:7]),
     .bot_op(net_6503[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_6593), .purst(purst), .slf_op(net_5915[0:7]),
     .pgate(pgate[303:288]), .bnr_op(net_6643[0:7]),
     .bnl_op(net_6475[0:7]), .tnr_op(net_6027[0:7]),
     .tnl_op(net_5859[0:7]));
ltile4rev I_12_17 ( .vdd_cntl(vdd_cntl[287:272]), .prog(prog),
     .carry_out(net_6649), .lft_op(net_6643[0:7]),
     .sp12_h_l(net_6543[0:23]), .sp4_h_l(net_6544[0:47]),
     .sp4_v_b(net_6547[0:47]), .sp12_v_b(net_5341[0:23]),
     .sp12_h_r(sp12_h_r_12_17[23:0]), .sp4_h_r(sp4_h_r_12_17[47:0]),
     .sp12_v_t(net_6657[0:23]), .sp4_v_t(net_6687[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_17[47:0]), .wl(wl[287:272]),
     .top_op(slf_op_12_18[7:0]), .rgt_op(rgt_op_12_17[7:0]),
     .bot_op(slf_op_12_16[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[287:272]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_6667), .purst(purst), .slf_op(slf_op_12_17[7:0]),
     .pgate(pgate[287:272]), .bnr_op(rgt_op_12_16[7:0]),
     .bnl_op(net_6615[0:7]), .tnr_op(rgt_op_12_18[7:0]),
     .tnl_op(net_5999[0:7]));
ltile4rev I_11_18 ( .vdd_cntl(vdd_cntl[303:288]), .prog(prog),
     .carry_out(net_6677), .lft_op(net_5915[0:7]),
     .sp12_h_l(net_6627[0:23]), .sp4_h_l(net_6628[0:47]),
     .sp4_v_b(net_6631[0:47]), .sp12_v_b(net_6545[0:23]),
     .sp12_h_r(net_6683[0:23]), .sp4_h_r(net_6684[0:47]),
     .sp12_v_t(net_6685[0:23]), .sp4_v_t(net_5987[0:47]),
     .sp4_r_v_b(net_6687[0:47]), .wl(wl[303:288]),
     .top_op(net_6027[0:7]), .rgt_op(slf_op_12_18[7:0]),
     .bot_op(net_6643[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[303:288]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_6537), .purst(purst), .slf_op(net_5999[0:7]),
     .pgate(pgate[303:288]), .bnr_op(slf_op_12_17[7:0]),
     .bnl_op(net_6503[0:7]), .tnr_op(slf_op_12_19[7:0]),
     .tnl_op(net_5887[0:7]));
ltile4rev I_11_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_6705), .lft_op(slf_op_10_11[7:0]),
     .sp12_h_l(net_6767[0:23]), .sp4_h_l(net_6768[0:47]),
     .sp4_v_b(sp4_v_b_11_11[47:0]), .sp12_v_b(sp12_v_b_11_11[23:0]),
     .sp12_h_r(net_6711[0:23]), .sp4_h_r(net_6712[0:47]),
     .sp12_v_t(net_6713[0:23]), .sp4_v_t(net_6799[0:47]),
     .sp4_r_v_b(sp4_v_b_12_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7427[0:7]), .rgt_op(slf_op_12_11[7:0]),
     .bot_op(bot_op_11_11[7:0]), .bl(bl[599:546]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(carry_in_11_11), .purst(purst),
     .slf_op(slf_op_11_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_11_11[7:0]), .bnl_op(bnl_op_11_11[7:0]),
     .tnr_op(slf_op_12_12[7:0]), .tnl_op(net_7343[0:7]));
ltile4rev I_12_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_7479), .lft_op(net_7427[0:7]),
     .sp12_h_l(net_6851[0:23]), .sp4_h_l(net_6852[0:47]),
     .sp4_v_b(net_6855[0:47]), .sp12_v_b(net_6825[0:23]),
     .sp12_h_r(sp12_h_r_12_12[23:0]), .sp4_h_r(sp4_h_r_12_12[47:0]),
     .sp12_v_t(net_6741[0:23]), .sp4_v_t(net_7359[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_12[47:0]), .wl(wl[207:192]),
     .top_op(slf_op_12_13[7:0]), .rgt_op(rgt_op_12_12[7:0]),
     .bot_op(slf_op_12_11[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_6817), .purst(purst), .slf_op(slf_op_12_12[7:0]),
     .pgate(pgate[207:192]), .bnr_op(rgt_op_12_11[7:0]),
     .bnl_op(slf_op_11_11[7:0]), .tnr_op(rgt_op_12_13[7:0]),
     .tnl_op(net_7455[0:7]));
ltile4rev I_10_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_6761), .lft_op(slf_op_09_11[7:0]),
     .sp12_h_l(net_4835[0:23]), .sp4_h_l(net_4836[0:47]),
     .sp4_v_b(sp4_v_b_10_11[47:0]), .sp12_v_b(sp12_v_b_10_11[23:0]),
     .sp12_h_r(net_6767[0:23]), .sp4_h_r(net_6768[0:47]),
     .sp12_v_t(net_6769[0:23]), .sp4_v_t(net_4811[0:47]),
     .sp4_r_v_b(sp4_v_b_11_11[47:0]), .wl(wl[191:176]),
     .top_op(net_7343[0:7]), .rgt_op(slf_op_11_11[7:0]),
     .bot_op(bot_op_10_11[7:0]), .bl(bl[545:492]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(carry_in_10_11), .purst(purst),
     .slf_op(slf_op_10_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_10_11[7:0]), .bnl_op(bnl_op_10_11[7:0]),
     .tnr_op(net_7427[0:7]), .tnl_op(net_7259[0:7]));
ltile4rev I_10_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_6789), .lft_op(net_7259[0:7]),
     .sp12_h_l(net_4807[0:23]), .sp4_h_l(net_4808[0:47]),
     .sp4_v_b(net_4811[0:47]), .sp12_v_b(net_6769[0:23]),
     .sp12_h_r(net_6795[0:23]), .sp4_h_r(net_6796[0:47]),
     .sp12_v_t(net_6797[0:23]), .sp4_v_t(net_7331[0:47]),
     .sp4_r_v_b(net_6799[0:47]), .wl(wl[207:192]),
     .top_op(net_7315[0:7]), .rgt_op(net_7427[0:7]),
     .bot_op(slf_op_10_11[7:0]), .bl(bl[545:492]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_6761), .purst(purst), .slf_op(net_7343[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_11_11[7:0]),
     .bnl_op(slf_op_09_11[7:0]), .tnr_op(net_7455[0:7]),
     .tnl_op(net_7287[0:7]));
ltile4rev I_12_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_6817), .lft_op(slf_op_11_11[7:0]),
     .sp12_h_l(net_6711[0:23]), .sp4_h_l(net_6712[0:47]),
     .sp4_v_b(sp4_v_b_12_11[47:0]), .sp12_v_b(sp12_v_b_12_11[23:0]),
     .sp12_h_r(sp12_h_r_12_11[23:0]), .sp4_h_r(sp4_h_r_12_11[47:0]),
     .sp12_v_t(net_6825[0:23]), .sp4_v_t(net_6855[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_11[47:0]), .wl(wl[191:176]),
     .top_op(slf_op_12_12[7:0]), .rgt_op(rgt_op_12_11[7:0]),
     .bot_op(bot_op_12_11[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(carry_in_12_11), .purst(purst),
     .slf_op(slf_op_12_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_12_11[7:0]), .bnl_op(bnl_op_12_11[7:0]),
     .tnr_op(rgt_op_12_12[7:0]), .tnl_op(net_7427[0:7]));
ltile4rev I_11_12 ( .vdd_cntl(vdd_cntl[207:192]), .prog(prog),
     .carry_out(net_6845), .lft_op(net_7343[0:7]),
     .sp12_h_l(net_6795[0:23]), .sp4_h_l(net_6796[0:47]),
     .sp4_v_b(net_6799[0:47]), .sp12_v_b(net_6713[0:23]),
     .sp12_h_r(net_6851[0:23]), .sp4_h_r(net_6852[0:47]),
     .sp12_v_t(net_6853[0:23]), .sp4_v_t(net_7415[0:47]),
     .sp4_r_v_b(net_6855[0:47]), .wl(wl[207:192]),
     .top_op(net_7455[0:7]), .rgt_op(slf_op_12_12[7:0]),
     .bot_op(slf_op_11_11[7:0]), .bl(bl[599:546]),
     .reset_b(reset_b[207:192]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_6705), .purst(purst), .slf_op(net_7427[0:7]),
     .pgate(pgate[207:192]), .bnr_op(slf_op_12_11[7:0]),
     .bnl_op(slf_op_10_11[7:0]), .tnr_op(slf_op_12_13[7:0]),
     .tnl_op(net_7315[0:7]));
ltile4rev I_02_11 ( .vdd_cntl(vdd_cntl[191:176]), .prog(prog),
     .carry_out(net_6873), .lft_op(slf_op_01_11[7:0]),
     .sp12_h_l(net_4695[0:23]), .sp4_h_l(net_4696[0:47]),
     .sp4_v_b(sp4_v_b_02_11[47:0]), .sp12_v_b(sp12_v_b_02_11[23:0]),
     .sp12_h_r(net_6879[0:23]), .sp4_h_r(net_6880[0:47]),
     .sp12_v_t(net_6881[0:23]), .sp4_v_t(net_4671[0:47]),
     .sp4_r_v_b(sp4_v_b_03_11[47:0]), .wl(wl[191:176]),
     .top_op(net_6923[0:7]), .rgt_op(slf_op_03_11[7:0]),
     .bot_op(bot_op_02_11[7:0]), .bl(bl[125:72]),
     .reset_b(reset_b[191:176]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(carry_in_02_11), .purst(purst),
     .slf_op(slf_op_02_11[7:0]), .pgate(pgate[191:176]),
     .bnr_op(bnr_op_02_11[7:0]), .bnl_op(bnl_op_02_11[7:0]),
     .tnr_op(net_7007[0:7]), .tnl_op(net_4701[0:7]));
ltile4rev I_01_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_6901), .lft_op({io_l_24[3], io_l_24[2], io_l_24[1],
     io_l_24[0], io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0]}),
     .sp12_h_l(net_4260[0:23]), .sp4_h_l(net_4259[0:47]),
     .sp4_v_b(net_4670[0:47]), .sp12_v_b(net_4669[0:23]),
     .sp12_h_r(net_6907[0:23]), .sp4_h_r(net_6908[0:47]),
     .sp12_v_t(net_6909[0:23]), .sp4_v_t(net_6910[0:47]),
     .sp4_r_v_b(net_6911[0:47]), .wl(wl[223:208]),
     .top_op(net_6913[0:7]), .rgt_op(net_6951[0:7]),
     .bot_op(net_4701[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_4661), .purst(purst), .slf_op(net_4673[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_6923[0:7]),
     .bnl_op({io_l_22[3], io_l_22[2], io_l_22[1], io_l_22[0],
     io_l_22[3], io_l_22[2], io_l_22[1], io_l_22[0]}),
     .tnr_op(net_5159[0:7]), .tnl_op({io_l_26[3], io_l_26[2],
     io_l_26[1], io_l_26[0], io_l_26[3], io_l_26[2], io_l_26[1],
     io_l_26[0]}));
ltile4rev I_01_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_6929), .lft_op({io_l_26[3], io_l_26[2], io_l_26[1],
     io_l_26[0], io_l_26[3], io_l_26[2], io_l_26[1], io_l_26[0]}),
     .sp12_h_l(net_4226[0:23]), .sp4_h_l(net_4225[0:47]),
     .sp4_v_b(net_6910[0:47]), .sp12_v_b(net_6909[0:23]),
     .sp12_h_r(net_6935[0:23]), .sp4_h_r(net_6936[0:47]),
     .sp12_v_t(net_6937[0:23]), .sp4_v_t(net_6938[0:47]),
     .sp4_r_v_b(net_6939[0:47]), .wl(wl[239:224]),
     .top_op(net_6941[0:7]), .rgt_op(net_5159[0:7]),
     .bot_op(net_4673[0:7]), .bl(bl[71:18]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_00[7:0]),
     .carry_in(net_6901), .purst(purst), .slf_op(net_6913[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_6951[0:7]),
     .bnl_op({io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0],
     io_l_24[3], io_l_24[2], io_l_24[1], io_l_24[0]}),
     .tnr_op(net_5131[0:7]), .tnl_op({io_l_28[3], io_l_28[2],
     io_l_28[1], io_l_28[0], io_l_28[3], io_l_28[2], io_l_28[1],
     io_l_28[0]}));
ltile4rev I_02_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_6957), .lft_op(net_6913[0:7]),
     .sp12_h_l(net_6935[0:23]), .sp4_h_l(net_6936[0:47]),
     .sp4_v_b(net_6939[0:47]), .sp12_v_b(net_6993[0:23]),
     .sp12_h_r(net_6963[0:23]), .sp4_h_r(net_6964[0:47]),
     .sp12_v_t(net_6965[0:23]), .sp4_v_t(net_5147[0:47]),
     .sp4_r_v_b(net_6967[0:47]), .wl(wl[239:224]),
     .top_op(net_5131[0:7]), .rgt_op(net_5075[0:7]),
     .bot_op(net_6951[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_6985), .purst(purst), .slf_op(net_5159[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_6979[0:7]),
     .bnl_op(net_4673[0:7]), .tnr_op(net_5103[0:7]),
     .tnl_op(net_6941[0:7]));
ltile4rev I_02_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_6985), .lft_op(net_4673[0:7]),
     .sp12_h_l(net_6907[0:23]), .sp4_h_l(net_6908[0:47]),
     .sp4_v_b(net_6911[0:47]), .sp12_v_b(net_4641[0:23]),
     .sp12_h_r(net_6991[0:23]), .sp4_h_r(net_6992[0:47]),
     .sp12_v_t(net_6993[0:23]), .sp4_v_t(net_6939[0:47]),
     .sp4_r_v_b(net_6995[0:47]), .wl(wl[223:208]),
     .top_op(net_5159[0:7]), .rgt_op(net_6979[0:7]),
     .bot_op(net_6923[0:7]), .bl(bl[125:72]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_01[7:0]),
     .carry_in(net_4633), .purst(purst), .slf_op(net_6951[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7007[0:7]),
     .bnl_op(net_4701[0:7]), .tnr_op(net_5075[0:7]),
     .tnl_op(net_6913[0:7]));
ltile4rev I_05_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7013), .lft_op(net_7119[0:7]),
     .sp12_h_l(net_7159[0:23]), .sp4_h_l(net_7160[0:47]),
     .sp4_v_b(net_7163[0:47]), .sp12_v_b(net_4473[0:23]),
     .sp12_h_r(net_7019[0:23]), .sp4_h_r(net_7020[0:47]),
     .sp12_v_t(net_7021[0:23]), .sp4_v_t(net_7135[0:47]),
     .sp4_r_v_b(net_7023[0:47]), .wl(wl[223:208]),
     .top_op(net_5019[0:7]), .rgt_op(net_7738[0:7]),
     .bot_op(net_7175[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_4465), .purst(purst), .slf_op(net_7147[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_4461[0:7]),
     .bnl_op(net_7091[0:7]), .tnr_op(net_7037[0:7]),
     .tnl_op(net_4935[0:7]));
ltile4rev I_05_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7041), .lft_op(net_4935[0:7]),
     .sp12_h_l(net_7131[0:23]), .sp4_h_l(net_7132[0:47]),
     .sp4_v_b(net_7135[0:47]), .sp12_v_b(net_7021[0:23]),
     .sp12_h_r(net_7047[0:23]), .sp4_h_r(net_7048[0:47]),
     .sp12_v_t(net_7049[0:23]), .sp4_v_t(net_5007[0:47]),
     .sp4_r_v_b(net_7051[0:47]), .wl(wl[239:224]),
     .top_op(net_4991[0:7]), .rgt_op(net_7037[0:7]),
     .bot_op(net_7147[0:7]), .bl(bl[287:234]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_04[7:0]),
     .carry_in(net_7013), .purst(purst), .slf_op(net_5019[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7738[0:7]),
     .bnl_op(net_7119[0:7]), .tnr_op(net_7688[0:7]),
     .tnl_op(net_4963[0:7]));
ltile4rev I_03_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7069), .lft_op(net_6951[0:7]),
     .sp12_h_l(net_6991[0:23]), .sp4_h_l(net_6992[0:47]),
     .sp4_v_b(net_6995[0:47]), .sp12_v_b(net_4529[0:23]),
     .sp12_h_r(net_7075[0:23]), .sp4_h_r(net_7076[0:47]),
     .sp12_v_t(net_7077[0:23]), .sp4_v_t(net_6967[0:47]),
     .sp4_r_v_b(net_7079[0:47]), .wl(wl[223:208]),
     .top_op(net_5075[0:7]), .rgt_op(net_7119[0:7]),
     .bot_op(net_7007[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_4521), .purst(purst), .slf_op(net_6979[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7091[0:7]),
     .bnl_op(net_6923[0:7]), .tnr_op(net_4935[0:7]),
     .tnl_op(net_5159[0:7]));
ltile4rev I_03_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7097), .lft_op(net_5159[0:7]),
     .sp12_h_l(net_6963[0:23]), .sp4_h_l(net_6964[0:47]),
     .sp4_v_b(net_6967[0:47]), .sp12_v_b(net_7077[0:23]),
     .sp12_h_r(net_7103[0:23]), .sp4_h_r(net_7104[0:47]),
     .sp12_v_t(net_7105[0:23]), .sp4_v_t(net_5063[0:47]),
     .sp4_r_v_b(net_7107[0:47]), .wl(wl[239:224]),
     .top_op(net_5103[0:7]), .rgt_op(net_4935[0:7]),
     .bot_op(net_6979[0:7]), .bl(bl[179:126]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_02[7:0]),
     .carry_in(net_7069), .purst(purst), .slf_op(net_5075[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7119[0:7]),
     .bnl_op(net_6951[0:7]), .tnr_op(net_4963[0:7]),
     .tnl_op(net_5131[0:7]));
ltile4rev I_04_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7125), .lft_op(net_5075[0:7]),
     .sp12_h_l(net_7103[0:23]), .sp4_h_l(net_7104[0:47]),
     .sp4_v_b(net_7107[0:47]), .sp12_v_b(net_7161[0:23]),
     .sp12_h_r(net_7131[0:23]), .sp4_h_r(net_7132[0:47]),
     .sp12_v_t(net_7133[0:23]), .sp4_v_t(net_4923[0:47]),
     .sp4_r_v_b(net_7135[0:47]), .wl(wl[239:224]),
     .top_op(net_4963[0:7]), .rgt_op(net_5019[0:7]),
     .bot_op(net_7119[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_7153), .purst(purst), .slf_op(net_4935[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7147[0:7]),
     .bnl_op(net_6979[0:7]), .tnr_op(net_4991[0:7]),
     .tnl_op(net_5103[0:7]));
ltile4rev I_04_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7153), .lft_op(net_6979[0:7]),
     .sp12_h_l(net_7075[0:23]), .sp4_h_l(net_7076[0:47]),
     .sp4_v_b(net_7079[0:47]), .sp12_v_b(net_4557[0:23]),
     .sp12_h_r(net_7159[0:23]), .sp4_h_r(net_7160[0:47]),
     .sp12_v_t(net_7161[0:23]), .sp4_v_t(net_7107[0:47]),
     .sp4_r_v_b(net_7163[0:47]), .wl(wl[223:208]),
     .top_op(net_4935[0:7]), .rgt_op(net_7147[0:7]),
     .bot_op(net_7091[0:7]), .bl(bl[233:180]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_03[7:0]),
     .carry_in(net_4549), .purst(purst), .slf_op(net_7119[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7175[0:7]),
     .bnl_op(net_7007[0:7]), .tnr_op(net_5019[0:7]),
     .tnl_op(net_5075[0:7]));
ltile4rev I_07_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7181), .lft_op(net_7037[0:7]),
     .sp12_h_l(net_7676[0:23]), .sp4_h_l(net_7679[0:47]),
     .sp4_v_b(net_7681[0:47]), .sp12_v_b(net_7217[0:23]),
     .sp12_h_r(net_7187[0:23]), .sp4_h_r(net_7188[0:47]),
     .sp12_v_t(net_7189[0:23]), .sp4_v_t(net_7645[0:47]),
     .sp4_r_v_b(net_7191[0:47]), .wl(wl[239:224]),
     .top_op(net_7193[0:7]), .rgt_op(net_7249[0:7]),
     .bot_op(net_4617[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_7209), .purst(purst), .slf_op(net_7221[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_4785[0:7]),
     .bnl_op(net_7738[0:7]), .tnr_op(net_7277[0:7]),
     .tnl_op(net_7688[0:7]));
ltile4rev I_07_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7209), .lft_op(net_7738[0:7]),
     .sp12_h_l(net_7677[0:23]), .sp4_h_l(net_7678[0:47]),
     .sp4_v_b(net_7682[0:47]), .sp12_v_b(net_4613[0:23]),
     .sp12_h_r(net_7215[0:23]), .sp4_h_r(net_7216[0:47]),
     .sp12_v_t(net_7217[0:23]), .sp4_v_t(net_7681[0:47]),
     .sp4_r_v_b(net_7219[0:47]), .wl(wl[223:208]),
     .top_op(net_7221[0:7]), .rgt_op(net_4785[0:7]),
     .bot_op(net_4729[0:7]), .bl(bl[383:330]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_06[7:0]),
     .carry_in(net_4605), .purst(purst), .slf_op(net_4617[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_4757[0:7]),
     .bnl_op(net_4461[0:7]), .tnr_op(net_7249[0:7]),
     .tnl_op(net_7037[0:7]));
ltile4rev I_08_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7237), .lft_op(net_4617[0:7]),
     .sp12_h_l(net_7215[0:23]), .sp4_h_l(net_7216[0:47]),
     .sp4_v_b(net_7219[0:47]), .sp12_v_b(net_4781[0:23]),
     .sp12_h_r(net_7243[0:23]), .sp4_h_r(net_7244[0:47]),
     .sp12_v_t(net_7245[0:23]), .sp4_v_t(net_7191[0:47]),
     .sp4_r_v_b(net_7247[0:47]), .wl(wl[223:208]),
     .top_op(net_7249[0:7]), .rgt_op(net_7287[0:7]),
     .bot_op(net_4757[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_4773), .purst(purst), .slf_op(net_4785[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7259[0:7]),
     .bnl_op(net_4729[0:7]), .tnr_op(net_5215[0:7]),
     .tnl_op(net_7221[0:7]));
ltile4rev I_08_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7265), .lft_op(net_7221[0:7]),
     .sp12_h_l(net_7187[0:23]), .sp4_h_l(net_7188[0:47]),
     .sp4_v_b(net_7191[0:47]), .sp12_v_b(net_7245[0:23]),
     .sp12_h_r(net_7271[0:23]), .sp4_h_r(net_7272[0:47]),
     .sp12_v_t(net_7273[0:23]), .sp4_v_t(net_5175[0:47]),
     .sp4_r_v_b(net_7275[0:47]), .wl(wl[239:224]),
     .top_op(net_7277[0:7]), .rgt_op(net_5215[0:7]),
     .bot_op(net_4785[0:7]), .bl(bl[437:384]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_07[7:0]),
     .carry_in(net_7237), .purst(purst), .slf_op(net_7249[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7287[0:7]),
     .bnl_op(net_4617[0:7]), .tnr_op(net_5243[0:7]),
     .tnl_op(net_7193[0:7]));
ltile4rev I_09_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7293), .lft_op(net_7249[0:7]),
     .sp12_h_l(net_7271[0:23]), .sp4_h_l(net_7272[0:47]),
     .sp4_v_b(net_7275[0:47]), .sp12_v_b(net_7329[0:23]),
     .sp12_h_r(net_7299[0:23]), .sp4_h_r(net_7300[0:47]),
     .sp12_v_t(net_7301[0:23]), .sp4_v_t(net_5203[0:47]),
     .sp4_r_v_b(net_7303[0:47]), .wl(wl[239:224]),
     .top_op(net_5243[0:7]), .rgt_op(net_5299[0:7]),
     .bot_op(net_7287[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_7321), .purst(purst), .slf_op(net_5215[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7315[0:7]),
     .bnl_op(net_4785[0:7]), .tnr_op(net_5271[0:7]),
     .tnl_op(net_7277[0:7]));
ltile4rev I_09_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7321), .lft_op(net_4785[0:7]),
     .sp12_h_l(net_7243[0:23]), .sp4_h_l(net_7244[0:47]),
     .sp4_v_b(net_7247[0:47]), .sp12_v_b(net_4809[0:23]),
     .sp12_h_r(net_7327[0:23]), .sp4_h_r(net_7328[0:47]),
     .sp12_v_t(net_7329[0:23]), .sp4_v_t(net_7275[0:47]),
     .sp4_r_v_b(net_7331[0:47]), .wl(wl[223:208]),
     .top_op(net_5215[0:7]), .rgt_op(net_7315[0:7]),
     .bot_op(net_7259[0:7]), .bl(bl[491:438]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_08[7:0]),
     .carry_in(net_4801), .purst(purst), .slf_op(net_7287[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7343[0:7]),
     .bnl_op(net_4757[0:7]), .tnr_op(net_5299[0:7]),
     .tnl_op(net_7249[0:7]));
ltile4rev I_11_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7349), .lft_op(net_7315[0:7]),
     .sp12_h_l(net_7411[0:23]), .sp4_h_l(net_7412[0:47]),
     .sp4_v_b(net_7415[0:47]), .sp12_v_b(net_6853[0:23]),
     .sp12_h_r(net_7355[0:23]), .sp4_h_r(net_7356[0:47]),
     .sp12_v_t(net_7357[0:23]), .sp4_v_t(net_7443[0:47]),
     .sp4_r_v_b(net_7359[0:47]), .wl(wl[223:208]),
     .top_op(net_5383[0:7]), .rgt_op(slf_op_12_13[7:0]),
     .bot_op(net_7427[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_6845), .purst(purst), .slf_op(net_7455[0:7]),
     .pgate(pgate[223:208]), .bnr_op(slf_op_12_12[7:0]),
     .bnl_op(net_7343[0:7]), .tnr_op(slf_op_12_14[7:0]),
     .tnl_op(net_5299[0:7]));
ltile4rev I_12_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7377), .lft_op(net_5383[0:7]),
     .sp12_h_l(net_7495[0:23]), .sp4_h_l(net_7496[0:47]),
     .sp4_v_b(net_7499[0:47]), .sp12_v_b(net_7469[0:23]),
     .sp12_h_r(sp12_h_r_12_14[23:0]), .sp4_h_r(sp4_h_r_12_14[47:0]),
     .sp12_v_t(net_7385[0:23]), .sp4_v_t(net_5315[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_14[47:0]), .wl(wl[239:224]),
     .top_op(slf_op_12_15[7:0]), .rgt_op(rgt_op_12_14[7:0]),
     .bot_op(slf_op_12_13[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_7461), .purst(purst), .slf_op(slf_op_12_14[7:0]),
     .pgate(pgate[239:224]), .bnr_op(rgt_op_12_13[7:0]),
     .bnl_op(net_7455[0:7]), .tnr_op(rgt_op_12_15[7:0]),
     .tnl_op(net_5411[0:7]));
ltile4rev I_10_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7405), .lft_op(net_7287[0:7]),
     .sp12_h_l(net_7327[0:23]), .sp4_h_l(net_7328[0:47]),
     .sp4_v_b(net_7331[0:47]), .sp12_v_b(net_6797[0:23]),
     .sp12_h_r(net_7411[0:23]), .sp4_h_r(net_7412[0:47]),
     .sp12_v_t(net_7413[0:23]), .sp4_v_t(net_7303[0:47]),
     .sp4_r_v_b(net_7415[0:47]), .wl(wl[223:208]),
     .top_op(net_5299[0:7]), .rgt_op(net_7455[0:7]),
     .bot_op(net_7343[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_6789), .purst(purst), .slf_op(net_7315[0:7]),
     .pgate(pgate[223:208]), .bnr_op(net_7427[0:7]),
     .bnl_op(net_7259[0:7]), .tnr_op(net_5383[0:7]),
     .tnl_op(net_5215[0:7]));
ltile4rev I_10_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7433), .lft_op(net_5215[0:7]),
     .sp12_h_l(net_7299[0:23]), .sp4_h_l(net_7300[0:47]),
     .sp4_v_b(net_7303[0:47]), .sp12_v_b(net_7413[0:23]),
     .sp12_h_r(net_7439[0:23]), .sp4_h_r(net_7440[0:47]),
     .sp12_v_t(net_7441[0:23]), .sp4_v_t(net_5287[0:47]),
     .sp4_r_v_b(net_7443[0:47]), .wl(wl[239:224]),
     .top_op(net_5271[0:7]), .rgt_op(net_5383[0:7]),
     .bot_op(net_7315[0:7]), .bl(bl[545:492]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_09[7:0]),
     .carry_in(net_7405), .purst(purst), .slf_op(net_5299[0:7]),
     .pgate(pgate[239:224]), .bnr_op(net_7455[0:7]),
     .bnl_op(net_7287[0:7]), .tnr_op(net_5411[0:7]),
     .tnl_op(net_5243[0:7]));
ltile4rev I_12_13 ( .vdd_cntl(vdd_cntl[223:208]), .prog(prog),
     .carry_out(net_7461), .lft_op(net_7455[0:7]),
     .sp12_h_l(net_7355[0:23]), .sp4_h_l(net_7356[0:47]),
     .sp4_v_b(net_7359[0:47]), .sp12_v_b(net_6741[0:23]),
     .sp12_h_r(sp12_h_r_12_13[23:0]), .sp4_h_r(sp4_h_r_12_13[47:0]),
     .sp12_v_t(net_7469[0:23]), .sp4_v_t(net_7499[0:47]),
     .sp4_r_v_b(sp4_r_v_b_12_13[47:0]), .wl(wl[223:208]),
     .top_op(slf_op_12_14[7:0]), .rgt_op(rgt_op_12_13[7:0]),
     .bot_op(slf_op_12_12[7:0]), .bl(bl[653:600]),
     .reset_b(reset_b[223:208]), .glb_netwk(glb_netwk_11[7:0]),
     .carry_in(net_7479), .purst(purst), .slf_op(slf_op_12_13[7:0]),
     .pgate(pgate[223:208]), .bnr_op(rgt_op_12_12[7:0]),
     .bnl_op(net_7427[0:7]), .tnr_op(rgt_op_12_14[7:0]),
     .tnl_op(net_5383[0:7]));
ltile4rev I_11_14 ( .vdd_cntl(vdd_cntl[239:224]), .prog(prog),
     .carry_out(net_7489), .lft_op(net_5299[0:7]),
     .sp12_h_l(net_7439[0:23]), .sp4_h_l(net_7440[0:47]),
     .sp4_v_b(net_7443[0:47]), .sp12_v_b(net_7357[0:23]),
     .sp12_h_r(net_7495[0:23]), .sp4_h_r(net_7496[0:47]),
     .sp12_v_t(net_7497[0:23]), .sp4_v_t(net_5371[0:47]),
     .sp4_r_v_b(net_7499[0:47]), .wl(wl[239:224]),
     .top_op(net_5411[0:7]), .rgt_op(slf_op_12_14[7:0]),
     .bot_op(net_7455[0:7]), .bl(bl[599:546]),
     .reset_b(reset_b[239:224]), .glb_netwk(glb_netwk_10[7:0]),
     .carry_in(net_7349), .purst(purst), .slf_op(net_5383[0:7]),
     .pgate(pgate[239:224]), .bnr_op(slf_op_12_13[7:0]),
     .bnl_op(net_7315[0:7]), .tnr_op(slf_op_12_15[7:0]),
     .tnl_op(net_5271[0:7]));
inv_hvt I1014 ( .A(net_7522), .Y(fabric_out_226));
inv_hvt I1016 ( .A(net_7520), .Y(fabric_out_228));
inv_hvt I1017 ( .A(net_8052), .Y(net_7520));
inv_hvt I1013 ( .A(net_8086), .Y(net_7522));
inv_hvt I1010 ( .A(padin_t[23]), .Y(net_7524));
inv_hvt I1007 ( .A(net_7525), .Y(fabric_out_30));
inv_hvt I1011 ( .A(net_7524), .Y(padin_226));
inv_hvt I1012 ( .A(net_7529), .Y(padin_30));
inv_hvt I1006 ( .A(net_7531), .Y(net_7525));
inv_hvt I1015 ( .A(padin_l[20]), .Y(net_7529));
clk_quad_bufx8 I_quad_driver ( .clko(net2col_drivers[7:0]),
     .clki(glb_in[7:0]));
bram_4kprouting_tbank I_bram0617 ( .glb_netwk(glb_netwk_05[7:0]),
     .vdd_cntl_bot(vdd_cntl[287:272]),
     .vdd_cntl_top(vdd_cntl[303:288]), .bm_sdo_o(net_7605),
     .bm_sdi_i(net_7607), .bm_sclkrw_i(net_7608), .bm_sdo_i(net_7543),
     .bm_sweb_i(net_7609), .bm_sdi_o(net_7545), .bm_sclkrw_o(net_7546),
     .bm_sweb_o(net_7547), .slf_op_top(net_6225[0:7]),
     .slf_op_bot(net_7614[0:7]), .wl_top(wl[303:288]),
     .wl_bot(wl[287:272]), .top_op_top(net_7552[0:7]),
     .tnl_op_top(net_5607[0:7]), .tnl_op_bot(net_5635[0:7]),
     .reset_b_top(reset_b[303:288]), .reset_b_bot(reset_b[287:272]),
     .prog(prog), .pgate_top(pgate[303:288]),
     .pgate_bot(pgate[287:272]), .lft_op_top(net_5635[0:7]),
     .lft_op_bot(net_6335[0:7]), .bm_wdummymux_en_i(net_7660),
     .bot_op_bot(net_6223[0:7]), .bnl_op_top(net_6335[0:7]),
     .bnl_op_bot(net_6363[0:7]), .sp12_v_t_top(net_7566[0:23]),
     .sp12_v_b_bot(net_7634[0:23]), .bm_init_i(net_7656),
     .sp12_h_l_top(net_6235[0:23]), .sp12_h_l_bot(net_6207[0:23]),
     .sp4_v_t_top(net_5483[0:47]), .sp4_v_b_top(net_6239[0:47]),
     .sp4_v_b_bot(net_6211[0:47]), .sp4_h_l_top(net_6236[0:47]),
     .sp4_h_l_bot(net_6208[0:47]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(net_7655), .bm_sa_i(net_7657[0:7]),
     .bm_sclk_i(net_7658), .bm_sreb_i(net_7659),
     .bm_rcapmux_en_o(net_7581), .bm_init_o(net_7582),
     .bm_sa_o(net_7583[0:7]), .bm_sclk_o(net_7584),
     .bm_sreb_o(net_7585), .bm_wdummymux_en_o(net_7586),
     .bnr_op_top(net_5037[0:7]), .rgt_op_top(net_6409[0:7]),
     .tnr_op_top(net_6381[0:7]), .tnr_op_bot(net_6409[0:7]),
     .sp12_h_r_top(net_7591[0:23]), .sp12_h_r_bot(net_7592[0:23]),
     .sp4_h_r_bot(net_7593[0:47]), .sp4_h_r_top(net_7594[0:47]),
     .rgt_op_bot(net_5037[0:7]), .sp4_r_v_b_top(net_7596[0:47]),
     .sp4_r_v_b_bot(net_7597[0:47]), .bnr_op_bot(net_5177[0:7]));
bram_4kprouting_tbank I_bram0615 ( .glb_netwk(glb_netwk_05[7:0]),
     .vdd_cntl_bot(vdd_cntl[255:240]),
     .vdd_cntl_top(vdd_cntl[271:256]), .bm_sdo_o(net_7667),
     .bm_sdi_i(net_7669), .bm_sclkrw_i(net_7670), .bm_sdo_i(net_7605),
     .bm_sweb_i(net_7671), .bm_sdi_o(net_7607), .bm_sclkrw_o(net_7608),
     .bm_sweb_o(net_7609), .slf_op_top(net_6223[0:7]),
     .slf_op_bot(net_7688[0:7]), .wl_top(wl[271:256]),
     .wl_bot(wl[255:240]), .top_op_top(net_7614[0:7]),
     .tnr_op_top(net_5037[0:7]), .tnr_op_bot(net_5177[0:7]),
     .tnl_op_top(net_6335[0:7]), .tnl_op_bot(net_6363[0:7]),
     .rgt_op_top(net_5177[0:7]), .rgt_op_bot(net_7193[0:7]),
     .reset_b_top(reset_b[271:256]), .reset_b_bot(reset_b[255:240]),
     .prog(prog), .pgate_top(pgate[271:256]),
     .pgate_bot(pgate[255:240]), .lft_op_top(net_6363[0:7]),
     .lft_op_bot(net_4991[0:7]), .bm_wdummymux_en_i(net_7722),
     .bot_op_bot(net_7037[0:7]), .bnr_op_top(net_7193[0:7]),
     .bnr_op_bot(net_7221[0:7]), .bnl_op_top(net_4991[0:7]),
     .bnl_op_bot(net_5019[0:7]), .sp12_v_t_top(net_7634[0:23]),
     .sp12_v_b_bot(net_7702[0:23]), .bm_init_i(net_7718),
     .sp12_h_r_top(net_7637[0:23]), .sp12_h_r_bot(net_7638[0:23]),
     .sp12_h_l_top(net_4891[0:23]), .sp12_h_l_bot(net_4863[0:23]),
     .sp4_v_t_top(net_6211[0:47]), .sp4_v_b_top(net_4895[0:47]),
     .sp4_v_b_bot(net_4867[0:47]), .sp4_r_v_b_top(net_7644[0:47]),
     .sp4_r_v_b_bot(net_7645[0:47]), .sp4_h_r_top(net_7646[0:47]),
     .sp4_h_r_bot(net_7647[0:47]), .sp4_h_l_top(net_4892[0:47]),
     .sp4_h_l_bot(net_4864[0:47]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(net_7717), .bm_sa_i(net_7719[0:7]),
     .bm_sclk_i(net_7720), .bm_sreb_i(net_7721),
     .bm_rcapmux_en_o(net_7655), .bm_init_o(net_7656),
     .bm_sa_o(net_7657[0:7]), .bm_sclk_o(net_7658),
     .bm_sreb_o(net_7659), .bm_wdummymux_en_o(net_7660));
bram_4kprouting_tbank I_bram0613 ( .glb_netwk(glb_netwk_05[7:0]),
     .vdd_cntl_bot(vdd_cntl[223:208]),
     .vdd_cntl_top(vdd_cntl[239:224]), .bm_sdo_o(net_7729),
     .bm_sdi_i(net_7731), .bm_sclkrw_i(net_7732), .bm_sdo_i(net_7667),
     .bm_sweb_i(net_7733), .bm_sdi_o(net_7669), .bm_sclkrw_o(net_7670),
     .bm_sweb_o(net_7671), .bnr_op_top(net_4617[0:7]),
     .rgt_op_top(net_7221[0:7]), .tnr_op_top(net_7193[0:7]),
     .tnr_op_bot(net_7221[0:7]), .sp12_h_r_top(net_7676[0:23]),
     .sp12_h_r_bot(net_7677[0:23]), .sp4_h_r_bot(net_7678[0:47]),
     .sp4_h_r_top(net_7679[0:47]), .rgt_op_bot(net_4617[0:7]),
     .sp4_r_v_b_top(net_7681[0:47]), .sp4_r_v_b_bot(net_7682[0:47]),
     .bnr_op_bot(net_4729[0:7]), .slf_op_top(net_7037[0:7]),
     .slf_op_bot(net_7738[0:7]), .wl_top(wl[239:224]),
     .wl_bot(wl[223:208]), .top_op_top(net_7688[0:7]),
     .tnl_op_top(net_4991[0:7]), .tnl_op_bot(net_5019[0:7]),
     .reset_b_top(reset_b[239:224]), .reset_b_bot(reset_b[223:208]),
     .prog(prog), .pgate_top(pgate[239:224]),
     .pgate_bot(pgate[223:208]), .lft_op_top(net_5019[0:7]),
     .lft_op_bot(net_7147[0:7]), .bm_wdummymux_en_i(net_7784),
     .bot_op_bot(net_4461[0:7]), .bnl_op_top(net_7147[0:7]),
     .bnl_op_bot(net_7175[0:7]), .sp12_v_t_top(net_7702[0:23]),
     .sp12_v_b_bot(net_7758[0:23]), .bm_init_i(net_7780),
     .sp12_h_l_top(net_7047[0:23]), .sp12_h_l_bot(net_7019[0:23]),
     .sp4_v_t_top(net_4867[0:47]), .sp4_v_b_top(net_7051[0:47]),
     .sp4_v_b_bot(net_7023[0:47]), .sp4_h_l_top(net_7048[0:47]),
     .sp4_h_l_bot(net_7020[0:47]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(net_7779), .bm_sa_i(net_7781[0:7]),
     .bm_sclk_i(net_7782), .bm_sreb_i(net_7783),
     .bm_rcapmux_en_o(net_7717), .bm_init_o(net_7718),
     .bm_sa_o(net_7719[0:7]), .bm_sclk_o(net_7720),
     .bm_sreb_o(net_7721), .bm_wdummymux_en_o(net_7722));
bram_4kprouting_tbankout I_bram0611 ( .glb_netwk(glb_netwk_05[7:0]),
     .vdd_cntl_bot(vdd_cntl[191:176]),
     .vdd_cntl_top(vdd_cntl[207:192]), .bm_sdo_o(bm_sdo_o),
     .bm_sdi_i(bm_sdi_i), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sdo_i(net_7729), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(net_7731),
     .bm_sclkrw_o(net_7732), .bm_sweb_o(net_7733),
     .slf_op_top(net_4461[0:7]), .slf_op_bot(slf_op_06_11[7:0]),
     .wl_top(wl[207:192]), .wl_bot(wl[191:176]),
     .top_op_top(net_7738[0:7]), .tnr_op_top(net_4617[0:7]),
     .tnr_op_bot(net_4729[0:7]), .tnl_op_top(net_7147[0:7]),
     .tnl_op_bot(net_7175[0:7]), .rgt_op_top(net_4729[0:7]),
     .rgt_op_bot(slf_op_07_11[7:0]), .reset_b_top(reset_b[207:192]),
     .reset_b_bot(reset_b[191:176]), .prog(prog),
     .pgate_top(pgate[207:192]), .pgate_bot(pgate[191:176]),
     .lft_op_top(net_7175[0:7]), .lft_op_bot(slf_op_05_11[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_06_11[7:0]), .bnr_op_top(slf_op_07_11[7:0]),
     .bnr_op_bot(bnr_op_06_11[7:0]), .bnl_op_top(slf_op_05_11[7:0]),
     .bnl_op_bot(bnl_op_06_11[7:0]), .sp12_v_t_top(net_7758[0:23]),
     .sp12_v_b_bot(sp12_v_b_06_11[23:0]), .bm_init_i(bm_init_i),
     .sp12_h_r_top(net_7761[0:23]), .sp12_h_r_bot(net_7762[0:23]),
     .sp12_h_l_top(net_4471[0:23]), .sp12_h_l_bot(net_4443[0:23]),
     .sp4_v_t_top(net_7023[0:47]), .sp4_v_b_top(net_4475[0:47]),
     .sp4_v_b_bot(sp4_v_b_06_11[47:0]), .sp4_r_v_b_top(net_7768[0:47]),
     .sp4_r_v_b_bot(sp4_v_b_07_11[47:0]), .sp4_h_r_top(net_7770[0:47]),
     .sp4_h_r_bot(net_7771[0:47]), .sp4_h_l_top(net_4472[0:47]),
     .sp4_h_l_bot(net_4444[0:47]), .bl(bl[329:288]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(net_7779), .bm_init_o(net_7780),
     .bm_sa_o(net_7781[0:7]), .bm_sclk_o(net_7782),
     .bm_sreb_o(net_7783), .bm_wdummymux_en_o(net_7784));
clk_colbufx8 I790 ( .clko(glb_netwk_07[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I798 ( .clko(glb_netwk_11[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I787 ( .clko(glb_netwk_03[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I791 ( .clko(glb_netwk_05[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I788 ( .clko(glb_netwk_02[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I800 ( .clko(glb_netwk_08[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I786 ( .clko(glb_netwk_01[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I789 ( .clko(glb_netwk_06[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I799 ( .clko(glb_netwk_09[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I797 ( .clko(glb_netwk_10[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I793 ( .clko(glb_netwk_io_l[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I792 ( .clko(glb_netwk_04[7:0]),
     .clki(net2col_drivers[7:0]));
clk_colbufx8 I785 ( .clko(glb_netwk_00[7:0]),
     .clki(net2col_drivers[7:0]));
io_col4 I_03_21_iot05 ( .ceb(net_04420), .cf(cf_t[71:48]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_7814), .sdo(net_7850), .sdi(net_7816),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[2]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[5:4]), .pado(pado_t[5:4]),
     .padeb(padeb_t[5:4]), .sp4_v_t(net_7874[0:15]),
     .sp4_h_l(net_7831[0:47]), .sp12_h_l(net_5565[0:23]), .prog(prog),
     .spi_ss_in_b(net_7834[0:1]), .tnl_op(net_8143[0:7]),
     .lft_op(net_7871[0:7]), .bnl_op(net_7837[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7840[0:15]), .wl(wl[351:336]), .bl({bl[127], bl[126],
     bl[165], bl[163], bl[154], bl[160], bl[159], bl[158], bl[157],
     bl[156], bl[137], bl[136], bl[135], bl[134], bl[133], bl[132],
     bl[167], bl[166]}), .slf_op(io_t_4[3:0]),
     .glb_netwk(glb_netwk_02[7:0]));
io_col4 I_02_21_iot03 ( .ceb(net_04420), .cf(cf_t[47:24]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_7848), .sdo(net_8122), .sdi(net_7850),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[1]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[3:2]), .pado(pado_t[3:2]),
     .padeb(padeb_t[3:2]), .sp4_v_t(net_8146[0:15]),
     .sp4_h_l(net_7865[0:47]), .sp12_h_l(net_5705[0:23]), .prog(prog),
     .spi_ss_in_b(net_7868[0:1]), .tnl_op(net_5765[0:7]),
     .lft_op(net_8143[0:7]), .bnl_op(net_7871[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7874[0:15]), .wl(wl[351:336]), .bl({bl[73], bl[72],
     bl[111], bl[109], bl[100], bl[106], bl[105], bl[104], bl[103],
     bl[102], bl[83], bl[82], bl[81], bl[80], bl[79], bl[78], bl[113],
     bl[112]}), .slf_op(io_t_2[3:0]), .glb_netwk(glb_netwk_01[7:0]));
io_col4 I_04_21_iot07 ( .ceb(net_04420), .cf(cf_t[95:72]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_7882), .sdo(net_7816), .sdi(net_7884),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[3]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[7:6]), .pado(pado_t[7:6]),
     .padeb(padeb_t[7:6]), .sp4_v_t(net_7840[0:15]),
     .sp4_h_l(net_7899[0:47]), .sp12_h_l(net_5593[0:23]), .prog(prog),
     .spi_ss_in_b(net_7902[0:1]), .tnl_op(net_7871[0:7]),
     .lft_op(net_7837[0:7]), .bnl_op(net_7905[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7908[0:15]), .wl(wl[351:336]), .bl({bl[181], bl[180],
     bl[219], bl[217], bl[208], bl[214], bl[213], bl[212], bl[211],
     bl[210], bl[191], bl[190], bl[189], bl[188], bl[187], bl[186],
     bl[221], bl[220]}), .slf_op(io_t_6[3:0]),
     .glb_netwk(glb_netwk_03[7:0]));
io_col4 I_07_21_iot13 ( .ceb(net_04420), .cf(cf_t[167:144]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_7916), .sdo(net_8190), .sdi(net_7918),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[6]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[13:12]), .pado(pado_t[13:12]),
     .padeb(padeb_t[13:12]), .sp4_v_t(net_8214[0:15]),
     .sp4_h_l(net_7933[0:47]), .sp12_h_l(net_5649[0:23]), .prog(prog),
     .spi_ss_in_b(net_7936[0:1]), .tnl_op(net_8177[0:7]),
     .lft_op(net_8211[0:7]), .bnl_op(net_7939[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7942[0:15]), .wl(wl[351:336]), .bl({bl[331], bl[330],
     bl[369], bl[367], bl[358], bl[364], bl[363], bl[362], bl[361],
     bl[360], bl[341], bl[340], bl[339], bl[338], bl[337], bl[336],
     bl[371], bl[370]}), .slf_op(io_t_12[3:0]),
     .glb_netwk(glb_netwk_06[7:0]));
io_col4 I_08_21_iot15 ( .ceb(net_04420), .cf(cf_t[191:168]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_7950), .sdo(net_7918), .sdi(net_7952),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[7]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[15:14]), .pado(pado_t[15:14]),
     .padeb(padeb_t[15:14]), .sp4_v_t(net_7942[0:15]),
     .sp4_h_l(net_7967[0:47]), .sp12_h_l(net_5845[0:23]), .prog(prog),
     .spi_ss_in_b(net_7970[0:1]), .tnl_op(net_8211[0:7]),
     .lft_op(net_7939[0:7]), .bnl_op(net_7973[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_7976[0:15]), .wl(wl[351:336]), .bl({bl[385], bl[384],
     bl[423], bl[421], bl[412], bl[418], bl[417], bl[416], bl[415],
     bl[414], bl[395], bl[394], bl[393], bl[392], bl[391], bl[390],
     bl[425], bl[424]}), .slf_op(io_t_14[3:0]),
     .glb_netwk(glb_netwk_07[7:0]));
io_col4 I_09_21_iot17 ( .ceb(net_04420), .cf(cf_t[215:192]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_7984), .sdo(net_7952), .sdi(net_7986),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[8]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[17:16]), .pado(pado_t[17:16]),
     .padeb(padeb_t[17:16]), .sp4_v_t(net_7976[0:15]),
     .sp4_h_l(net_8001[0:47]), .sp12_h_l(net_5873[0:23]), .prog(prog),
     .spi_ss_in_b(net_8004[0:1]), .tnl_op(net_7939[0:7]),
     .lft_op(net_7973[0:7]), .bnl_op(net_8007[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8010[0:15]), .wl(wl[351:336]), .bl({bl[439], bl[438],
     bl[477], bl[475], bl[466], bl[472], bl[471], bl[470], bl[469],
     bl[468], bl[449], bl[448], bl[447], bl[446], bl[445], bl[444],
     bl[479], bl[478]}), .slf_op(io_t_16[3:0]),
     .glb_netwk(glb_netwk_08[7:0]));
io_col4 I_10_21_iot19 ( .ceb(net_04420), .cf(cf_t[239:216]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_8018), .sdo(net_7986), .sdi(net_8020),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[9]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[19:18]), .pado(pado_t[19:18]),
     .padeb(padeb_t[19:18]), .sp4_v_t(net_8010[0:15]),
     .sp4_h_l(net_8035[0:47]), .sp12_h_l(net_6013[0:23]), .prog(prog),
     .spi_ss_in_b(net_8038[0:1]), .tnl_op(net_7973[0:7]),
     .lft_op(net_8007[0:7]), .bnl_op(net_8041[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8044[0:15]), .wl(wl[351:336]), .bl({bl[493], bl[492],
     bl[531], bl[529], bl[520], bl[526], bl[525], bl[524], bl[523],
     bl[522], bl[503], bl[502], bl[501], bl[500], bl[499], bl[498],
     bl[533], bl[532]}), .slf_op(io_t_18[3:0]),
     .glb_netwk(glb_netwk_09[7:0]));
io_col4 I_11_21_iot21 ( .ceb(net_04420), .cf(cf_t[263:240]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_8052), .sdo(net_8020), .sdi(net_8054),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[10]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[21:20]), .pado(pado_t[21:20]),
     .padeb(padeb_t[21:20]), .sp4_v_t(net_8044[0:15]),
     .sp4_h_l(net_8069[0:47]), .sp12_h_l(net_6069[0:23]), .prog(prog),
     .spi_ss_in_b(net_8072[0:1]), .tnl_op(net_8007[0:7]),
     .lft_op(net_8041[0:7]), .bnl_op(slf_op_12_20[7:0]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8078[0:15]), .wl(wl[351:336]), .bl({bl[547], bl[546],
     bl[585], bl[583], bl[574], bl[580], bl[579], bl[578], bl[577],
     bl[576], bl[557], bl[556], bl[555], bl[554], bl[553], bl[552],
     bl[587], bl[586]}), .slf_op(io_t_20[3:0]),
     .glb_netwk(glb_netwk_10[7:0]));
io_col4 I_12_21_iot23 ( .ceb(net_04420), .cf(cf_t[287:264]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_8086), .sdo(net_8054), .sdi(net_8088),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[11]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[23:22]), .pado(pado_t[23:22]),
     .padeb(padeb_t[23:22]), .sp4_v_t(net_8078[0:15]),
     .sp4_h_l(net_8103[0:47]), .sp12_h_l(net_5957[0:23]), .prog(prog),
     .spi_ss_in_b(net_8106[0:1]), .tnl_op(net_8041[0:7]),
     .lft_op(slf_op_12_20[7:0]), .bnl_op(rgt_op_12_20[7:0]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(sp4_h_r_12_21[15:0]), .wl(wl[351:336]), .bl({bl[601],
     bl[600], bl[639], bl[637], bl[628], bl[634], bl[633], bl[632],
     bl[631], bl[630], bl[611], bl[610], bl[609], bl[608], bl[607],
     bl[606], bl[641], bl[640]}), .slf_op(slf_op_12_21[3:0]),
     .glb_netwk(glb_netwk_11[7:0]));
io_col4 I_01_21_iot01 ( .ceb(net_04420), .cf(cf_t[23:0]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_8120), .sdo(net_4405), .sdi(net_8122),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[0]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[1:0]), .pado(pado_t[1:0]),
     .padeb(padeb_t[1:0]), .sp4_v_t(net_4020[0:15]),
     .sp4_h_l(net_8137[0:47]), .sp12_h_l(net_5733[0:23]), .prog(prog),
     .spi_ss_in_b(net_8140[0:1]), .tnl_op({io_l_38[3], io_l_38[2],
     io_l_38[1], io_l_38[0], io_l_38[3], io_l_38[2], io_l_38[1],
     io_l_38[0]}), .lft_op(net_5765[0:7]), .bnl_op(net_8143[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8146[0:15]), .wl(wl[351:336]), .bl({bl[19], bl[18],
     bl[57], bl[55], bl[46], bl[52], bl[51], bl[50], bl[49], bl[48],
     bl[29], bl[28], bl[27], bl[26], bl[25], bl[24], bl[59], bl[58]}),
     .slf_op(io_t_0[3:0]), .glb_netwk(glb_netwk_00[7:0]));
io_col4 I_05_21_iot09 ( .ceb(net_04420), .cf(cf_t[119:96]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_8154), .sdo(net_7884), .sdi(net_8156),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[4]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[9:8]), .pado(pado_t[9:8]),
     .padeb(padeb_t[9:8]), .sp4_v_t(net_7908[0:15]),
     .sp4_h_l(net_8171[0:47]), .sp12_h_l(net_5509[0:23]), .prog(prog),
     .spi_ss_in_b(net_8174[0:1]), .tnl_op(net_7837[0:7]),
     .lft_op(net_7905[0:7]), .bnl_op(net_8177[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8180[0:15]), .wl(wl[351:336]), .bl({bl[235], bl[234],
     bl[273], bl[271], bl[262], bl[268], bl[267], bl[266], bl[265],
     bl[264], bl[245], bl[244], bl[243], bl[242], bl[241], bl[240],
     bl[275], bl[274]}), .slf_op(io_t_8[3:0]),
     .glb_netwk(glb_netwk_04[7:0]));
io_col4 I_06_21_iot11 ( .ceb(net_04420), .cf(cf_t[143:120]),
     .vdd_cntl(vdd_cntl[351:336]), .hold(hold_t_l),
     .fabric_out(net_8188), .sdo(net_8156), .sdi(net_8190),
     .spiout({tiegnd, tiegnd}), .cdone_in(end_of_startup_top_l[5]),
     .spioeb({tievdd, tievdd}), .mode(net_4415), .shift(net_4429),
     .hiz_b(net_4433), .r(net_4419), .bs_en(net_4427), .tclk(net_4407),
     .update(net_4431), .padin(padin_t[11:10]), .pado(pado_t[11:10]),
     .padeb(padeb_t[11:10]), .sp4_v_t(net_8180[0:15]),
     .sp4_h_l(net_4383[0:47]), .sp12_h_l(net_4376[0:23]), .prog(prog),
     .spi_ss_in_b(net_8208[0:1]), .tnl_op(net_7905[0:7]),
     .lft_op(net_8177[0:7]), .bnl_op(net_8211[0:7]),
     .pgate(pgate[351:336]), .reset(reset_b[351:336]),
     .sp4_v_b(net_8214[0:15]), .wl(wl[351:336]), .bl({bl[289], bl[288],
     bl[315], bl[313], bl[304], bl[310], bl[309], bl[308], bl[307],
     bl[306], bl[299], bl[298], bl[297], bl[296], bl[295], bl[294],
     bl[317], bl[316]}), .slf_op(io_t_10[3:0]),
     .glb_netwk(glb_netwk_05[7:0]));

endmodule
// Library - leafcell, Cell - bram_bufferx16_2inv, View - schematic
// LAST TIME SAVED: Aug  4 12:31:20 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module bram_bufferx16_2inv ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - misc, Cell - smc_and_jtag_ice4frr, View - schematic
// LAST TIME SAVED: Apr  8 13:57:07 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module smc_and_jtag_ice4frr ( bm_bank_sdi, bm_banksel, bm_clk, bm_init,
     bm_rcapmux_en, bm_sa, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_banksel, cm_clk, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2, cm_sdi_u3, data_muxsel, data_muxsel1,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0, j_hiz_b,
     j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck, j_tdi,
     j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, psdo, rst_b,
     smc_load_nvcm_bstream, smc_osc_fsel, smc_oscoff_b, smc_podt_off,
     smc_podt_rst, smc_read, smc_row_inc, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rsr_rst, smc_rwl_en, smc_seq_rst,
     smc_wcram_rst, smc_wdis_dclk, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, tdo_oe_pad, tdo_pad,
     bm_bank_sdo, boot, bp0, bschain_sdo, cdone_in, cm_last_rsr,
     cm_monitor_cell, cm_sdo_u0, cm_sdo_u1, cm_sdo_u2, cm_sdo_u3,
     cnt_podt_out, coldboot_sel, creset_b, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b, osc_clk, por_b,
     psdi, spi_clk_in, spi_sdi, spi_ss_in_b, tck_pad, tdi_pad, tms_pad,
     trst_pad, warmboot_sel );
output  bm_clk, bm_init, bm_rcapmux_en, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_clk, data_muxsel,
     data_muxsel1, en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0,
     j_hiz_b, j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck,
     j_tdi, j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, rst_b,
     smc_load_nvcm_bstream, smc_oscoff_b, smc_podt_off, smc_podt_rst,
     smc_read, smc_row_inc, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rsr_rst, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_wdis_dclk, smc_write, smc_wset_prec, smc_wset_precgnd,
     smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_oe_pad, tdo_pad;

input  boot, bp0, bschain_sdo, cdone_in, cm_last_rsr, cnt_podt_out,
     creset_b, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, osc_clk, por_b, spi_clk_in, spi_sdi,
     spi_ss_in_b, tck_pad, tdi_pad, tms_pad, trst_pad;

output [1:0]  cm_sdi_u3;
output [7:0]  bm_sa;
output [1:0]  cm_sdi_u0;
output [1:0]  cm_sdi_u1;
output [3:0]  bm_banksel;
output [1:0]  smc_osc_fsel;
output [7:1]  psdo;
output [1:0]  cm_sdi_u2;
output [3:0]  bm_bank_sdi;
output [3:0]  cm_banksel;

input [1:0]  cm_sdo_u2;
input [1:0]  coldboot_sel;
input [1:0]  cm_sdo_u0;
input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdo_u3;
input [3:0]  cm_monitor_cell;
input [7:1]  psdi;
input [1:0]  warmboot_sel;
input [3:0]  bm_bank_sdo;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - leafcell, Cell - bram_hbuffer_2xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:01:06 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module bram_hbuffer_2xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;
output [3:0]  bm_sdi_o;
output [3:0]  bm_sdo_o;
output [3:0]  bm_banksel_o;

input [3:0]  bm_sdi_i;
input [3:0]  bm_banksel_i;
input [3:0]  bm_sdo_i;
input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx16_2inv I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_3_ ( .in(bm_sdo_i[3]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I2_2_ ( .in(bm_sdo_i[2]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_3_ ( .in(bm_banksel_i[3]),
     .out(bm_banksel_o[3]));
bram_bufferx16_2inv I13_2_ ( .in(bm_banksel_i[2]),
     .out(bm_banksel_o[2]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_icg, View - schematic
// LAST TIME SAVED: Jun 25 14:02:00 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module bram_icg ( clkout, clk, en );
output  clkout;

input  clk, en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(net027), .Y(net014), .B(c));
inv_tri_2_hvt I7 ( .Tb(cn), .T(c), .A(net027), .Y(net023));
inv_tri_2_hvt I5 ( .Tb(c), .T(cn), .A(en), .Y(net023));
inv_hvt I391 ( .A(net014), .Y(clkout));
inv_hvt I6 ( .A(net023), .Y(net027));
inv_hvt I4 ( .A(cn), .Y(c));
inv_hvt I3 ( .A(clk), .Y(cn));

endmodule
// Library - leafcell, Cell - bram_hbuffer_dff_2xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:02:56 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module bram_hbuffer_dff_2xbank ( bm_banksel_o, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclkrw_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [3:0]  bm_sdi_o;
output [3:0]  bm_banksel_o;
output [1:0]  bm_sclk_o;
output [7:0]  bm_sa_o;
output [3:0]  bm_sdo_o;

input [7:0]  bm_sa_i;
input [3:0]  bm_sdo_i;
input [3:0]  bm_banksel_i;
input [3:0]  bm_sdi_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net102;

wire  [0:3]  net103;



tielo I23 ( .tielo(net057));
bram_icg I47 ( .en(net74), .clk(bm_sclk_i), .clkout(net61));
bram_icg I19 ( .en(net72), .clk(bm_sclk_i), .clkout(net64));
bram_bufferx16_2inv I16_3_ ( .in(net103[0]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I16_2_ ( .in(net103[1]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I16_1_ ( .in(net103[2]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I16_0_ ( .in(net103[3]), .out(bm_sdo_o[0]));
bram_bufferx4 I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx4 I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx4 I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx4 I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx4 I22 ( .in(net64), .out(bm_sclk_o[1]));
bram_bufferx4 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx4 I13_3_ ( .in(bm_banksel_i[3]), .out(bm_banksel_o[3]));
bram_bufferx4 I13_2_ ( .in(bm_banksel_i[2]), .out(bm_banksel_o[2]));
bram_bufferx4 I13_1_ ( .in(bm_banksel_i[1]), .out(bm_banksel_o[1]));
bram_bufferx4 I13_0_ ( .in(bm_banksel_i[0]), .out(bm_banksel_o[0]));
bram_bufferx4 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx4 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx4 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx4 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx4 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx4 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx4 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx4 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx4 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx4 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx4 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx4 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx4 I18 ( .in(net61), .out(bm_sclk_o[0]));
bram_bufferx4 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));
leafcell_ml_dff_schematic I48_3_ ( .R(net057), .D(bm_sdo_i[3]),
     .CLK(bm_sclk_i), .QN(net102[0]), .Q(net103[0]));
leafcell_ml_dff_schematic I48_2_ ( .R(net057), .D(bm_sdo_i[2]),
     .CLK(bm_sclk_i), .QN(net102[1]), .Q(net103[1]));
leafcell_ml_dff_schematic I48_1_ ( .R(net057), .D(bm_sdo_i[1]),
     .CLK(bm_sclk_i), .QN(net102[2]), .Q(net103[2]));
leafcell_ml_dff_schematic I48_0_ ( .R(net057), .D(bm_sdo_i[0]),
     .CLK(bm_sclk_i), .QN(net102[3]), .Q(net103[3]));
nor2_hvt I20 ( .A(bm_banksel_i[2]), .B(bm_banksel_i[3]), .Y(net67));
nor2_hvt I49 ( .A(bm_banksel_i[0]), .B(bm_banksel_i[1]), .Y(net70));
inv_hvt I21 ( .A(net67), .Y(net72));
inv_hvt I17 ( .A(net70), .Y(net74));

endmodule
// Library - leafcell, Cell - bram_hbuffer_1xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:50:36 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module bram_hbuffer_1xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_banksel_o;
output [1:0]  bm_sdo_o;

input [1:0]  bm_sdo_i;
input [1:0]  bm_banksel_i;
input [1:0]  bm_sdi_i;
input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_bufferx2e, View - schematic
// LAST TIME SAVED: Jun 25 13:54:30 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module bram_bufferx2e ( out, en, in );
output  out;

input  en, in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net7), .Y(out));
nand2_hvt I193 ( .A(en), .Y(net7), .B(in));

endmodule
// Library - leafcell, Cell - bram_bank_logic_bot, View - schematic
// LAST TIME SAVED: Aug 31 18:48:17 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module bram_bank_logic_bot ( bm_sclkrw_o, bm_sdo_o, bm_sweb_o,
     bm_banksel_i, bm_sclk_i, bm_sclkrw_i, bm_sdo_i, bm_sweb_i );

input  bm_sclk_i, bm_sclkrw_i, bm_sweb_i;

output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sclkrw_o;

input [1:0]  bm_banksel_i;
input [1:0]  bm_sdo_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net25;

wire  [1:0]  net26;



bram_bufferx16_2inv I51_1_ ( .in(net26[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I51_0_ ( .in(net26[0]), .out(bm_sdo_o[0]));
leafcell_ml_dff_schematic I52_1_ ( .R(net020), .D(bm_sdo_i[1]),
     .CLK(bm_sclk_i), .QN(net25[0]), .Q(net26[1]));
leafcell_ml_dff_schematic I52_0_ ( .R(net020), .D(bm_sdo_i[0]),
     .CLK(bm_sclk_i), .QN(net25[1]), .Q(net26[0]));
bram_bufferx2e I54_1_ ( .in(bm_sweb_i), .en(bm_banksel_i[1]),
     .out(bm_sweb_o[1]));
bram_bufferx2e I54_0_ ( .in(bm_sweb_i), .en(bm_banksel_i[0]),
     .out(bm_sweb_o[0]));
bram_bufferx2e I48_1_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[1]),
     .out(bm_sclkrw_o[1]));
bram_bufferx2e I48_0_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[0]),
     .out(bm_sclkrw_o[0]));
tielo I55 ( .tielo(net020));

endmodule
// Library - xpmem, Cell - cram2x2x2, View - schematic
// LAST TIME SAVED: Apr 14 10:40:03 2008
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module cram2x2x2 ( q, q_b, bl, pgate_l, pgate_r, r_gnd_l, r_gnd_r,
     reset_b_l, reset_b_r, wl_l, wl_r );



output [7:0]  q_b;
output [7:0]  q;

inout [3:0]  bl;

input [1:0]  wl_r;
input [1:0]  r_gnd_r;
input [1:0]  reset_b_r;
input [1:0]  pgate_l;
input [1:0]  pgate_r;
input [1:0]  wl_l;
input [1:0]  r_gnd_l;
input [1:0]  reset_b_l;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imrgt ( .bl(bl[3:2]), .q_b(q_b[7:4]), .reset(reset_b_r[1:0]),
     .q(q[7:4]), .wl(wl_r[1:0]), .r_vdd(r_gnd_r[1:0]),
     .pgate(pgate_r[1:0]));
cram2x2 Imleft ( .reset(reset_b_l[1:0]), .r_vdd(r_gnd_l[1:0]),
     .pgate(pgate_l[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl_l[1:0]));

endmodule
// Library - xpmem, Cell - cramrow174bl4, View - schematic
// LAST TIME SAVED: Sep 25 20:58:33 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module cramrow174bl4 ( bl, pgate_l, pgate_r, reset_l, reset_r,
     vdd_cntl_l, vdd_cntl_r, wl_l, wl_r );


inout [3:0]  bl;

input [173:0]  vdd_cntl_l;
input [173:0]  reset_r;
input [173:0]  vdd_cntl_r;
input [173:0]  wl_r;
input [173:0]  pgate_r;
input [173:0]  pgate_l;
input [173:0]  wl_l;
input [173:0]  reset_l;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net073;

wire  [0:7]  net61;

wire  [0:687]  net036;

wire  [0:687]  net032;

wire  [173:0]  r_vdd;

wire  [173:0]  r_vdd_r;



cram2x2x2 xcram_85_ ( .pgate_l(pgate_l[171:170]), .wl_l(wl_l[171:170]),
     .reset_b_l(reset_l[171:170]), .r_gnd_l(r_vdd[171:170]),
     .r_gnd_r(r_vdd_r[171:170]), .pgate_r(pgate_r[171:170]),
     .wl_r(wl_r[171:170]), .reset_b_r(reset_r[171:170]),
     .q(net032[0:7]), .q_b(net036[0:7]), .bl(bl[3:0]));
cram2x2x2 xcram_84_ ( .pgate_l(pgate_l[169:168]), .wl_l(wl_l[169:168]),
     .reset_b_l(reset_l[169:168]), .r_gnd_l(r_vdd[169:168]),
     .r_gnd_r(r_vdd_r[169:168]), .pgate_r(pgate_r[169:168]),
     .wl_r(wl_r[169:168]), .reset_b_r(reset_r[169:168]),
     .q(net032[8:15]), .q_b(net036[8:15]), .bl(bl[3:0]));
cram2x2x2 xcram_83_ ( .pgate_l(pgate_l[167:166]), .wl_l(wl_l[167:166]),
     .reset_b_l(reset_l[167:166]), .r_gnd_l(r_vdd[167:166]),
     .r_gnd_r(r_vdd_r[167:166]), .pgate_r(pgate_r[167:166]),
     .wl_r(wl_r[167:166]), .reset_b_r(reset_r[167:166]),
     .q(net032[16:23]), .q_b(net036[16:23]), .bl(bl[3:0]));
cram2x2x2 xcram_82_ ( .pgate_l(pgate_l[165:164]), .wl_l(wl_l[165:164]),
     .reset_b_l(reset_l[165:164]), .r_gnd_l(r_vdd[165:164]),
     .r_gnd_r(r_vdd_r[165:164]), .pgate_r(pgate_r[165:164]),
     .wl_r(wl_r[165:164]), .reset_b_r(reset_r[165:164]),
     .q(net032[24:31]), .q_b(net036[24:31]), .bl(bl[3:0]));
cram2x2x2 xcram_81_ ( .pgate_l(pgate_l[163:162]), .wl_l(wl_l[163:162]),
     .reset_b_l(reset_l[163:162]), .r_gnd_l(r_vdd[163:162]),
     .r_gnd_r(r_vdd_r[163:162]), .pgate_r(pgate_r[163:162]),
     .wl_r(wl_r[163:162]), .reset_b_r(reset_r[163:162]),
     .q(net032[32:39]), .q_b(net036[32:39]), .bl(bl[3:0]));
cram2x2x2 xcram_80_ ( .pgate_l(pgate_l[161:160]), .wl_l(wl_l[161:160]),
     .reset_b_l(reset_l[161:160]), .r_gnd_l(r_vdd[161:160]),
     .r_gnd_r(r_vdd_r[161:160]), .pgate_r(pgate_r[161:160]),
     .wl_r(wl_r[161:160]), .reset_b_r(reset_r[161:160]),
     .q(net032[40:47]), .q_b(net036[40:47]), .bl(bl[3:0]));
cram2x2x2 xcram_79_ ( .pgate_l(pgate_l[159:158]), .wl_l(wl_l[159:158]),
     .reset_b_l(reset_l[159:158]), .r_gnd_l(r_vdd[159:158]),
     .r_gnd_r(r_vdd_r[159:158]), .pgate_r(pgate_r[159:158]),
     .wl_r(wl_r[159:158]), .reset_b_r(reset_r[159:158]),
     .q(net032[48:55]), .q_b(net036[48:55]), .bl(bl[3:0]));
cram2x2x2 xcram_78_ ( .pgate_l(pgate_l[157:156]), .wl_l(wl_l[157:156]),
     .reset_b_l(reset_l[157:156]), .r_gnd_l(r_vdd[157:156]),
     .r_gnd_r(r_vdd_r[157:156]), .pgate_r(pgate_r[157:156]),
     .wl_r(wl_r[157:156]), .reset_b_r(reset_r[157:156]),
     .q(net032[56:63]), .q_b(net036[56:63]), .bl(bl[3:0]));
cram2x2x2 xcram_77_ ( .pgate_l(pgate_l[155:154]), .wl_l(wl_l[155:154]),
     .reset_b_l(reset_l[155:154]), .r_gnd_l(r_vdd[155:154]),
     .r_gnd_r(r_vdd_r[155:154]), .pgate_r(pgate_r[155:154]),
     .wl_r(wl_r[155:154]), .reset_b_r(reset_r[155:154]),
     .q(net032[64:71]), .q_b(net036[64:71]), .bl(bl[3:0]));
cram2x2x2 xcram_76_ ( .pgate_l(pgate_l[153:152]), .wl_l(wl_l[153:152]),
     .reset_b_l(reset_l[153:152]), .r_gnd_l(r_vdd[153:152]),
     .r_gnd_r(r_vdd_r[153:152]), .pgate_r(pgate_r[153:152]),
     .wl_r(wl_r[153:152]), .reset_b_r(reset_r[153:152]),
     .q(net032[72:79]), .q_b(net036[72:79]), .bl(bl[3:0]));
cram2x2x2 xcram_75_ ( .pgate_l(pgate_l[151:150]), .wl_l(wl_l[151:150]),
     .reset_b_l(reset_l[151:150]), .r_gnd_l(r_vdd[151:150]),
     .r_gnd_r(r_vdd_r[151:150]), .pgate_r(pgate_r[151:150]),
     .wl_r(wl_r[151:150]), .reset_b_r(reset_r[151:150]),
     .q(net032[80:87]), .q_b(net036[80:87]), .bl(bl[3:0]));
cram2x2x2 xcram_74_ ( .pgate_l(pgate_l[149:148]), .wl_l(wl_l[149:148]),
     .reset_b_l(reset_l[149:148]), .r_gnd_l(r_vdd[149:148]),
     .r_gnd_r(r_vdd_r[149:148]), .pgate_r(pgate_r[149:148]),
     .wl_r(wl_r[149:148]), .reset_b_r(reset_r[149:148]),
     .q(net032[88:95]), .q_b(net036[88:95]), .bl(bl[3:0]));
cram2x2x2 xcram_73_ ( .pgate_l(pgate_l[147:146]), .wl_l(wl_l[147:146]),
     .reset_b_l(reset_l[147:146]), .r_gnd_l(r_vdd[147:146]),
     .r_gnd_r(r_vdd_r[147:146]), .pgate_r(pgate_r[147:146]),
     .wl_r(wl_r[147:146]), .reset_b_r(reset_r[147:146]),
     .q(net032[96:103]), .q_b(net036[96:103]), .bl(bl[3:0]));
cram2x2x2 xcram_72_ ( .pgate_l(pgate_l[145:144]), .wl_l(wl_l[145:144]),
     .reset_b_l(reset_l[145:144]), .r_gnd_l(r_vdd[145:144]),
     .r_gnd_r(r_vdd_r[145:144]), .pgate_r(pgate_r[145:144]),
     .wl_r(wl_r[145:144]), .reset_b_r(reset_r[145:144]),
     .q(net032[104:111]), .q_b(net036[104:111]), .bl(bl[3:0]));
cram2x2x2 xcram_71_ ( .pgate_l(pgate_l[143:142]), .wl_l(wl_l[143:142]),
     .reset_b_l(reset_l[143:142]), .r_gnd_l(r_vdd[143:142]),
     .r_gnd_r(r_vdd_r[143:142]), .pgate_r(pgate_r[143:142]),
     .wl_r(wl_r[143:142]), .reset_b_r(reset_r[143:142]),
     .q(net032[112:119]), .q_b(net036[112:119]), .bl(bl[3:0]));
cram2x2x2 xcram_70_ ( .pgate_l(pgate_l[141:140]), .wl_l(wl_l[141:140]),
     .reset_b_l(reset_l[141:140]), .r_gnd_l(r_vdd[141:140]),
     .r_gnd_r(r_vdd_r[141:140]), .pgate_r(pgate_r[141:140]),
     .wl_r(wl_r[141:140]), .reset_b_r(reset_r[141:140]),
     .q(net032[120:127]), .q_b(net036[120:127]), .bl(bl[3:0]));
cram2x2x2 xcram_69_ ( .pgate_l(pgate_l[139:138]), .wl_l(wl_l[139:138]),
     .reset_b_l(reset_l[139:138]), .r_gnd_l(r_vdd[139:138]),
     .r_gnd_r(r_vdd_r[139:138]), .pgate_r(pgate_r[139:138]),
     .wl_r(wl_r[139:138]), .reset_b_r(reset_r[139:138]),
     .q(net032[128:135]), .q_b(net036[128:135]), .bl(bl[3:0]));
cram2x2x2 xcram_68_ ( .pgate_l(pgate_l[137:136]), .wl_l(wl_l[137:136]),
     .reset_b_l(reset_l[137:136]), .r_gnd_l(r_vdd[137:136]),
     .r_gnd_r(r_vdd_r[137:136]), .pgate_r(pgate_r[137:136]),
     .wl_r(wl_r[137:136]), .reset_b_r(reset_r[137:136]),
     .q(net032[136:143]), .q_b(net036[136:143]), .bl(bl[3:0]));
cram2x2x2 xcram_67_ ( .pgate_l(pgate_l[135:134]), .wl_l(wl_l[135:134]),
     .reset_b_l(reset_l[135:134]), .r_gnd_l(r_vdd[135:134]),
     .r_gnd_r(r_vdd_r[135:134]), .pgate_r(pgate_r[135:134]),
     .wl_r(wl_r[135:134]), .reset_b_r(reset_r[135:134]),
     .q(net032[144:151]), .q_b(net036[144:151]), .bl(bl[3:0]));
cram2x2x2 xcram_66_ ( .pgate_l(pgate_l[133:132]), .wl_l(wl_l[133:132]),
     .reset_b_l(reset_l[133:132]), .r_gnd_l(r_vdd[133:132]),
     .r_gnd_r(r_vdd_r[133:132]), .pgate_r(pgate_r[133:132]),
     .wl_r(wl_r[133:132]), .reset_b_r(reset_r[133:132]),
     .q(net032[152:159]), .q_b(net036[152:159]), .bl(bl[3:0]));
cram2x2x2 xcram_65_ ( .pgate_l(pgate_l[131:130]), .wl_l(wl_l[131:130]),
     .reset_b_l(reset_l[131:130]), .r_gnd_l(r_vdd[131:130]),
     .r_gnd_r(r_vdd_r[131:130]), .pgate_r(pgate_r[131:130]),
     .wl_r(wl_r[131:130]), .reset_b_r(reset_r[131:130]),
     .q(net032[160:167]), .q_b(net036[160:167]), .bl(bl[3:0]));
cram2x2x2 xcram_64_ ( .pgate_l(pgate_l[129:128]), .wl_l(wl_l[129:128]),
     .reset_b_l(reset_l[129:128]), .r_gnd_l(r_vdd[129:128]),
     .r_gnd_r(r_vdd_r[129:128]), .pgate_r(pgate_r[129:128]),
     .wl_r(wl_r[129:128]), .reset_b_r(reset_r[129:128]),
     .q(net032[168:175]), .q_b(net036[168:175]), .bl(bl[3:0]));
cram2x2x2 xcram_63_ ( .pgate_l(pgate_l[127:126]), .wl_l(wl_l[127:126]),
     .reset_b_l(reset_l[127:126]), .r_gnd_l(r_vdd[127:126]),
     .r_gnd_r(r_vdd_r[127:126]), .pgate_r(pgate_r[127:126]),
     .wl_r(wl_r[127:126]), .reset_b_r(reset_r[127:126]),
     .q(net032[176:183]), .q_b(net036[176:183]), .bl(bl[3:0]));
cram2x2x2 xcram_62_ ( .pgate_l(pgate_l[125:124]), .wl_l(wl_l[125:124]),
     .reset_b_l(reset_l[125:124]), .r_gnd_l(r_vdd[125:124]),
     .r_gnd_r(r_vdd_r[125:124]), .pgate_r(pgate_r[125:124]),
     .wl_r(wl_r[125:124]), .reset_b_r(reset_r[125:124]),
     .q(net032[184:191]), .q_b(net036[184:191]), .bl(bl[3:0]));
cram2x2x2 xcram_61_ ( .pgate_l(pgate_l[123:122]), .wl_l(wl_l[123:122]),
     .reset_b_l(reset_l[123:122]), .r_gnd_l(r_vdd[123:122]),
     .r_gnd_r(r_vdd_r[123:122]), .pgate_r(pgate_r[123:122]),
     .wl_r(wl_r[123:122]), .reset_b_r(reset_r[123:122]),
     .q(net032[192:199]), .q_b(net036[192:199]), .bl(bl[3:0]));
cram2x2x2 xcram_60_ ( .pgate_l(pgate_l[121:120]), .wl_l(wl_l[121:120]),
     .reset_b_l(reset_l[121:120]), .r_gnd_l(r_vdd[121:120]),
     .r_gnd_r(r_vdd_r[121:120]), .pgate_r(pgate_r[121:120]),
     .wl_r(wl_r[121:120]), .reset_b_r(reset_r[121:120]),
     .q(net032[200:207]), .q_b(net036[200:207]), .bl(bl[3:0]));
cram2x2x2 xcram_59_ ( .pgate_l(pgate_l[119:118]), .wl_l(wl_l[119:118]),
     .reset_b_l(reset_l[119:118]), .r_gnd_l(r_vdd[119:118]),
     .r_gnd_r(r_vdd_r[119:118]), .pgate_r(pgate_r[119:118]),
     .wl_r(wl_r[119:118]), .reset_b_r(reset_r[119:118]),
     .q(net032[208:215]), .q_b(net036[208:215]), .bl(bl[3:0]));
cram2x2x2 xcram_58_ ( .pgate_l(pgate_l[117:116]), .wl_l(wl_l[117:116]),
     .reset_b_l(reset_l[117:116]), .r_gnd_l(r_vdd[117:116]),
     .r_gnd_r(r_vdd_r[117:116]), .pgate_r(pgate_r[117:116]),
     .wl_r(wl_r[117:116]), .reset_b_r(reset_r[117:116]),
     .q(net032[216:223]), .q_b(net036[216:223]), .bl(bl[3:0]));
cram2x2x2 xcram_57_ ( .pgate_l(pgate_l[115:114]), .wl_l(wl_l[115:114]),
     .reset_b_l(reset_l[115:114]), .r_gnd_l(r_vdd[115:114]),
     .r_gnd_r(r_vdd_r[115:114]), .pgate_r(pgate_r[115:114]),
     .wl_r(wl_r[115:114]), .reset_b_r(reset_r[115:114]),
     .q(net032[224:231]), .q_b(net036[224:231]), .bl(bl[3:0]));
cram2x2x2 xcram_56_ ( .pgate_l(pgate_l[113:112]), .wl_l(wl_l[113:112]),
     .reset_b_l(reset_l[113:112]), .r_gnd_l(r_vdd[113:112]),
     .r_gnd_r(r_vdd_r[113:112]), .pgate_r(pgate_r[113:112]),
     .wl_r(wl_r[113:112]), .reset_b_r(reset_r[113:112]),
     .q(net032[232:239]), .q_b(net036[232:239]), .bl(bl[3:0]));
cram2x2x2 xcram_55_ ( .pgate_l(pgate_l[111:110]), .wl_l(wl_l[111:110]),
     .reset_b_l(reset_l[111:110]), .r_gnd_l(r_vdd[111:110]),
     .r_gnd_r(r_vdd_r[111:110]), .pgate_r(pgate_r[111:110]),
     .wl_r(wl_r[111:110]), .reset_b_r(reset_r[111:110]),
     .q(net032[240:247]), .q_b(net036[240:247]), .bl(bl[3:0]));
cram2x2x2 xcram_54_ ( .pgate_l(pgate_l[109:108]), .wl_l(wl_l[109:108]),
     .reset_b_l(reset_l[109:108]), .r_gnd_l(r_vdd[109:108]),
     .r_gnd_r(r_vdd_r[109:108]), .pgate_r(pgate_r[109:108]),
     .wl_r(wl_r[109:108]), .reset_b_r(reset_r[109:108]),
     .q(net032[248:255]), .q_b(net036[248:255]), .bl(bl[3:0]));
cram2x2x2 xcram_53_ ( .pgate_l(pgate_l[107:106]), .wl_l(wl_l[107:106]),
     .reset_b_l(reset_l[107:106]), .r_gnd_l(r_vdd[107:106]),
     .r_gnd_r(r_vdd_r[107:106]), .pgate_r(pgate_r[107:106]),
     .wl_r(wl_r[107:106]), .reset_b_r(reset_r[107:106]),
     .q(net032[256:263]), .q_b(net036[256:263]), .bl(bl[3:0]));
cram2x2x2 xcram_52_ ( .pgate_l(pgate_l[105:104]), .wl_l(wl_l[105:104]),
     .reset_b_l(reset_l[105:104]), .r_gnd_l(r_vdd[105:104]),
     .r_gnd_r(r_vdd_r[105:104]), .pgate_r(pgate_r[105:104]),
     .wl_r(wl_r[105:104]), .reset_b_r(reset_r[105:104]),
     .q(net032[264:271]), .q_b(net036[264:271]), .bl(bl[3:0]));
cram2x2x2 xcram_51_ ( .pgate_l(pgate_l[103:102]), .wl_l(wl_l[103:102]),
     .reset_b_l(reset_l[103:102]), .r_gnd_l(r_vdd[103:102]),
     .r_gnd_r(r_vdd_r[103:102]), .pgate_r(pgate_r[103:102]),
     .wl_r(wl_r[103:102]), .reset_b_r(reset_r[103:102]),
     .q(net032[272:279]), .q_b(net036[272:279]), .bl(bl[3:0]));
cram2x2x2 xcram_50_ ( .pgate_l(pgate_l[101:100]), .wl_l(wl_l[101:100]),
     .reset_b_l(reset_l[101:100]), .r_gnd_l(r_vdd[101:100]),
     .r_gnd_r(r_vdd_r[101:100]), .pgate_r(pgate_r[101:100]),
     .wl_r(wl_r[101:100]), .reset_b_r(reset_r[101:100]),
     .q(net032[280:287]), .q_b(net036[280:287]), .bl(bl[3:0]));
cram2x2x2 xcram_49_ ( .pgate_l(pgate_l[99:98]), .wl_l(wl_l[99:98]),
     .reset_b_l(reset_l[99:98]), .r_gnd_l(r_vdd[99:98]),
     .r_gnd_r(r_vdd_r[99:98]), .pgate_r(pgate_r[99:98]),
     .wl_r(wl_r[99:98]), .reset_b_r(reset_r[99:98]),
     .q(net032[288:295]), .q_b(net036[288:295]), .bl(bl[3:0]));
cram2x2x2 xcram_48_ ( .pgate_l(pgate_l[97:96]), .wl_l(wl_l[97:96]),
     .reset_b_l(reset_l[97:96]), .r_gnd_l(r_vdd[97:96]),
     .r_gnd_r(r_vdd_r[97:96]), .pgate_r(pgate_r[97:96]),
     .wl_r(wl_r[97:96]), .reset_b_r(reset_r[97:96]),
     .q(net032[296:303]), .q_b(net036[296:303]), .bl(bl[3:0]));
cram2x2x2 xcram_47_ ( .pgate_l(pgate_l[95:94]), .wl_l(wl_l[95:94]),
     .reset_b_l(reset_l[95:94]), .r_gnd_l(r_vdd[95:94]),
     .r_gnd_r(r_vdd_r[95:94]), .pgate_r(pgate_r[95:94]),
     .wl_r(wl_r[95:94]), .reset_b_r(reset_r[95:94]),
     .q(net032[304:311]), .q_b(net036[304:311]), .bl(bl[3:0]));
cram2x2x2 xcram_46_ ( .pgate_l(pgate_l[93:92]), .wl_l(wl_l[93:92]),
     .reset_b_l(reset_l[93:92]), .r_gnd_l(r_vdd[93:92]),
     .r_gnd_r(r_vdd_r[93:92]), .pgate_r(pgate_r[93:92]),
     .wl_r(wl_r[93:92]), .reset_b_r(reset_r[93:92]),
     .q(net032[312:319]), .q_b(net036[312:319]), .bl(bl[3:0]));
cram2x2x2 xcram_45_ ( .pgate_l(pgate_l[91:90]), .wl_l(wl_l[91:90]),
     .reset_b_l(reset_l[91:90]), .r_gnd_l(r_vdd[91:90]),
     .r_gnd_r(r_vdd_r[91:90]), .pgate_r(pgate_r[91:90]),
     .wl_r(wl_r[91:90]), .reset_b_r(reset_r[91:90]),
     .q(net032[320:327]), .q_b(net036[320:327]), .bl(bl[3:0]));
cram2x2x2 xcram_44_ ( .pgate_l(pgate_l[89:88]), .wl_l(wl_l[89:88]),
     .reset_b_l(reset_l[89:88]), .r_gnd_l(r_vdd[89:88]),
     .r_gnd_r(r_vdd_r[89:88]), .pgate_r(pgate_r[89:88]),
     .wl_r(wl_r[89:88]), .reset_b_r(reset_r[89:88]),
     .q(net032[328:335]), .q_b(net036[328:335]), .bl(bl[3:0]));
cram2x2x2 xcram_43_ ( .pgate_l(pgate_l[87:86]), .wl_l(wl_l[87:86]),
     .reset_b_l(reset_l[87:86]), .r_gnd_l(r_vdd[87:86]),
     .r_gnd_r(r_vdd_r[87:86]), .pgate_r(pgate_r[87:86]),
     .wl_r(wl_r[87:86]), .reset_b_r(reset_r[87:86]),
     .q(net032[336:343]), .q_b(net036[336:343]), .bl(bl[3:0]));
cram2x2x2 xcram_42_ ( .pgate_l(pgate_l[85:84]), .wl_l(wl_l[85:84]),
     .reset_b_l(reset_l[85:84]), .r_gnd_l(r_vdd[85:84]),
     .r_gnd_r(r_vdd_r[85:84]), .pgate_r(pgate_r[85:84]),
     .wl_r(wl_r[85:84]), .reset_b_r(reset_r[85:84]),
     .q(net032[344:351]), .q_b(net036[344:351]), .bl(bl[3:0]));
cram2x2x2 xcram_41_ ( .pgate_l(pgate_l[83:82]), .wl_l(wl_l[83:82]),
     .reset_b_l(reset_l[83:82]), .r_gnd_l(r_vdd[83:82]),
     .r_gnd_r(r_vdd_r[83:82]), .pgate_r(pgate_r[83:82]),
     .wl_r(wl_r[83:82]), .reset_b_r(reset_r[83:82]),
     .q(net032[352:359]), .q_b(net036[352:359]), .bl(bl[3:0]));
cram2x2x2 xcram_40_ ( .pgate_l(pgate_l[81:80]), .wl_l(wl_l[81:80]),
     .reset_b_l(reset_l[81:80]), .r_gnd_l(r_vdd[81:80]),
     .r_gnd_r(r_vdd_r[81:80]), .pgate_r(pgate_r[81:80]),
     .wl_r(wl_r[81:80]), .reset_b_r(reset_r[81:80]),
     .q(net032[360:367]), .q_b(net036[360:367]), .bl(bl[3:0]));
cram2x2x2 xcram_39_ ( .pgate_l(pgate_l[79:78]), .wl_l(wl_l[79:78]),
     .reset_b_l(reset_l[79:78]), .r_gnd_l(r_vdd[79:78]),
     .r_gnd_r(r_vdd_r[79:78]), .pgate_r(pgate_r[79:78]),
     .wl_r(wl_r[79:78]), .reset_b_r(reset_r[79:78]),
     .q(net032[368:375]), .q_b(net036[368:375]), .bl(bl[3:0]));
cram2x2x2 xcram_38_ ( .pgate_l(pgate_l[77:76]), .wl_l(wl_l[77:76]),
     .reset_b_l(reset_l[77:76]), .r_gnd_l(r_vdd[77:76]),
     .r_gnd_r(r_vdd_r[77:76]), .pgate_r(pgate_r[77:76]),
     .wl_r(wl_r[77:76]), .reset_b_r(reset_r[77:76]),
     .q(net032[376:383]), .q_b(net036[376:383]), .bl(bl[3:0]));
cram2x2x2 xcram_37_ ( .pgate_l(pgate_l[75:74]), .wl_l(wl_l[75:74]),
     .reset_b_l(reset_l[75:74]), .r_gnd_l(r_vdd[75:74]),
     .r_gnd_r(r_vdd_r[75:74]), .pgate_r(pgate_r[75:74]),
     .wl_r(wl_r[75:74]), .reset_b_r(reset_r[75:74]),
     .q(net032[384:391]), .q_b(net036[384:391]), .bl(bl[3:0]));
cram2x2x2 xcram_36_ ( .pgate_l(pgate_l[73:72]), .wl_l(wl_l[73:72]),
     .reset_b_l(reset_l[73:72]), .r_gnd_l(r_vdd[73:72]),
     .r_gnd_r(r_vdd_r[73:72]), .pgate_r(pgate_r[73:72]),
     .wl_r(wl_r[73:72]), .reset_b_r(reset_r[73:72]),
     .q(net032[392:399]), .q_b(net036[392:399]), .bl(bl[3:0]));
cram2x2x2 xcram_35_ ( .pgate_l(pgate_l[71:70]), .wl_l(wl_l[71:70]),
     .reset_b_l(reset_l[71:70]), .r_gnd_l(r_vdd[71:70]),
     .r_gnd_r(r_vdd_r[71:70]), .pgate_r(pgate_r[71:70]),
     .wl_r(wl_r[71:70]), .reset_b_r(reset_r[71:70]),
     .q(net032[400:407]), .q_b(net036[400:407]), .bl(bl[3:0]));
cram2x2x2 xcram_34_ ( .pgate_l(pgate_l[69:68]), .wl_l(wl_l[69:68]),
     .reset_b_l(reset_l[69:68]), .r_gnd_l(r_vdd[69:68]),
     .r_gnd_r(r_vdd_r[69:68]), .pgate_r(pgate_r[69:68]),
     .wl_r(wl_r[69:68]), .reset_b_r(reset_r[69:68]),
     .q(net032[408:415]), .q_b(net036[408:415]), .bl(bl[3:0]));
cram2x2x2 xcram_33_ ( .pgate_l(pgate_l[67:66]), .wl_l(wl_l[67:66]),
     .reset_b_l(reset_l[67:66]), .r_gnd_l(r_vdd[67:66]),
     .r_gnd_r(r_vdd_r[67:66]), .pgate_r(pgate_r[67:66]),
     .wl_r(wl_r[67:66]), .reset_b_r(reset_r[67:66]),
     .q(net032[416:423]), .q_b(net036[416:423]), .bl(bl[3:0]));
cram2x2x2 xcram_32_ ( .pgate_l(pgate_l[65:64]), .wl_l(wl_l[65:64]),
     .reset_b_l(reset_l[65:64]), .r_gnd_l(r_vdd[65:64]),
     .r_gnd_r(r_vdd_r[65:64]), .pgate_r(pgate_r[65:64]),
     .wl_r(wl_r[65:64]), .reset_b_r(reset_r[65:64]),
     .q(net032[424:431]), .q_b(net036[424:431]), .bl(bl[3:0]));
cram2x2x2 xcram_31_ ( .pgate_l(pgate_l[63:62]), .wl_l(wl_l[63:62]),
     .reset_b_l(reset_l[63:62]), .r_gnd_l(r_vdd[63:62]),
     .r_gnd_r(r_vdd_r[63:62]), .pgate_r(pgate_r[63:62]),
     .wl_r(wl_r[63:62]), .reset_b_r(reset_r[63:62]),
     .q(net032[432:439]), .q_b(net036[432:439]), .bl(bl[3:0]));
cram2x2x2 xcram_30_ ( .pgate_l(pgate_l[61:60]), .wl_l(wl_l[61:60]),
     .reset_b_l(reset_l[61:60]), .r_gnd_l(r_vdd[61:60]),
     .r_gnd_r(r_vdd_r[61:60]), .pgate_r(pgate_r[61:60]),
     .wl_r(wl_r[61:60]), .reset_b_r(reset_r[61:60]),
     .q(net032[440:447]), .q_b(net036[440:447]), .bl(bl[3:0]));
cram2x2x2 xcram_29_ ( .pgate_l(pgate_l[59:58]), .wl_l(wl_l[59:58]),
     .reset_b_l(reset_l[59:58]), .r_gnd_l(r_vdd[59:58]),
     .r_gnd_r(r_vdd_r[59:58]), .pgate_r(pgate_r[59:58]),
     .wl_r(wl_r[59:58]), .reset_b_r(reset_r[59:58]),
     .q(net032[448:455]), .q_b(net036[448:455]), .bl(bl[3:0]));
cram2x2x2 xcram_28_ ( .pgate_l(pgate_l[57:56]), .wl_l(wl_l[57:56]),
     .reset_b_l(reset_l[57:56]), .r_gnd_l(r_vdd[57:56]),
     .r_gnd_r(r_vdd_r[57:56]), .pgate_r(pgate_r[57:56]),
     .wl_r(wl_r[57:56]), .reset_b_r(reset_r[57:56]),
     .q(net032[456:463]), .q_b(net036[456:463]), .bl(bl[3:0]));
cram2x2x2 xcram_27_ ( .pgate_l(pgate_l[55:54]), .wl_l(wl_l[55:54]),
     .reset_b_l(reset_l[55:54]), .r_gnd_l(r_vdd[55:54]),
     .r_gnd_r(r_vdd_r[55:54]), .pgate_r(pgate_r[55:54]),
     .wl_r(wl_r[55:54]), .reset_b_r(reset_r[55:54]),
     .q(net032[464:471]), .q_b(net036[464:471]), .bl(bl[3:0]));
cram2x2x2 xcram_26_ ( .pgate_l(pgate_l[53:52]), .wl_l(wl_l[53:52]),
     .reset_b_l(reset_l[53:52]), .r_gnd_l(r_vdd[53:52]),
     .r_gnd_r(r_vdd_r[53:52]), .pgate_r(pgate_r[53:52]),
     .wl_r(wl_r[53:52]), .reset_b_r(reset_r[53:52]),
     .q(net032[472:479]), .q_b(net036[472:479]), .bl(bl[3:0]));
cram2x2x2 xcram_25_ ( .pgate_l(pgate_l[51:50]), .wl_l(wl_l[51:50]),
     .reset_b_l(reset_l[51:50]), .r_gnd_l(r_vdd[51:50]),
     .r_gnd_r(r_vdd_r[51:50]), .pgate_r(pgate_r[51:50]),
     .wl_r(wl_r[51:50]), .reset_b_r(reset_r[51:50]),
     .q(net032[480:487]), .q_b(net036[480:487]), .bl(bl[3:0]));
cram2x2x2 xcram_24_ ( .pgate_l(pgate_l[49:48]), .wl_l(wl_l[49:48]),
     .reset_b_l(reset_l[49:48]), .r_gnd_l(r_vdd[49:48]),
     .r_gnd_r(r_vdd_r[49:48]), .pgate_r(pgate_r[49:48]),
     .wl_r(wl_r[49:48]), .reset_b_r(reset_r[49:48]),
     .q(net032[488:495]), .q_b(net036[488:495]), .bl(bl[3:0]));
cram2x2x2 xcram_23_ ( .pgate_l(pgate_l[47:46]), .wl_l(wl_l[47:46]),
     .reset_b_l(reset_l[47:46]), .r_gnd_l(r_vdd[47:46]),
     .r_gnd_r(r_vdd_r[47:46]), .pgate_r(pgate_r[47:46]),
     .wl_r(wl_r[47:46]), .reset_b_r(reset_r[47:46]),
     .q(net032[496:503]), .q_b(net036[496:503]), .bl(bl[3:0]));
cram2x2x2 xcram_22_ ( .pgate_l(pgate_l[45:44]), .wl_l(wl_l[45:44]),
     .reset_b_l(reset_l[45:44]), .r_gnd_l(r_vdd[45:44]),
     .r_gnd_r(r_vdd_r[45:44]), .pgate_r(pgate_r[45:44]),
     .wl_r(wl_r[45:44]), .reset_b_r(reset_r[45:44]),
     .q(net032[504:511]), .q_b(net036[504:511]), .bl(bl[3:0]));
cram2x2x2 xcram_21_ ( .pgate_l(pgate_l[43:42]), .wl_l(wl_l[43:42]),
     .reset_b_l(reset_l[43:42]), .r_gnd_l(r_vdd[43:42]),
     .r_gnd_r(r_vdd_r[43:42]), .pgate_r(pgate_r[43:42]),
     .wl_r(wl_r[43:42]), .reset_b_r(reset_r[43:42]),
     .q(net032[512:519]), .q_b(net036[512:519]), .bl(bl[3:0]));
cram2x2x2 xcram_20_ ( .pgate_l(pgate_l[41:40]), .wl_l(wl_l[41:40]),
     .reset_b_l(reset_l[41:40]), .r_gnd_l(r_vdd[41:40]),
     .r_gnd_r(r_vdd_r[41:40]), .pgate_r(pgate_r[41:40]),
     .wl_r(wl_r[41:40]), .reset_b_r(reset_r[41:40]),
     .q(net032[520:527]), .q_b(net036[520:527]), .bl(bl[3:0]));
cram2x2x2 xcram_19_ ( .pgate_l(pgate_l[39:38]), .wl_l(wl_l[39:38]),
     .reset_b_l(reset_l[39:38]), .r_gnd_l(r_vdd[39:38]),
     .r_gnd_r(r_vdd_r[39:38]), .pgate_r(pgate_r[39:38]),
     .wl_r(wl_r[39:38]), .reset_b_r(reset_r[39:38]),
     .q(net032[528:535]), .q_b(net036[528:535]), .bl(bl[3:0]));
cram2x2x2 xcram_18_ ( .pgate_l(pgate_l[37:36]), .wl_l(wl_l[37:36]),
     .reset_b_l(reset_l[37:36]), .r_gnd_l(r_vdd[37:36]),
     .r_gnd_r(r_vdd_r[37:36]), .pgate_r(pgate_r[37:36]),
     .wl_r(wl_r[37:36]), .reset_b_r(reset_r[37:36]),
     .q(net032[536:543]), .q_b(net036[536:543]), .bl(bl[3:0]));
cram2x2x2 xcram_17_ ( .pgate_l(pgate_l[35:34]), .wl_l(wl_l[35:34]),
     .reset_b_l(reset_l[35:34]), .r_gnd_l(r_vdd[35:34]),
     .r_gnd_r(r_vdd_r[35:34]), .pgate_r(pgate_r[35:34]),
     .wl_r(wl_r[35:34]), .reset_b_r(reset_r[35:34]),
     .q(net032[544:551]), .q_b(net036[544:551]), .bl(bl[3:0]));
cram2x2x2 xcram_16_ ( .pgate_l(pgate_l[33:32]), .wl_l(wl_l[33:32]),
     .reset_b_l(reset_l[33:32]), .r_gnd_l(r_vdd[33:32]),
     .r_gnd_r(r_vdd_r[33:32]), .pgate_r(pgate_r[33:32]),
     .wl_r(wl_r[33:32]), .reset_b_r(reset_r[33:32]),
     .q(net032[552:559]), .q_b(net036[552:559]), .bl(bl[3:0]));
cram2x2x2 xcram_15_ ( .pgate_l(pgate_l[31:30]), .wl_l(wl_l[31:30]),
     .reset_b_l(reset_l[31:30]), .r_gnd_l(r_vdd[31:30]),
     .r_gnd_r(r_vdd_r[31:30]), .pgate_r(pgate_r[31:30]),
     .wl_r(wl_r[31:30]), .reset_b_r(reset_r[31:30]),
     .q(net032[560:567]), .q_b(net036[560:567]), .bl(bl[3:0]));
cram2x2x2 xcram_14_ ( .pgate_l(pgate_l[29:28]), .wl_l(wl_l[29:28]),
     .reset_b_l(reset_l[29:28]), .r_gnd_l(r_vdd[29:28]),
     .r_gnd_r(r_vdd_r[29:28]), .pgate_r(pgate_r[29:28]),
     .wl_r(wl_r[29:28]), .reset_b_r(reset_r[29:28]),
     .q(net032[568:575]), .q_b(net036[568:575]), .bl(bl[3:0]));
cram2x2x2 xcram_13_ ( .pgate_l(pgate_l[27:26]), .wl_l(wl_l[27:26]),
     .reset_b_l(reset_l[27:26]), .r_gnd_l(r_vdd[27:26]),
     .r_gnd_r(r_vdd_r[27:26]), .pgate_r(pgate_r[27:26]),
     .wl_r(wl_r[27:26]), .reset_b_r(reset_r[27:26]),
     .q(net032[576:583]), .q_b(net036[576:583]), .bl(bl[3:0]));
cram2x2x2 xcram_12_ ( .pgate_l(pgate_l[25:24]), .wl_l(wl_l[25:24]),
     .reset_b_l(reset_l[25:24]), .r_gnd_l(r_vdd[25:24]),
     .r_gnd_r(r_vdd_r[25:24]), .pgate_r(pgate_r[25:24]),
     .wl_r(wl_r[25:24]), .reset_b_r(reset_r[25:24]),
     .q(net032[584:591]), .q_b(net036[584:591]), .bl(bl[3:0]));
cram2x2x2 xcram_11_ ( .pgate_l(pgate_l[23:22]), .wl_l(wl_l[23:22]),
     .reset_b_l(reset_l[23:22]), .r_gnd_l(r_vdd[23:22]),
     .r_gnd_r(r_vdd_r[23:22]), .pgate_r(pgate_r[23:22]),
     .wl_r(wl_r[23:22]), .reset_b_r(reset_r[23:22]),
     .q(net032[592:599]), .q_b(net036[592:599]), .bl(bl[3:0]));
cram2x2x2 xcram_10_ ( .pgate_l(pgate_l[21:20]), .wl_l(wl_l[21:20]),
     .reset_b_l(reset_l[21:20]), .r_gnd_l(r_vdd[21:20]),
     .r_gnd_r(r_vdd_r[21:20]), .pgate_r(pgate_r[21:20]),
     .wl_r(wl_r[21:20]), .reset_b_r(reset_r[21:20]),
     .q(net032[600:607]), .q_b(net036[600:607]), .bl(bl[3:0]));
cram2x2x2 xcram_9_ ( .pgate_l(pgate_l[19:18]), .wl_l(wl_l[19:18]),
     .reset_b_l(reset_l[19:18]), .r_gnd_l(r_vdd[19:18]),
     .r_gnd_r(r_vdd_r[19:18]), .pgate_r(pgate_r[19:18]),
     .wl_r(wl_r[19:18]), .reset_b_r(reset_r[19:18]),
     .q(net032[608:615]), .q_b(net036[608:615]), .bl(bl[3:0]));
cram2x2x2 xcram_8_ ( .pgate_l(pgate_l[17:16]), .wl_l(wl_l[17:16]),
     .reset_b_l(reset_l[17:16]), .r_gnd_l(r_vdd[17:16]),
     .r_gnd_r(r_vdd_r[17:16]), .pgate_r(pgate_r[17:16]),
     .wl_r(wl_r[17:16]), .reset_b_r(reset_r[17:16]),
     .q(net032[616:623]), .q_b(net036[616:623]), .bl(bl[3:0]));
cram2x2x2 xcram_7_ ( .pgate_l(pgate_l[15:14]), .wl_l(wl_l[15:14]),
     .reset_b_l(reset_l[15:14]), .r_gnd_l(r_vdd[15:14]),
     .r_gnd_r(r_vdd_r[15:14]), .pgate_r(pgate_r[15:14]),
     .wl_r(wl_r[15:14]), .reset_b_r(reset_r[15:14]),
     .q(net032[624:631]), .q_b(net036[624:631]), .bl(bl[3:0]));
cram2x2x2 xcram_6_ ( .pgate_l(pgate_l[13:12]), .wl_l(wl_l[13:12]),
     .reset_b_l(reset_l[13:12]), .r_gnd_l(r_vdd[13:12]),
     .r_gnd_r(r_vdd_r[13:12]), .pgate_r(pgate_r[13:12]),
     .wl_r(wl_r[13:12]), .reset_b_r(reset_r[13:12]),
     .q(net032[632:639]), .q_b(net036[632:639]), .bl(bl[3:0]));
cram2x2x2 xcram_5_ ( .pgate_l(pgate_l[11:10]), .wl_l(wl_l[11:10]),
     .reset_b_l(reset_l[11:10]), .r_gnd_l(r_vdd[11:10]),
     .r_gnd_r(r_vdd_r[11:10]), .pgate_r(pgate_r[11:10]),
     .wl_r(wl_r[11:10]), .reset_b_r(reset_r[11:10]),
     .q(net032[640:647]), .q_b(net036[640:647]), .bl(bl[3:0]));
cram2x2x2 xcram_4_ ( .pgate_l(pgate_l[9:8]), .wl_l(wl_l[9:8]),
     .reset_b_l(reset_l[9:8]), .r_gnd_l(r_vdd[9:8]),
     .r_gnd_r(r_vdd_r[9:8]), .pgate_r(pgate_r[9:8]), .wl_r(wl_r[9:8]),
     .reset_b_r(reset_r[9:8]), .q(net032[648:655]),
     .q_b(net036[648:655]), .bl(bl[3:0]));
cram2x2x2 xcram_3_ ( .pgate_l(pgate_l[7:6]), .wl_l(wl_l[7:6]),
     .reset_b_l(reset_l[7:6]), .r_gnd_l(r_vdd[7:6]),
     .r_gnd_r(r_vdd_r[7:6]), .pgate_r(pgate_r[7:6]), .wl_r(wl_r[7:6]),
     .reset_b_r(reset_r[7:6]), .q(net032[656:663]),
     .q_b(net036[656:663]), .bl(bl[3:0]));
cram2x2x2 xcram_2_ ( .pgate_l(pgate_l[5:4]), .wl_l(wl_l[5:4]),
     .reset_b_l(reset_l[5:4]), .r_gnd_l(r_vdd[5:4]),
     .r_gnd_r(r_vdd_r[5:4]), .pgate_r(pgate_r[5:4]), .wl_r(wl_r[5:4]),
     .reset_b_r(reset_r[5:4]), .q(net032[664:671]),
     .q_b(net036[664:671]), .bl(bl[3:0]));
cram2x2x2 xcram_1_ ( .pgate_l(pgate_l[3:2]), .wl_l(wl_l[3:2]),
     .reset_b_l(reset_l[3:2]), .r_gnd_l(r_vdd[3:2]),
     .r_gnd_r(r_vdd_r[3:2]), .pgate_r(pgate_r[3:2]), .wl_r(wl_r[3:2]),
     .reset_b_r(reset_r[3:2]), .q(net032[672:679]),
     .q_b(net036[672:679]), .bl(bl[3:0]));
cram2x2x2 xcram_0_ ( .pgate_l(pgate_l[1:0]), .wl_l(wl_l[1:0]),
     .reset_b_l(reset_l[1:0]), .r_gnd_l(r_vdd[1:0]),
     .r_gnd_r(r_vdd_r[1:0]), .pgate_r(pgate_r[1:0]), .wl_r(wl_r[1:0]),
     .reset_b_r(reset_r[1:0]), .q(net032[680:687]),
     .q_b(net036[680:687]), .bl(bl[3:0]));
cram2x2x2 I299 ( .pgate_l(pgate_l[173:172]), .wl_l(wl_l[173:172]),
     .reset_b_l(reset_l[173:172]), .r_gnd_l(r_vdd[173:172]),
     .r_gnd_r(r_vdd_r[173:172]), .pgate_r(pgate_r[173:172]),
     .wl_r(wl_r[173:172]), .reset_b_r(reset_r[173:172]),
     .q(net073[0:7]), .q_b(net61[0:7]), .bl(bl[3:0]));
pch_hvt  M0_173_ ( .D(r_vdd_r[173]), .B(vdd_), .G(vdd_cntl_r[173]),
     .S(vdd_));
pch_hvt  M0_172_ ( .D(r_vdd_r[172]), .B(vdd_), .G(vdd_cntl_r[172]),
     .S(vdd_));
pch_hvt  M0_171_ ( .D(r_vdd_r[171]), .B(vdd_), .G(vdd_cntl_r[171]),
     .S(vdd_));
pch_hvt  M0_170_ ( .D(r_vdd_r[170]), .B(vdd_), .G(vdd_cntl_r[170]),
     .S(vdd_));
pch_hvt  M0_169_ ( .D(r_vdd_r[169]), .B(vdd_), .G(vdd_cntl_r[169]),
     .S(vdd_));
pch_hvt  M0_168_ ( .D(r_vdd_r[168]), .B(vdd_), .G(vdd_cntl_r[168]),
     .S(vdd_));
pch_hvt  M0_167_ ( .D(r_vdd_r[167]), .B(vdd_), .G(vdd_cntl_r[167]),
     .S(vdd_));
pch_hvt  M0_166_ ( .D(r_vdd_r[166]), .B(vdd_), .G(vdd_cntl_r[166]),
     .S(vdd_));
pch_hvt  M0_165_ ( .D(r_vdd_r[165]), .B(vdd_), .G(vdd_cntl_r[165]),
     .S(vdd_));
pch_hvt  M0_164_ ( .D(r_vdd_r[164]), .B(vdd_), .G(vdd_cntl_r[164]),
     .S(vdd_));
pch_hvt  M0_163_ ( .D(r_vdd_r[163]), .B(vdd_), .G(vdd_cntl_r[163]),
     .S(vdd_));
pch_hvt  M0_162_ ( .D(r_vdd_r[162]), .B(vdd_), .G(vdd_cntl_r[162]),
     .S(vdd_));
pch_hvt  M0_161_ ( .D(r_vdd_r[161]), .B(vdd_), .G(vdd_cntl_r[161]),
     .S(vdd_));
pch_hvt  M0_160_ ( .D(r_vdd_r[160]), .B(vdd_), .G(vdd_cntl_r[160]),
     .S(vdd_));
pch_hvt  M0_159_ ( .D(r_vdd_r[159]), .B(vdd_), .G(vdd_cntl_r[159]),
     .S(vdd_));
pch_hvt  M0_158_ ( .D(r_vdd_r[158]), .B(vdd_), .G(vdd_cntl_r[158]),
     .S(vdd_));
pch_hvt  M0_157_ ( .D(r_vdd_r[157]), .B(vdd_), .G(vdd_cntl_r[157]),
     .S(vdd_));
pch_hvt  M0_156_ ( .D(r_vdd_r[156]), .B(vdd_), .G(vdd_cntl_r[156]),
     .S(vdd_));
pch_hvt  M0_155_ ( .D(r_vdd_r[155]), .B(vdd_), .G(vdd_cntl_r[155]),
     .S(vdd_));
pch_hvt  M0_154_ ( .D(r_vdd_r[154]), .B(vdd_), .G(vdd_cntl_r[154]),
     .S(vdd_));
pch_hvt  M0_153_ ( .D(r_vdd_r[153]), .B(vdd_), .G(vdd_cntl_r[153]),
     .S(vdd_));
pch_hvt  M0_152_ ( .D(r_vdd_r[152]), .B(vdd_), .G(vdd_cntl_r[152]),
     .S(vdd_));
pch_hvt  M0_151_ ( .D(r_vdd_r[151]), .B(vdd_), .G(vdd_cntl_r[151]),
     .S(vdd_));
pch_hvt  M0_150_ ( .D(r_vdd_r[150]), .B(vdd_), .G(vdd_cntl_r[150]),
     .S(vdd_));
pch_hvt  M0_149_ ( .D(r_vdd_r[149]), .B(vdd_), .G(vdd_cntl_r[149]),
     .S(vdd_));
pch_hvt  M0_148_ ( .D(r_vdd_r[148]), .B(vdd_), .G(vdd_cntl_r[148]),
     .S(vdd_));
pch_hvt  M0_147_ ( .D(r_vdd_r[147]), .B(vdd_), .G(vdd_cntl_r[147]),
     .S(vdd_));
pch_hvt  M0_146_ ( .D(r_vdd_r[146]), .B(vdd_), .G(vdd_cntl_r[146]),
     .S(vdd_));
pch_hvt  M0_145_ ( .D(r_vdd_r[145]), .B(vdd_), .G(vdd_cntl_r[145]),
     .S(vdd_));
pch_hvt  M0_144_ ( .D(r_vdd_r[144]), .B(vdd_), .G(vdd_cntl_r[144]),
     .S(vdd_));
pch_hvt  M0_143_ ( .D(r_vdd_r[143]), .B(vdd_), .G(vdd_cntl_r[143]),
     .S(vdd_));
pch_hvt  M0_142_ ( .D(r_vdd_r[142]), .B(vdd_), .G(vdd_cntl_r[142]),
     .S(vdd_));
pch_hvt  M0_141_ ( .D(r_vdd_r[141]), .B(vdd_), .G(vdd_cntl_r[141]),
     .S(vdd_));
pch_hvt  M0_140_ ( .D(r_vdd_r[140]), .B(vdd_), .G(vdd_cntl_r[140]),
     .S(vdd_));
pch_hvt  M0_139_ ( .D(r_vdd_r[139]), .B(vdd_), .G(vdd_cntl_r[139]),
     .S(vdd_));
pch_hvt  M0_138_ ( .D(r_vdd_r[138]), .B(vdd_), .G(vdd_cntl_r[138]),
     .S(vdd_));
pch_hvt  M0_137_ ( .D(r_vdd_r[137]), .B(vdd_), .G(vdd_cntl_r[137]),
     .S(vdd_));
pch_hvt  M0_136_ ( .D(r_vdd_r[136]), .B(vdd_), .G(vdd_cntl_r[136]),
     .S(vdd_));
pch_hvt  M0_135_ ( .D(r_vdd_r[135]), .B(vdd_), .G(vdd_cntl_r[135]),
     .S(vdd_));
pch_hvt  M0_134_ ( .D(r_vdd_r[134]), .B(vdd_), .G(vdd_cntl_r[134]),
     .S(vdd_));
pch_hvt  M0_133_ ( .D(r_vdd_r[133]), .B(vdd_), .G(vdd_cntl_r[133]),
     .S(vdd_));
pch_hvt  M0_132_ ( .D(r_vdd_r[132]), .B(vdd_), .G(vdd_cntl_r[132]),
     .S(vdd_));
pch_hvt  M0_131_ ( .D(r_vdd_r[131]), .B(vdd_), .G(vdd_cntl_r[131]),
     .S(vdd_));
pch_hvt  M0_130_ ( .D(r_vdd_r[130]), .B(vdd_), .G(vdd_cntl_r[130]),
     .S(vdd_));
pch_hvt  M0_129_ ( .D(r_vdd_r[129]), .B(vdd_), .G(vdd_cntl_r[129]),
     .S(vdd_));
pch_hvt  M0_128_ ( .D(r_vdd_r[128]), .B(vdd_), .G(vdd_cntl_r[128]),
     .S(vdd_));
pch_hvt  M0_127_ ( .D(r_vdd_r[127]), .B(vdd_), .G(vdd_cntl_r[127]),
     .S(vdd_));
pch_hvt  M0_126_ ( .D(r_vdd_r[126]), .B(vdd_), .G(vdd_cntl_r[126]),
     .S(vdd_));
pch_hvt  M0_125_ ( .D(r_vdd_r[125]), .B(vdd_), .G(vdd_cntl_r[125]),
     .S(vdd_));
pch_hvt  M0_124_ ( .D(r_vdd_r[124]), .B(vdd_), .G(vdd_cntl_r[124]),
     .S(vdd_));
pch_hvt  M0_123_ ( .D(r_vdd_r[123]), .B(vdd_), .G(vdd_cntl_r[123]),
     .S(vdd_));
pch_hvt  M0_122_ ( .D(r_vdd_r[122]), .B(vdd_), .G(vdd_cntl_r[122]),
     .S(vdd_));
pch_hvt  M0_121_ ( .D(r_vdd_r[121]), .B(vdd_), .G(vdd_cntl_r[121]),
     .S(vdd_));
pch_hvt  M0_120_ ( .D(r_vdd_r[120]), .B(vdd_), .G(vdd_cntl_r[120]),
     .S(vdd_));
pch_hvt  M0_119_ ( .D(r_vdd_r[119]), .B(vdd_), .G(vdd_cntl_r[119]),
     .S(vdd_));
pch_hvt  M0_118_ ( .D(r_vdd_r[118]), .B(vdd_), .G(vdd_cntl_r[118]),
     .S(vdd_));
pch_hvt  M0_117_ ( .D(r_vdd_r[117]), .B(vdd_), .G(vdd_cntl_r[117]),
     .S(vdd_));
pch_hvt  M0_116_ ( .D(r_vdd_r[116]), .B(vdd_), .G(vdd_cntl_r[116]),
     .S(vdd_));
pch_hvt  M0_115_ ( .D(r_vdd_r[115]), .B(vdd_), .G(vdd_cntl_r[115]),
     .S(vdd_));
pch_hvt  M0_114_ ( .D(r_vdd_r[114]), .B(vdd_), .G(vdd_cntl_r[114]),
     .S(vdd_));
pch_hvt  M0_113_ ( .D(r_vdd_r[113]), .B(vdd_), .G(vdd_cntl_r[113]),
     .S(vdd_));
pch_hvt  M0_112_ ( .D(r_vdd_r[112]), .B(vdd_), .G(vdd_cntl_r[112]),
     .S(vdd_));
pch_hvt  M0_111_ ( .D(r_vdd_r[111]), .B(vdd_), .G(vdd_cntl_r[111]),
     .S(vdd_));
pch_hvt  M0_110_ ( .D(r_vdd_r[110]), .B(vdd_), .G(vdd_cntl_r[110]),
     .S(vdd_));
pch_hvt  M0_109_ ( .D(r_vdd_r[109]), .B(vdd_), .G(vdd_cntl_r[109]),
     .S(vdd_));
pch_hvt  M0_108_ ( .D(r_vdd_r[108]), .B(vdd_), .G(vdd_cntl_r[108]),
     .S(vdd_));
pch_hvt  M0_107_ ( .D(r_vdd_r[107]), .B(vdd_), .G(vdd_cntl_r[107]),
     .S(vdd_));
pch_hvt  M0_106_ ( .D(r_vdd_r[106]), .B(vdd_), .G(vdd_cntl_r[106]),
     .S(vdd_));
pch_hvt  M0_105_ ( .D(r_vdd_r[105]), .B(vdd_), .G(vdd_cntl_r[105]),
     .S(vdd_));
pch_hvt  M0_104_ ( .D(r_vdd_r[104]), .B(vdd_), .G(vdd_cntl_r[104]),
     .S(vdd_));
pch_hvt  M0_103_ ( .D(r_vdd_r[103]), .B(vdd_), .G(vdd_cntl_r[103]),
     .S(vdd_));
pch_hvt  M0_102_ ( .D(r_vdd_r[102]), .B(vdd_), .G(vdd_cntl_r[102]),
     .S(vdd_));
pch_hvt  M0_101_ ( .D(r_vdd_r[101]), .B(vdd_), .G(vdd_cntl_r[101]),
     .S(vdd_));
pch_hvt  M0_100_ ( .D(r_vdd_r[100]), .B(vdd_), .G(vdd_cntl_r[100]),
     .S(vdd_));
pch_hvt  M0_99_ ( .D(r_vdd_r[99]), .B(vdd_), .G(vdd_cntl_r[99]),
     .S(vdd_));
pch_hvt  M0_98_ ( .D(r_vdd_r[98]), .B(vdd_), .G(vdd_cntl_r[98]),
     .S(vdd_));
pch_hvt  M0_97_ ( .D(r_vdd_r[97]), .B(vdd_), .G(vdd_cntl_r[97]),
     .S(vdd_));
pch_hvt  M0_96_ ( .D(r_vdd_r[96]), .B(vdd_), .G(vdd_cntl_r[96]),
     .S(vdd_));
pch_hvt  M0_95_ ( .D(r_vdd_r[95]), .B(vdd_), .G(vdd_cntl_r[95]),
     .S(vdd_));
pch_hvt  M0_94_ ( .D(r_vdd_r[94]), .B(vdd_), .G(vdd_cntl_r[94]),
     .S(vdd_));
pch_hvt  M0_93_ ( .D(r_vdd_r[93]), .B(vdd_), .G(vdd_cntl_r[93]),
     .S(vdd_));
pch_hvt  M0_92_ ( .D(r_vdd_r[92]), .B(vdd_), .G(vdd_cntl_r[92]),
     .S(vdd_));
pch_hvt  M0_91_ ( .D(r_vdd_r[91]), .B(vdd_), .G(vdd_cntl_r[91]),
     .S(vdd_));
pch_hvt  M0_90_ ( .D(r_vdd_r[90]), .B(vdd_), .G(vdd_cntl_r[90]),
     .S(vdd_));
pch_hvt  M0_89_ ( .D(r_vdd_r[89]), .B(vdd_), .G(vdd_cntl_r[89]),
     .S(vdd_));
pch_hvt  M0_88_ ( .D(r_vdd_r[88]), .B(vdd_), .G(vdd_cntl_r[88]),
     .S(vdd_));
pch_hvt  M0_87_ ( .D(r_vdd_r[87]), .B(vdd_), .G(vdd_cntl_r[87]),
     .S(vdd_));
pch_hvt  M0_86_ ( .D(r_vdd_r[86]), .B(vdd_), .G(vdd_cntl_r[86]),
     .S(vdd_));
pch_hvt  M0_85_ ( .D(r_vdd_r[85]), .B(vdd_), .G(vdd_cntl_r[85]),
     .S(vdd_));
pch_hvt  M0_84_ ( .D(r_vdd_r[84]), .B(vdd_), .G(vdd_cntl_r[84]),
     .S(vdd_));
pch_hvt  M0_83_ ( .D(r_vdd_r[83]), .B(vdd_), .G(vdd_cntl_r[83]),
     .S(vdd_));
pch_hvt  M0_82_ ( .D(r_vdd_r[82]), .B(vdd_), .G(vdd_cntl_r[82]),
     .S(vdd_));
pch_hvt  M0_81_ ( .D(r_vdd_r[81]), .B(vdd_), .G(vdd_cntl_r[81]),
     .S(vdd_));
pch_hvt  M0_80_ ( .D(r_vdd_r[80]), .B(vdd_), .G(vdd_cntl_r[80]),
     .S(vdd_));
pch_hvt  M0_79_ ( .D(r_vdd_r[79]), .B(vdd_), .G(vdd_cntl_r[79]),
     .S(vdd_));
pch_hvt  M0_78_ ( .D(r_vdd_r[78]), .B(vdd_), .G(vdd_cntl_r[78]),
     .S(vdd_));
pch_hvt  M0_77_ ( .D(r_vdd_r[77]), .B(vdd_), .G(vdd_cntl_r[77]),
     .S(vdd_));
pch_hvt  M0_76_ ( .D(r_vdd_r[76]), .B(vdd_), .G(vdd_cntl_r[76]),
     .S(vdd_));
pch_hvt  M0_75_ ( .D(r_vdd_r[75]), .B(vdd_), .G(vdd_cntl_r[75]),
     .S(vdd_));
pch_hvt  M0_74_ ( .D(r_vdd_r[74]), .B(vdd_), .G(vdd_cntl_r[74]),
     .S(vdd_));
pch_hvt  M0_73_ ( .D(r_vdd_r[73]), .B(vdd_), .G(vdd_cntl_r[73]),
     .S(vdd_));
pch_hvt  M0_72_ ( .D(r_vdd_r[72]), .B(vdd_), .G(vdd_cntl_r[72]),
     .S(vdd_));
pch_hvt  M0_71_ ( .D(r_vdd_r[71]), .B(vdd_), .G(vdd_cntl_r[71]),
     .S(vdd_));
pch_hvt  M0_70_ ( .D(r_vdd_r[70]), .B(vdd_), .G(vdd_cntl_r[70]),
     .S(vdd_));
pch_hvt  M0_69_ ( .D(r_vdd_r[69]), .B(vdd_), .G(vdd_cntl_r[69]),
     .S(vdd_));
pch_hvt  M0_68_ ( .D(r_vdd_r[68]), .B(vdd_), .G(vdd_cntl_r[68]),
     .S(vdd_));
pch_hvt  M0_67_ ( .D(r_vdd_r[67]), .B(vdd_), .G(vdd_cntl_r[67]),
     .S(vdd_));
pch_hvt  M0_66_ ( .D(r_vdd_r[66]), .B(vdd_), .G(vdd_cntl_r[66]),
     .S(vdd_));
pch_hvt  M0_65_ ( .D(r_vdd_r[65]), .B(vdd_), .G(vdd_cntl_r[65]),
     .S(vdd_));
pch_hvt  M0_64_ ( .D(r_vdd_r[64]), .B(vdd_), .G(vdd_cntl_r[64]),
     .S(vdd_));
pch_hvt  M0_63_ ( .D(r_vdd_r[63]), .B(vdd_), .G(vdd_cntl_r[63]),
     .S(vdd_));
pch_hvt  M0_62_ ( .D(r_vdd_r[62]), .B(vdd_), .G(vdd_cntl_r[62]),
     .S(vdd_));
pch_hvt  M0_61_ ( .D(r_vdd_r[61]), .B(vdd_), .G(vdd_cntl_r[61]),
     .S(vdd_));
pch_hvt  M0_60_ ( .D(r_vdd_r[60]), .B(vdd_), .G(vdd_cntl_r[60]),
     .S(vdd_));
pch_hvt  M0_59_ ( .D(r_vdd_r[59]), .B(vdd_), .G(vdd_cntl_r[59]),
     .S(vdd_));
pch_hvt  M0_58_ ( .D(r_vdd_r[58]), .B(vdd_), .G(vdd_cntl_r[58]),
     .S(vdd_));
pch_hvt  M0_57_ ( .D(r_vdd_r[57]), .B(vdd_), .G(vdd_cntl_r[57]),
     .S(vdd_));
pch_hvt  M0_56_ ( .D(r_vdd_r[56]), .B(vdd_), .G(vdd_cntl_r[56]),
     .S(vdd_));
pch_hvt  M0_55_ ( .D(r_vdd_r[55]), .B(vdd_), .G(vdd_cntl_r[55]),
     .S(vdd_));
pch_hvt  M0_54_ ( .D(r_vdd_r[54]), .B(vdd_), .G(vdd_cntl_r[54]),
     .S(vdd_));
pch_hvt  M0_53_ ( .D(r_vdd_r[53]), .B(vdd_), .G(vdd_cntl_r[53]),
     .S(vdd_));
pch_hvt  M0_52_ ( .D(r_vdd_r[52]), .B(vdd_), .G(vdd_cntl_r[52]),
     .S(vdd_));
pch_hvt  M0_51_ ( .D(r_vdd_r[51]), .B(vdd_), .G(vdd_cntl_r[51]),
     .S(vdd_));
pch_hvt  M0_50_ ( .D(r_vdd_r[50]), .B(vdd_), .G(vdd_cntl_r[50]),
     .S(vdd_));
pch_hvt  M0_49_ ( .D(r_vdd_r[49]), .B(vdd_), .G(vdd_cntl_r[49]),
     .S(vdd_));
pch_hvt  M0_48_ ( .D(r_vdd_r[48]), .B(vdd_), .G(vdd_cntl_r[48]),
     .S(vdd_));
pch_hvt  M0_47_ ( .D(r_vdd_r[47]), .B(vdd_), .G(vdd_cntl_r[47]),
     .S(vdd_));
pch_hvt  M0_46_ ( .D(r_vdd_r[46]), .B(vdd_), .G(vdd_cntl_r[46]),
     .S(vdd_));
pch_hvt  M0_45_ ( .D(r_vdd_r[45]), .B(vdd_), .G(vdd_cntl_r[45]),
     .S(vdd_));
pch_hvt  M0_44_ ( .D(r_vdd_r[44]), .B(vdd_), .G(vdd_cntl_r[44]),
     .S(vdd_));
pch_hvt  M0_43_ ( .D(r_vdd_r[43]), .B(vdd_), .G(vdd_cntl_r[43]),
     .S(vdd_));
pch_hvt  M0_42_ ( .D(r_vdd_r[42]), .B(vdd_), .G(vdd_cntl_r[42]),
     .S(vdd_));
pch_hvt  M0_41_ ( .D(r_vdd_r[41]), .B(vdd_), .G(vdd_cntl_r[41]),
     .S(vdd_));
pch_hvt  M0_40_ ( .D(r_vdd_r[40]), .B(vdd_), .G(vdd_cntl_r[40]),
     .S(vdd_));
pch_hvt  M0_39_ ( .D(r_vdd_r[39]), .B(vdd_), .G(vdd_cntl_r[39]),
     .S(vdd_));
pch_hvt  M0_38_ ( .D(r_vdd_r[38]), .B(vdd_), .G(vdd_cntl_r[38]),
     .S(vdd_));
pch_hvt  M0_37_ ( .D(r_vdd_r[37]), .B(vdd_), .G(vdd_cntl_r[37]),
     .S(vdd_));
pch_hvt  M0_36_ ( .D(r_vdd_r[36]), .B(vdd_), .G(vdd_cntl_r[36]),
     .S(vdd_));
pch_hvt  M0_35_ ( .D(r_vdd_r[35]), .B(vdd_), .G(vdd_cntl_r[35]),
     .S(vdd_));
pch_hvt  M0_34_ ( .D(r_vdd_r[34]), .B(vdd_), .G(vdd_cntl_r[34]),
     .S(vdd_));
pch_hvt  M0_33_ ( .D(r_vdd_r[33]), .B(vdd_), .G(vdd_cntl_r[33]),
     .S(vdd_));
pch_hvt  M0_32_ ( .D(r_vdd_r[32]), .B(vdd_), .G(vdd_cntl_r[32]),
     .S(vdd_));
pch_hvt  M0_31_ ( .D(r_vdd_r[31]), .B(vdd_), .G(vdd_cntl_r[31]),
     .S(vdd_));
pch_hvt  M0_30_ ( .D(r_vdd_r[30]), .B(vdd_), .G(vdd_cntl_r[30]),
     .S(vdd_));
pch_hvt  M0_29_ ( .D(r_vdd_r[29]), .B(vdd_), .G(vdd_cntl_r[29]),
     .S(vdd_));
pch_hvt  M0_28_ ( .D(r_vdd_r[28]), .B(vdd_), .G(vdd_cntl_r[28]),
     .S(vdd_));
pch_hvt  M0_27_ ( .D(r_vdd_r[27]), .B(vdd_), .G(vdd_cntl_r[27]),
     .S(vdd_));
pch_hvt  M0_26_ ( .D(r_vdd_r[26]), .B(vdd_), .G(vdd_cntl_r[26]),
     .S(vdd_));
pch_hvt  M0_25_ ( .D(r_vdd_r[25]), .B(vdd_), .G(vdd_cntl_r[25]),
     .S(vdd_));
pch_hvt  M0_24_ ( .D(r_vdd_r[24]), .B(vdd_), .G(vdd_cntl_r[24]),
     .S(vdd_));
pch_hvt  M0_23_ ( .D(r_vdd_r[23]), .B(vdd_), .G(vdd_cntl_r[23]),
     .S(vdd_));
pch_hvt  M0_22_ ( .D(r_vdd_r[22]), .B(vdd_), .G(vdd_cntl_r[22]),
     .S(vdd_));
pch_hvt  M0_21_ ( .D(r_vdd_r[21]), .B(vdd_), .G(vdd_cntl_r[21]),
     .S(vdd_));
pch_hvt  M0_20_ ( .D(r_vdd_r[20]), .B(vdd_), .G(vdd_cntl_r[20]),
     .S(vdd_));
pch_hvt  M0_19_ ( .D(r_vdd_r[19]), .B(vdd_), .G(vdd_cntl_r[19]),
     .S(vdd_));
pch_hvt  M0_18_ ( .D(r_vdd_r[18]), .B(vdd_), .G(vdd_cntl_r[18]),
     .S(vdd_));
pch_hvt  M0_17_ ( .D(r_vdd_r[17]), .B(vdd_), .G(vdd_cntl_r[17]),
     .S(vdd_));
pch_hvt  M0_16_ ( .D(r_vdd_r[16]), .B(vdd_), .G(vdd_cntl_r[16]),
     .S(vdd_));
pch_hvt  M0_15_ ( .D(r_vdd_r[15]), .B(vdd_), .G(vdd_cntl_r[15]),
     .S(vdd_));
pch_hvt  M0_14_ ( .D(r_vdd_r[14]), .B(vdd_), .G(vdd_cntl_r[14]),
     .S(vdd_));
pch_hvt  M0_13_ ( .D(r_vdd_r[13]), .B(vdd_), .G(vdd_cntl_r[13]),
     .S(vdd_));
pch_hvt  M0_12_ ( .D(r_vdd_r[12]), .B(vdd_), .G(vdd_cntl_r[12]),
     .S(vdd_));
pch_hvt  M0_11_ ( .D(r_vdd_r[11]), .B(vdd_), .G(vdd_cntl_r[11]),
     .S(vdd_));
pch_hvt  M0_10_ ( .D(r_vdd_r[10]), .B(vdd_), .G(vdd_cntl_r[10]),
     .S(vdd_));
pch_hvt  M0_9_ ( .D(r_vdd_r[9]), .B(vdd_), .G(vdd_cntl_r[9]),
     .S(vdd_));
pch_hvt  M0_8_ ( .D(r_vdd_r[8]), .B(vdd_), .G(vdd_cntl_r[8]),
     .S(vdd_));
pch_hvt  M0_7_ ( .D(r_vdd_r[7]), .B(vdd_), .G(vdd_cntl_r[7]),
     .S(vdd_));
pch_hvt  M0_6_ ( .D(r_vdd_r[6]), .B(vdd_), .G(vdd_cntl_r[6]),
     .S(vdd_));
pch_hvt  M0_5_ ( .D(r_vdd_r[5]), .B(vdd_), .G(vdd_cntl_r[5]),
     .S(vdd_));
pch_hvt  M0_4_ ( .D(r_vdd_r[4]), .B(vdd_), .G(vdd_cntl_r[4]),
     .S(vdd_));
pch_hvt  M0_3_ ( .D(r_vdd_r[3]), .B(vdd_), .G(vdd_cntl_r[3]),
     .S(vdd_));
pch_hvt  M0_2_ ( .D(r_vdd_r[2]), .B(vdd_), .G(vdd_cntl_r[2]),
     .S(vdd_));
pch_hvt  M0_1_ ( .D(r_vdd_r[1]), .B(vdd_), .G(vdd_cntl_r[1]),
     .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd_r[0]), .B(vdd_), .G(vdd_cntl_r[0]),
     .S(vdd_));
pch_hvt  vdd_cntrl_173_ ( .D(r_vdd[173]), .B(vdd_),
     .G(vdd_cntl_l[173]), .S(vdd_));
pch_hvt  vdd_cntrl_172_ ( .D(r_vdd[172]), .B(vdd_),
     .G(vdd_cntl_l[172]), .S(vdd_));
pch_hvt  vdd_cntrl_171_ ( .D(r_vdd[171]), .B(vdd_),
     .G(vdd_cntl_l[171]), .S(vdd_));
pch_hvt  vdd_cntrl_170_ ( .D(r_vdd[170]), .B(vdd_),
     .G(vdd_cntl_l[170]), .S(vdd_));
pch_hvt  vdd_cntrl_169_ ( .D(r_vdd[169]), .B(vdd_),
     .G(vdd_cntl_l[169]), .S(vdd_));
pch_hvt  vdd_cntrl_168_ ( .D(r_vdd[168]), .B(vdd_),
     .G(vdd_cntl_l[168]), .S(vdd_));
pch_hvt  vdd_cntrl_167_ ( .D(r_vdd[167]), .B(vdd_),
     .G(vdd_cntl_l[167]), .S(vdd_));
pch_hvt  vdd_cntrl_166_ ( .D(r_vdd[166]), .B(vdd_),
     .G(vdd_cntl_l[166]), .S(vdd_));
pch_hvt  vdd_cntrl_165_ ( .D(r_vdd[165]), .B(vdd_),
     .G(vdd_cntl_l[165]), .S(vdd_));
pch_hvt  vdd_cntrl_164_ ( .D(r_vdd[164]), .B(vdd_),
     .G(vdd_cntl_l[164]), .S(vdd_));
pch_hvt  vdd_cntrl_163_ ( .D(r_vdd[163]), .B(vdd_),
     .G(vdd_cntl_l[163]), .S(vdd_));
pch_hvt  vdd_cntrl_162_ ( .D(r_vdd[162]), .B(vdd_),
     .G(vdd_cntl_l[162]), .S(vdd_));
pch_hvt  vdd_cntrl_161_ ( .D(r_vdd[161]), .B(vdd_),
     .G(vdd_cntl_l[161]), .S(vdd_));
pch_hvt  vdd_cntrl_160_ ( .D(r_vdd[160]), .B(vdd_),
     .G(vdd_cntl_l[160]), .S(vdd_));
pch_hvt  vdd_cntrl_159_ ( .D(r_vdd[159]), .B(vdd_),
     .G(vdd_cntl_l[159]), .S(vdd_));
pch_hvt  vdd_cntrl_158_ ( .D(r_vdd[158]), .B(vdd_),
     .G(vdd_cntl_l[158]), .S(vdd_));
pch_hvt  vdd_cntrl_157_ ( .D(r_vdd[157]), .B(vdd_),
     .G(vdd_cntl_l[157]), .S(vdd_));
pch_hvt  vdd_cntrl_156_ ( .D(r_vdd[156]), .B(vdd_),
     .G(vdd_cntl_l[156]), .S(vdd_));
pch_hvt  vdd_cntrl_155_ ( .D(r_vdd[155]), .B(vdd_),
     .G(vdd_cntl_l[155]), .S(vdd_));
pch_hvt  vdd_cntrl_154_ ( .D(r_vdd[154]), .B(vdd_),
     .G(vdd_cntl_l[154]), .S(vdd_));
pch_hvt  vdd_cntrl_153_ ( .D(r_vdd[153]), .B(vdd_),
     .G(vdd_cntl_l[153]), .S(vdd_));
pch_hvt  vdd_cntrl_152_ ( .D(r_vdd[152]), .B(vdd_),
     .G(vdd_cntl_l[152]), .S(vdd_));
pch_hvt  vdd_cntrl_151_ ( .D(r_vdd[151]), .B(vdd_),
     .G(vdd_cntl_l[151]), .S(vdd_));
pch_hvt  vdd_cntrl_150_ ( .D(r_vdd[150]), .B(vdd_),
     .G(vdd_cntl_l[150]), .S(vdd_));
pch_hvt  vdd_cntrl_149_ ( .D(r_vdd[149]), .B(vdd_),
     .G(vdd_cntl_l[149]), .S(vdd_));
pch_hvt  vdd_cntrl_148_ ( .D(r_vdd[148]), .B(vdd_),
     .G(vdd_cntl_l[148]), .S(vdd_));
pch_hvt  vdd_cntrl_147_ ( .D(r_vdd[147]), .B(vdd_),
     .G(vdd_cntl_l[147]), .S(vdd_));
pch_hvt  vdd_cntrl_146_ ( .D(r_vdd[146]), .B(vdd_),
     .G(vdd_cntl_l[146]), .S(vdd_));
pch_hvt  vdd_cntrl_145_ ( .D(r_vdd[145]), .B(vdd_),
     .G(vdd_cntl_l[145]), .S(vdd_));
pch_hvt  vdd_cntrl_144_ ( .D(r_vdd[144]), .B(vdd_),
     .G(vdd_cntl_l[144]), .S(vdd_));
pch_hvt  vdd_cntrl_143_ ( .D(r_vdd[143]), .B(vdd_),
     .G(vdd_cntl_l[143]), .S(vdd_));
pch_hvt  vdd_cntrl_142_ ( .D(r_vdd[142]), .B(vdd_),
     .G(vdd_cntl_l[142]), .S(vdd_));
pch_hvt  vdd_cntrl_141_ ( .D(r_vdd[141]), .B(vdd_),
     .G(vdd_cntl_l[141]), .S(vdd_));
pch_hvt  vdd_cntrl_140_ ( .D(r_vdd[140]), .B(vdd_),
     .G(vdd_cntl_l[140]), .S(vdd_));
pch_hvt  vdd_cntrl_139_ ( .D(r_vdd[139]), .B(vdd_),
     .G(vdd_cntl_l[139]), .S(vdd_));
pch_hvt  vdd_cntrl_138_ ( .D(r_vdd[138]), .B(vdd_),
     .G(vdd_cntl_l[138]), .S(vdd_));
pch_hvt  vdd_cntrl_137_ ( .D(r_vdd[137]), .B(vdd_),
     .G(vdd_cntl_l[137]), .S(vdd_));
pch_hvt  vdd_cntrl_136_ ( .D(r_vdd[136]), .B(vdd_),
     .G(vdd_cntl_l[136]), .S(vdd_));
pch_hvt  vdd_cntrl_135_ ( .D(r_vdd[135]), .B(vdd_),
     .G(vdd_cntl_l[135]), .S(vdd_));
pch_hvt  vdd_cntrl_134_ ( .D(r_vdd[134]), .B(vdd_),
     .G(vdd_cntl_l[134]), .S(vdd_));
pch_hvt  vdd_cntrl_133_ ( .D(r_vdd[133]), .B(vdd_),
     .G(vdd_cntl_l[133]), .S(vdd_));
pch_hvt  vdd_cntrl_132_ ( .D(r_vdd[132]), .B(vdd_),
     .G(vdd_cntl_l[132]), .S(vdd_));
pch_hvt  vdd_cntrl_131_ ( .D(r_vdd[131]), .B(vdd_),
     .G(vdd_cntl_l[131]), .S(vdd_));
pch_hvt  vdd_cntrl_130_ ( .D(r_vdd[130]), .B(vdd_),
     .G(vdd_cntl_l[130]), .S(vdd_));
pch_hvt  vdd_cntrl_129_ ( .D(r_vdd[129]), .B(vdd_),
     .G(vdd_cntl_l[129]), .S(vdd_));
pch_hvt  vdd_cntrl_128_ ( .D(r_vdd[128]), .B(vdd_),
     .G(vdd_cntl_l[128]), .S(vdd_));
pch_hvt  vdd_cntrl_127_ ( .D(r_vdd[127]), .B(vdd_),
     .G(vdd_cntl_l[127]), .S(vdd_));
pch_hvt  vdd_cntrl_126_ ( .D(r_vdd[126]), .B(vdd_),
     .G(vdd_cntl_l[126]), .S(vdd_));
pch_hvt  vdd_cntrl_125_ ( .D(r_vdd[125]), .B(vdd_),
     .G(vdd_cntl_l[125]), .S(vdd_));
pch_hvt  vdd_cntrl_124_ ( .D(r_vdd[124]), .B(vdd_),
     .G(vdd_cntl_l[124]), .S(vdd_));
pch_hvt  vdd_cntrl_123_ ( .D(r_vdd[123]), .B(vdd_),
     .G(vdd_cntl_l[123]), .S(vdd_));
pch_hvt  vdd_cntrl_122_ ( .D(r_vdd[122]), .B(vdd_),
     .G(vdd_cntl_l[122]), .S(vdd_));
pch_hvt  vdd_cntrl_121_ ( .D(r_vdd[121]), .B(vdd_),
     .G(vdd_cntl_l[121]), .S(vdd_));
pch_hvt  vdd_cntrl_120_ ( .D(r_vdd[120]), .B(vdd_),
     .G(vdd_cntl_l[120]), .S(vdd_));
pch_hvt  vdd_cntrl_119_ ( .D(r_vdd[119]), .B(vdd_),
     .G(vdd_cntl_l[119]), .S(vdd_));
pch_hvt  vdd_cntrl_118_ ( .D(r_vdd[118]), .B(vdd_),
     .G(vdd_cntl_l[118]), .S(vdd_));
pch_hvt  vdd_cntrl_117_ ( .D(r_vdd[117]), .B(vdd_),
     .G(vdd_cntl_l[117]), .S(vdd_));
pch_hvt  vdd_cntrl_116_ ( .D(r_vdd[116]), .B(vdd_),
     .G(vdd_cntl_l[116]), .S(vdd_));
pch_hvt  vdd_cntrl_115_ ( .D(r_vdd[115]), .B(vdd_),
     .G(vdd_cntl_l[115]), .S(vdd_));
pch_hvt  vdd_cntrl_114_ ( .D(r_vdd[114]), .B(vdd_),
     .G(vdd_cntl_l[114]), .S(vdd_));
pch_hvt  vdd_cntrl_113_ ( .D(r_vdd[113]), .B(vdd_),
     .G(vdd_cntl_l[113]), .S(vdd_));
pch_hvt  vdd_cntrl_112_ ( .D(r_vdd[112]), .B(vdd_),
     .G(vdd_cntl_l[112]), .S(vdd_));
pch_hvt  vdd_cntrl_111_ ( .D(r_vdd[111]), .B(vdd_),
     .G(vdd_cntl_l[111]), .S(vdd_));
pch_hvt  vdd_cntrl_110_ ( .D(r_vdd[110]), .B(vdd_),
     .G(vdd_cntl_l[110]), .S(vdd_));
pch_hvt  vdd_cntrl_109_ ( .D(r_vdd[109]), .B(vdd_),
     .G(vdd_cntl_l[109]), .S(vdd_));
pch_hvt  vdd_cntrl_108_ ( .D(r_vdd[108]), .B(vdd_),
     .G(vdd_cntl_l[108]), .S(vdd_));
pch_hvt  vdd_cntrl_107_ ( .D(r_vdd[107]), .B(vdd_),
     .G(vdd_cntl_l[107]), .S(vdd_));
pch_hvt  vdd_cntrl_106_ ( .D(r_vdd[106]), .B(vdd_),
     .G(vdd_cntl_l[106]), .S(vdd_));
pch_hvt  vdd_cntrl_105_ ( .D(r_vdd[105]), .B(vdd_),
     .G(vdd_cntl_l[105]), .S(vdd_));
pch_hvt  vdd_cntrl_104_ ( .D(r_vdd[104]), .B(vdd_),
     .G(vdd_cntl_l[104]), .S(vdd_));
pch_hvt  vdd_cntrl_103_ ( .D(r_vdd[103]), .B(vdd_),
     .G(vdd_cntl_l[103]), .S(vdd_));
pch_hvt  vdd_cntrl_102_ ( .D(r_vdd[102]), .B(vdd_),
     .G(vdd_cntl_l[102]), .S(vdd_));
pch_hvt  vdd_cntrl_101_ ( .D(r_vdd[101]), .B(vdd_),
     .G(vdd_cntl_l[101]), .S(vdd_));
pch_hvt  vdd_cntrl_100_ ( .D(r_vdd[100]), .B(vdd_),
     .G(vdd_cntl_l[100]), .S(vdd_));
pch_hvt  vdd_cntrl_99_ ( .D(r_vdd[99]), .B(vdd_), .G(vdd_cntl_l[99]),
     .S(vdd_));
pch_hvt  vdd_cntrl_98_ ( .D(r_vdd[98]), .B(vdd_), .G(vdd_cntl_l[98]),
     .S(vdd_));
pch_hvt  vdd_cntrl_97_ ( .D(r_vdd[97]), .B(vdd_), .G(vdd_cntl_l[97]),
     .S(vdd_));
pch_hvt  vdd_cntrl_96_ ( .D(r_vdd[96]), .B(vdd_), .G(vdd_cntl_l[96]),
     .S(vdd_));
pch_hvt  vdd_cntrl_95_ ( .D(r_vdd[95]), .B(vdd_), .G(vdd_cntl_l[95]),
     .S(vdd_));
pch_hvt  vdd_cntrl_94_ ( .D(r_vdd[94]), .B(vdd_), .G(vdd_cntl_l[94]),
     .S(vdd_));
pch_hvt  vdd_cntrl_93_ ( .D(r_vdd[93]), .B(vdd_), .G(vdd_cntl_l[93]),
     .S(vdd_));
pch_hvt  vdd_cntrl_92_ ( .D(r_vdd[92]), .B(vdd_), .G(vdd_cntl_l[92]),
     .S(vdd_));
pch_hvt  vdd_cntrl_91_ ( .D(r_vdd[91]), .B(vdd_), .G(vdd_cntl_l[91]),
     .S(vdd_));
pch_hvt  vdd_cntrl_90_ ( .D(r_vdd[90]), .B(vdd_), .G(vdd_cntl_l[90]),
     .S(vdd_));
pch_hvt  vdd_cntrl_89_ ( .D(r_vdd[89]), .B(vdd_), .G(vdd_cntl_l[89]),
     .S(vdd_));
pch_hvt  vdd_cntrl_88_ ( .D(r_vdd[88]), .B(vdd_), .G(vdd_cntl_l[88]),
     .S(vdd_));
pch_hvt  vdd_cntrl_87_ ( .D(r_vdd[87]), .B(vdd_), .G(vdd_cntl_l[87]),
     .S(vdd_));
pch_hvt  vdd_cntrl_86_ ( .D(r_vdd[86]), .B(vdd_), .G(vdd_cntl_l[86]),
     .S(vdd_));
pch_hvt  vdd_cntrl_85_ ( .D(r_vdd[85]), .B(vdd_), .G(vdd_cntl_l[85]),
     .S(vdd_));
pch_hvt  vdd_cntrl_84_ ( .D(r_vdd[84]), .B(vdd_), .G(vdd_cntl_l[84]),
     .S(vdd_));
pch_hvt  vdd_cntrl_83_ ( .D(r_vdd[83]), .B(vdd_), .G(vdd_cntl_l[83]),
     .S(vdd_));
pch_hvt  vdd_cntrl_82_ ( .D(r_vdd[82]), .B(vdd_), .G(vdd_cntl_l[82]),
     .S(vdd_));
pch_hvt  vdd_cntrl_81_ ( .D(r_vdd[81]), .B(vdd_), .G(vdd_cntl_l[81]),
     .S(vdd_));
pch_hvt  vdd_cntrl_80_ ( .D(r_vdd[80]), .B(vdd_), .G(vdd_cntl_l[80]),
     .S(vdd_));
pch_hvt  vdd_cntrl_79_ ( .D(r_vdd[79]), .B(vdd_), .G(vdd_cntl_l[79]),
     .S(vdd_));
pch_hvt  vdd_cntrl_78_ ( .D(r_vdd[78]), .B(vdd_), .G(vdd_cntl_l[78]),
     .S(vdd_));
pch_hvt  vdd_cntrl_77_ ( .D(r_vdd[77]), .B(vdd_), .G(vdd_cntl_l[77]),
     .S(vdd_));
pch_hvt  vdd_cntrl_76_ ( .D(r_vdd[76]), .B(vdd_), .G(vdd_cntl_l[76]),
     .S(vdd_));
pch_hvt  vdd_cntrl_75_ ( .D(r_vdd[75]), .B(vdd_), .G(vdd_cntl_l[75]),
     .S(vdd_));
pch_hvt  vdd_cntrl_74_ ( .D(r_vdd[74]), .B(vdd_), .G(vdd_cntl_l[74]),
     .S(vdd_));
pch_hvt  vdd_cntrl_73_ ( .D(r_vdd[73]), .B(vdd_), .G(vdd_cntl_l[73]),
     .S(vdd_));
pch_hvt  vdd_cntrl_72_ ( .D(r_vdd[72]), .B(vdd_), .G(vdd_cntl_l[72]),
     .S(vdd_));
pch_hvt  vdd_cntrl_71_ ( .D(r_vdd[71]), .B(vdd_), .G(vdd_cntl_l[71]),
     .S(vdd_));
pch_hvt  vdd_cntrl_70_ ( .D(r_vdd[70]), .B(vdd_), .G(vdd_cntl_l[70]),
     .S(vdd_));
pch_hvt  vdd_cntrl_69_ ( .D(r_vdd[69]), .B(vdd_), .G(vdd_cntl_l[69]),
     .S(vdd_));
pch_hvt  vdd_cntrl_68_ ( .D(r_vdd[68]), .B(vdd_), .G(vdd_cntl_l[68]),
     .S(vdd_));
pch_hvt  vdd_cntrl_67_ ( .D(r_vdd[67]), .B(vdd_), .G(vdd_cntl_l[67]),
     .S(vdd_));
pch_hvt  vdd_cntrl_66_ ( .D(r_vdd[66]), .B(vdd_), .G(vdd_cntl_l[66]),
     .S(vdd_));
pch_hvt  vdd_cntrl_65_ ( .D(r_vdd[65]), .B(vdd_), .G(vdd_cntl_l[65]),
     .S(vdd_));
pch_hvt  vdd_cntrl_64_ ( .D(r_vdd[64]), .B(vdd_), .G(vdd_cntl_l[64]),
     .S(vdd_));
pch_hvt  vdd_cntrl_63_ ( .D(r_vdd[63]), .B(vdd_), .G(vdd_cntl_l[63]),
     .S(vdd_));
pch_hvt  vdd_cntrl_62_ ( .D(r_vdd[62]), .B(vdd_), .G(vdd_cntl_l[62]),
     .S(vdd_));
pch_hvt  vdd_cntrl_61_ ( .D(r_vdd[61]), .B(vdd_), .G(vdd_cntl_l[61]),
     .S(vdd_));
pch_hvt  vdd_cntrl_60_ ( .D(r_vdd[60]), .B(vdd_), .G(vdd_cntl_l[60]),
     .S(vdd_));
pch_hvt  vdd_cntrl_59_ ( .D(r_vdd[59]), .B(vdd_), .G(vdd_cntl_l[59]),
     .S(vdd_));
pch_hvt  vdd_cntrl_58_ ( .D(r_vdd[58]), .B(vdd_), .G(vdd_cntl_l[58]),
     .S(vdd_));
pch_hvt  vdd_cntrl_57_ ( .D(r_vdd[57]), .B(vdd_), .G(vdd_cntl_l[57]),
     .S(vdd_));
pch_hvt  vdd_cntrl_56_ ( .D(r_vdd[56]), .B(vdd_), .G(vdd_cntl_l[56]),
     .S(vdd_));
pch_hvt  vdd_cntrl_55_ ( .D(r_vdd[55]), .B(vdd_), .G(vdd_cntl_l[55]),
     .S(vdd_));
pch_hvt  vdd_cntrl_54_ ( .D(r_vdd[54]), .B(vdd_), .G(vdd_cntl_l[54]),
     .S(vdd_));
pch_hvt  vdd_cntrl_53_ ( .D(r_vdd[53]), .B(vdd_), .G(vdd_cntl_l[53]),
     .S(vdd_));
pch_hvt  vdd_cntrl_52_ ( .D(r_vdd[52]), .B(vdd_), .G(vdd_cntl_l[52]),
     .S(vdd_));
pch_hvt  vdd_cntrl_51_ ( .D(r_vdd[51]), .B(vdd_), .G(vdd_cntl_l[51]),
     .S(vdd_));
pch_hvt  vdd_cntrl_50_ ( .D(r_vdd[50]), .B(vdd_), .G(vdd_cntl_l[50]),
     .S(vdd_));
pch_hvt  vdd_cntrl_49_ ( .D(r_vdd[49]), .B(vdd_), .G(vdd_cntl_l[49]),
     .S(vdd_));
pch_hvt  vdd_cntrl_48_ ( .D(r_vdd[48]), .B(vdd_), .G(vdd_cntl_l[48]),
     .S(vdd_));
pch_hvt  vdd_cntrl_47_ ( .D(r_vdd[47]), .B(vdd_), .G(vdd_cntl_l[47]),
     .S(vdd_));
pch_hvt  vdd_cntrl_46_ ( .D(r_vdd[46]), .B(vdd_), .G(vdd_cntl_l[46]),
     .S(vdd_));
pch_hvt  vdd_cntrl_45_ ( .D(r_vdd[45]), .B(vdd_), .G(vdd_cntl_l[45]),
     .S(vdd_));
pch_hvt  vdd_cntrl_44_ ( .D(r_vdd[44]), .B(vdd_), .G(vdd_cntl_l[44]),
     .S(vdd_));
pch_hvt  vdd_cntrl_43_ ( .D(r_vdd[43]), .B(vdd_), .G(vdd_cntl_l[43]),
     .S(vdd_));
pch_hvt  vdd_cntrl_42_ ( .D(r_vdd[42]), .B(vdd_), .G(vdd_cntl_l[42]),
     .S(vdd_));
pch_hvt  vdd_cntrl_41_ ( .D(r_vdd[41]), .B(vdd_), .G(vdd_cntl_l[41]),
     .S(vdd_));
pch_hvt  vdd_cntrl_40_ ( .D(r_vdd[40]), .B(vdd_), .G(vdd_cntl_l[40]),
     .S(vdd_));
pch_hvt  vdd_cntrl_39_ ( .D(r_vdd[39]), .B(vdd_), .G(vdd_cntl_l[39]),
     .S(vdd_));
pch_hvt  vdd_cntrl_38_ ( .D(r_vdd[38]), .B(vdd_), .G(vdd_cntl_l[38]),
     .S(vdd_));
pch_hvt  vdd_cntrl_37_ ( .D(r_vdd[37]), .B(vdd_), .G(vdd_cntl_l[37]),
     .S(vdd_));
pch_hvt  vdd_cntrl_36_ ( .D(r_vdd[36]), .B(vdd_), .G(vdd_cntl_l[36]),
     .S(vdd_));
pch_hvt  vdd_cntrl_35_ ( .D(r_vdd[35]), .B(vdd_), .G(vdd_cntl_l[35]),
     .S(vdd_));
pch_hvt  vdd_cntrl_34_ ( .D(r_vdd[34]), .B(vdd_), .G(vdd_cntl_l[34]),
     .S(vdd_));
pch_hvt  vdd_cntrl_33_ ( .D(r_vdd[33]), .B(vdd_), .G(vdd_cntl_l[33]),
     .S(vdd_));
pch_hvt  vdd_cntrl_32_ ( .D(r_vdd[32]), .B(vdd_), .G(vdd_cntl_l[32]),
     .S(vdd_));
pch_hvt  vdd_cntrl_31_ ( .D(r_vdd[31]), .B(vdd_), .G(vdd_cntl_l[31]),
     .S(vdd_));
pch_hvt  vdd_cntrl_30_ ( .D(r_vdd[30]), .B(vdd_), .G(vdd_cntl_l[30]),
     .S(vdd_));
pch_hvt  vdd_cntrl_29_ ( .D(r_vdd[29]), .B(vdd_), .G(vdd_cntl_l[29]),
     .S(vdd_));
pch_hvt  vdd_cntrl_28_ ( .D(r_vdd[28]), .B(vdd_), .G(vdd_cntl_l[28]),
     .S(vdd_));
pch_hvt  vdd_cntrl_27_ ( .D(r_vdd[27]), .B(vdd_), .G(vdd_cntl_l[27]),
     .S(vdd_));
pch_hvt  vdd_cntrl_26_ ( .D(r_vdd[26]), .B(vdd_), .G(vdd_cntl_l[26]),
     .S(vdd_));
pch_hvt  vdd_cntrl_25_ ( .D(r_vdd[25]), .B(vdd_), .G(vdd_cntl_l[25]),
     .S(vdd_));
pch_hvt  vdd_cntrl_24_ ( .D(r_vdd[24]), .B(vdd_), .G(vdd_cntl_l[24]),
     .S(vdd_));
pch_hvt  vdd_cntrl_23_ ( .D(r_vdd[23]), .B(vdd_), .G(vdd_cntl_l[23]),
     .S(vdd_));
pch_hvt  vdd_cntrl_22_ ( .D(r_vdd[22]), .B(vdd_), .G(vdd_cntl_l[22]),
     .S(vdd_));
pch_hvt  vdd_cntrl_21_ ( .D(r_vdd[21]), .B(vdd_), .G(vdd_cntl_l[21]),
     .S(vdd_));
pch_hvt  vdd_cntrl_20_ ( .D(r_vdd[20]), .B(vdd_), .G(vdd_cntl_l[20]),
     .S(vdd_));
pch_hvt  vdd_cntrl_19_ ( .D(r_vdd[19]), .B(vdd_), .G(vdd_cntl_l[19]),
     .S(vdd_));
pch_hvt  vdd_cntrl_18_ ( .D(r_vdd[18]), .B(vdd_), .G(vdd_cntl_l[18]),
     .S(vdd_));
pch_hvt  vdd_cntrl_17_ ( .D(r_vdd[17]), .B(vdd_), .G(vdd_cntl_l[17]),
     .S(vdd_));
pch_hvt  vdd_cntrl_16_ ( .D(r_vdd[16]), .B(vdd_), .G(vdd_cntl_l[16]),
     .S(vdd_));
pch_hvt  vdd_cntrl_15_ ( .D(r_vdd[15]), .B(vdd_), .G(vdd_cntl_l[15]),
     .S(vdd_));
pch_hvt  vdd_cntrl_14_ ( .D(r_vdd[14]), .B(vdd_), .G(vdd_cntl_l[14]),
     .S(vdd_));
pch_hvt  vdd_cntrl_13_ ( .D(r_vdd[13]), .B(vdd_), .G(vdd_cntl_l[13]),
     .S(vdd_));
pch_hvt  vdd_cntrl_12_ ( .D(r_vdd[12]), .B(vdd_), .G(vdd_cntl_l[12]),
     .S(vdd_));
pch_hvt  vdd_cntrl_11_ ( .D(r_vdd[11]), .B(vdd_), .G(vdd_cntl_l[11]),
     .S(vdd_));
pch_hvt  vdd_cntrl_10_ ( .D(r_vdd[10]), .B(vdd_), .G(vdd_cntl_l[10]),
     .S(vdd_));
pch_hvt  vdd_cntrl_9_ ( .D(r_vdd[9]), .B(vdd_), .G(vdd_cntl_l[9]),
     .S(vdd_));
pch_hvt  vdd_cntrl_8_ ( .D(r_vdd[8]), .B(vdd_), .G(vdd_cntl_l[8]),
     .S(vdd_));
pch_hvt  vdd_cntrl_7_ ( .D(r_vdd[7]), .B(vdd_), .G(vdd_cntl_l[7]),
     .S(vdd_));
pch_hvt  vdd_cntrl_6_ ( .D(r_vdd[6]), .B(vdd_), .G(vdd_cntl_l[6]),
     .S(vdd_));
pch_hvt  vdd_cntrl_5_ ( .D(r_vdd[5]), .B(vdd_), .G(vdd_cntl_l[5]),
     .S(vdd_));
pch_hvt  vdd_cntrl_4_ ( .D(r_vdd[4]), .B(vdd_), .G(vdd_cntl_l[4]),
     .S(vdd_));
pch_hvt  vdd_cntrl_3_ ( .D(r_vdd[3]), .B(vdd_), .G(vdd_cntl_l[3]),
     .S(vdd_));
pch_hvt  vdd_cntrl_2_ ( .D(r_vdd[2]), .B(vdd_), .G(vdd_cntl_l[2]),
     .S(vdd_));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));

endmodule
// Library - leafcell, Cell - clk_mux2to1, View - schematic
// LAST TIME SAVED: Jul 24 18:58:03 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module clk_mux2to1 ( clk, cbit, cbitb, min, prog );
output  clk;

input  cbit, cbitb, prog;

input [1:0]  min;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I289 ( .A(net29), .Y(clk));
inv_hvt I288 ( .A(prog), .Y(net27));
nand2_hvt I287 ( .A(net27), .Y(net29), .B(st2));
txgate_hvt I249 ( .in(min[1]), .out(st2), .pp(cbitb), .nn(cbit));
txgate_hvt I248 ( .in(min[0]), .out(st2), .pp(cbit), .nn(cbitb));

endmodule
// Library - leafcell, Cell - clk_mux2to1x4, View - schematic
// LAST TIME SAVED: Sep 26 10:53:26 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module clk_mux2to1x4 ( gnet, bl, min0, min1, min2, min3, pgate_l,
     pgate_r, prog, reset_l, reset_r, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r );


input  prog;

output [3:0]  gnet;

inout [3:0]  bl;

input [1:0]  min1;
input [1:0]  vdd_cntl_l;
input [1:0]  vdd_cntl_r;
input [1:0]  pgate_r;
input [1:0]  min3;
input [1:0]  wl_r;
input [1:0]  min0;
input [1:0]  pgate_l;
input [1:0]  reset_r;
input [1:0]  reset_l;
input [1:0]  min2;
input [1:0]  wl_l;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [7:0]  cbitb;

wire  [7:0]  cbit;

wire  [0:1]  l_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(l_vdd[0]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(l_vdd[1]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl_r[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl_r[0]), .S(vdd_));
cram2x2 I292 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset_l[1:0]),
     .q(cbit[3:0]), .wl(wl_l[1:0]), .r_vdd(l_vdd[0:1]),
     .pgate(pgate_l[1:0]));
cram2x2 I298 ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset_r[1:0]),
     .q(cbit[7:4]), .wl(wl_r[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate_r[1:0]));
clk_mux2to1 I295 ( .prog(prog), .cbit(cbit[3]), .cbitb(cbitb[3]),
     .min(min3[1:0]), .clk(gnet[3]));
clk_mux2to1 I293 ( .prog(prog), .cbit(cbit[1]), .cbitb(cbitb[1]),
     .min(min1[1:0]), .clk(gnet[1]));
clk_mux2to1 I294 ( .prog(prog), .cbit(cbit[2]), .cbitb(cbitb[2]),
     .min(min2[1:0]), .clk(gnet[2]));
clk_mux2to1 I291 ( .prog(prog), .cbit(cbit[0]), .cbitb(cbitb[0]),
     .min(min0[1:0]), .clk(gnet[0]));

endmodule
// Library - ice4chip, Cell - CHIP_route_right_ice4f_guc, View -
//schematic
// LAST TIME SAVED: Apr 21 19:24:04 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module CHIP_route_right_ice4f_guc ( bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bldld, cm_banksel_bltrd1_3_,
     cm_clk_blbrd, cm_clk_bltrd1, cm_sdi_u0, cm_sdi_u1, cm_sdi_u2d,
     cm_sdi_u3d2, core_por_b0, core_por_b1, core_por_b_rowu2,
     core_por_b_rowu3, core_por_bb, cram_pgateoff, cram_prec,
     cram_prec_blbrd, cram_prec_bltrd1, cram_pullup_b,
     .cram_pullup_b_blbrd(cram_pullup_b_bldrd), cram_pullup_b_bltrd1,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, cram_write_blbrd,
     cram_write_bltrd1, data_muxsel, data_muxsel1, data_muxsel1_blbrd,
     data_muxsel1_bltrd1, data_muxsel_blbrd, data_muxsel_bltrd1,
     .en_8bcibfig_b_bltrd1(en_8bconfig_b_bltrd1), en_8bconfig_b,
     en_8bconfig_b_blbrd, end_of_startup, gint_hz, gsr, hiz_b0,
     j_rst_b, j_tck, j_tdi, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr, md_spi_b, mode0,
     nvcm_spi_sdi, nvcm_spi_ss_b, pgate_r, psdo, reset_b_r, row_test0,
     rst_b, sdo_enable, shift0, smc_clk_out, smc_load_nvcm_bstream,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk, smc_wdis_dclk_blbrd,
     smc_wdis_dclk_bltrd1, smc_write0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, totdopad, update0, vdd_cntl_r, wl_r,
     bm_sdo_o, bp0, cdone_in, cf_r, cm_sdo_u0d1, cm_sdo_u1d3,
     cm_sdo_u2d1, cm_sdo_u3, crst_filterout, fabric_out_122,
     fabric_out_126, fabric_out_136, fromsdo, last_rsr3,
     monitor_celld4, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, smc_core_por_bottom1, smc_core_por_bottom2,
     spi_ss_in_bbank, spi_ss_in_r, tck_pad, tdi_pad, tms_pad, trst_pad,
     vddio_rightbank );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bltrd1_3_, cm_clk_blbrd,
     cm_clk_bltrd1, core_por_b0, core_por_b1, core_por_b_rowu2,
     core_por_b_rowu3, core_por_bb, cram_pgateoff, cram_prec,
     cram_prec_blbrd, cram_prec_bltrd1, cram_pullup_b,
     cram_pullup_b_bldrd, cram_pullup_b_bltrd1, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, cram_write_blbrd, cram_write_bltrd1,
     data_muxsel, data_muxsel1, data_muxsel1_blbrd,
     data_muxsel1_bltrd1, data_muxsel_blbrd, data_muxsel_bltrd1,
     en_8bconfig_b_bltrd1, en_8bconfig_b, en_8bconfig_b_blbrd,
     end_of_startup, gint_hz, gsr, hiz_b0, j_rst_b, j_tck, j_tdi,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, nvcm_spi_sdi, nvcm_spi_ss_b, row_test0, rst_b, sdo_enable,
     shift0, smc_clk_out, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk, smc_wdis_dclk_blbrd,
     smc_wdis_dclk_bltrd1, smc_write0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, totdopad, update0;

input  bp0, cdone_in, crst_filterout, fabric_out_122, fabric_out_126,
     fabric_out_136, fromsdo, last_rsr3, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, tck_pad, tdi_pad,
     tms_pad, trst_pad, vddio_rightbank;

output [351:0]  wl_r;
output [351:0]  vdd_cntl_r;
output [3:0]  bm_sdi_i;
output [7:1]  psdo;
output [351:0]  pgate_r;
output [1:0]  cm_sdi_u2d;
output [1:0]  cm_sdi_u0;
output [351:0]  reset_b_r;
output [1:0]  cm_sdi_u3d2;
output [1:0]  last_rsr;
output [1:0]  cm_sdi_u1;
output [3:0]  bm_banksel_i;
output [1:0]  cm_banksel_bldld;
output [7:0]  bm_sa_i;

input [1:0]  cm_sdo_u2d1;
input [3:0]  bm_sdo_o;
input [1:0]  cf_r;
input [1:0]  cm_sdo_u0d1;
input [1:0]  monitor_celld4;
input [1:0]  cm_sdo_u1d3;
input [4:0]  spi_ss_in_bbank;
input [1:0]  cm_sdo_u3;
input [7:1]  spi_ss_in_r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdi_u3;

wire  [1:0]  smc_osco_fsel;

wire  [1:0]  cm_sdi_u2;

wire  [7:1]  spi_ss_in_rd;

wire  [3:2]  monitor_celldd;

wire  [1:0]  cm_sdo_u3d1;

wire  [3:0]  cm_banksel;

wire  [1:0]  u1_in;

wire  [1:0]  u0_in;



CHIP_route_right0smc I462 ( .vddio_rightbank(vddio_rightbank),
     .spi_ss_in_r(spi_ss_in_r[7:1]), .last_rsr(last_rsr[1:0]),
     .cm_banksel_bltrd1_3_(cm_banksel_bltrd1_3_),
     .crst_filterout(crst_filterout), .cm_sdo_u3(cm_sdo_u3[1:0]),
     .vdd_cntl_r(vdd_cntl_r[351:0]),
     .smc_wdis_dclk_bltrd1(smc_wdis_dclk_bltrd1),
     .reset_b_r(reset_b_r[351:0]),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd_2_),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .j_tck(j_tck), .en_8bcibfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel1_bltrd1(data_muxsel1_bltrd1),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1), .core_por_b1(core_por_b1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .cm_clk_bltrd1(cm_clk_bltrd1),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1), .wl_r(wl_r[351:0]),
     .cm_sdi_u2(cm_sdi_u2[1:0]), .cm_sdi_u3(cm_sdi_u3[1:0]),
     .smc_podt_rst(smc_podt_rst), .smc_osco_fsel(smc_osco_fsel[1:0]),
     .smc_oscoff_b(smc_oscoff_b), .smc_podt_off(smc_podt_off),
     .cnt_podt_out(cnt_podt_out), .osc_clk(osc_clk),
     .u1_in(u1_in[1:0]), .u0_in(u0_in[1:0]),
     .spi_ss_in_rd(spi_ss_in_rd[7:1]), .cm_sdo_u3d1(cm_sdo_u3d1[1:0]),
     .cm_banksel(cm_banksel[3:0]),
     .smc_row_inc_fromsmc(smc_row_inc_fromsmc),
     .smc_rsr_rst_fromsmc(smc_rsr_rst_fromsmc),
     .smc_wwlwrt_en(smc_wwlwrt_en),
     .smc_wset_precgnd(smc_wset_precgnd), .smc_seq_rst(smc_seq_rst),
     .smc_write(smc_write0), .smc_rwl_en(smc_rwl_en),
     .smc_wcram_rst(smc_wcram_rst), .smc_wset_prec(smc_wset_prec),
     .smc_rrst_pullwlen(smc_rrst_pullwlen), .smc_read(net355),
     .smc_rprec(smc_rprec), .smc_rpull_b(smc_rpull_b),
     .smc_clk(cm_clk), .smc_write0(smc_write0), .cf_r(cf_r[1:0]),
     .core_por_b_rowu2(core_por_b_rowu2), .core_por_b0(core_por_b0),
     .row_test0(row_test0), .smc_row_inc(smc_row_inc),
     .cram_pgateoff(cram_pgateoff), .core_por_bb(core_por_bb),
     .smc_wwlwrt_dis(smc_wwlwrt_dis), .cram_wl_en(cram_wl_en),
     .cram_vddoff(cram_vddoff), .cram_rst(cram_rst),
     .smc_rsr_rst(smc_rsr_rst), .j_rst_b(j_rst_b),
     .cram_prec_blbrd(cram_prec_blbrd),
     .cram_pullup_b_blbrd(cram_pullup_b_bldrd),
     .cram_write_blbrd(cram_write_blbrd),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .cm_clk_blbrd(cm_clk_blbrd),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk(smc_wdis_dclk), .smc_clk_out(smc_clk_out),
     .en_8bconfig_b(en_8bconfig_b), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel), .cram_write(cram_write),
     .cram_prec(cram_prec), .cram_pullup_b(cram_pullup_b),
     .core_por_b_rowu3(core_por_b_rowu3), .pgate_r(pgate_r[351:0]),
     .cm_banksel_bldld(cm_banksel_bldld[1:0]),
     .monitor_celldd(monitor_celldd[3:2]), .smc_por_b0(smc_por_b0));
// smc_and_jtag_ice4frr I_smc_and_jtag (
smc_and_jtag I_smc_and_jtag (
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot), .bp0(bp0),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_spi_ss_b(nvcm_spi_ss_b), .nvcm_spi_sdi(nvcm_spi_sdi),
     .j_shift0(shift0), .j_ceb0(ceb0), .warmboot_sel({fabric_out_126,
     fabric_out_122}), .trst_pad(trst_pad), .tms_pad(tms_pad),
     .tdi_pad(tdi_pad), .tck_pad(tck_pad),
     .spi_ss_in_b(spi_ss_in_bbank[4]), .spi_sdi(spi_ss_in_bbank[2]),
     .spi_clk_in(spi_ss_in_bbank[3]), .psdi(spi_ss_in_rd[7:1]),
     .por_b(smc_por_b0), .osc_clk(osc_clk), .creset_b(crst_filterout),
     .coldboot_sel(spi_ss_in_bbank[1:0]), .cnt_podt_out(cnt_podt_out),
     .cm_sdo_u3(cm_sdo_u3d1[1:0]), .cm_sdo_u2(cm_sdo_u2d1[1:0]),
     .cm_sdo_u1(cm_sdo_u1d3[1:0]), .cm_sdo_u0(cm_sdo_u0d1[1:0]),
     .cm_monitor_cell({monitor_celldd[3:2], monitor_celld4[1:0]}),
     .cm_last_rsr(last_rsr3), .cdone_in(cdone_in),
     .bschain_sdo(fromsdo), .boot(fabric_out_136),
     .bm_bank_sdo(bm_sdo_o[3:0]), .tdo_pad(totdopad),
     .tdo_oe_pad(sdo_enable), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .spi_clk_out(spi_clk_out), .smc_wwlwrt_en(smc_wwlwrt_en),
     .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wdis_dclk(smc_wdis_dclk), .smc_wcram_rst(smc_wcram_rst),
     .smc_seq_rst(smc_seq_rst), .smc_rwl_en(smc_rwl_en),
     .smc_rsr_rst(smc_rsr_rst_fromsmc),
     .smc_rrst_pullwlen(smc_rrst_pullwlen), .smc_rpull_b(smc_rpull_b),
     .smc_rprec(smc_rprec), .smc_row_inc(smc_row_inc_fromsmc),
     .cm_clk(cm_clk), .smc_read(net355), .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]), .psdo(psdo[7:1]),
     .md_spi_b(md_spi_b), .j_upd_dr(update0), .j_tdi(j_tdi),
     .j_tck(j_tck), .j_sft_dr(shiftfromsmc), .j_rst_b(j_rst_b),
     .j_row_test(row_test0), .j_mode(mode0), .j_hiz_b(hiz_b0),
     .gsr(gsr), .gint_hz(gint_hz), .end_of_startup(end_of_startup),
     .en_8bconfig_b(en_8bconfig_b), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel), .cm_sdi_u3(cm_sdi_u3[1:0]),
     .cm_sdi_u2(cm_sdi_u2[1:0]), .cm_sdi_u1(u1_in[1:0]),
     .cm_sdi_u0(u0_in[1:0]), .cm_banksel(cm_banksel[3:0]),
     .cdone_out(cdone_out), .bs_en(bs_en0),
     .bm_wdummymux_en(bm_wdummymux_en_i), .bm_sreb(bm_sreb_i),
     .bm_sclkrw(bm_sclkrw_i), .bm_sa(bm_sa_i[7:0]),
     .bm_rcapmux_en(bm_rcapmux_en_i), .bm_init(bm_init_i),
     .bm_clk(bm_sclk_i), .bm_banksel(bm_banksel_i[3:0]),
     .bm_bank_sdi(bm_sdi_i[3:0]), .bm_sweb(bm_sweb_i));

endmodule
// Library - leafcell, Cell - QUAD_x4, View - schematic
// LAST TIME SAVED: Feb  8 14:15:23 2008
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module QUAD_x4 ( bm_sdo_o, cf_b, cf_l, cf_r, cf_t, fabric_out_122,
     fabric_out_126, fabric_out_136, padeb_b, padeb_l, padeb_r,
     padeb_t, pado_b, pado_l, pado_r, pado_t, sdo_pad, spi_ss_in_b,
     spi_ss_in_lft_b, spi_ss_in_r, bl_bot, bl_top, bm_banksel_i,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en,
     cdone_in_bot_r, ceb, end_of_startup_l, end_of_startup_r,
     end_of_startup_t, hiz_b, mode, padin_b, padin_l, padin_r, padin_t,
     pgate_l, pgate_r, prog, purst, r, reset_b_l, reset_b_r, sdi_pad,
     shift, spioeb_b, spioeb_lft_b, spiout_b, spiout_lft_b, spiout_r,
     tclk, tiegnd, tievdd, update, vdd_cntl_l, vdd_cntl_r, wl_l, wl_r
     );
output  fabric_out_122, fabric_out_126, fabric_out_136, sdo_pad;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb, hiz_b, mode, prog,
     purst, r, sdi_pad, shift, tclk, tiegnd, tievdd, update;

output [47:24]  spi_ss_in_b;
output [19:0]  spi_ss_in_lft_b;
output [47:0]  padeb_t;
output [479:0]  cf_l;
output [39:0]  padeb_l;
output [479:0]  cf_r;
output [47:0]  pado_b;
output [3:0]  bm_sdo_o;
output [39:0]  pado_l;
output [47:0]  padeb_b;
output [575:0]  cf_b;
output [39:0]  pado_r;
output [47:0]  pado_t;
output [39:0]  padeb_r;
output [39:0]  spi_ss_in_r;
output [575:0]  cf_t;

inout [1311:0]  bl_bot;
inout [1311:0]  bl_top;

input [19:0]  spiout_r;
input [19:0]  spioeb_lft_b;
input [7:0]  bm_sa_i;
input [3:0]  bm_sdi_i;
input [47:24]  spioeb_b;
input [39:0]  padin_r;
input [19:0]  spiout_lft_b;
input [3:0]  bm_banksel_i;
input [47:24]  spiout_b;
input [19:0]  end_of_startup_r;
input [351:0]  wl_l;
input [23:0]  end_of_startup_t;
input [39:0]  padin_l;
input [351:0]  pgate_r;
input [351:0]  wl_r;
input [47:0]  padin_t;
input [19:0]  end_of_startup_l;
input [351:0]  vdd_cntl_r;
input [351:0]  pgate_l;
input [351:0]  vdd_cntl_l;
input [351:0]  reset_b_l;
input [11:0]  cdone_in_bot_r;
input [351:0]  reset_b_r;
input [47:0]  padin_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net1235;

wire  [0:47]  net1417;

wire  [0:23]  net1499;

wire  [0:23]  net1318;

wire  [0:7]  net810;

wire  [0:7]  net1296;

wire  [0:23]  net965;

wire  [0:7]  net1333;

wire  [0:47]  net1322;

wire  [0:7]  net1029;

wire  [0:7]  net815;

wire  [0:47]  net1405;

wire  [0:47]  net1421;

wire  [0:7]  net1207;

wire  [0:23]  net1500;

wire  [0:7]  net1027;

wire  [0:7]  net1339;

wire  [0:7]  net1552;

wire  [0:47]  net1416;

wire  [0:23]  net1320;

wire  [0:23]  net1390;

wire  [0:15]  net1508;

wire  [0:7]  net1327;

wire  [0:23]  net966;

wire  [0:47]  net1616;

wire  [0:7]  net1654;

wire  [0:7]  net1344;

wire  [0:23]  net1503;

wire  [0:23]  net1391;

wire  [0:7]  net1700;

wire  [0:47]  net1398;

wire  [0:1]  net1698;

wire  [0:47]  net1603;

wire  [0:47]  net984;

wire  [0:7]  net1354;

wire  [0:47]  net1420;

wire  [0:7]  net1332;

wire  [0:23]  net1315;

wire  [0:47]  net1350;

wire  [0:23]  net960;

wire  [0:23]  net1392;

wire  [0:47]  net1611;

wire  [0:7]  net809;

wire  [3:0]  slf_op_13_21;

wire  [0:7]  net1515;

wire  [0:7]  net1559;

wire  [0:23]  net1501;

wire  [0:47]  net1396;

wire  [0:7]  net1556;

wire  [0:1]  net1292;

wire  [0:7]  net1522;

wire  [0:47]  net988;

wire  [0:1]  net1289;

wire  [0:23]  net1313;

wire  [0:47]  net1615;

wire  [0:7]  net817;

wire  [0:23]  net962;

wire  [0:47]  net1403;

wire  [0:7]  net1233;

wire  [0:7]  net1331;

wire  [0:23]  net1384;

wire  [0:7]  net1517;

wire  [0:23]  net1314;

wire  [0:7]  net1514;

wire  [3:0]  slf_op_12_00;

wire  [0:1]  net1379;

wire  [0:47]  net1411;

wire  [0:23]  net961;

wire  [0:7]  net1342;

wire  [1:0]  bm_bank10_banksel_o;

wire  [0:47]  net1422;

wire  [0:7]  net1352;

wire  [0:47]  net1612;

wire  [0:7]  net1678;

wire  [0:1]  net1716;

wire  [0:7]  net1553;

wire  [0:47]  net981;

wire  [3:0]  slf_op_13_00;

wire  [0:47]  net1610;

wire  [0:7]  net1037;

wire  [0:23]  net1381;

wire  [0:7]  net1032;

wire  [0:23]  net1386;

wire  [0:7]  net1554;

wire  [0:3]  net1667;

wire  [3:0]  slf_op_12_21;

wire  [0:47]  net1410;

wire  [0:1]  net1294;

wire  [0:3]  net1671;

wire  [0:7]  net1031;

wire  [0:47]  net1618;

wire  [7:0]  glb_net;

wire  [0:23]  net969;

wire  [0:47]  net1614;

wire  [0:23]  net1383;

wire  [0:7]  net1338;

wire  [0:7]  net1558;

wire  [0:3]  net1666;

wire  [0:7]  net1034;

wire  [0:23]  net1382;

wire  [0:7]  net816;

wire  [0:7]  net1345;

wire  [0:47]  net1617;

wire  [0:23]  net963;

wire  [0:23]  net1317;

wire  [0:7]  net1231;

wire  [0:7]  net1035;

wire  [0:7]  net1028;

wire  [0:7]  net1551;

wire  [0:47]  net1409;

wire  [0:7]  net1537;

wire  [3:0]  slf_op_00_11;

wire  [0:7]  net819;

wire  [0:7]  net1340;

wire  [0:47]  net1600;

wire  [0:23]  net1385;

wire  [0:47]  net991;

wire  [0:7]  net1343;

wire  [0:47]  net987;

wire  [0:23]  net1504;

wire  [1:0]  bm_sweb_b2_o;

wire  [0:47]  net990;

wire  [0:47]  net983;

wire  [0:7]  net1229;

wire  [0:1]  net1721;

wire  [0:7]  net1360;

wire  [0:15]  net1299;

wire  [1:0]  bm_sdi_b2_o;

wire  [0:7]  net1334;

wire  [0:23]  net1388;

wire  [0:7]  net1359;

wire  [0:47]  net1401;

wire  [0:47]  net1419;

wire  [0:7]  net820;

wire  [0:7]  net1426;

wire  [0:47]  net980;

wire  [0:7]  net1227;

wire  [0:47]  net1394;

wire  [0:7]  net1357;

wire  [0:23]  net1312;

wire  [0:7]  net1330;

wire  [0:47]  net1395;

wire  [0:7]  net1518;

wire  [0:7]  net813;

wire  [0:23]  net1505;

wire  [0:47]  net986;

wire  [0:7]  net1033;

wire  [0:7]  net811;

wire  [3:0]  slf_op_00_10;

wire  [0:47]  net1601;

wire  [0:47]  net1606;

wire  [0:47]  net1404;

wire  [0:23]  net1389;

wire  [0:7]  net1341;

wire  [0:7]  net1321;

wire  [0:7]  net1232;

wire  [0:23]  net959;

wire  [0:7]  net1328;

wire  [0:23]  net1387;

wire  [0:47]  net1605;

wire  [0:23]  net968;

wire  [0:7]  net1234;

wire  [3:0]  slf_op_25_10;

wire  [0:7]  net1310;

wire  [0:23]  net964;

wire  [0:7]  net858;

wire  [0:7]  net1516;

wire  [0:47]  net985;

wire  [0:23]  net1506;

wire  [0:7]  net1548;

wire  [0:7]  net1520;

wire  [0:23]  net1507;

wire  [0:23]  net1316;

wire  [0:47]  net989;

wire  [0:7]  net1230;

wire  [0:47]  net1609;

wire  [1:0]  bm_sclkrw_b2_o;

wire  [0:7]  net1284;

wire  [0:47]  net1408;

wire  [0:7]  net1415;

wire  [0:23]  net958;

wire  [0:47]  net1414;

wire  [0:47]  net1400;

wire  [0:23]  net967;

wire  [0:7]  net1329;

wire  [0:7]  net1335;

wire  [0:47]  net1613;

wire  [0:1]  net1715;

wire  [0:7]  net812;

wire  [0:7]  net1519;

wire  [0:1]  net869;

wire  [0:47]  net1413;

wire  [0:7]  net1353;

wire  [0:47]  net1418;

wire  [0:7]  net1325;

wire  [0:23]  net1498;

wire  [0:47]  net1402;

wire  [0:7]  net1355;

wire  [0:7]  net1326;

wire  [0:7]  net1555;

wire  [0:47]  net1412;

wire  [0:3]  net1024;

wire  [0:7]  net1521;

wire  [0:47]  net1602;

wire  [3:0]  bm_bank30_banksel_o;

wire  [0:47]  net1607;

wire  [1:0]  bm_bank30_sclk_o;

wire  [0:47]  net982;

wire  [0:15]  net884;

wire  [0:47]  net1393;

wire  [0:47]  net1323;

wire  [0:47]  net1604;

wire  [0:23]  net1502;

wire  [0:7]  net1356;

wire  [0:7]  net1236;

wire  [0:15]  net1324;

wire  [1:0]  bm_sweb_b0_o;

wire  [0:47]  net1407;

wire  [0:1]  net866;

wire  [0:47]  net1397;

wire  [0:23]  net1319;

wire  [0:47]  net1399;

wire  [0:7]  net1036;

wire  [0:7]  net1030;

wire  [0:7]  net1557;

wire  [3:0]  bm_bank30_sdi_o;

wire  [0:47]  net1406;

wire  [3:0]  bm_bank30_sdo_i;

wire  [0:1]  net867;

wire  [7:0]  bm_sa_b1_o;

wire  [0:23]  net1311;

wire  [0:47]  net1599;

wire  [0:7]  net814;

wire  [1:0]  bm_sdi_b0_o;

wire  [1:0]  bm_sclkrw_b0_o;

wire  [0:7]  net1228;

wire  [0:7]  net1358;



QUAD_BR I_BR ( .ceb_mi(ceb), .ceb_o(net01027), .ceb_i(net01230),
     .tnr_op_24_10(net1024[0:3]), .bnl_op_13_01(slf_op_12_00[3:0]),
     .tiegnd(tiegnd), .tnl_op_24_10(net809[0:7]),
     .tnl_op_25_10(net810[0:7]), .tnl_op_21_10(net811[0:7]),
     .tnl_op_20_10(net812[0:7]), .tnl_op_19_10(net813[0:7]),
     .tnl_op_18_10(net814[0:7]), .tnl_op_17_10(net815[0:7]),
     .tnl_op_16_10(net816[0:7]), .tnl_op_15_10(net817[0:7]),
     .tnl_op_14_10(net1310[0:7]), .tnl_op_23_10(net819[0:7]),
     .tnl_op_22_10(net820[0:7]), .tnr_op_23_10(net810[0:7]),
     .tnr_op_22_10(net809[0:7]), .tnr_op_21_10(net819[0:7]),
     .tnr_op_20_10(net820[0:7]), .tnr_op_19_10(net811[0:7]),
     .tnr_op_18_10(net812[0:7]), .tnr_op_17_10(net813[0:7]),
     .tnr_op_16_10(net814[0:7]), .tnr_op_15_10(net815[0:7]),
     .tnr_op_14_10(net816[0:7]), .tnr_op_13_10(net817[0:7]),
     .hiz_b_o(net832), .bs_en_o(net833), .r_o(net834),
     .update_o(net835), .mode_o(net836), .tclk_o(net837),
     .tclk_mi(tclk), .bs_en_mi(bs_en), .r_mi(r), .hiz_b_mi(hiz_b),
     .update_mi(update), .shift_mi(shift), .update_i(net1265),
     .mode_i(net1264), .shift_o(net846), .shift_i(net1261),
     .r_i(net1262), .hiz_b_i(net1263), .mode_mi(mode),
     .bs_en_i(net1260), .tclk_i(net1266), .bm_sdi_o(bm_sdi_b2_o[1:0]),
     .bm_sweb_o(bm_sweb_b2_o[1:0]), .bm_sreb_o(net855),
     .bm_sclkrw_o(bm_sclkrw_b2_o[1:0]), .bm_sclk_o(net857),
     .bm_sa_o(net858[0:7]), .bm_init_o(net859), .bm_sdo_i({bm_sdo_b3_o,
     bm_sdi_b2_o[0]}), .bm_rcapmux_en_o(net861),
     .bm_wdummymux_en_o(net862), .bm_sdi_i(bm_bank30_sdi_o[3:2]),
     .bm_rcapmux_en_i(net1681), .bm_wdummymux_en_i(net1682),
     .bm_sdo_o(net866[0:1]), .bm_sweb_i(net867[0:1]),
     .bm_sreb_i(net1675), .bm_sclkrw_i(net869[0:1]),
     .bm_sclk_i(bm_bank30_sclk_o[1]), .bm_sa_i(net1678[0:7]),
     .bm_init_i(net1679), .cdone_in_rgt_b(end_of_startup_r[9:0]),
     .cdone_in_bot_r(cdone_in_bot_r[11:0]), .vdd_cntl({vdd_cntl_r[174],
     vdd_cntl_r[175], vdd_cntl_r[172], vdd_cntl_r[173],
     vdd_cntl_r[170], vdd_cntl_r[171], vdd_cntl_r[168],
     vdd_cntl_r[169], vdd_cntl_r[166], vdd_cntl_r[167],
     vdd_cntl_r[164], vdd_cntl_r[165], vdd_cntl_r[162],
     vdd_cntl_r[163], vdd_cntl_r[160], vdd_cntl_r[161],
     vdd_cntl_r[158], vdd_cntl_r[159], vdd_cntl_r[156],
     vdd_cntl_r[157], vdd_cntl_r[154], vdd_cntl_r[155],
     vdd_cntl_r[152], vdd_cntl_r[153], vdd_cntl_r[150],
     vdd_cntl_r[151], vdd_cntl_r[148], vdd_cntl_r[149],
     vdd_cntl_r[146], vdd_cntl_r[147], vdd_cntl_r[144],
     vdd_cntl_r[145], vdd_cntl_r[142], vdd_cntl_r[143],
     vdd_cntl_r[140], vdd_cntl_r[141], vdd_cntl_r[138],
     vdd_cntl_r[139], vdd_cntl_r[136], vdd_cntl_r[137],
     vdd_cntl_r[134], vdd_cntl_r[135], vdd_cntl_r[132],
     vdd_cntl_r[133], vdd_cntl_r[130], vdd_cntl_r[131],
     vdd_cntl_r[128], vdd_cntl_r[129], vdd_cntl_r[126],
     vdd_cntl_r[127], vdd_cntl_r[124], vdd_cntl_r[125],
     vdd_cntl_r[122], vdd_cntl_r[123], vdd_cntl_r[120],
     vdd_cntl_r[121], vdd_cntl_r[118], vdd_cntl_r[119],
     vdd_cntl_r[116], vdd_cntl_r[117], vdd_cntl_r[114],
     vdd_cntl_r[115], vdd_cntl_r[112], vdd_cntl_r[113],
     vdd_cntl_r[110], vdd_cntl_r[111], vdd_cntl_r[108],
     vdd_cntl_r[109], vdd_cntl_r[106], vdd_cntl_r[107],
     vdd_cntl_r[104], vdd_cntl_r[105], vdd_cntl_r[102],
     vdd_cntl_r[103], vdd_cntl_r[100], vdd_cntl_r[101], vdd_cntl_r[98],
     vdd_cntl_r[99], vdd_cntl_r[96], vdd_cntl_r[97], vdd_cntl_r[94],
     vdd_cntl_r[95], vdd_cntl_r[92], vdd_cntl_r[93], vdd_cntl_r[90],
     vdd_cntl_r[91], vdd_cntl_r[88], vdd_cntl_r[89], vdd_cntl_r[86],
     vdd_cntl_r[87], vdd_cntl_r[84], vdd_cntl_r[85], vdd_cntl_r[82],
     vdd_cntl_r[83], vdd_cntl_r[80], vdd_cntl_r[81], vdd_cntl_r[78],
     vdd_cntl_r[79], vdd_cntl_r[76], vdd_cntl_r[77], vdd_cntl_r[74],
     vdd_cntl_r[75], vdd_cntl_r[72], vdd_cntl_r[73], vdd_cntl_r[70],
     vdd_cntl_r[71], vdd_cntl_r[68], vdd_cntl_r[69], vdd_cntl_r[66],
     vdd_cntl_r[67], vdd_cntl_r[64], vdd_cntl_r[65], vdd_cntl_r[62],
     vdd_cntl_r[63], vdd_cntl_r[60], vdd_cntl_r[61], vdd_cntl_r[58],
     vdd_cntl_r[59], vdd_cntl_r[56], vdd_cntl_r[57], vdd_cntl_r[54],
     vdd_cntl_r[55], vdd_cntl_r[52], vdd_cntl_r[53], vdd_cntl_r[50],
     vdd_cntl_r[51], vdd_cntl_r[48], vdd_cntl_r[49], vdd_cntl_r[46],
     vdd_cntl_r[47], vdd_cntl_r[44], vdd_cntl_r[45], vdd_cntl_r[42],
     vdd_cntl_r[43], vdd_cntl_r[40], vdd_cntl_r[41], vdd_cntl_r[38],
     vdd_cntl_r[39], vdd_cntl_r[36], vdd_cntl_r[37], vdd_cntl_r[34],
     vdd_cntl_r[35], vdd_cntl_r[32], vdd_cntl_r[33], vdd_cntl_r[30],
     vdd_cntl_r[31], vdd_cntl_r[28], vdd_cntl_r[29], vdd_cntl_r[26],
     vdd_cntl_r[27], vdd_cntl_r[24], vdd_cntl_r[25], vdd_cntl_r[22],
     vdd_cntl_r[23], vdd_cntl_r[20], vdd_cntl_r[21], vdd_cntl_r[18],
     vdd_cntl_r[19], vdd_cntl_r[16], vdd_cntl_r[17], vdd_cntl_r[0],
     vdd_cntl_r[1], vdd_cntl_r[3], vdd_cntl_r[2], vdd_cntl_r[4],
     vdd_cntl_r[5], vdd_cntl_r[7], vdd_cntl_r[6], vdd_cntl_r[8],
     vdd_cntl_r[9], vdd_cntl_r[11], vdd_cntl_r[10], vdd_cntl_r[12],
     vdd_cntl_r[13], vdd_cntl_r[15], vdd_cntl_r[14]}),
     .cf_r(cf_r[239:0]), .cf_b(cf_b[575:288]),
     .hold_b_r(bank_cntl_bottom), .hold_r_b(bank_cntl_right),
     .padin_94(padin_94), .padin_162(padin_162), .glb_in(glb_net[7:0]),
     .slf_op_13_00(slf_op_13_00[3:0]), .sp4_v_t_25_10(net884[0:15]),
     .spioeb_b(spioeb_b[47:24]), .padeb_b(padeb_b[47:24]),
     .pado_b(pado_b[47:24]), .padin_b(padin_b[47:24]),
     .spi_ss_in_b(spi_ss_in_b[47:24]), .top_op_24_10(net810[0:7]),
     .top_op_23_10(net809[0:7]), .top_op_22_10(net819[0:7]),
     .top_op_21_10(net820[0:7]), .top_op_20_10(net811[0:7]),
     .top_op_19_10(net812[0:7]), .top_op_18_10(net813[0:7]),
     .top_op_17_10(net814[0:7]), .top_op_16_10(net815[0:7]),
     .top_op_15_10(net816[0:7]), .top_op_14_10(net817[0:7]),
     .top_op_13_10(net1310[0:7]), .fabric_out_94(fabric_out_94),
     .tnl_op_13_10(net1415[0:7]), .spiout_r(spiout_r[19:0]),
     .spiout_b(spiout_b[47:24]), .spioeb_r({tievdd, tievdd, tiegnd,
     tievdd, tiegnd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tiegnd}), .sdi_pad(sdi_pad), .padin_r(padin_r[19:0]),
     .fabric_out_98(bank_cntl_bottom), .lft_op_13_10(net1537[0:7]),
     .lft_op_13_09(net1352[0:7]), .lft_op_13_08(net1353[0:7]),
     .lft_op_13_07(net1354[0:7]), .lft_op_13_06(net1355[0:7]),
     .lft_op_13_05(net1356[0:7]), .lft_op_13_04(net1357[0:7]),
     .lft_op_13_03(net1426[0:7]), .lft_op_13_02(net1358[0:7]),
     .lft_op_13_01(net1359[0:7]), .slf_op_25_10(slf_op_25_10[3:0]),
     .fabric_out_162(fabric_out_162), .spi_ss_in_r(spi_ss_in_r[19:0]),
     .slf_op_24_10(net1027[0:7]), .slf_op_23_10(net1028[0:7]),
     .slf_op_22_10(net1029[0:7]), .slf_op_21_10(net1030[0:7]),
     .slf_op_20_10(net1031[0:7]), .slf_op_19_10(net1032[0:7]),
     .slf_op_18_10(net1033[0:7]), .slf_op_17_10(net1034[0:7]),
     .slf_op_16_10(net1035[0:7]), .slf_op_15_10(net1036[0:7]),
     .slf_op_14_10(net1037[0:7]), .slf_op_13_10(net1548[0:7]),
     .slf_op_13_09(net1338[0:7]), .slf_op_13_08(net1339[0:7]),
     .slf_op_13_07(net1321[0:7]), .slf_op_13_06(net1340[0:7]),
     .slf_op_13_05(net1341[0:7]), .slf_op_13_04(net1342[0:7]),
     .slf_op_13_03(net1343[0:7]), .slf_op_13_02(net1344[0:7]),
     .slf_op_13_01(net1345[0:7]), .sdo_pad(sdo_pad),
     .pado_r(pado_r[19:0]), .padeb_r(padeb_r[19:0]),
     .fabric_out_136(fabric_out_136), .carry_out_24_10(net948),
     .carry_out_23_10(net949), .carry_out_22_10(net950),
     .carry_out_21_10(net951), .carry_out_20_10(net952),
     .carry_out_18_10(net953), .carry_out_15_10(net954),
     .carry_out_17_10(net955), .carry_out_16_10(net956),
     .carry_out_14_10(net957), .sp12_v_t_24_10(net958[0:23]),
     .sp12_v_t_23_10(net959[0:23]), .sp12_v_t_22_10(net960[0:23]),
     .sp12_v_t_21_10(net961[0:23]), .sp12_v_t_20_10(net962[0:23]),
     .sp12_v_t_19_10(net963[0:23]), .sp12_v_t_18_10(net964[0:23]),
     .sp12_v_t_17_10(net965[0:23]), .sp12_v_t_16_10(net966[0:23]),
     .sp12_v_t_15_10(net967[0:23]), .sp12_v_t_14_10(net968[0:23]),
     .sp12_v_t_13_10(net969[0:23]), .sp12_h_l_13_10(net1319[0:23]),
     .sp12_h_l_13_09(net1320[0:23]), .sp12_h_l_13_08(net1316[0:23]),
     .sp12_h_l_13_07(net1317[0:23]), .sp12_h_l_13_06(net1318[0:23]),
     .sp12_h_l_13_05(net1315[0:23]), .sp12_h_l_13_04(net1311[0:23]),
     .sp12_h_l_13_03(net1314[0:23]), .sp12_h_l_13_02(net1313[0:23]),
     .sp12_h_l_13_01(net1312[0:23]), .sp4_v_t_24_10(net980[0:47]),
     .sp4_v_t_23_10(net981[0:47]), .sp4_v_t_22_10(net982[0:47]),
     .sp4_v_t_21_10(net983[0:47]), .sp4_v_t_20_10(net984[0:47]),
     .sp4_v_t_19_10(net985[0:47]), .sp4_v_t_18_10(net986[0:47]),
     .sp4_v_t_17_10(net987[0:47]), .sp4_v_t_16_10(net988[0:47]),
     .sp4_v_t_15_10(net989[0:47]), .sp4_v_t_14_10(net990[0:47]),
     .sp4_v_t_13_10(net991[0:47]), .sp4_v_b_13_10(net1405[0:47]),
     .sp4_v_b_13_09(net1406[0:47]), .sp4_v_b_13_08(net1407[0:47]),
     .sp4_v_b_13_07(net1408[0:47]), .sp4_v_b_13_06(net1409[0:47]),
     .sp4_v_b_13_05(net1410[0:47]), .sp4_v_b_13_04(net1411[0:47]),
     .sp4_v_b_13_03(net1412[0:47]), .sp4_v_b_13_02(net1413[0:47]),
     .sp4_v_b_13_01(net1414[0:47]), .sp4_h_l_13_10(net1416[0:47]),
     .sp4_h_l_13_09(net1417[0:47]), .sp4_h_l_13_08(net1322[0:47]),
     .sp4_h_l_13_07(net1323[0:47]), .sp4_h_l_13_06(net1418[0:47]),
     .sp4_h_l_13_05(net1419[0:47]), .sp4_h_l_13_04(net1420[0:47]),
     .sp4_h_l_13_03(net1350[0:47]), .sp4_h_l_13_02(net1421[0:47]),
     .sp4_h_l_13_01(net1422[0:47]), .sp4_h_l_13_00(net1299[0:15]),
     .bl({bl_bot[1297], bl_bot[1296], bl_bot[1295], bl_bot[1294],
     bl_bot[1303], bl_bot[1302], bl_bot[1301], bl_bot[1300],
     bl_bot[1299], bl_bot[1298], bl_bot[1309], bl_bot[1308],
     bl_bot[1307], bl_bot[1306], bl_bot[1305], bl_bot[1304],
     bl_bot[1311], bl_bot[1310], bl_bot[1243], bl_bot[1242],
     bl_bot[1241], bl_bot[1240], bl_bot[1253], bl_bot[1252],
     bl_bot[1251], bl_bot[1250], bl_bot[1249], bl_bot[1248],
     bl_bot[1247], bl_bot[1246], bl_bot[1245], bl_bot[1244],
     bl_bot[1265], bl_bot[1264], bl_bot[1263], bl_bot[1262],
     bl_bot[1261], bl_bot[1260], bl_bot[1259], bl_bot[1258],
     bl_bot[1257], bl_bot[1256], bl_bot[1255], bl_bot[1254],
     bl_bot[1293], bl_bot[1292], bl_bot[1291], bl_bot[1290],
     bl_bot[1289], bl_bot[1288], bl_bot[1287], bl_bot[1286],
     bl_bot[1285], bl_bot[1284], bl_bot[1283], bl_bot[1282],
     bl_bot[1281], bl_bot[1280], bl_bot[1279], bl_bot[1278],
     bl_bot[1277], bl_bot[1276], bl_bot[1275], bl_bot[1274],
     bl_bot[1273], bl_bot[1272], bl_bot[1271], bl_bot[1270],
     bl_bot[1269], bl_bot[1268], bl_bot[1267], bl_bot[1266],
     bl_bot[1189], bl_bot[1188], bl_bot[1187], bl_bot[1186],
     bl_bot[1199], bl_bot[1198], bl_bot[1197], bl_bot[1196],
     bl_bot[1195], bl_bot[1194], bl_bot[1193], bl_bot[1192],
     bl_bot[1191], bl_bot[1190], bl_bot[1211], bl_bot[1210],
     bl_bot[1209], bl_bot[1208], bl_bot[1207], bl_bot[1206],
     bl_bot[1205], bl_bot[1204], bl_bot[1203], bl_bot[1202],
     bl_bot[1201], bl_bot[1200], bl_bot[1239], bl_bot[1238],
     bl_bot[1237], bl_bot[1236], bl_bot[1235], bl_bot[1234],
     bl_bot[1233], bl_bot[1232], bl_bot[1231], bl_bot[1230],
     bl_bot[1229], bl_bot[1228], bl_bot[1227], bl_bot[1226],
     bl_bot[1225], bl_bot[1224], bl_bot[1223], bl_bot[1222],
     bl_bot[1221], bl_bot[1220], bl_bot[1219], bl_bot[1218],
     bl_bot[1217], bl_bot[1216], bl_bot[1215], bl_bot[1214],
     bl_bot[1213], bl_bot[1212], bl_bot[1135], bl_bot[1134],
     bl_bot[1133], bl_bot[1132], bl_bot[1145], bl_bot[1144],
     bl_bot[1143], bl_bot[1142], bl_bot[1141], bl_bot[1140],
     bl_bot[1139], bl_bot[1138], bl_bot[1137], bl_bot[1136],
     bl_bot[1157], bl_bot[1156], bl_bot[1155], bl_bot[1154],
     bl_bot[1153], bl_bot[1152], bl_bot[1151], bl_bot[1150],
     bl_bot[1149], bl_bot[1148], bl_bot[1147], bl_bot[1146],
     bl_bot[1185], bl_bot[1184], bl_bot[1183], bl_bot[1182],
     bl_bot[1181], bl_bot[1180], bl_bot[1179], bl_bot[1178],
     bl_bot[1177], bl_bot[1176], bl_bot[1175], bl_bot[1174],
     bl_bot[1173], bl_bot[1172], bl_bot[1171], bl_bot[1170],
     bl_bot[1169], bl_bot[1168], bl_bot[1167], bl_bot[1166],
     bl_bot[1165], bl_bot[1164], bl_bot[1163], bl_bot[1162],
     bl_bot[1161], bl_bot[1160], bl_bot[1159], bl_bot[1158],
     bl_bot[1081], bl_bot[1080], bl_bot[1079], bl_bot[1078],
     bl_bot[1091], bl_bot[1090], bl_bot[1089], bl_bot[1088],
     bl_bot[1087], bl_bot[1086], bl_bot[1085], bl_bot[1084],
     bl_bot[1083], bl_bot[1082], bl_bot[1103], bl_bot[1102],
     bl_bot[1101], bl_bot[1100], bl_bot[1099], bl_bot[1098],
     bl_bot[1097], bl_bot[1096], bl_bot[1095], bl_bot[1094],
     bl_bot[1093], bl_bot[1092], bl_bot[1131], bl_bot[1130],
     bl_bot[1129], bl_bot[1128], bl_bot[1127], bl_bot[1126],
     bl_bot[1125], bl_bot[1124], bl_bot[1123], bl_bot[1122],
     bl_bot[1121], bl_bot[1120], bl_bot[1119], bl_bot[1118],
     bl_bot[1117], bl_bot[1116], bl_bot[1115], bl_bot[1114],
     bl_bot[1113], bl_bot[1112], bl_bot[1111], bl_bot[1110],
     bl_bot[1109], bl_bot[1108], bl_bot[1107], bl_bot[1106],
     bl_bot[1105], bl_bot[1104], bl_bot[1027], bl_bot[1026],
     bl_bot[1025], bl_bot[1024], bl_bot[1037], bl_bot[1036],
     bl_bot[1035], bl_bot[1034], bl_bot[1033], bl_bot[1032],
     bl_bot[1031], bl_bot[1030], bl_bot[1029], bl_bot[1028],
     bl_bot[1049], bl_bot[1048], bl_bot[1047], bl_bot[1046],
     bl_bot[1045], bl_bot[1044], bl_bot[1043], bl_bot[1042],
     bl_bot[1041], bl_bot[1040], bl_bot[1039], bl_bot[1038],
     bl_bot[1077], bl_bot[1076], bl_bot[1075], bl_bot[1074],
     bl_bot[1073], bl_bot[1072], bl_bot[1071], bl_bot[1070],
     bl_bot[1069], bl_bot[1068], bl_bot[1067], bl_bot[1066],
     bl_bot[1065], bl_bot[1064], bl_bot[1063], bl_bot[1062],
     bl_bot[1061], bl_bot[1060], bl_bot[1059], bl_bot[1058],
     bl_bot[1057], bl_bot[1056], bl_bot[1055], bl_bot[1054],
     bl_bot[1053], bl_bot[1052], bl_bot[1051], bl_bot[1050],
     bl_bot[985], bl_bot[984], bl_bot[983], bl_bot[982], bl_bot[995],
     bl_bot[994], bl_bot[993], bl_bot[992], bl_bot[991], bl_bot[990],
     bl_bot[989], bl_bot[988], bl_bot[987], bl_bot[986], bl_bot[1007],
     bl_bot[1006], bl_bot[1005], bl_bot[1004], bl_bot[1003],
     bl_bot[1002], bl_bot[1001], bl_bot[1000], bl_bot[999],
     bl_bot[998], bl_bot[997], bl_bot[996], bl_bot[1023], bl_bot[1022],
     bl_bot[1021], bl_bot[1020], bl_bot[1019], bl_bot[1018],
     bl_bot[1017], bl_bot[1016], bl_bot[1015], bl_bot[1014],
     bl_bot[1013], bl_bot[1012], bl_bot[1011], bl_bot[1010],
     bl_bot[1009], bl_bot[1008], bl_bot[931], bl_bot[930], bl_bot[929],
     bl_bot[928], bl_bot[941], bl_bot[940], bl_bot[939], bl_bot[938],
     bl_bot[937], bl_bot[936], bl_bot[935], bl_bot[934], bl_bot[933],
     bl_bot[932], bl_bot[953], bl_bot[952], bl_bot[951], bl_bot[950],
     bl_bot[949], bl_bot[948], bl_bot[947], bl_bot[946], bl_bot[945],
     bl_bot[944], bl_bot[943], bl_bot[942], bl_bot[981], bl_bot[980],
     bl_bot[979], bl_bot[978], bl_bot[977], bl_bot[976], bl_bot[975],
     bl_bot[974], bl_bot[973], bl_bot[972], bl_bot[971], bl_bot[970],
     bl_bot[969], bl_bot[968], bl_bot[967], bl_bot[966], bl_bot[965],
     bl_bot[964], bl_bot[963], bl_bot[962], bl_bot[961], bl_bot[960],
     bl_bot[959], bl_bot[958], bl_bot[957], bl_bot[956], bl_bot[955],
     bl_bot[954], bl_bot[877], bl_bot[876], bl_bot[875], bl_bot[874],
     bl_bot[887], bl_bot[886], bl_bot[885], bl_bot[884], bl_bot[883],
     bl_bot[882], bl_bot[881], bl_bot[880], bl_bot[879], bl_bot[878],
     bl_bot[899], bl_bot[898], bl_bot[897], bl_bot[896], bl_bot[895],
     bl_bot[894], bl_bot[893], bl_bot[892], bl_bot[891], bl_bot[890],
     bl_bot[889], bl_bot[888], bl_bot[927], bl_bot[926], bl_bot[925],
     bl_bot[924], bl_bot[923], bl_bot[922], bl_bot[921], bl_bot[920],
     bl_bot[919], bl_bot[918], bl_bot[917], bl_bot[916], bl_bot[915],
     bl_bot[914], bl_bot[913], bl_bot[912], bl_bot[911], bl_bot[910],
     bl_bot[909], bl_bot[908], bl_bot[907], bl_bot[906], bl_bot[905],
     bl_bot[904], bl_bot[903], bl_bot[902], bl_bot[901], bl_bot[900],
     bl_bot[823], bl_bot[822], bl_bot[821], bl_bot[820], bl_bot[833],
     bl_bot[832], bl_bot[831], bl_bot[830], bl_bot[829], bl_bot[828],
     bl_bot[827], bl_bot[826], bl_bot[825], bl_bot[824], bl_bot[845],
     bl_bot[844], bl_bot[843], bl_bot[842], bl_bot[841], bl_bot[840],
     bl_bot[839], bl_bot[838], bl_bot[837], bl_bot[836], bl_bot[835],
     bl_bot[834], bl_bot[873], bl_bot[872], bl_bot[871], bl_bot[870],
     bl_bot[869], bl_bot[868], bl_bot[867], bl_bot[866], bl_bot[865],
     bl_bot[864], bl_bot[863], bl_bot[862], bl_bot[861], bl_bot[860],
     bl_bot[859], bl_bot[858], bl_bot[857], bl_bot[856], bl_bot[855],
     bl_bot[854], bl_bot[853], bl_bot[852], bl_bot[851], bl_bot[850],
     bl_bot[849], bl_bot[848], bl_bot[847], bl_bot[846], bl_bot[769],
     bl_bot[768], bl_bot[767], bl_bot[766], bl_bot[779], bl_bot[778],
     bl_bot[777], bl_bot[776], bl_bot[775], bl_bot[774], bl_bot[773],
     bl_bot[772], bl_bot[771], bl_bot[770], bl_bot[791], bl_bot[790],
     bl_bot[789], bl_bot[788], bl_bot[787], bl_bot[786], bl_bot[785],
     bl_bot[784], bl_bot[783], bl_bot[782], bl_bot[781], bl_bot[780],
     bl_bot[819], bl_bot[818], bl_bot[817], bl_bot[816], bl_bot[815],
     bl_bot[814], bl_bot[813], bl_bot[812], bl_bot[811], bl_bot[810],
     bl_bot[809], bl_bot[808], bl_bot[807], bl_bot[806], bl_bot[805],
     bl_bot[804], bl_bot[803], bl_bot[802], bl_bot[801], bl_bot[800],
     bl_bot[799], bl_bot[798], bl_bot[797], bl_bot[796], bl_bot[795],
     bl_bot[794], bl_bot[793], bl_bot[792], bl_bot[715], bl_bot[714],
     bl_bot[713], bl_bot[712], bl_bot[725], bl_bot[724], bl_bot[723],
     bl_bot[722], bl_bot[721], bl_bot[720], bl_bot[719], bl_bot[718],
     bl_bot[717], bl_bot[716], bl_bot[737], bl_bot[736], bl_bot[735],
     bl_bot[734], bl_bot[733], bl_bot[732], bl_bot[731], bl_bot[730],
     bl_bot[729], bl_bot[728], bl_bot[727], bl_bot[726], bl_bot[765],
     bl_bot[764], bl_bot[763], bl_bot[762], bl_bot[761], bl_bot[760],
     bl_bot[759], bl_bot[758], bl_bot[757], bl_bot[756], bl_bot[755],
     bl_bot[754], bl_bot[753], bl_bot[752], bl_bot[751], bl_bot[750],
     bl_bot[749], bl_bot[748], bl_bot[747], bl_bot[746], bl_bot[745],
     bl_bot[744], bl_bot[743], bl_bot[742], bl_bot[741], bl_bot[740],
     bl_bot[739], bl_bot[738], bl_bot[661], bl_bot[660], bl_bot[659],
     bl_bot[658], bl_bot[671], bl_bot[670], bl_bot[669], bl_bot[668],
     bl_bot[667], bl_bot[666], bl_bot[665], bl_bot[664], bl_bot[663],
     bl_bot[662], bl_bot[683], bl_bot[682], bl_bot[681], bl_bot[680],
     bl_bot[679], bl_bot[678], bl_bot[677], bl_bot[676], bl_bot[675],
     bl_bot[674], bl_bot[673], bl_bot[672], bl_bot[711], bl_bot[710],
     bl_bot[709], bl_bot[708], bl_bot[707], bl_bot[706], bl_bot[705],
     bl_bot[704], bl_bot[703], bl_bot[702], bl_bot[701], bl_bot[700],
     bl_bot[699], bl_bot[698], bl_bot[697], bl_bot[696], bl_bot[695],
     bl_bot[694], bl_bot[693], bl_bot[692], bl_bot[691], bl_bot[690],
     bl_bot[689], bl_bot[688], bl_bot[687], bl_bot[686], bl_bot[685],
     bl_bot[684]}), .fabric_out_122(fabric_out_122),
     .carry_out_13_10(net1015), .fabric_out_126(fabric_out_126),
     .sdi(net1361), .purst(purst), .prog(prog), .sdo(net1066),
     .wl({wl_r[174], wl_r[175], wl_r[172], wl_r[173], wl_r[170],
     wl_r[171], wl_r[168], wl_r[169], wl_r[166], wl_r[167], wl_r[164],
     wl_r[165], wl_r[162], wl_r[163], wl_r[160], wl_r[161], wl_r[158],
     wl_r[159], wl_r[156], wl_r[157], wl_r[154], wl_r[155], wl_r[152],
     wl_r[153], wl_r[150], wl_r[151], wl_r[148], wl_r[149], wl_r[146],
     wl_r[147], wl_r[144], wl_r[145], wl_r[142], wl_r[143], wl_r[140],
     wl_r[141], wl_r[138], wl_r[139], wl_r[136], wl_r[137], wl_r[134],
     wl_r[135], wl_r[132], wl_r[133], wl_r[130], wl_r[131], wl_r[128],
     wl_r[129], wl_r[126], wl_r[127], wl_r[124], wl_r[125], wl_r[122],
     wl_r[123], wl_r[120], wl_r[121], wl_r[118], wl_r[119], wl_r[116],
     wl_r[117], wl_r[114], wl_r[115], wl_r[112], wl_r[113], wl_r[110],
     wl_r[111], wl_r[108], wl_r[109], wl_r[106], wl_r[107], wl_r[104],
     wl_r[105], wl_r[102], wl_r[103], wl_r[100], wl_r[101], wl_r[98],
     wl_r[99], wl_r[96], wl_r[97], wl_r[94], wl_r[95], wl_r[92],
     wl_r[93], wl_r[90], wl_r[91], wl_r[88], wl_r[89], wl_r[86],
     wl_r[87], wl_r[84], wl_r[85], wl_r[82], wl_r[83], wl_r[80],
     wl_r[81], wl_r[78], wl_r[79], wl_r[76], wl_r[77], wl_r[74],
     wl_r[75], wl_r[72], wl_r[73], wl_r[70], wl_r[71], wl_r[68],
     wl_r[69], wl_r[66], wl_r[67], wl_r[64], wl_r[65], wl_r[62],
     wl_r[63], wl_r[60], wl_r[61], wl_r[58], wl_r[59], wl_r[56],
     wl_r[57], wl_r[54], wl_r[55], wl_r[52], wl_r[53], wl_r[50],
     wl_r[51], wl_r[48], wl_r[49], wl_r[46], wl_r[47], wl_r[44],
     wl_r[45], wl_r[42], wl_r[43], wl_r[40], wl_r[41], wl_r[38],
     wl_r[39], wl_r[36], wl_r[37], wl_r[34], wl_r[35], wl_r[32],
     wl_r[33], wl_r[30], wl_r[31], wl_r[28], wl_r[29], wl_r[26],
     wl_r[27], wl_r[24], wl_r[25], wl_r[22], wl_r[23], wl_r[20],
     wl_r[21], wl_r[18], wl_r[19], wl_r[16], wl_r[17], wl_r[0],
     wl_r[1], wl_r[3], wl_r[2], wl_r[4], wl_r[5], wl_r[7], wl_r[6],
     wl_r[8], wl_r[9], wl_r[11], wl_r[10], wl_r[12], wl_r[13],
     wl_r[15], wl_r[14]}), .reset_b({reset_b_r[174], reset_b_r[175],
     reset_b_r[172], reset_b_r[173], reset_b_r[170], reset_b_r[171],
     reset_b_r[168], reset_b_r[169], reset_b_r[166], reset_b_r[167],
     reset_b_r[164], reset_b_r[165], reset_b_r[162], reset_b_r[163],
     reset_b_r[160], reset_b_r[161], reset_b_r[158], reset_b_r[159],
     reset_b_r[156], reset_b_r[157], reset_b_r[154], reset_b_r[155],
     reset_b_r[152], reset_b_r[153], reset_b_r[150], reset_b_r[151],
     reset_b_r[148], reset_b_r[149], reset_b_r[146], reset_b_r[147],
     reset_b_r[144], reset_b_r[145], reset_b_r[142], reset_b_r[143],
     reset_b_r[140], reset_b_r[141], reset_b_r[138], reset_b_r[139],
     reset_b_r[136], reset_b_r[137], reset_b_r[134], reset_b_r[135],
     reset_b_r[132], reset_b_r[133], reset_b_r[130], reset_b_r[131],
     reset_b_r[128], reset_b_r[129], reset_b_r[126], reset_b_r[127],
     reset_b_r[124], reset_b_r[125], reset_b_r[122], reset_b_r[123],
     reset_b_r[120], reset_b_r[121], reset_b_r[118], reset_b_r[119],
     reset_b_r[116], reset_b_r[117], reset_b_r[114], reset_b_r[115],
     reset_b_r[112], reset_b_r[113], reset_b_r[110], reset_b_r[111],
     reset_b_r[108], reset_b_r[109], reset_b_r[106], reset_b_r[107],
     reset_b_r[104], reset_b_r[105], reset_b_r[102], reset_b_r[103],
     reset_b_r[100], reset_b_r[101], reset_b_r[98], reset_b_r[99],
     reset_b_r[96], reset_b_r[97], reset_b_r[94], reset_b_r[95],
     reset_b_r[92], reset_b_r[93], reset_b_r[90], reset_b_r[91],
     reset_b_r[88], reset_b_r[89], reset_b_r[86], reset_b_r[87],
     reset_b_r[84], reset_b_r[85], reset_b_r[82], reset_b_r[83],
     reset_b_r[80], reset_b_r[81], reset_b_r[78], reset_b_r[79],
     reset_b_r[76], reset_b_r[77], reset_b_r[74], reset_b_r[75],
     reset_b_r[72], reset_b_r[73], reset_b_r[70], reset_b_r[71],
     reset_b_r[68], reset_b_r[69], reset_b_r[66], reset_b_r[67],
     reset_b_r[64], reset_b_r[65], reset_b_r[62], reset_b_r[63],
     reset_b_r[60], reset_b_r[61], reset_b_r[58], reset_b_r[59],
     reset_b_r[56], reset_b_r[57], reset_b_r[54], reset_b_r[55],
     reset_b_r[52], reset_b_r[53], reset_b_r[50], reset_b_r[51],
     reset_b_r[48], reset_b_r[49], reset_b_r[46], reset_b_r[47],
     reset_b_r[44], reset_b_r[45], reset_b_r[42], reset_b_r[43],
     reset_b_r[40], reset_b_r[41], reset_b_r[38], reset_b_r[39],
     reset_b_r[36], reset_b_r[37], reset_b_r[34], reset_b_r[35],
     reset_b_r[32], reset_b_r[33], reset_b_r[30], reset_b_r[31],
     reset_b_r[28], reset_b_r[29], reset_b_r[26], reset_b_r[27],
     reset_b_r[24], reset_b_r[25], reset_b_r[22], reset_b_r[23],
     reset_b_r[20], reset_b_r[21], reset_b_r[18], reset_b_r[19],
     reset_b_r[16], reset_b_r[17], reset_b_r[0], reset_b_r[1],
     reset_b_r[3], reset_b_r[2], reset_b_r[4], reset_b_r[5],
     reset_b_r[7], reset_b_r[6], reset_b_r[8], reset_b_r[9],
     reset_b_r[11], reset_b_r[10], reset_b_r[12], reset_b_r[13],
     reset_b_r[15], reset_b_r[14]}), .pgate({pgate_r[174],
     pgate_r[175], pgate_r[172], pgate_r[173], pgate_r[170],
     pgate_r[171], pgate_r[168], pgate_r[169], pgate_r[166],
     pgate_r[167], pgate_r[164], pgate_r[165], pgate_r[162],
     pgate_r[163], pgate_r[160], pgate_r[161], pgate_r[158],
     pgate_r[159], pgate_r[156], pgate_r[157], pgate_r[154],
     pgate_r[155], pgate_r[152], pgate_r[153], pgate_r[150],
     pgate_r[151], pgate_r[148], pgate_r[149], pgate_r[146],
     pgate_r[147], pgate_r[144], pgate_r[145], pgate_r[142],
     pgate_r[143], pgate_r[140], pgate_r[141], pgate_r[138],
     pgate_r[139], pgate_r[136], pgate_r[137], pgate_r[134],
     pgate_r[135], pgate_r[132], pgate_r[133], pgate_r[130],
     pgate_r[131], pgate_r[128], pgate_r[129], pgate_r[126],
     pgate_r[127], pgate_r[124], pgate_r[125], pgate_r[122],
     pgate_r[123], pgate_r[120], pgate_r[121], pgate_r[118],
     pgate_r[119], pgate_r[116], pgate_r[117], pgate_r[114],
     pgate_r[115], pgate_r[112], pgate_r[113], pgate_r[110],
     pgate_r[111], pgate_r[108], pgate_r[109], pgate_r[106],
     pgate_r[107], pgate_r[104], pgate_r[105], pgate_r[102],
     pgate_r[103], pgate_r[100], pgate_r[101], pgate_r[98],
     pgate_r[99], pgate_r[96], pgate_r[97], pgate_r[94], pgate_r[95],
     pgate_r[92], pgate_r[93], pgate_r[90], pgate_r[91], pgate_r[88],
     pgate_r[89], pgate_r[86], pgate_r[87], pgate_r[84], pgate_r[85],
     pgate_r[82], pgate_r[83], pgate_r[80], pgate_r[81], pgate_r[78],
     pgate_r[79], pgate_r[76], pgate_r[77], pgate_r[74], pgate_r[75],
     pgate_r[72], pgate_r[73], pgate_r[70], pgate_r[71], pgate_r[68],
     pgate_r[69], pgate_r[66], pgate_r[67], pgate_r[64], pgate_r[65],
     pgate_r[62], pgate_r[63], pgate_r[60], pgate_r[61], pgate_r[58],
     pgate_r[59], pgate_r[56], pgate_r[57], pgate_r[54], pgate_r[55],
     pgate_r[52], pgate_r[53], pgate_r[50], pgate_r[51], pgate_r[48],
     pgate_r[49], pgate_r[46], pgate_r[47], pgate_r[44], pgate_r[45],
     pgate_r[42], pgate_r[43], pgate_r[40], pgate_r[41], pgate_r[38],
     pgate_r[39], pgate_r[36], pgate_r[37], pgate_r[34], pgate_r[35],
     pgate_r[32], pgate_r[33], pgate_r[30], pgate_r[31], pgate_r[28],
     pgate_r[29], pgate_r[26], pgate_r[27], pgate_r[24], pgate_r[25],
     pgate_r[22], pgate_r[23], pgate_r[20], pgate_r[21], pgate_r[18],
     pgate_r[19], pgate_r[16], pgate_r[17], pgate_r[0], pgate_r[1],
     pgate_r[3], pgate_r[2], pgate_r[4], pgate_r[5], pgate_r[7],
     pgate_r[6], pgate_r[8], pgate_r[9], pgate_r[11], pgate_r[10],
     pgate_r[12], pgate_r[13], pgate_r[15], pgate_r[14]}));
QUAD_TR I_TR ( .ceb_i(net01027), .ceb_o(net01435),
     .io_r_00_24_11(net1024[0:3]), .tnl_op_13_20(slf_op_12_21[3:0]),
     .bnl_op_25_11(net1027[0:7]), .bnr_op_23_11(net1027[0:7]),
     .bnr_op_22_11(net1028[0:7]), .bnr_op_21_11(net1029[0:7]),
     .bnr_op_20_11(net1030[0:7]), .bnr_op_19_11(net1031[0:7]),
     .bnr_op_18_11(net1032[0:7]), .bnr_op_17_11(net1033[0:7]),
     .bnr_op_16_11(net1034[0:7]), .bnr_op_15_11(net1035[0:7]),
     .bnr_op_14_11(net1036[0:7]), .bnr_op_13_11(net1037[0:7]),
     .bnl_op_24_11(net1028[0:7]), .bnl_op_23_11(net1029[0:7]),
     .bnl_op_22_11(net1030[0:7]), .bnl_op_21_11(net1031[0:7]),
     .bnl_op_20_11(net1032[0:7]), .bnl_op_19_11(net1033[0:7]),
     .bnl_op_18_11(net1034[0:7]), .bnl_op_17_11(net1035[0:7]),
     .bnl_op_16_11(net1036[0:7]), .bnl_op_15_11(net1037[0:7]),
     .bnl_op_14_11(net1548[0:7]), .hiz_b_i(net832), .bs_en_i(net833),
     .shift_i(net846), .r_i(net834), .tclk_i(net837),
     .update_i(net835), .mode_i(net836), .mode_o(net1459),
     .shift_o(net1460), .update_o(net1461), .hiz_b_o(net1462),
     .r_o(net1463), .bs_en_o(net1464), .tclk_o(net1465),
     .tiegnd(tiegnd), .tievdd(tievdd), .wl({wl_r[351], wl_r[350],
     wl_r[348], wl_r[349], wl_r[347], wl_r[346], wl_r[344], wl_r[345],
     wl_r[343], wl_r[342], wl_r[340], wl_r[341], wl_r[339], wl_r[338],
     wl_r[336], wl_r[337], wl_r[334], wl_r[335], wl_r[332], wl_r[333],
     wl_r[330], wl_r[331], wl_r[328], wl_r[329], wl_r[326], wl_r[327],
     wl_r[324], wl_r[325], wl_r[322], wl_r[323], wl_r[320], wl_r[321],
     wl_r[318], wl_r[319], wl_r[316], wl_r[317], wl_r[314], wl_r[315],
     wl_r[312], wl_r[313], wl_r[310], wl_r[311], wl_r[308], wl_r[309],
     wl_r[306], wl_r[307], wl_r[304], wl_r[305], wl_r[302], wl_r[303],
     wl_r[300], wl_r[301], wl_r[298], wl_r[299], wl_r[296], wl_r[297],
     wl_r[294], wl_r[295], wl_r[292], wl_r[293], wl_r[290], wl_r[291],
     wl_r[288], wl_r[289], wl_r[286], wl_r[287], wl_r[284], wl_r[285],
     wl_r[282], wl_r[283], wl_r[280], wl_r[281], wl_r[278], wl_r[279],
     wl_r[276], wl_r[277], wl_r[274], wl_r[275], wl_r[272], wl_r[273],
     wl_r[270], wl_r[271], wl_r[268], wl_r[269], wl_r[266], wl_r[267],
     wl_r[264], wl_r[265], wl_r[262], wl_r[263], wl_r[260], wl_r[261],
     wl_r[258], wl_r[259], wl_r[256], wl_r[257], wl_r[254], wl_r[255],
     wl_r[252], wl_r[253], wl_r[250], wl_r[251], wl_r[248], wl_r[249],
     wl_r[246], wl_r[247], wl_r[244], wl_r[245], wl_r[242], wl_r[243],
     wl_r[240], wl_r[241], wl_r[238], wl_r[239], wl_r[236], wl_r[237],
     wl_r[234], wl_r[235], wl_r[232], wl_r[233], wl_r[230], wl_r[231],
     wl_r[228], wl_r[229], wl_r[226], wl_r[227], wl_r[224], wl_r[225],
     wl_r[222], wl_r[223], wl_r[220], wl_r[221], wl_r[218], wl_r[219],
     wl_r[216], wl_r[217], wl_r[214], wl_r[215], wl_r[212], wl_r[213],
     wl_r[210], wl_r[211], wl_r[208], wl_r[209], wl_r[206], wl_r[207],
     wl_r[204], wl_r[205], wl_r[202], wl_r[203], wl_r[200], wl_r[201],
     wl_r[198], wl_r[199], wl_r[196], wl_r[197], wl_r[194], wl_r[195],
     wl_r[192], wl_r[193], wl_r[190], wl_r[191], wl_r[188], wl_r[189],
     wl_r[186], wl_r[187], wl_r[184], wl_r[185], wl_r[182], wl_r[183],
     wl_r[180], wl_r[181], wl_r[178], wl_r[179], wl_r[176],
     wl_r[177]}), .sdi(net1066), .reset_b({reset_b_r[351],
     reset_b_r[350], reset_b_r[348], reset_b_r[349], reset_b_r[347],
     reset_b_r[346], reset_b_r[344], reset_b_r[345], reset_b_r[343],
     reset_b_r[342], reset_b_r[340], reset_b_r[341], reset_b_r[339],
     reset_b_r[338], reset_b_r[336], reset_b_r[337], reset_b_r[334],
     reset_b_r[335], reset_b_r[332], reset_b_r[333], reset_b_r[330],
     reset_b_r[331], reset_b_r[328], reset_b_r[329], reset_b_r[326],
     reset_b_r[327], reset_b_r[324], reset_b_r[325], reset_b_r[322],
     reset_b_r[323], reset_b_r[320], reset_b_r[321], reset_b_r[318],
     reset_b_r[319], reset_b_r[316], reset_b_r[317], reset_b_r[314],
     reset_b_r[315], reset_b_r[312], reset_b_r[313], reset_b_r[310],
     reset_b_r[311], reset_b_r[308], reset_b_r[309], reset_b_r[306],
     reset_b_r[307], reset_b_r[304], reset_b_r[305], reset_b_r[302],
     reset_b_r[303], reset_b_r[300], reset_b_r[301], reset_b_r[298],
     reset_b_r[299], reset_b_r[296], reset_b_r[297], reset_b_r[294],
     reset_b_r[295], reset_b_r[292], reset_b_r[293], reset_b_r[290],
     reset_b_r[291], reset_b_r[288], reset_b_r[289], reset_b_r[286],
     reset_b_r[287], reset_b_r[284], reset_b_r[285], reset_b_r[282],
     reset_b_r[283], reset_b_r[280], reset_b_r[281], reset_b_r[278],
     reset_b_r[279], reset_b_r[276], reset_b_r[277], reset_b_r[274],
     reset_b_r[275], reset_b_r[272], reset_b_r[273], reset_b_r[270],
     reset_b_r[271], reset_b_r[268], reset_b_r[269], reset_b_r[266],
     reset_b_r[267], reset_b_r[264], reset_b_r[265], reset_b_r[262],
     reset_b_r[263], reset_b_r[260], reset_b_r[261], reset_b_r[258],
     reset_b_r[259], reset_b_r[256], reset_b_r[257], reset_b_r[254],
     reset_b_r[255], reset_b_r[252], reset_b_r[253], reset_b_r[250],
     reset_b_r[251], reset_b_r[248], reset_b_r[249], reset_b_r[246],
     reset_b_r[247], reset_b_r[244], reset_b_r[245], reset_b_r[242],
     reset_b_r[243], reset_b_r[240], reset_b_r[241], reset_b_r[238],
     reset_b_r[239], reset_b_r[236], reset_b_r[237], reset_b_r[234],
     reset_b_r[235], reset_b_r[232], reset_b_r[233], reset_b_r[230],
     reset_b_r[231], reset_b_r[228], reset_b_r[229], reset_b_r[226],
     reset_b_r[227], reset_b_r[224], reset_b_r[225], reset_b_r[222],
     reset_b_r[223], reset_b_r[220], reset_b_r[221], reset_b_r[218],
     reset_b_r[219], reset_b_r[216], reset_b_r[217], reset_b_r[214],
     reset_b_r[215], reset_b_r[212], reset_b_r[213], reset_b_r[210],
     reset_b_r[211], reset_b_r[208], reset_b_r[209], reset_b_r[206],
     reset_b_r[207], reset_b_r[204], reset_b_r[205], reset_b_r[202],
     reset_b_r[203], reset_b_r[200], reset_b_r[201], reset_b_r[198],
     reset_b_r[199], reset_b_r[196], reset_b_r[197], reset_b_r[194],
     reset_b_r[195], reset_b_r[192], reset_b_r[193], reset_b_r[190],
     reset_b_r[191], reset_b_r[188], reset_b_r[189], reset_b_r[186],
     reset_b_r[187], reset_b_r[184], reset_b_r[185], reset_b_r[182],
     reset_b_r[183], reset_b_r[180], reset_b_r[181], reset_b_r[178],
     reset_b_r[179], reset_b_r[176], reset_b_r[177]}), .purst(purst),
     .prog(prog), .pgate({pgate_r[351], pgate_r[350], pgate_r[348],
     pgate_r[349], pgate_r[347], pgate_r[346], pgate_r[344],
     pgate_r[345], pgate_r[343], pgate_r[342], pgate_r[340],
     pgate_r[341], pgate_r[339], pgate_r[338], pgate_r[336],
     pgate_r[337], pgate_r[334], pgate_r[335], pgate_r[332],
     pgate_r[333], pgate_r[330], pgate_r[331], pgate_r[328],
     pgate_r[329], pgate_r[326], pgate_r[327], pgate_r[324],
     pgate_r[325], pgate_r[322], pgate_r[323], pgate_r[320],
     pgate_r[321], pgate_r[318], pgate_r[319], pgate_r[316],
     pgate_r[317], pgate_r[314], pgate_r[315], pgate_r[312],
     pgate_r[313], pgate_r[310], pgate_r[311], pgate_r[308],
     pgate_r[309], pgate_r[306], pgate_r[307], pgate_r[304],
     pgate_r[305], pgate_r[302], pgate_r[303], pgate_r[300],
     pgate_r[301], pgate_r[298], pgate_r[299], pgate_r[296],
     pgate_r[297], pgate_r[294], pgate_r[295], pgate_r[292],
     pgate_r[293], pgate_r[290], pgate_r[291], pgate_r[288],
     pgate_r[289], pgate_r[286], pgate_r[287], pgate_r[284],
     pgate_r[285], pgate_r[282], pgate_r[283], pgate_r[280],
     pgate_r[281], pgate_r[278], pgate_r[279], pgate_r[276],
     pgate_r[277], pgate_r[274], pgate_r[275], pgate_r[272],
     pgate_r[273], pgate_r[270], pgate_r[271], pgate_r[268],
     pgate_r[269], pgate_r[266], pgate_r[267], pgate_r[264],
     pgate_r[265], pgate_r[262], pgate_r[263], pgate_r[260],
     pgate_r[261], pgate_r[258], pgate_r[259], pgate_r[256],
     pgate_r[257], pgate_r[254], pgate_r[255], pgate_r[252],
     pgate_r[253], pgate_r[250], pgate_r[251], pgate_r[248],
     pgate_r[249], pgate_r[246], pgate_r[247], pgate_r[244],
     pgate_r[245], pgate_r[242], pgate_r[243], pgate_r[240],
     pgate_r[241], pgate_r[238], pgate_r[239], pgate_r[236],
     pgate_r[237], pgate_r[234], pgate_r[235], pgate_r[232],
     pgate_r[233], pgate_r[230], pgate_r[231], pgate_r[228],
     pgate_r[229], pgate_r[226], pgate_r[227], pgate_r[224],
     pgate_r[225], pgate_r[222], pgate_r[223], pgate_r[220],
     pgate_r[221], pgate_r[218], pgate_r[219], pgate_r[216],
     pgate_r[217], pgate_r[214], pgate_r[215], pgate_r[212],
     pgate_r[213], pgate_r[210], pgate_r[211], pgate_r[208],
     pgate_r[209], pgate_r[206], pgate_r[207], pgate_r[204],
     pgate_r[205], pgate_r[202], pgate_r[203], pgate_r[200],
     pgate_r[201], pgate_r[198], pgate_r[199], pgate_r[196],
     pgate_r[197], pgate_r[194], pgate_r[195], pgate_r[192],
     pgate_r[193], pgate_r[190], pgate_r[191], pgate_r[188],
     pgate_r[189], pgate_r[186], pgate_r[187], pgate_r[184],
     pgate_r[185], pgate_r[182], pgate_r[183], pgate_r[180],
     pgate_r[181], pgate_r[178], pgate_r[179], pgate_r[176],
     pgate_r[177]}), .padin_r(padin_r[39:20]),
     .sp4_h_l_13_21(net1508[0:15]), .sp4_v_b_25_11(net884[0:15]),
     .lft_op_13_10(net1551[0:7]), .lft_op_13_09(net1552[0:7]),
     .lft_op_13_08(net1553[0:7]), .lft_op_13_07(net1554[0:7]),
     .lft_op_13_06(net1555[0:7]), .lft_op_13_05(net1556[0:7]),
     .lft_op_13_04(net1557[0:7]), .lft_op_13_03(net1558[0:7]),
     .lft_op_13_02(net1559[0:7]), .lft_op_13_01(net1415[0:7]),
     .carry_in_24_11(net948), .carry_in_23_11(net949),
     .carry_in_22_11(net950), .carry_in_21_11(net951),
     .carry_in_20_11(net952), .carry_in_18_11(net953),
     .carry_in_17_11(net955), .carry_in_16_11(net956),
     .carry_in_15_11(net954), .carry_in_14_11(net957),
     .carry_in_13_11(net1015), .bot_op_24_11(net1027[0:7]),
     .bot_op_23_11(net1028[0:7]), .bot_op_22_11(net1029[0:7]),
     .bot_op_21_11(net1030[0:7]), .bot_op_20_11(net1031[0:7]),
     .bot_op_19_11(net1032[0:7]), .bot_op_18_11(net1033[0:7]),
     .bot_op_17_11(net1034[0:7]), .bot_op_16_11(net1035[0:7]),
     .bot_op_15_11(net1036[0:7]), .bot_op_14_11(net1037[0:7]),
     .bot_op_13_11(net1548[0:7]), .bnr_op_24_11({slf_op_25_10[3],
     slf_op_25_10[2], slf_op_25_10[1], slf_op_25_10[0],
     slf_op_25_10[3], slf_op_25_10[2], slf_op_25_10[1],
     slf_op_25_10[0]}), .bnl_op_13_11(net1537[0:7]),
     .spi_ss_in_r(spi_ss_in_r[39:20]), .slf_op_24_11(net810[0:7]),
     .slf_op_23_11(net809[0:7]), .slf_op_22_11(net819[0:7]),
     .slf_op_21_11(net820[0:7]), .slf_op_20_11(net811[0:7]),
     .slf_op_19_11(net812[0:7]), .slf_op_18_11(net813[0:7]),
     .slf_op_17_11(net814[0:7]), .slf_op_16_11(net815[0:7]),
     .slf_op_15_11(net816[0:7]), .slf_op_14_11(net817[0:7]),
     .slf_op_13_11(net1310[0:7]), .slf_op_13_10(net1514[0:7]),
     .slf_op_13_09(net1515[0:7]), .slf_op_13_08(net1516[0:7]),
     .slf_op_13_07(net1517[0:7]), .slf_op_13_06(net1518[0:7]),
     .slf_op_13_05(net1519[0:7]), .slf_op_13_04(net1520[0:7]),
     .slf_op_13_03(net1521[0:7]), .slf_op_13_02(net1522[0:7]),
     .sdo(net1623), .pado_r(pado_r[39:20]), .padeb_r(padeb_r[39:20]),
     .vdd_cntl({vdd_cntl_r[351], vdd_cntl_r[350], vdd_cntl_r[348],
     vdd_cntl_r[349], vdd_cntl_r[347], vdd_cntl_r[346],
     vdd_cntl_r[344], vdd_cntl_r[345], vdd_cntl_r[343],
     vdd_cntl_r[342], vdd_cntl_r[340], vdd_cntl_r[341],
     vdd_cntl_r[339], vdd_cntl_r[338], vdd_cntl_r[336],
     vdd_cntl_r[337], vdd_cntl_r[334], vdd_cntl_r[335],
     vdd_cntl_r[332], vdd_cntl_r[333], vdd_cntl_r[330],
     vdd_cntl_r[331], vdd_cntl_r[328], vdd_cntl_r[329],
     vdd_cntl_r[326], vdd_cntl_r[327], vdd_cntl_r[324],
     vdd_cntl_r[325], vdd_cntl_r[322], vdd_cntl_r[323],
     vdd_cntl_r[320], vdd_cntl_r[321], vdd_cntl_r[318],
     vdd_cntl_r[319], vdd_cntl_r[316], vdd_cntl_r[317],
     vdd_cntl_r[314], vdd_cntl_r[315], vdd_cntl_r[312],
     vdd_cntl_r[313], vdd_cntl_r[310], vdd_cntl_r[311],
     vdd_cntl_r[308], vdd_cntl_r[309], vdd_cntl_r[306],
     vdd_cntl_r[307], vdd_cntl_r[304], vdd_cntl_r[305],
     vdd_cntl_r[302], vdd_cntl_r[303], vdd_cntl_r[300],
     vdd_cntl_r[301], vdd_cntl_r[298], vdd_cntl_r[299],
     vdd_cntl_r[296], vdd_cntl_r[297], vdd_cntl_r[294],
     vdd_cntl_r[295], vdd_cntl_r[292], vdd_cntl_r[293],
     vdd_cntl_r[290], vdd_cntl_r[291], vdd_cntl_r[288],
     vdd_cntl_r[289], vdd_cntl_r[286], vdd_cntl_r[287],
     vdd_cntl_r[284], vdd_cntl_r[285], vdd_cntl_r[282],
     vdd_cntl_r[283], vdd_cntl_r[280], vdd_cntl_r[281],
     vdd_cntl_r[278], vdd_cntl_r[279], vdd_cntl_r[276],
     vdd_cntl_r[277], vdd_cntl_r[274], vdd_cntl_r[275],
     vdd_cntl_r[272], vdd_cntl_r[273], vdd_cntl_r[270],
     vdd_cntl_r[271], vdd_cntl_r[268], vdd_cntl_r[269],
     vdd_cntl_r[266], vdd_cntl_r[267], vdd_cntl_r[264],
     vdd_cntl_r[265], vdd_cntl_r[262], vdd_cntl_r[263],
     vdd_cntl_r[260], vdd_cntl_r[261], vdd_cntl_r[258],
     vdd_cntl_r[259], vdd_cntl_r[256], vdd_cntl_r[257],
     vdd_cntl_r[254], vdd_cntl_r[255], vdd_cntl_r[252],
     vdd_cntl_r[253], vdd_cntl_r[250], vdd_cntl_r[251],
     vdd_cntl_r[248], vdd_cntl_r[249], vdd_cntl_r[246],
     vdd_cntl_r[247], vdd_cntl_r[244], vdd_cntl_r[245],
     vdd_cntl_r[242], vdd_cntl_r[243], vdd_cntl_r[240],
     vdd_cntl_r[241], vdd_cntl_r[238], vdd_cntl_r[239],
     vdd_cntl_r[236], vdd_cntl_r[237], vdd_cntl_r[234],
     vdd_cntl_r[235], vdd_cntl_r[232], vdd_cntl_r[233],
     vdd_cntl_r[230], vdd_cntl_r[231], vdd_cntl_r[228],
     vdd_cntl_r[229], vdd_cntl_r[226], vdd_cntl_r[227],
     vdd_cntl_r[224], vdd_cntl_r[225], vdd_cntl_r[222],
     vdd_cntl_r[223], vdd_cntl_r[220], vdd_cntl_r[221],
     vdd_cntl_r[218], vdd_cntl_r[219], vdd_cntl_r[216],
     vdd_cntl_r[217], vdd_cntl_r[214], vdd_cntl_r[215],
     vdd_cntl_r[212], vdd_cntl_r[213], vdd_cntl_r[210],
     vdd_cntl_r[211], vdd_cntl_r[208], vdd_cntl_r[209],
     vdd_cntl_r[206], vdd_cntl_r[207], vdd_cntl_r[204],
     vdd_cntl_r[205], vdd_cntl_r[202], vdd_cntl_r[203],
     vdd_cntl_r[200], vdd_cntl_r[201], vdd_cntl_r[198],
     vdd_cntl_r[199], vdd_cntl_r[196], vdd_cntl_r[197],
     vdd_cntl_r[194], vdd_cntl_r[195], vdd_cntl_r[192],
     vdd_cntl_r[193], vdd_cntl_r[190], vdd_cntl_r[191],
     vdd_cntl_r[188], vdd_cntl_r[189], vdd_cntl_r[186],
     vdd_cntl_r[187], vdd_cntl_r[184], vdd_cntl_r[185],
     vdd_cntl_r[182], vdd_cntl_r[183], vdd_cntl_r[180],
     vdd_cntl_r[181], vdd_cntl_r[178], vdd_cntl_r[179],
     vdd_cntl_r[176], vdd_cntl_r[177]}),
     .slf_op_13_21(slf_op_13_21[3:0]), .fabric_out_223(fabric_out_223),
     .fabric_out_168(bank_cntl_right), .fabric_out_163(fabric_out_163),
     .sp12_v_b_24_11(net958[0:23]), .sp12_v_b_23_11(net959[0:23]),
     .sp12_v_b_22_11(net960[0:23]), .sp12_v_b_21_11(net961[0:23]),
     .sp12_v_b_20_11(net962[0:23]), .sp12_v_b_19_11(net963[0:23]),
     .sp12_v_b_18_11(net964[0:23]), .sp12_v_b_17_11(net965[0:23]),
     .sp12_v_b_16_11(net966[0:23]), .sp12_v_b_15_11(net967[0:23]),
     .sp12_v_b_14_11(net968[0:23]), .sp12_v_b_13_11(net969[0:23]),
     .sp12_h_l_13_10(net1501[0:23]), .sp12_h_l_13_09(net1502[0:23]),
     .sp12_h_l_13_08(net1503[0:23]), .sp12_h_l_13_07(net1504[0:23]),
     .sp12_h_l_13_06(net1505[0:23]), .sp12_h_l_13_05(net1506[0:23]),
     .sp12_h_l_13_04(net1507[0:23]), .sp12_h_l_13_03(net1498[0:23]),
     .sp12_h_l_13_02(net1500[0:23]), .sp12_h_l_13_01(net1499[0:23]),
     .sp4_v_b_24_11(net980[0:47]), .sp4_v_b_23_11(net981[0:47]),
     .sp4_v_b_22_11(net982[0:47]), .sp4_v_b_21_11(net983[0:47]),
     .sp4_v_b_20_11(net984[0:47]), .sp4_v_b_19_11(net985[0:47]),
     .sp4_v_b_18_11(net986[0:47]), .sp4_v_b_17_11(net987[0:47]),
     .sp4_v_b_16_11(net988[0:47]), .sp4_v_b_15_11(net989[0:47]),
     .sp4_v_b_14_11(net990[0:47]), .sp4_v_b_13_11(net991[0:47]),
     .sp4_v_b_13_10(net1599[0:47]), .sp4_v_b_13_09(net1600[0:47]),
     .sp4_v_b_13_08(net1601[0:47]), .sp4_v_b_13_07(net1602[0:47]),
     .sp4_v_b_13_06(net1603[0:47]), .sp4_v_b_13_05(net1604[0:47]),
     .sp4_v_b_13_04(net1605[0:47]), .sp4_v_b_13_03(net1606[0:47]),
     .sp4_v_b_13_02(net1607[0:47]), .sp4_h_l_13_10(net1609[0:47]),
     .sp4_h_l_13_09(net1610[0:47]), .sp4_h_l_13_08(net1611[0:47]),
     .sp4_h_l_13_07(net1612[0:47]), .sp4_h_l_13_06(net1613[0:47]),
     .sp4_h_l_13_05(net1614[0:47]), .sp4_h_l_13_04(net1615[0:47]),
     .sp4_h_l_13_03(net1616[0:47]), .sp4_h_l_13_02(net1617[0:47]),
     .sp4_h_l_13_01(net1618[0:47]), .bl({bl_top[1297], bl_top[1296],
     bl_top[1295], bl_top[1294], bl_top[1303], bl_top[1302],
     bl_top[1301], bl_top[1300], bl_top[1299], bl_top[1298],
     bl_top[1309], bl_top[1308], bl_top[1307], bl_top[1306],
     bl_top[1305], bl_top[1304], bl_top[1311], bl_top[1310],
     bl_top[1243], bl_top[1242], bl_top[1241], bl_top[1240],
     bl_top[1253], bl_top[1252], bl_top[1251], bl_top[1250],
     bl_top[1249], bl_top[1248], bl_top[1247], bl_top[1246],
     bl_top[1245], bl_top[1244], bl_top[1265], bl_top[1264],
     bl_top[1263], bl_top[1262], bl_top[1261], bl_top[1260],
     bl_top[1259], bl_top[1258], bl_top[1257], bl_top[1256],
     bl_top[1255], bl_top[1254], bl_top[1293], bl_top[1292],
     bl_top[1291], bl_top[1290], bl_top[1289], bl_top[1288],
     bl_top[1287], bl_top[1286], bl_top[1285], bl_top[1284],
     bl_top[1283], bl_top[1282], bl_top[1281], bl_top[1280],
     bl_top[1279], bl_top[1278], bl_top[1277], bl_top[1276],
     bl_top[1275], bl_top[1274], bl_top[1273], bl_top[1272],
     bl_top[1271], bl_top[1270], bl_top[1269], bl_top[1268],
     bl_top[1267], bl_top[1266], bl_top[1189], bl_top[1188],
     bl_top[1187], bl_top[1186], bl_top[1199], bl_top[1198],
     bl_top[1197], bl_top[1196], bl_top[1195], bl_top[1194],
     bl_top[1193], bl_top[1192], bl_top[1191], bl_top[1190],
     bl_top[1211], bl_top[1210], bl_top[1209], bl_top[1208],
     bl_top[1207], bl_top[1206], bl_top[1205], bl_top[1204],
     bl_top[1203], bl_top[1202], bl_top[1201], bl_top[1200],
     bl_top[1239], bl_top[1238], bl_top[1237], bl_top[1236],
     bl_top[1235], bl_top[1234], bl_top[1233], bl_top[1232],
     bl_top[1231], bl_top[1230], bl_top[1229], bl_top[1228],
     bl_top[1227], bl_top[1226], bl_top[1225], bl_top[1224],
     bl_top[1223], bl_top[1222], bl_top[1221], bl_top[1220],
     bl_top[1219], bl_top[1218], bl_top[1217], bl_top[1216],
     bl_top[1215], bl_top[1214], bl_top[1213], bl_top[1212],
     bl_top[1135], bl_top[1134], bl_top[1133], bl_top[1132],
     bl_top[1145], bl_top[1144], bl_top[1143], bl_top[1142],
     bl_top[1141], bl_top[1140], bl_top[1139], bl_top[1138],
     bl_top[1137], bl_top[1136], bl_top[1157], bl_top[1156],
     bl_top[1155], bl_top[1154], bl_top[1153], bl_top[1152],
     bl_top[1151], bl_top[1150], bl_top[1149], bl_top[1148],
     bl_top[1147], bl_top[1146], bl_top[1185], bl_top[1184],
     bl_top[1183], bl_top[1182], bl_top[1181], bl_top[1180],
     bl_top[1179], bl_top[1178], bl_top[1177], bl_top[1176],
     bl_top[1175], bl_top[1174], bl_top[1173], bl_top[1172],
     bl_top[1171], bl_top[1170], bl_top[1169], bl_top[1168],
     bl_top[1167], bl_top[1166], bl_top[1165], bl_top[1164],
     bl_top[1163], bl_top[1162], bl_top[1161], bl_top[1160],
     bl_top[1159], bl_top[1158], bl_top[1081], bl_top[1080],
     bl_top[1079], bl_top[1078], bl_top[1091], bl_top[1090],
     bl_top[1089], bl_top[1088], bl_top[1087], bl_top[1086],
     bl_top[1085], bl_top[1084], bl_top[1083], bl_top[1082],
     bl_top[1103], bl_top[1102], bl_top[1101], bl_top[1100],
     bl_top[1099], bl_top[1098], bl_top[1097], bl_top[1096],
     bl_top[1095], bl_top[1094], bl_top[1093], bl_top[1092],
     bl_top[1131], bl_top[1130], bl_top[1129], bl_top[1128],
     bl_top[1127], bl_top[1126], bl_top[1125], bl_top[1124],
     bl_top[1123], bl_top[1122], bl_top[1121], bl_top[1120],
     bl_top[1119], bl_top[1118], bl_top[1117], bl_top[1116],
     bl_top[1115], bl_top[1114], bl_top[1113], bl_top[1112],
     bl_top[1111], bl_top[1110], bl_top[1109], bl_top[1108],
     bl_top[1107], bl_top[1106], bl_top[1105], bl_top[1104],
     bl_top[1027], bl_top[1026], bl_top[1025], bl_top[1024],
     bl_top[1037], bl_top[1036], bl_top[1035], bl_top[1034],
     bl_top[1033], bl_top[1032], bl_top[1031], bl_top[1030],
     bl_top[1029], bl_top[1028], bl_top[1049], bl_top[1048],
     bl_top[1047], bl_top[1046], bl_top[1045], bl_top[1044],
     bl_top[1043], bl_top[1042], bl_top[1041], bl_top[1040],
     bl_top[1039], bl_top[1038], bl_top[1077], bl_top[1076],
     bl_top[1075], bl_top[1074], bl_top[1073], bl_top[1072],
     bl_top[1071], bl_top[1070], bl_top[1069], bl_top[1068],
     bl_top[1067], bl_top[1066], bl_top[1065], bl_top[1064],
     bl_top[1063], bl_top[1062], bl_top[1061], bl_top[1060],
     bl_top[1059], bl_top[1058], bl_top[1057], bl_top[1056],
     bl_top[1055], bl_top[1054], bl_top[1053], bl_top[1052],
     bl_top[1051], bl_top[1050], bl_top[985], bl_top[984], bl_top[983],
     bl_top[982], bl_top[995], bl_top[994], bl_top[993], bl_top[992],
     bl_top[991], bl_top[990], bl_top[989], bl_top[988], bl_top[987],
     bl_top[986], bl_top[1007], bl_top[1006], bl_top[1005],
     bl_top[1004], bl_top[1003], bl_top[1002], bl_top[1001],
     bl_top[1000], bl_top[999], bl_top[998], bl_top[997], bl_top[996],
     bl_top[1023], bl_top[1022], bl_top[1021], bl_top[1020],
     bl_top[1019], bl_top[1018], bl_top[1017], bl_top[1016],
     bl_top[1015], bl_top[1014], bl_top[1013], bl_top[1012],
     bl_top[1011], bl_top[1010], bl_top[1009], bl_top[1008],
     bl_top[931], bl_top[930], bl_top[929], bl_top[928], bl_top[941],
     bl_top[940], bl_top[939], bl_top[938], bl_top[937], bl_top[936],
     bl_top[935], bl_top[934], bl_top[933], bl_top[932], bl_top[953],
     bl_top[952], bl_top[951], bl_top[950], bl_top[949], bl_top[948],
     bl_top[947], bl_top[946], bl_top[945], bl_top[944], bl_top[943],
     bl_top[942], bl_top[981], bl_top[980], bl_top[979], bl_top[978],
     bl_top[977], bl_top[976], bl_top[975], bl_top[974], bl_top[973],
     bl_top[972], bl_top[971], bl_top[970], bl_top[969], bl_top[968],
     bl_top[967], bl_top[966], bl_top[965], bl_top[964], bl_top[963],
     bl_top[962], bl_top[961], bl_top[960], bl_top[959], bl_top[958],
     bl_top[957], bl_top[956], bl_top[955], bl_top[954], bl_top[877],
     bl_top[876], bl_top[875], bl_top[874], bl_top[887], bl_top[886],
     bl_top[885], bl_top[884], bl_top[883], bl_top[882], bl_top[881],
     bl_top[880], bl_top[879], bl_top[878], bl_top[899], bl_top[898],
     bl_top[897], bl_top[896], bl_top[895], bl_top[894], bl_top[893],
     bl_top[892], bl_top[891], bl_top[890], bl_top[889], bl_top[888],
     bl_top[927], bl_top[926], bl_top[925], bl_top[924], bl_top[923],
     bl_top[922], bl_top[921], bl_top[920], bl_top[919], bl_top[918],
     bl_top[917], bl_top[916], bl_top[915], bl_top[914], bl_top[913],
     bl_top[912], bl_top[911], bl_top[910], bl_top[909], bl_top[908],
     bl_top[907], bl_top[906], bl_top[905], bl_top[904], bl_top[903],
     bl_top[902], bl_top[901], bl_top[900], bl_top[823], bl_top[822],
     bl_top[821], bl_top[820], bl_top[833], bl_top[832], bl_top[831],
     bl_top[830], bl_top[829], bl_top[828], bl_top[827], bl_top[826],
     bl_top[825], bl_top[824], bl_top[845], bl_top[844], bl_top[843],
     bl_top[842], bl_top[841], bl_top[840], bl_top[839], bl_top[838],
     bl_top[837], bl_top[836], bl_top[835], bl_top[834], bl_top[873],
     bl_top[872], bl_top[871], bl_top[870], bl_top[869], bl_top[868],
     bl_top[867], bl_top[866], bl_top[865], bl_top[864], bl_top[863],
     bl_top[862], bl_top[861], bl_top[860], bl_top[859], bl_top[858],
     bl_top[857], bl_top[856], bl_top[855], bl_top[854], bl_top[853],
     bl_top[852], bl_top[851], bl_top[850], bl_top[849], bl_top[848],
     bl_top[847], bl_top[846], bl_top[769], bl_top[768], bl_top[767],
     bl_top[766], bl_top[779], bl_top[778], bl_top[777], bl_top[776],
     bl_top[775], bl_top[774], bl_top[773], bl_top[772], bl_top[771],
     bl_top[770], bl_top[791], bl_top[790], bl_top[789], bl_top[788],
     bl_top[787], bl_top[786], bl_top[785], bl_top[784], bl_top[783],
     bl_top[782], bl_top[781], bl_top[780], bl_top[819], bl_top[818],
     bl_top[817], bl_top[816], bl_top[815], bl_top[814], bl_top[813],
     bl_top[812], bl_top[811], bl_top[810], bl_top[809], bl_top[808],
     bl_top[807], bl_top[806], bl_top[805], bl_top[804], bl_top[803],
     bl_top[802], bl_top[801], bl_top[800], bl_top[799], bl_top[798],
     bl_top[797], bl_top[796], bl_top[795], bl_top[794], bl_top[793],
     bl_top[792], bl_top[715], bl_top[714], bl_top[713], bl_top[712],
     bl_top[725], bl_top[724], bl_top[723], bl_top[722], bl_top[721],
     bl_top[720], bl_top[719], bl_top[718], bl_top[717], bl_top[716],
     bl_top[737], bl_top[736], bl_top[735], bl_top[734], bl_top[733],
     bl_top[732], bl_top[731], bl_top[730], bl_top[729], bl_top[728],
     bl_top[727], bl_top[726], bl_top[765], bl_top[764], bl_top[763],
     bl_top[762], bl_top[761], bl_top[760], bl_top[759], bl_top[758],
     bl_top[757], bl_top[756], bl_top[755], bl_top[754], bl_top[753],
     bl_top[752], bl_top[751], bl_top[750], bl_top[749], bl_top[748],
     bl_top[747], bl_top[746], bl_top[745], bl_top[744], bl_top[743],
     bl_top[742], bl_top[741], bl_top[740], bl_top[739], bl_top[738],
     bl_top[661], bl_top[660], bl_top[659], bl_top[658], bl_top[671],
     bl_top[670], bl_top[669], bl_top[668], bl_top[667], bl_top[666],
     bl_top[665], bl_top[664], bl_top[663], bl_top[662], bl_top[683],
     bl_top[682], bl_top[681], bl_top[680], bl_top[679], bl_top[678],
     bl_top[677], bl_top[676], bl_top[675], bl_top[674], bl_top[673],
     bl_top[672], bl_top[711], bl_top[710], bl_top[709], bl_top[708],
     bl_top[707], bl_top[706], bl_top[705], bl_top[704], bl_top[703],
     bl_top[702], bl_top[701], bl_top[700], bl_top[699], bl_top[698],
     bl_top[697], bl_top[696], bl_top[695], bl_top[694], bl_top[693],
     bl_top[692], bl_top[691], bl_top[690], bl_top[689], bl_top[688],
     bl_top[687], bl_top[686], bl_top[685], bl_top[684]}),
     .end_of_startup_r(end_of_startup_r[19:10]), .cf_t(cf_t[575:288]),
     .cf_r(cf_r[479:240]), .hold_t_r(bank_cntl_top),
     .hold_r_t(bank_cntl_right), .padin_223(padin_223),
     .padin_163(padin_163), .glb_in(glb_net[7:0]),
     .pado_t(pado_t[47:24]), .padeb_t(padeb_t[47:24]),
     .padin_t(padin_t[47:24]),
     .end_of_startup_top_r(end_of_startup_t[23:12]),
     .bm_sreb_o(net1205), .bm_sclk_o(net1206), .bm_sa_o(net1207[0:7]),
     .bm_init_o(net1208), .bm_rcapmux_en_o(net1209),
     .bm_wdummymux_en_o(net1210), .bm_rcapmux_en_i(net861),
     .bm_wdummymux_en_i(net862), .bm_sreb_i(net855),
     .bm_sclk_i(net857), .bm_sa_i(net858[0:7]), .bm_init_i(net859),
     .bm_sclkrw_i(bm_sclkrw_b2_o[1]), .bm_sdi_i(bm_sdi_b2_o[1]),
     .bm_sweb_i(bm_sweb_b2_o[1]), .bm_sdo_o(bm_sdo_b3_o),
     .bm_sdo_i(net1223), .bm_sweb_o(net1222), .bm_sdi_o(net1223),
     .bm_sclkrw_o(net1224));
QUAD_BL I_BL ( net1285, net1287, net1284[0:7], net1283,
     bm_sclkrw_b0_o[1:0], bm_sdi_b0_o[1:0], net1379[0:1], net1281,
     bm_sweb_b0_o[1:0], net1288, net1260, net1378, net1377, net1376,
     net1375, net1374, net1373, net1372, net1371, net1370, net1369,
     net1368, net01230, cf_b[287:0], cf_l[239:0], fabric_out_34,
     bank_cntl_left, fabric_out_93, net1263, net1264, padeb_b[23:0],
     padeb_l[19:0], padin_34, padin_93, pado_b[23:0], pado_l[19:0],
     net1262, net1361, net1261, slf_op_00_10[3:0], net1227[0:7],
     net1228[0:7], net1229[0:7], net1230[0:7], net1231[0:7],
     net1360[0:7], net1232[0:7], net1233[0:7], net1234[0:7],
     net1235[0:7], net1236[0:7], slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0], net1359[0:7], net1358[0:7],
     net1426[0:7], net1357[0:7], net1356[0:7], net1355[0:7],
     net1354[0:7], net1353[0:7], net1352[0:7], net1537[0:7],
     spi_ss_in_lft_b[19:0], net1266, net1265, {bl_bot[603],
     bl_bot[602], bl_bot[601], bl_bot[600], bl_bot[613], bl_bot[612],
     bl_bot[611], bl_bot[610], bl_bot[609], bl_bot[608], bl_bot[607],
     bl_bot[606], bl_bot[605], bl_bot[604], bl_bot[625], bl_bot[624],
     bl_bot[623], bl_bot[622], bl_bot[621], bl_bot[620], bl_bot[619],
     bl_bot[618], bl_bot[617], bl_bot[616], bl_bot[615], bl_bot[614],
     bl_bot[653], bl_bot[652], bl_bot[651], bl_bot[650], bl_bot[649],
     bl_bot[648], bl_bot[647], bl_bot[646], bl_bot[645], bl_bot[644],
     bl_bot[643], bl_bot[642], bl_bot[641], bl_bot[640], bl_bot[639],
     bl_bot[638], bl_bot[637], bl_bot[636], bl_bot[635], bl_bot[634],
     bl_bot[633], bl_bot[632], bl_bot[631], bl_bot[630], bl_bot[629],
     bl_bot[628], bl_bot[627], bl_bot[626], bl_bot[549], bl_bot[548],
     bl_bot[547], bl_bot[546], bl_bot[559], bl_bot[558], bl_bot[557],
     bl_bot[556], bl_bot[555], bl_bot[554], bl_bot[553], bl_bot[552],
     bl_bot[551], bl_bot[550], bl_bot[571], bl_bot[570], bl_bot[569],
     bl_bot[568], bl_bot[567], bl_bot[566], bl_bot[565], bl_bot[564],
     bl_bot[563], bl_bot[562], bl_bot[561], bl_bot[560], bl_bot[599],
     bl_bot[598], bl_bot[597], bl_bot[596], bl_bot[595], bl_bot[594],
     bl_bot[593], bl_bot[592], bl_bot[591], bl_bot[590], bl_bot[589],
     bl_bot[588], bl_bot[587], bl_bot[586], bl_bot[585], bl_bot[584],
     bl_bot[583], bl_bot[582], bl_bot[581], bl_bot[580], bl_bot[579],
     bl_bot[578], bl_bot[577], bl_bot[576], bl_bot[575], bl_bot[574],
     bl_bot[573], bl_bot[572], bl_bot[495], bl_bot[494], bl_bot[493],
     bl_bot[492], bl_bot[505], bl_bot[504], bl_bot[503], bl_bot[502],
     bl_bot[501], bl_bot[500], bl_bot[499], bl_bot[498], bl_bot[497],
     bl_bot[496], bl_bot[517], bl_bot[516], bl_bot[515], bl_bot[514],
     bl_bot[513], bl_bot[512], bl_bot[511], bl_bot[510], bl_bot[509],
     bl_bot[508], bl_bot[507], bl_bot[506], bl_bot[545], bl_bot[544],
     bl_bot[543], bl_bot[542], bl_bot[541], bl_bot[540], bl_bot[539],
     bl_bot[538], bl_bot[537], bl_bot[536], bl_bot[535], bl_bot[534],
     bl_bot[533], bl_bot[532], bl_bot[531], bl_bot[530], bl_bot[529],
     bl_bot[528], bl_bot[527], bl_bot[526], bl_bot[525], bl_bot[524],
     bl_bot[523], bl_bot[522], bl_bot[521], bl_bot[520], bl_bot[519],
     bl_bot[518], bl_bot[441], bl_bot[440], bl_bot[439], bl_bot[438],
     bl_bot[451], bl_bot[450], bl_bot[449], bl_bot[448], bl_bot[447],
     bl_bot[446], bl_bot[445], bl_bot[444], bl_bot[443], bl_bot[442],
     bl_bot[463], bl_bot[462], bl_bot[461], bl_bot[460], bl_bot[459],
     bl_bot[458], bl_bot[457], bl_bot[456], bl_bot[455], bl_bot[454],
     bl_bot[453], bl_bot[452], bl_bot[491], bl_bot[490], bl_bot[489],
     bl_bot[488], bl_bot[487], bl_bot[486], bl_bot[485], bl_bot[484],
     bl_bot[483], bl_bot[482], bl_bot[481], bl_bot[480], bl_bot[479],
     bl_bot[478], bl_bot[477], bl_bot[476], bl_bot[475], bl_bot[474],
     bl_bot[473], bl_bot[472], bl_bot[471], bl_bot[470], bl_bot[469],
     bl_bot[468], bl_bot[467], bl_bot[466], bl_bot[465], bl_bot[464],
     bl_bot[387], bl_bot[386], bl_bot[385], bl_bot[384], bl_bot[397],
     bl_bot[396], bl_bot[395], bl_bot[394], bl_bot[393], bl_bot[392],
     bl_bot[391], bl_bot[390], bl_bot[389], bl_bot[388], bl_bot[409],
     bl_bot[408], bl_bot[407], bl_bot[406], bl_bot[405], bl_bot[404],
     bl_bot[403], bl_bot[402], bl_bot[401], bl_bot[400], bl_bot[399],
     bl_bot[398], bl_bot[437], bl_bot[436], bl_bot[435], bl_bot[434],
     bl_bot[433], bl_bot[432], bl_bot[431], bl_bot[430], bl_bot[429],
     bl_bot[428], bl_bot[427], bl_bot[426], bl_bot[425], bl_bot[424],
     bl_bot[423], bl_bot[422], bl_bot[421], bl_bot[420], bl_bot[419],
     bl_bot[418], bl_bot[417], bl_bot[416], bl_bot[415], bl_bot[414],
     bl_bot[413], bl_bot[412], bl_bot[411], bl_bot[410], bl_bot[333],
     bl_bot[332], bl_bot[331], bl_bot[330], bl_bot[343], bl_bot[342],
     bl_bot[341], bl_bot[340], bl_bot[339], bl_bot[338], bl_bot[337],
     bl_bot[336], bl_bot[335], bl_bot[334], bl_bot[355], bl_bot[354],
     bl_bot[353], bl_bot[352], bl_bot[351], bl_bot[350], bl_bot[349],
     bl_bot[348], bl_bot[347], bl_bot[346], bl_bot[345], bl_bot[344],
     bl_bot[383], bl_bot[382], bl_bot[381], bl_bot[380], bl_bot[379],
     bl_bot[378], bl_bot[377], bl_bot[376], bl_bot[375], bl_bot[374],
     bl_bot[373], bl_bot[372], bl_bot[371], bl_bot[370], bl_bot[369],
     bl_bot[368], bl_bot[367], bl_bot[366], bl_bot[365], bl_bot[364],
     bl_bot[363], bl_bot[362], bl_bot[361], bl_bot[360], bl_bot[359],
     bl_bot[358], bl_bot[357], bl_bot[356], bl_bot[291], bl_bot[290],
     bl_bot[289], bl_bot[288], bl_bot[301], bl_bot[300], bl_bot[299],
     bl_bot[298], bl_bot[297], bl_bot[296], bl_bot[295], bl_bot[294],
     bl_bot[293], bl_bot[292], bl_bot[313], bl_bot[312], bl_bot[311],
     bl_bot[310], bl_bot[309], bl_bot[308], bl_bot[307], bl_bot[306],
     bl_bot[305], bl_bot[304], bl_bot[303], bl_bot[302], bl_bot[329],
     bl_bot[328], bl_bot[327], bl_bot[326], bl_bot[325], bl_bot[324],
     bl_bot[323], bl_bot[322], bl_bot[321], bl_bot[320], bl_bot[319],
     bl_bot[318], bl_bot[317], bl_bot[316], bl_bot[315], bl_bot[314],
     bl_bot[237], bl_bot[236], bl_bot[235], bl_bot[234], bl_bot[247],
     bl_bot[246], bl_bot[245], bl_bot[244], bl_bot[243], bl_bot[242],
     bl_bot[241], bl_bot[240], bl_bot[239], bl_bot[238], bl_bot[259],
     bl_bot[258], bl_bot[257], bl_bot[256], bl_bot[255], bl_bot[254],
     bl_bot[253], bl_bot[252], bl_bot[251], bl_bot[250], bl_bot[249],
     bl_bot[248], bl_bot[287], bl_bot[286], bl_bot[285], bl_bot[284],
     bl_bot[283], bl_bot[282], bl_bot[281], bl_bot[280], bl_bot[279],
     bl_bot[278], bl_bot[277], bl_bot[276], bl_bot[275], bl_bot[274],
     bl_bot[273], bl_bot[272], bl_bot[271], bl_bot[270], bl_bot[269],
     bl_bot[268], bl_bot[267], bl_bot[266], bl_bot[265], bl_bot[264],
     bl_bot[263], bl_bot[262], bl_bot[261], bl_bot[260], bl_bot[183],
     bl_bot[182], bl_bot[181], bl_bot[180], bl_bot[193], bl_bot[192],
     bl_bot[191], bl_bot[190], bl_bot[189], bl_bot[188], bl_bot[187],
     bl_bot[186], bl_bot[185], bl_bot[184], bl_bot[205], bl_bot[204],
     bl_bot[203], bl_bot[202], bl_bot[201], bl_bot[200], bl_bot[199],
     bl_bot[198], bl_bot[197], bl_bot[196], bl_bot[195], bl_bot[194],
     bl_bot[233], bl_bot[232], bl_bot[231], bl_bot[230], bl_bot[229],
     bl_bot[228], bl_bot[227], bl_bot[226], bl_bot[225], bl_bot[224],
     bl_bot[223], bl_bot[222], bl_bot[221], bl_bot[220], bl_bot[219],
     bl_bot[218], bl_bot[217], bl_bot[216], bl_bot[215], bl_bot[214],
     bl_bot[213], bl_bot[212], bl_bot[211], bl_bot[210], bl_bot[209],
     bl_bot[208], bl_bot[207], bl_bot[206], bl_bot[129], bl_bot[128],
     bl_bot[127], bl_bot[126], bl_bot[139], bl_bot[138], bl_bot[137],
     bl_bot[136], bl_bot[135], bl_bot[134], bl_bot[133], bl_bot[132],
     bl_bot[131], bl_bot[130], bl_bot[151], bl_bot[150], bl_bot[149],
     bl_bot[148], bl_bot[147], bl_bot[146], bl_bot[145], bl_bot[144],
     bl_bot[143], bl_bot[142], bl_bot[141], bl_bot[140], bl_bot[179],
     bl_bot[178], bl_bot[177], bl_bot[176], bl_bot[175], bl_bot[174],
     bl_bot[173], bl_bot[172], bl_bot[171], bl_bot[170], bl_bot[169],
     bl_bot[168], bl_bot[167], bl_bot[166], bl_bot[165], bl_bot[164],
     bl_bot[163], bl_bot[162], bl_bot[161], bl_bot[160], bl_bot[159],
     bl_bot[158], bl_bot[157], bl_bot[156], bl_bot[155], bl_bot[154],
     bl_bot[153], bl_bot[152], bl_bot[75], bl_bot[74], bl_bot[73],
     bl_bot[72], bl_bot[85], bl_bot[84], bl_bot[83], bl_bot[82],
     bl_bot[81], bl_bot[80], bl_bot[79], bl_bot[78], bl_bot[77],
     bl_bot[76], bl_bot[97], bl_bot[96], bl_bot[95], bl_bot[94],
     bl_bot[93], bl_bot[92], bl_bot[91], bl_bot[90], bl_bot[89],
     bl_bot[88], bl_bot[87], bl_bot[86], bl_bot[125], bl_bot[124],
     bl_bot[123], bl_bot[122], bl_bot[121], bl_bot[120], bl_bot[119],
     bl_bot[118], bl_bot[117], bl_bot[116], bl_bot[115], bl_bot[114],
     bl_bot[113], bl_bot[112], bl_bot[111], bl_bot[110], bl_bot[109],
     bl_bot[108], bl_bot[107], bl_bot[106], bl_bot[105], bl_bot[104],
     bl_bot[103], bl_bot[102], bl_bot[101], bl_bot[100], bl_bot[99],
     bl_bot[98], bl_bot[21], bl_bot[20], bl_bot[19], bl_bot[18],
     bl_bot[31], bl_bot[30], bl_bot[29], bl_bot[28], bl_bot[27],
     bl_bot[26], bl_bot[25], bl_bot[24], bl_bot[23], bl_bot[22],
     bl_bot[43], bl_bot[42], bl_bot[41], bl_bot[40], bl_bot[39],
     bl_bot[38], bl_bot[37], bl_bot[36], bl_bot[35], bl_bot[34],
     bl_bot[33], bl_bot[32], bl_bot[71], bl_bot[70], bl_bot[69],
     bl_bot[68], bl_bot[67], bl_bot[66], bl_bot[65], bl_bot[64],
     bl_bot[63], bl_bot[62], bl_bot[61], bl_bot[60], bl_bot[59],
     bl_bot[58], bl_bot[57], bl_bot[56], bl_bot[55], bl_bot[54],
     bl_bot[53], bl_bot[52], bl_bot[51], bl_bot[50], bl_bot[49],
     bl_bot[48], bl_bot[47], bl_bot[46], bl_bot[45], bl_bot[44],
     bl_bot[14], bl_bot[15], bl_bot[16], bl_bot[17], bl_bot[8],
     bl_bot[9], bl_bot[10], bl_bot[11], bl_bot[12], bl_bot[13],
     bl_bot[2], bl_bot[3], bl_bot[4], bl_bot[5], bl_bot[6], bl_bot[7],
     bl_bot[0], bl_bot[1]}, {pgate_l[174], pgate_l[175], pgate_l[172],
     pgate_l[173], pgate_l[170], pgate_l[171], pgate_l[168],
     pgate_l[169], pgate_l[166], pgate_l[167], pgate_l[164],
     pgate_l[165], pgate_l[162], pgate_l[163], pgate_l[160],
     pgate_l[161], pgate_l[158], pgate_l[159], pgate_l[156],
     pgate_l[157], pgate_l[154], pgate_l[155], pgate_l[152],
     pgate_l[153], pgate_l[150], pgate_l[151], pgate_l[148],
     pgate_l[149], pgate_l[146], pgate_l[147], pgate_l[144],
     pgate_l[145], pgate_l[142], pgate_l[143], pgate_l[140],
     pgate_l[141], pgate_l[138], pgate_l[139], pgate_l[136],
     pgate_l[137], pgate_l[134], pgate_l[135], pgate_l[132],
     pgate_l[133], pgate_l[130], pgate_l[131], pgate_l[128],
     pgate_l[129], pgate_l[126], pgate_l[127], pgate_l[124],
     pgate_l[125], pgate_l[122], pgate_l[123], pgate_l[120],
     pgate_l[121], pgate_l[118], pgate_l[119], pgate_l[116],
     pgate_l[117], pgate_l[114], pgate_l[115], pgate_l[112],
     pgate_l[113], pgate_l[110], pgate_l[111], pgate_l[108],
     pgate_l[109], pgate_l[106], pgate_l[107], pgate_l[104],
     pgate_l[105], pgate_l[102], pgate_l[103], pgate_l[100],
     pgate_l[101], pgate_l[98], pgate_l[99], pgate_l[96], pgate_l[97],
     pgate_l[94], pgate_l[95], pgate_l[92], pgate_l[93], pgate_l[90],
     pgate_l[91], pgate_l[88], pgate_l[89], pgate_l[86], pgate_l[87],
     pgate_l[84], pgate_l[85], pgate_l[82], pgate_l[83], pgate_l[80],
     pgate_l[81], pgate_l[78], pgate_l[79], pgate_l[76], pgate_l[77],
     pgate_l[74], pgate_l[75], pgate_l[72], pgate_l[73], pgate_l[70],
     pgate_l[71], pgate_l[68], pgate_l[69], pgate_l[66], pgate_l[67],
     pgate_l[64], pgate_l[65], pgate_l[62], pgate_l[63], pgate_l[60],
     pgate_l[61], pgate_l[58], pgate_l[59], pgate_l[56], pgate_l[57],
     pgate_l[54], pgate_l[55], pgate_l[52], pgate_l[53], pgate_l[50],
     pgate_l[51], pgate_l[48], pgate_l[49], pgate_l[46], pgate_l[47],
     pgate_l[44], pgate_l[45], pgate_l[42], pgate_l[43], pgate_l[40],
     pgate_l[41], pgate_l[38], pgate_l[39], pgate_l[36], pgate_l[37],
     pgate_l[34], pgate_l[35], pgate_l[32], pgate_l[33], pgate_l[30],
     pgate_l[31], pgate_l[28], pgate_l[29], pgate_l[26], pgate_l[27],
     pgate_l[24], pgate_l[25], pgate_l[22], pgate_l[23], pgate_l[20],
     pgate_l[21], pgate_l[18], pgate_l[19], pgate_l[16], pgate_l[17],
     pgate_l[0], pgate_l[1], pgate_l[3], pgate_l[2], pgate_l[4],
     pgate_l[5], pgate_l[7], pgate_l[6], pgate_l[8], pgate_l[9],
     pgate_l[11], pgate_l[10], pgate_l[12], pgate_l[13], pgate_l[15],
     pgate_l[14]}, {reset_b_l[174], reset_b_l[175], reset_b_l[172],
     reset_b_l[173], reset_b_l[170], reset_b_l[171], reset_b_l[168],
     reset_b_l[169], reset_b_l[166], reset_b_l[167], reset_b_l[164],
     reset_b_l[165], reset_b_l[162], reset_b_l[163], reset_b_l[160],
     reset_b_l[161], reset_b_l[158], reset_b_l[159], reset_b_l[156],
     reset_b_l[157], reset_b_l[154], reset_b_l[155], reset_b_l[152],
     reset_b_l[153], reset_b_l[150], reset_b_l[151], reset_b_l[148],
     reset_b_l[149], reset_b_l[146], reset_b_l[147], reset_b_l[144],
     reset_b_l[145], reset_b_l[142], reset_b_l[143], reset_b_l[140],
     reset_b_l[141], reset_b_l[138], reset_b_l[139], reset_b_l[136],
     reset_b_l[137], reset_b_l[134], reset_b_l[135], reset_b_l[132],
     reset_b_l[133], reset_b_l[130], reset_b_l[131], reset_b_l[128],
     reset_b_l[129], reset_b_l[126], reset_b_l[127], reset_b_l[124],
     reset_b_l[125], reset_b_l[122], reset_b_l[123], reset_b_l[120],
     reset_b_l[121], reset_b_l[118], reset_b_l[119], reset_b_l[116],
     reset_b_l[117], reset_b_l[114], reset_b_l[115], reset_b_l[112],
     reset_b_l[113], reset_b_l[110], reset_b_l[111], reset_b_l[108],
     reset_b_l[109], reset_b_l[106], reset_b_l[107], reset_b_l[104],
     reset_b_l[105], reset_b_l[102], reset_b_l[103], reset_b_l[100],
     reset_b_l[101], reset_b_l[98], reset_b_l[99], reset_b_l[96],
     reset_b_l[97], reset_b_l[94], reset_b_l[95], reset_b_l[92],
     reset_b_l[93], reset_b_l[90], reset_b_l[91], reset_b_l[88],
     reset_b_l[89], reset_b_l[86], reset_b_l[87], reset_b_l[84],
     reset_b_l[85], reset_b_l[82], reset_b_l[83], reset_b_l[80],
     reset_b_l[81], reset_b_l[78], reset_b_l[79], reset_b_l[76],
     reset_b_l[77], reset_b_l[74], reset_b_l[75], reset_b_l[72],
     reset_b_l[73], reset_b_l[70], reset_b_l[71], reset_b_l[68],
     reset_b_l[69], reset_b_l[66], reset_b_l[67], reset_b_l[64],
     reset_b_l[65], reset_b_l[62], reset_b_l[63], reset_b_l[60],
     reset_b_l[61], reset_b_l[58], reset_b_l[59], reset_b_l[56],
     reset_b_l[57], reset_b_l[54], reset_b_l[55], reset_b_l[52],
     reset_b_l[53], reset_b_l[50], reset_b_l[51], reset_b_l[48],
     reset_b_l[49], reset_b_l[46], reset_b_l[47], reset_b_l[44],
     reset_b_l[45], reset_b_l[42], reset_b_l[43], reset_b_l[40],
     reset_b_l[41], reset_b_l[38], reset_b_l[39], reset_b_l[36],
     reset_b_l[37], reset_b_l[34], reset_b_l[35], reset_b_l[32],
     reset_b_l[33], reset_b_l[30], reset_b_l[31], reset_b_l[28],
     reset_b_l[29], reset_b_l[26], reset_b_l[27], reset_b_l[24],
     reset_b_l[25], reset_b_l[22], reset_b_l[23], reset_b_l[20],
     reset_b_l[21], reset_b_l[18], reset_b_l[19], reset_b_l[16],
     reset_b_l[17], reset_b_l[0], reset_b_l[1], reset_b_l[3],
     reset_b_l[2], reset_b_l[4], reset_b_l[5], reset_b_l[7],
     reset_b_l[6], reset_b_l[8], reset_b_l[9], reset_b_l[11],
     reset_b_l[10], reset_b_l[12], reset_b_l[13], reset_b_l[15],
     reset_b_l[14]}, net1299[0:15], net1422[0:47], net1421[0:47],
     net1350[0:47], net1420[0:47], net1419[0:47], net1418[0:47],
     net1323[0:47], net1322[0:47], net1417[0:47], net1416[0:47],
     net1414[0:47], net1413[0:47], net1412[0:47], net1411[0:47],
     net1410[0:47], net1409[0:47], net1408[0:47], net1407[0:47],
     net1406[0:47], net1405[0:47], net1324[0:15], net1404[0:47],
     net1403[0:47], net1402[0:47], net1401[0:47], net1400[0:47],
     net1399[0:47], net1398[0:47], net1397[0:47], net1396[0:47],
     net1395[0:47], net1394[0:47], net1393[0:47], net1312[0:23],
     net1313[0:23], net1314[0:23], net1311[0:23], net1315[0:23],
     net1318[0:23], net1317[0:23], net1316[0:23], net1320[0:23],
     net1319[0:23], net1392[0:23], net1391[0:23], net1390[0:23],
     net1389[0:23], net1388[0:23], net1387[0:23], net1386[0:23],
     net1385[0:23], net1384[0:23], net1383[0:23], net1382[0:23],
     net1381[0:23], {vdd_cntl_l[174], vdd_cntl_l[175], vdd_cntl_l[172],
     vdd_cntl_l[173], vdd_cntl_l[170], vdd_cntl_l[171],
     vdd_cntl_l[168], vdd_cntl_l[169], vdd_cntl_l[166],
     vdd_cntl_l[167], vdd_cntl_l[164], vdd_cntl_l[165],
     vdd_cntl_l[162], vdd_cntl_l[163], vdd_cntl_l[160],
     vdd_cntl_l[161], vdd_cntl_l[158], vdd_cntl_l[159],
     vdd_cntl_l[156], vdd_cntl_l[157], vdd_cntl_l[154],
     vdd_cntl_l[155], vdd_cntl_l[152], vdd_cntl_l[153],
     vdd_cntl_l[150], vdd_cntl_l[151], vdd_cntl_l[148],
     vdd_cntl_l[149], vdd_cntl_l[146], vdd_cntl_l[147],
     vdd_cntl_l[144], vdd_cntl_l[145], vdd_cntl_l[142],
     vdd_cntl_l[143], vdd_cntl_l[140], vdd_cntl_l[141],
     vdd_cntl_l[138], vdd_cntl_l[139], vdd_cntl_l[136],
     vdd_cntl_l[137], vdd_cntl_l[134], vdd_cntl_l[135],
     vdd_cntl_l[132], vdd_cntl_l[133], vdd_cntl_l[130],
     vdd_cntl_l[131], vdd_cntl_l[128], vdd_cntl_l[129],
     vdd_cntl_l[126], vdd_cntl_l[127], vdd_cntl_l[124],
     vdd_cntl_l[125], vdd_cntl_l[122], vdd_cntl_l[123],
     vdd_cntl_l[120], vdd_cntl_l[121], vdd_cntl_l[118],
     vdd_cntl_l[119], vdd_cntl_l[116], vdd_cntl_l[117],
     vdd_cntl_l[114], vdd_cntl_l[115], vdd_cntl_l[112],
     vdd_cntl_l[113], vdd_cntl_l[110], vdd_cntl_l[111],
     vdd_cntl_l[108], vdd_cntl_l[109], vdd_cntl_l[106],
     vdd_cntl_l[107], vdd_cntl_l[104], vdd_cntl_l[105],
     vdd_cntl_l[102], vdd_cntl_l[103], vdd_cntl_l[100],
     vdd_cntl_l[101], vdd_cntl_l[98], vdd_cntl_l[99], vdd_cntl_l[96],
     vdd_cntl_l[97], vdd_cntl_l[94], vdd_cntl_l[95], vdd_cntl_l[92],
     vdd_cntl_l[93], vdd_cntl_l[90], vdd_cntl_l[91], vdd_cntl_l[88],
     vdd_cntl_l[89], vdd_cntl_l[86], vdd_cntl_l[87], vdd_cntl_l[84],
     vdd_cntl_l[85], vdd_cntl_l[82], vdd_cntl_l[83], vdd_cntl_l[80],
     vdd_cntl_l[81], vdd_cntl_l[78], vdd_cntl_l[79], vdd_cntl_l[76],
     vdd_cntl_l[77], vdd_cntl_l[74], vdd_cntl_l[75], vdd_cntl_l[72],
     vdd_cntl_l[73], vdd_cntl_l[70], vdd_cntl_l[71], vdd_cntl_l[68],
     vdd_cntl_l[69], vdd_cntl_l[66], vdd_cntl_l[67], vdd_cntl_l[64],
     vdd_cntl_l[65], vdd_cntl_l[62], vdd_cntl_l[63], vdd_cntl_l[60],
     vdd_cntl_l[61], vdd_cntl_l[58], vdd_cntl_l[59], vdd_cntl_l[56],
     vdd_cntl_l[57], vdd_cntl_l[54], vdd_cntl_l[55], vdd_cntl_l[52],
     vdd_cntl_l[53], vdd_cntl_l[50], vdd_cntl_l[51], vdd_cntl_l[48],
     vdd_cntl_l[49], vdd_cntl_l[46], vdd_cntl_l[47], vdd_cntl_l[44],
     vdd_cntl_l[45], vdd_cntl_l[42], vdd_cntl_l[43], vdd_cntl_l[40],
     vdd_cntl_l[41], vdd_cntl_l[38], vdd_cntl_l[39], vdd_cntl_l[36],
     vdd_cntl_l[37], vdd_cntl_l[34], vdd_cntl_l[35], vdd_cntl_l[32],
     vdd_cntl_l[33], vdd_cntl_l[30], vdd_cntl_l[31], vdd_cntl_l[28],
     vdd_cntl_l[29], vdd_cntl_l[26], vdd_cntl_l[27], vdd_cntl_l[24],
     vdd_cntl_l[25], vdd_cntl_l[22], vdd_cntl_l[23], vdd_cntl_l[20],
     vdd_cntl_l[21], vdd_cntl_l[18], vdd_cntl_l[19], vdd_cntl_l[16],
     vdd_cntl_l[17], vdd_cntl_l[0], vdd_cntl_l[1], vdd_cntl_l[3],
     vdd_cntl_l[2], vdd_cntl_l[4], vdd_cntl_l[5], vdd_cntl_l[7],
     vdd_cntl_l[6], vdd_cntl_l[8], vdd_cntl_l[9], vdd_cntl_l[11],
     vdd_cntl_l[10], vdd_cntl_l[12], vdd_cntl_l[13], vdd_cntl_l[15],
     vdd_cntl_l[14]}, {wl_l[174], wl_l[175], wl_l[172], wl_l[173],
     wl_l[170], wl_l[171], wl_l[168], wl_l[169], wl_l[166], wl_l[167],
     wl_l[164], wl_l[165], wl_l[162], wl_l[163], wl_l[160], wl_l[161],
     wl_l[158], wl_l[159], wl_l[156], wl_l[157], wl_l[154], wl_l[155],
     wl_l[152], wl_l[153], wl_l[150], wl_l[151], wl_l[148], wl_l[149],
     wl_l[146], wl_l[147], wl_l[144], wl_l[145], wl_l[142], wl_l[143],
     wl_l[140], wl_l[141], wl_l[138], wl_l[139], wl_l[136], wl_l[137],
     wl_l[134], wl_l[135], wl_l[132], wl_l[133], wl_l[130], wl_l[131],
     wl_l[128], wl_l[129], wl_l[126], wl_l[127], wl_l[124], wl_l[125],
     wl_l[122], wl_l[123], wl_l[120], wl_l[121], wl_l[118], wl_l[119],
     wl_l[116], wl_l[117], wl_l[114], wl_l[115], wl_l[112], wl_l[113],
     wl_l[110], wl_l[111], wl_l[108], wl_l[109], wl_l[106], wl_l[107],
     wl_l[104], wl_l[105], wl_l[102], wl_l[103], wl_l[100], wl_l[101],
     wl_l[98], wl_l[99], wl_l[96], wl_l[97], wl_l[94], wl_l[95],
     wl_l[92], wl_l[93], wl_l[90], wl_l[91], wl_l[88], wl_l[89],
     wl_l[86], wl_l[87], wl_l[84], wl_l[85], wl_l[82], wl_l[83],
     wl_l[80], wl_l[81], wl_l[78], wl_l[79], wl_l[76], wl_l[77],
     wl_l[74], wl_l[75], wl_l[72], wl_l[73], wl_l[70], wl_l[71],
     wl_l[68], wl_l[69], wl_l[66], wl_l[67], wl_l[64], wl_l[65],
     wl_l[62], wl_l[63], wl_l[60], wl_l[61], wl_l[58], wl_l[59],
     wl_l[56], wl_l[57], wl_l[54], wl_l[55], wl_l[52], wl_l[53],
     wl_l[50], wl_l[51], wl_l[48], wl_l[49], wl_l[46], wl_l[47],
     wl_l[44], wl_l[45], wl_l[42], wl_l[43], wl_l[40], wl_l[41],
     wl_l[38], wl_l[39], wl_l[36], wl_l[37], wl_l[34], wl_l[35],
     wl_l[32], wl_l[33], wl_l[30], wl_l[31], wl_l[28], wl_l[29],
     wl_l[26], wl_l[27], wl_l[24], wl_l[25], wl_l[22], wl_l[23],
     wl_l[20], wl_l[21], wl_l[18], wl_l[19], wl_l[16], wl_l[17],
     wl_l[0], wl_l[1], wl_l[3], wl_l[2], wl_l[4], wl_l[5], wl_l[7],
     wl_l[6], wl_l[8], wl_l[9], wl_l[11], wl_l[10], wl_l[12], wl_l[13],
     wl_l[15], wl_l[14]}, net1297, net1290, net1296[0:7], net1295,
     net1294[0:1], net1289[0:1], {bm_sdo_b1_o, bm_sdi_b0_o[0]},
     net1293, net1292[0:1], net1291, slf_op_13_00[3:0], net1272,
     net01436, end_of_startup_l[9:0], glb_net[7:0], net1270,
     bank_cntl_bottom, bank_cntl_left, net1267, padin_b[23:0],
     padin_l[19:0], prog, purst, net1271, net1345[0:7], net1344[0:7],
     net1343[0:7], net1342[0:7], net1341[0:7], net1340[0:7],
     net1321[0:7], net1339[0:7], net1338[0:7], net1548[0:7], net1336,
     net1268, spioeb_lft_b[19:0], spiout_lft_b[19:0], net1273, tiegnd,
     tievdd, net1334[0:7], {slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0], slf_op_00_11[3],
     slf_op_00_11[2], slf_op_00_11[1], slf_op_00_11[0]}, net1334[0:7],
     net1331[0:7], net1332[0:7], net1335[0:7], net1330[0:7],
     net1325[0:7], net1333[0:7], net1328[0:7], net1327[0:7],
     net1329[0:7], net1326[0:7], net1331[0:7], net1332[0:7],
     net1335[0:7], net1330[0:7], net1325[0:7], net1333[0:7],
     net1328[0:7], net1327[0:7], net1329[0:7], net1326[0:7],
     net1415[0:7], net1310[0:7], net1334[0:7], net1331[0:7],
     net1332[0:7], net1335[0:7], net1330[0:7], net1325[0:7],
     net1333[0:7], net1328[0:7], net1327[0:7], net1329[0:7],
     net1326[0:7], net1415[0:7], net1269);
QUAD_TL I_TL ( .ceb_i(net01435), .ceb_o(net01436),
     .tnr_op_12_20(slf_op_13_21[3:0]), .bnr_op_11_11(net1537[0:7]),
     .bnr_op_10_11(net1236[0:7]), .bnr_op_09_11(net1235[0:7]),
     .bnr_op_08_11(net1234[0:7]), .bnr_op_07_11(net1233[0:7]),
     .bnr_op_06_11(net1232[0:7]), .bnr_op_05_11(net1360[0:7]),
     .bnr_op_04_11(net1231[0:7]), .bnr_op_03_11(net1230[0:7]),
     .bnr_op_02_11(net1229[0:7]), .bnr_op_01_11(net1228[0:7]),
     .bnr_op_00_11(net1227[0:7]), .bnl_op_12_11(net1236[0:7]),
     .bnl_op_11_11(net1235[0:7]), .bnl_op_10_11(net1234[0:7]),
     .bnl_op_09_11(net1233[0:7]), .bnl_op_08_11(net1232[0:7]),
     .bnl_op_07_11(net1360[0:7]), .bnl_op_06_11(net1231[0:7]),
     .bnl_op_05_11(net1230[0:7]), .bnl_op_04_11(net1229[0:7]),
     .bnl_op_03_11(net1228[0:7]), .bnl_op_02_11(net1227[0:7]),
     .shift_o(net1268), .hiz_b_o(net1270), .bs_en_o(net1272),
     .r_o(net1271), .tclk_o(net1273), .update_o(net1269),
     .mode_o(net1267), .mode_i(net1459), .shift_i(net1460),
     .update_i(net1461), .hiz_b_i(net1462), .r_i(net1463),
     .bs_en_i(net1464), .tclk_i(net1465), .tiegnd(tiegnd),
     .tievdd(tievdd), .bm_sdi_o(bm_sdo_b1_i), .bm_sweb_o(bm_sweb_b1_o),
     .bm_sreb_o(bm_sreb_b1_o), .bm_sclkrw_o(bm_sclkrw_b1_o),
     .bm_sclk_o(bm_sclk_b1_o), .bm_sa_o(bm_sa_b1_o[7:0]),
     .bm_init_o(bm_init_b1_o), .bm_sdo_i(bm_sdo_b1_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_b1_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_b1_o),
     .bm_sdi_i(bm_sdi_b0_o[1]), .bm_rcapmux_en_i(net1287),
     .bm_wdummymux_en_i(net1288), .bm_sdo_o(bm_sdo_b1_o),
     .bm_sweb_i(bm_sweb_b0_o[1]), .bm_sreb_i(net1281),
     .bm_sclkrw_i(bm_sclkrw_b0_o[1]), .bm_sclk_i(net1283),
     .bm_sa_i(net1284[0:7]), .bm_init_i(net1285),
     .end_of_startup_top_l(end_of_startup_t[11:0]),
     .end_of_startup_lft_t(end_of_startup_l[19:10]),
     .vdd_cntl({vdd_cntl_l[351], vdd_cntl_l[350], vdd_cntl_l[348],
     vdd_cntl_l[349], vdd_cntl_l[347], vdd_cntl_l[346],
     vdd_cntl_l[344], vdd_cntl_l[345], vdd_cntl_l[343],
     vdd_cntl_l[342], vdd_cntl_l[340], vdd_cntl_l[341],
     vdd_cntl_l[339], vdd_cntl_l[338], vdd_cntl_l[336],
     vdd_cntl_l[337], vdd_cntl_l[334], vdd_cntl_l[335],
     vdd_cntl_l[332], vdd_cntl_l[333], vdd_cntl_l[330],
     vdd_cntl_l[331], vdd_cntl_l[328], vdd_cntl_l[329],
     vdd_cntl_l[326], vdd_cntl_l[327], vdd_cntl_l[324],
     vdd_cntl_l[325], vdd_cntl_l[322], vdd_cntl_l[323],
     vdd_cntl_l[320], vdd_cntl_l[321], vdd_cntl_l[318],
     vdd_cntl_l[319], vdd_cntl_l[316], vdd_cntl_l[317],
     vdd_cntl_l[314], vdd_cntl_l[315], vdd_cntl_l[312],
     vdd_cntl_l[313], vdd_cntl_l[310], vdd_cntl_l[311],
     vdd_cntl_l[308], vdd_cntl_l[309], vdd_cntl_l[306],
     vdd_cntl_l[307], vdd_cntl_l[304], vdd_cntl_l[305],
     vdd_cntl_l[302], vdd_cntl_l[303], vdd_cntl_l[300],
     vdd_cntl_l[301], vdd_cntl_l[298], vdd_cntl_l[299],
     vdd_cntl_l[296], vdd_cntl_l[297], vdd_cntl_l[294],
     vdd_cntl_l[295], vdd_cntl_l[292], vdd_cntl_l[293],
     vdd_cntl_l[290], vdd_cntl_l[291], vdd_cntl_l[288],
     vdd_cntl_l[289], vdd_cntl_l[286], vdd_cntl_l[287],
     vdd_cntl_l[284], vdd_cntl_l[285], vdd_cntl_l[282],
     vdd_cntl_l[283], vdd_cntl_l[280], vdd_cntl_l[281],
     vdd_cntl_l[278], vdd_cntl_l[279], vdd_cntl_l[276],
     vdd_cntl_l[277], vdd_cntl_l[274], vdd_cntl_l[275],
     vdd_cntl_l[272], vdd_cntl_l[273], vdd_cntl_l[270],
     vdd_cntl_l[271], vdd_cntl_l[268], vdd_cntl_l[269],
     vdd_cntl_l[266], vdd_cntl_l[267], vdd_cntl_l[264],
     vdd_cntl_l[265], vdd_cntl_l[262], vdd_cntl_l[263],
     vdd_cntl_l[260], vdd_cntl_l[261], vdd_cntl_l[258],
     vdd_cntl_l[259], vdd_cntl_l[256], vdd_cntl_l[257],
     vdd_cntl_l[254], vdd_cntl_l[255], vdd_cntl_l[252],
     vdd_cntl_l[253], vdd_cntl_l[250], vdd_cntl_l[251],
     vdd_cntl_l[248], vdd_cntl_l[249], vdd_cntl_l[246],
     vdd_cntl_l[247], vdd_cntl_l[244], vdd_cntl_l[245],
     vdd_cntl_l[242], vdd_cntl_l[243], vdd_cntl_l[240],
     vdd_cntl_l[241], vdd_cntl_l[238], vdd_cntl_l[239],
     vdd_cntl_l[236], vdd_cntl_l[237], vdd_cntl_l[234],
     vdd_cntl_l[235], vdd_cntl_l[232], vdd_cntl_l[233],
     vdd_cntl_l[230], vdd_cntl_l[231], vdd_cntl_l[228],
     vdd_cntl_l[229], vdd_cntl_l[226], vdd_cntl_l[227],
     vdd_cntl_l[224], vdd_cntl_l[225], vdd_cntl_l[222],
     vdd_cntl_l[223], vdd_cntl_l[220], vdd_cntl_l[221],
     vdd_cntl_l[218], vdd_cntl_l[219], vdd_cntl_l[216],
     vdd_cntl_l[217], vdd_cntl_l[214], vdd_cntl_l[215],
     vdd_cntl_l[212], vdd_cntl_l[213], vdd_cntl_l[210],
     vdd_cntl_l[211], vdd_cntl_l[208], vdd_cntl_l[209],
     vdd_cntl_l[206], vdd_cntl_l[207], vdd_cntl_l[204],
     vdd_cntl_l[205], vdd_cntl_l[202], vdd_cntl_l[203],
     vdd_cntl_l[200], vdd_cntl_l[201], vdd_cntl_l[198],
     vdd_cntl_l[199], vdd_cntl_l[196], vdd_cntl_l[197],
     vdd_cntl_l[194], vdd_cntl_l[195], vdd_cntl_l[192],
     vdd_cntl_l[193], vdd_cntl_l[190], vdd_cntl_l[191],
     vdd_cntl_l[188], vdd_cntl_l[189], vdd_cntl_l[186],
     vdd_cntl_l[187], vdd_cntl_l[184], vdd_cntl_l[185],
     vdd_cntl_l[182], vdd_cntl_l[183], vdd_cntl_l[180],
     vdd_cntl_l[181], vdd_cntl_l[178], vdd_cntl_l[179],
     vdd_cntl_l[176], vdd_cntl_l[177]}), .cf_l(cf_l[479:240]),
     .cf_t(cf_t[287:0]), .hold_l_t(bank_cntl_left),
     .hold_t_l(bank_cntl_top), .padin_30(padin_30),
     .padin_226(padin_226), .glb_in(glb_net[7:0]),
     .sp12_h_r_12_13(net1498[0:23]), .sp12_h_r_12_11(net1499[0:23]),
     .sp12_h_r_12_12(net1500[0:23]), .sp12_h_r_12_20(net1501[0:23]),
     .sp12_h_r_12_19(net1502[0:23]), .sp12_h_r_12_18(net1503[0:23]),
     .sp12_h_r_12_17(net1504[0:23]), .sp12_h_r_12_16(net1505[0:23]),
     .sp12_h_r_12_15(net1506[0:23]), .sp12_h_r_12_14(net1507[0:23]),
     .sp4_h_r_12_21(net1508[0:15]), .sp4_v_b_00_11(net1324[0:15]),
     .bot_op_06_11(net1360[0:7]), .sp12_v_b_06_11(net1387[0:23]),
     .sp4_v_b_06_11(net1399[0:47]), .sp4_v_b_08_11(net1397[0:47]),
     .rgt_op_12_20(net1514[0:7]), .rgt_op_12_19(net1515[0:7]),
     .rgt_op_12_18(net1516[0:7]), .rgt_op_12_17(net1517[0:7]),
     .rgt_op_12_16(net1518[0:7]), .rgt_op_12_15(net1519[0:7]),
     .rgt_op_12_14(net1520[0:7]), .rgt_op_12_13(net1521[0:7]),
     .rgt_op_12_12(net1522[0:7]), .rgt_op_12_11(net1310[0:7]),
     .padin_t(padin_t[23:0]), .padin_l(padin_l[39:20]),
     .carry_in_12_11(net1368), .carry_in_11_11(net1369),
     .carry_in_10_11(net1370), .carry_in_09_11(net1371),
     .carry_in_08_11(net1372), .carry_in_07_11(net1373),
     .carry_in_05_11(net1374), .carry_in_04_11(net1375),
     .carry_in_03_11(net1376), .carry_in_02_11(net1377),
     .carry_in_01_11(net1378), .bot_op_12_11(net1537[0:7]),
     .bot_op_11_11(net1236[0:7]), .bot_op_10_11(net1235[0:7]),
     .bot_op_09_11(net1234[0:7]), .bot_op_08_11(net1233[0:7]),
     .bot_op_07_11(net1232[0:7]), .bot_op_05_11(net1231[0:7]),
     .bot_op_04_11(net1230[0:7]), .bot_op_03_11(net1229[0:7]),
     .bot_op_02_11(net1228[0:7]), .bot_op_01_11(net1227[0:7]),
     .bnr_op_12_11(net1548[0:7]), .bnl_op_01_11({slf_op_00_10[3],
     slf_op_00_10[2], slf_op_00_10[1], slf_op_00_10[0],
     slf_op_00_10[3], slf_op_00_10[2], slf_op_00_10[1],
     slf_op_00_10[0]}), .slf_op_12_21(slf_op_12_21[3:0]),
     .slf_op_12_20(net1551[0:7]), .slf_op_12_19(net1552[0:7]),
     .slf_op_12_18(net1553[0:7]), .slf_op_12_17(net1554[0:7]),
     .slf_op_12_16(net1555[0:7]), .slf_op_12_15(net1556[0:7]),
     .slf_op_12_14(net1557[0:7]), .slf_op_12_13(net1558[0:7]),
     .slf_op_12_12(net1559[0:7]), .slf_op_12_11(net1415[0:7]),
     .slf_op_11_11(net1326[0:7]), .slf_op_10_11(net1329[0:7]),
     .slf_op_09_11(net1327[0:7]), .slf_op_08_11(net1328[0:7]),
     .slf_op_07_11(net1333[0:7]), .slf_op_06_11(net1325[0:7]),
     .slf_op_05_11(net1330[0:7]), .slf_op_04_11(net1335[0:7]),
     .slf_op_03_11(net1332[0:7]), .slf_op_02_11(net1331[0:7]),
     .slf_op_01_11(net1334[0:7]), .slf_op_00_11(slf_op_00_11[3:0]),
     .pado_t(pado_t[23:0]), .pado_l(pado_l[39:20]),
     .padeb_t(padeb_t[23:0]), .padeb_l(padeb_l[39:20]),
     .fabric_out_30(fabric_out_30), .sp12_v_b_12_11(net1381[0:23]),
     .sp12_v_b_11_11(net1382[0:23]), .sp12_v_b_10_11(net1383[0:23]),
     .sp12_v_b_09_11(net1384[0:23]), .sp12_v_b_08_11(net1385[0:23]),
     .sp12_v_b_07_11(net1386[0:23]), .sp12_v_b_05_11(net1388[0:23]),
     .sp12_v_b_04_11(net1389[0:23]), .sp12_v_b_03_11(net1390[0:23]),
     .sp12_v_b_02_11(net1391[0:23]), .sp12_v_b_01_11(net1392[0:23]),
     .sp4_v_b_12_11(net1393[0:47]), .sp4_v_b_11_11(net1394[0:47]),
     .sp4_v_b_10_11(net1395[0:47]), .sp4_v_b_09_11(net1396[0:47]),
     .sp4_v_b_07_11(net1398[0:47]), .sp4_v_b_05_11(net1400[0:47]),
     .sp4_v_b_04_11(net1401[0:47]), .sp4_v_b_03_11(net1402[0:47]),
     .sp4_v_b_02_11(net1403[0:47]), .sp4_v_b_01_11(net1404[0:47]),
     .sp4_r_v_b_12_20(net1599[0:47]), .sp4_r_v_b_12_19(net1600[0:47]),
     .sp4_r_v_b_12_18(net1601[0:47]), .sp4_r_v_b_12_17(net1602[0:47]),
     .sp4_r_v_b_12_16(net1603[0:47]), .sp4_r_v_b_12_15(net1604[0:47]),
     .sp4_r_v_b_12_14(net1605[0:47]), .sp4_r_v_b_12_13(net1606[0:47]),
     .sp4_r_v_b_12_12(net1607[0:47]), .sp4_r_v_b_12_11(net991[0:47]),
     .sp4_h_r_12_20(net1609[0:47]), .sp4_h_r_12_19(net1610[0:47]),
     .sp4_h_r_12_18(net1611[0:47]), .sp4_h_r_12_17(net1612[0:47]),
     .sp4_h_r_12_16(net1613[0:47]), .sp4_h_r_12_15(net1614[0:47]),
     .sp4_h_r_12_14(net1615[0:47]), .sp4_h_r_12_13(net1616[0:47]),
     .sp4_h_r_12_12(net1617[0:47]), .sp4_h_r_12_11(net1618[0:47]),
     .bl({bl_top[603], bl_top[602], bl_top[601], bl_top[600],
     bl_top[613], bl_top[612], bl_top[611], bl_top[610], bl_top[609],
     bl_top[608], bl_top[607], bl_top[606], bl_top[605], bl_top[604],
     bl_top[625], bl_top[624], bl_top[623], bl_top[622], bl_top[621],
     bl_top[620], bl_top[619], bl_top[618], bl_top[617], bl_top[616],
     bl_top[615], bl_top[614], bl_top[653], bl_top[652], bl_top[651],
     bl_top[650], bl_top[649], bl_top[648], bl_top[647], bl_top[646],
     bl_top[645], bl_top[644], bl_top[643], bl_top[642], bl_top[641],
     bl_top[640], bl_top[639], bl_top[638], bl_top[637], bl_top[636],
     bl_top[635], bl_top[634], bl_top[633], bl_top[632], bl_top[631],
     bl_top[630], bl_top[629], bl_top[628], bl_top[627], bl_top[626],
     bl_top[549], bl_top[548], bl_top[547], bl_top[546], bl_top[559],
     bl_top[558], bl_top[557], bl_top[556], bl_top[555], bl_top[554],
     bl_top[553], bl_top[552], bl_top[551], bl_top[550], bl_top[571],
     bl_top[570], bl_top[569], bl_top[568], bl_top[567], bl_top[566],
     bl_top[565], bl_top[564], bl_top[563], bl_top[562], bl_top[561],
     bl_top[560], bl_top[599], bl_top[598], bl_top[597], bl_top[596],
     bl_top[595], bl_top[594], bl_top[593], bl_top[592], bl_top[591],
     bl_top[590], bl_top[589], bl_top[588], bl_top[587], bl_top[586],
     bl_top[585], bl_top[584], bl_top[583], bl_top[582], bl_top[581],
     bl_top[580], bl_top[579], bl_top[578], bl_top[577], bl_top[576],
     bl_top[575], bl_top[574], bl_top[573], bl_top[572], bl_top[495],
     bl_top[494], bl_top[493], bl_top[492], bl_top[505], bl_top[504],
     bl_top[503], bl_top[502], bl_top[501], bl_top[500], bl_top[499],
     bl_top[498], bl_top[497], bl_top[496], bl_top[517], bl_top[516],
     bl_top[515], bl_top[514], bl_top[513], bl_top[512], bl_top[511],
     bl_top[510], bl_top[509], bl_top[508], bl_top[507], bl_top[506],
     bl_top[545], bl_top[544], bl_top[543], bl_top[542], bl_top[541],
     bl_top[540], bl_top[539], bl_top[538], bl_top[537], bl_top[536],
     bl_top[535], bl_top[534], bl_top[533], bl_top[532], bl_top[531],
     bl_top[530], bl_top[529], bl_top[528], bl_top[527], bl_top[526],
     bl_top[525], bl_top[524], bl_top[523], bl_top[522], bl_top[521],
     bl_top[520], bl_top[519], bl_top[518], bl_top[441], bl_top[440],
     bl_top[439], bl_top[438], bl_top[451], bl_top[450], bl_top[449],
     bl_top[448], bl_top[447], bl_top[446], bl_top[445], bl_top[444],
     bl_top[443], bl_top[442], bl_top[463], bl_top[462], bl_top[461],
     bl_top[460], bl_top[459], bl_top[458], bl_top[457], bl_top[456],
     bl_top[455], bl_top[454], bl_top[453], bl_top[452], bl_top[491],
     bl_top[490], bl_top[489], bl_top[488], bl_top[487], bl_top[486],
     bl_top[485], bl_top[484], bl_top[483], bl_top[482], bl_top[481],
     bl_top[480], bl_top[479], bl_top[478], bl_top[477], bl_top[476],
     bl_top[475], bl_top[474], bl_top[473], bl_top[472], bl_top[471],
     bl_top[470], bl_top[469], bl_top[468], bl_top[467], bl_top[466],
     bl_top[465], bl_top[464], bl_top[387], bl_top[386], bl_top[385],
     bl_top[384], bl_top[397], bl_top[396], bl_top[395], bl_top[394],
     bl_top[393], bl_top[392], bl_top[391], bl_top[390], bl_top[389],
     bl_top[388], bl_top[409], bl_top[408], bl_top[407], bl_top[406],
     bl_top[405], bl_top[404], bl_top[403], bl_top[402], bl_top[401],
     bl_top[400], bl_top[399], bl_top[398], bl_top[437], bl_top[436],
     bl_top[435], bl_top[434], bl_top[433], bl_top[432], bl_top[431],
     bl_top[430], bl_top[429], bl_top[428], bl_top[427], bl_top[426],
     bl_top[425], bl_top[424], bl_top[423], bl_top[422], bl_top[421],
     bl_top[420], bl_top[419], bl_top[418], bl_top[417], bl_top[416],
     bl_top[415], bl_top[414], bl_top[413], bl_top[412], bl_top[411],
     bl_top[410], bl_top[333], bl_top[332], bl_top[331], bl_top[330],
     bl_top[343], bl_top[342], bl_top[341], bl_top[340], bl_top[339],
     bl_top[338], bl_top[337], bl_top[336], bl_top[335], bl_top[334],
     bl_top[355], bl_top[354], bl_top[353], bl_top[352], bl_top[351],
     bl_top[350], bl_top[349], bl_top[348], bl_top[347], bl_top[346],
     bl_top[345], bl_top[344], bl_top[383], bl_top[382], bl_top[381],
     bl_top[380], bl_top[379], bl_top[378], bl_top[377], bl_top[376],
     bl_top[375], bl_top[374], bl_top[373], bl_top[372], bl_top[371],
     bl_top[370], bl_top[369], bl_top[368], bl_top[367], bl_top[366],
     bl_top[365], bl_top[364], bl_top[363], bl_top[362], bl_top[361],
     bl_top[360], bl_top[359], bl_top[358], bl_top[357], bl_top[356],
     bl_top[291], bl_top[290], bl_top[289], bl_top[288], bl_top[301],
     bl_top[300], bl_top[299], bl_top[298], bl_top[297], bl_top[296],
     bl_top[295], bl_top[294], bl_top[293], bl_top[292], bl_top[313],
     bl_top[312], bl_top[311], bl_top[310], bl_top[309], bl_top[308],
     bl_top[307], bl_top[306], bl_top[305], bl_top[304], bl_top[303],
     bl_top[302], bl_top[329], bl_top[328], bl_top[327], bl_top[326],
     bl_top[325], bl_top[324], bl_top[323], bl_top[322], bl_top[321],
     bl_top[320], bl_top[319], bl_top[318], bl_top[317], bl_top[316],
     bl_top[315], bl_top[314], bl_top[237], bl_top[236], bl_top[235],
     bl_top[234], bl_top[247], bl_top[246], bl_top[245], bl_top[244],
     bl_top[243], bl_top[242], bl_top[241], bl_top[240], bl_top[239],
     bl_top[238], bl_top[259], bl_top[258], bl_top[257], bl_top[256],
     bl_top[255], bl_top[254], bl_top[253], bl_top[252], bl_top[251],
     bl_top[250], bl_top[249], bl_top[248], bl_top[287], bl_top[286],
     bl_top[285], bl_top[284], bl_top[283], bl_top[282], bl_top[281],
     bl_top[280], bl_top[279], bl_top[278], bl_top[277], bl_top[276],
     bl_top[275], bl_top[274], bl_top[273], bl_top[272], bl_top[271],
     bl_top[270], bl_top[269], bl_top[268], bl_top[267], bl_top[266],
     bl_top[265], bl_top[264], bl_top[263], bl_top[262], bl_top[261],
     bl_top[260], bl_top[183], bl_top[182], bl_top[181], bl_top[180],
     bl_top[193], bl_top[192], bl_top[191], bl_top[190], bl_top[189],
     bl_top[188], bl_top[187], bl_top[186], bl_top[185], bl_top[184],
     bl_top[205], bl_top[204], bl_top[203], bl_top[202], bl_top[201],
     bl_top[200], bl_top[199], bl_top[198], bl_top[197], bl_top[196],
     bl_top[195], bl_top[194], bl_top[233], bl_top[232], bl_top[231],
     bl_top[230], bl_top[229], bl_top[228], bl_top[227], bl_top[226],
     bl_top[225], bl_top[224], bl_top[223], bl_top[222], bl_top[221],
     bl_top[220], bl_top[219], bl_top[218], bl_top[217], bl_top[216],
     bl_top[215], bl_top[214], bl_top[213], bl_top[212], bl_top[211],
     bl_top[210], bl_top[209], bl_top[208], bl_top[207], bl_top[206],
     bl_top[129], bl_top[128], bl_top[127], bl_top[126], bl_top[139],
     bl_top[138], bl_top[137], bl_top[136], bl_top[135], bl_top[134],
     bl_top[133], bl_top[132], bl_top[131], bl_top[130], bl_top[151],
     bl_top[150], bl_top[149], bl_top[148], bl_top[147], bl_top[146],
     bl_top[145], bl_top[144], bl_top[143], bl_top[142], bl_top[141],
     bl_top[140], bl_top[179], bl_top[178], bl_top[177], bl_top[176],
     bl_top[175], bl_top[174], bl_top[173], bl_top[172], bl_top[171],
     bl_top[170], bl_top[169], bl_top[168], bl_top[167], bl_top[166],
     bl_top[165], bl_top[164], bl_top[163], bl_top[162], bl_top[161],
     bl_top[160], bl_top[159], bl_top[158], bl_top[157], bl_top[156],
     bl_top[155], bl_top[154], bl_top[153], bl_top[152], bl_top[75],
     bl_top[74], bl_top[73], bl_top[72], bl_top[85], bl_top[84],
     bl_top[83], bl_top[82], bl_top[81], bl_top[80], bl_top[79],
     bl_top[78], bl_top[77], bl_top[76], bl_top[97], bl_top[96],
     bl_top[95], bl_top[94], bl_top[93], bl_top[92], bl_top[91],
     bl_top[90], bl_top[89], bl_top[88], bl_top[87], bl_top[86],
     bl_top[125], bl_top[124], bl_top[123], bl_top[122], bl_top[121],
     bl_top[120], bl_top[119], bl_top[118], bl_top[117], bl_top[116],
     bl_top[115], bl_top[114], bl_top[113], bl_top[112], bl_top[111],
     bl_top[110], bl_top[109], bl_top[108], bl_top[107], bl_top[106],
     bl_top[105], bl_top[104], bl_top[103], bl_top[102], bl_top[101],
     bl_top[100], bl_top[99], bl_top[98], bl_top[21], bl_top[20],
     bl_top[19], bl_top[18], bl_top[31], bl_top[30], bl_top[29],
     bl_top[28], bl_top[27], bl_top[26], bl_top[25], bl_top[24],
     bl_top[23], bl_top[22], bl_top[43], bl_top[42], bl_top[41],
     bl_top[40], bl_top[39], bl_top[38], bl_top[37], bl_top[36],
     bl_top[35], bl_top[34], bl_top[33], bl_top[32], bl_top[71],
     bl_top[70], bl_top[69], bl_top[68], bl_top[67], bl_top[66],
     bl_top[65], bl_top[64], bl_top[63], bl_top[62], bl_top[61],
     bl_top[60], bl_top[59], bl_top[58], bl_top[57], bl_top[56],
     bl_top[55], bl_top[54], bl_top[53], bl_top[52], bl_top[51],
     bl_top[50], bl_top[49], bl_top[48], bl_top[47], bl_top[46],
     bl_top[45], bl_top[44], bl_top[14], bl_top[15], bl_top[16],
     bl_top[17], bl_top[8], bl_top[9], bl_top[10], bl_top[11],
     bl_top[12], bl_top[13], bl_top[2], bl_top[3], bl_top[4],
     bl_top[5], bl_top[6], bl_top[7], bl_top[0], bl_top[1]}),
     .fabric_out_226(fabric_out_226), .fabric_out_228(bank_cntl_top),
     .wl({wl_l[351], wl_l[350], wl_l[348], wl_l[349], wl_l[347],
     wl_l[346], wl_l[344], wl_l[345], wl_l[343], wl_l[342], wl_l[340],
     wl_l[341], wl_l[339], wl_l[338], wl_l[336], wl_l[337], wl_l[334],
     wl_l[335], wl_l[332], wl_l[333], wl_l[330], wl_l[331], wl_l[328],
     wl_l[329], wl_l[326], wl_l[327], wl_l[324], wl_l[325], wl_l[322],
     wl_l[323], wl_l[320], wl_l[321], wl_l[318], wl_l[319], wl_l[316],
     wl_l[317], wl_l[314], wl_l[315], wl_l[312], wl_l[313], wl_l[310],
     wl_l[311], wl_l[308], wl_l[309], wl_l[306], wl_l[307], wl_l[304],
     wl_l[305], wl_l[302], wl_l[303], wl_l[300], wl_l[301], wl_l[298],
     wl_l[299], wl_l[296], wl_l[297], wl_l[294], wl_l[295], wl_l[292],
     wl_l[293], wl_l[290], wl_l[291], wl_l[288], wl_l[289], wl_l[286],
     wl_l[287], wl_l[284], wl_l[285], wl_l[282], wl_l[283], wl_l[280],
     wl_l[281], wl_l[278], wl_l[279], wl_l[276], wl_l[277], wl_l[274],
     wl_l[275], wl_l[272], wl_l[273], wl_l[270], wl_l[271], wl_l[268],
     wl_l[269], wl_l[266], wl_l[267], wl_l[264], wl_l[265], wl_l[262],
     wl_l[263], wl_l[260], wl_l[261], wl_l[258], wl_l[259], wl_l[256],
     wl_l[257], wl_l[254], wl_l[255], wl_l[252], wl_l[253], wl_l[250],
     wl_l[251], wl_l[248], wl_l[249], wl_l[246], wl_l[247], wl_l[244],
     wl_l[245], wl_l[242], wl_l[243], wl_l[240], wl_l[241], wl_l[238],
     wl_l[239], wl_l[236], wl_l[237], wl_l[234], wl_l[235], wl_l[232],
     wl_l[233], wl_l[230], wl_l[231], wl_l[228], wl_l[229], wl_l[226],
     wl_l[227], wl_l[224], wl_l[225], wl_l[222], wl_l[223], wl_l[220],
     wl_l[221], wl_l[218], wl_l[219], wl_l[216], wl_l[217], wl_l[214],
     wl_l[215], wl_l[212], wl_l[213], wl_l[210], wl_l[211], wl_l[208],
     wl_l[209], wl_l[206], wl_l[207], wl_l[204], wl_l[205], wl_l[202],
     wl_l[203], wl_l[200], wl_l[201], wl_l[198], wl_l[199], wl_l[196],
     wl_l[197], wl_l[194], wl_l[195], wl_l[192], wl_l[193], wl_l[190],
     wl_l[191], wl_l[188], wl_l[189], wl_l[186], wl_l[187], wl_l[184],
     wl_l[185], wl_l[182], wl_l[183], wl_l[180], wl_l[181], wl_l[178],
     wl_l[179], wl_l[176], wl_l[177]}), .sdi(net1623),
     .reset_b({reset_b_l[351], reset_b_l[350], reset_b_l[348],
     reset_b_l[349], reset_b_l[347], reset_b_l[346], reset_b_l[344],
     reset_b_l[345], reset_b_l[343], reset_b_l[342], reset_b_l[340],
     reset_b_l[341], reset_b_l[339], reset_b_l[338], reset_b_l[336],
     reset_b_l[337], reset_b_l[334], reset_b_l[335], reset_b_l[332],
     reset_b_l[333], reset_b_l[330], reset_b_l[331], reset_b_l[328],
     reset_b_l[329], reset_b_l[326], reset_b_l[327], reset_b_l[324],
     reset_b_l[325], reset_b_l[322], reset_b_l[323], reset_b_l[320],
     reset_b_l[321], reset_b_l[318], reset_b_l[319], reset_b_l[316],
     reset_b_l[317], reset_b_l[314], reset_b_l[315], reset_b_l[312],
     reset_b_l[313], reset_b_l[310], reset_b_l[311], reset_b_l[308],
     reset_b_l[309], reset_b_l[306], reset_b_l[307], reset_b_l[304],
     reset_b_l[305], reset_b_l[302], reset_b_l[303], reset_b_l[300],
     reset_b_l[301], reset_b_l[298], reset_b_l[299], reset_b_l[296],
     reset_b_l[297], reset_b_l[294], reset_b_l[295], reset_b_l[292],
     reset_b_l[293], reset_b_l[290], reset_b_l[291], reset_b_l[288],
     reset_b_l[289], reset_b_l[286], reset_b_l[287], reset_b_l[284],
     reset_b_l[285], reset_b_l[282], reset_b_l[283], reset_b_l[280],
     reset_b_l[281], reset_b_l[278], reset_b_l[279], reset_b_l[276],
     reset_b_l[277], reset_b_l[274], reset_b_l[275], reset_b_l[272],
     reset_b_l[273], reset_b_l[270], reset_b_l[271], reset_b_l[268],
     reset_b_l[269], reset_b_l[266], reset_b_l[267], reset_b_l[264],
     reset_b_l[265], reset_b_l[262], reset_b_l[263], reset_b_l[260],
     reset_b_l[261], reset_b_l[258], reset_b_l[259], reset_b_l[256],
     reset_b_l[257], reset_b_l[254], reset_b_l[255], reset_b_l[252],
     reset_b_l[253], reset_b_l[250], reset_b_l[251], reset_b_l[248],
     reset_b_l[249], reset_b_l[246], reset_b_l[247], reset_b_l[244],
     reset_b_l[245], reset_b_l[242], reset_b_l[243], reset_b_l[240],
     reset_b_l[241], reset_b_l[238], reset_b_l[239], reset_b_l[236],
     reset_b_l[237], reset_b_l[234], reset_b_l[235], reset_b_l[232],
     reset_b_l[233], reset_b_l[230], reset_b_l[231], reset_b_l[228],
     reset_b_l[229], reset_b_l[226], reset_b_l[227], reset_b_l[224],
     reset_b_l[225], reset_b_l[222], reset_b_l[223], reset_b_l[220],
     reset_b_l[221], reset_b_l[218], reset_b_l[219], reset_b_l[216],
     reset_b_l[217], reset_b_l[214], reset_b_l[215], reset_b_l[212],
     reset_b_l[213], reset_b_l[210], reset_b_l[211], reset_b_l[208],
     reset_b_l[209], reset_b_l[206], reset_b_l[207], reset_b_l[204],
     reset_b_l[205], reset_b_l[202], reset_b_l[203], reset_b_l[200],
     reset_b_l[201], reset_b_l[198], reset_b_l[199], reset_b_l[196],
     reset_b_l[197], reset_b_l[194], reset_b_l[195], reset_b_l[192],
     reset_b_l[193], reset_b_l[190], reset_b_l[191], reset_b_l[188],
     reset_b_l[189], reset_b_l[186], reset_b_l[187], reset_b_l[184],
     reset_b_l[185], reset_b_l[182], reset_b_l[183], reset_b_l[180],
     reset_b_l[181], reset_b_l[178], reset_b_l[179], reset_b_l[176],
     reset_b_l[177]}), .purst(purst), .prog(prog),
     .pgate({pgate_l[351], pgate_l[350], pgate_l[348], pgate_l[349],
     pgate_l[347], pgate_l[346], pgate_l[344], pgate_l[345],
     pgate_l[343], pgate_l[342], pgate_l[340], pgate_l[341],
     pgate_l[339], pgate_l[338], pgate_l[336], pgate_l[337],
     pgate_l[334], pgate_l[335], pgate_l[332], pgate_l[333],
     pgate_l[330], pgate_l[331], pgate_l[328], pgate_l[329],
     pgate_l[326], pgate_l[327], pgate_l[324], pgate_l[325],
     pgate_l[322], pgate_l[323], pgate_l[320], pgate_l[321],
     pgate_l[318], pgate_l[319], pgate_l[316], pgate_l[317],
     pgate_l[314], pgate_l[315], pgate_l[312], pgate_l[313],
     pgate_l[310], pgate_l[311], pgate_l[308], pgate_l[309],
     pgate_l[306], pgate_l[307], pgate_l[304], pgate_l[305],
     pgate_l[302], pgate_l[303], pgate_l[300], pgate_l[301],
     pgate_l[298], pgate_l[299], pgate_l[296], pgate_l[297],
     pgate_l[294], pgate_l[295], pgate_l[292], pgate_l[293],
     pgate_l[290], pgate_l[291], pgate_l[288], pgate_l[289],
     pgate_l[286], pgate_l[287], pgate_l[284], pgate_l[285],
     pgate_l[282], pgate_l[283], pgate_l[280], pgate_l[281],
     pgate_l[278], pgate_l[279], pgate_l[276], pgate_l[277],
     pgate_l[274], pgate_l[275], pgate_l[272], pgate_l[273],
     pgate_l[270], pgate_l[271], pgate_l[268], pgate_l[269],
     pgate_l[266], pgate_l[267], pgate_l[264], pgate_l[265],
     pgate_l[262], pgate_l[263], pgate_l[260], pgate_l[261],
     pgate_l[258], pgate_l[259], pgate_l[256], pgate_l[257],
     pgate_l[254], pgate_l[255], pgate_l[252], pgate_l[253],
     pgate_l[250], pgate_l[251], pgate_l[248], pgate_l[249],
     pgate_l[246], pgate_l[247], pgate_l[244], pgate_l[245],
     pgate_l[242], pgate_l[243], pgate_l[240], pgate_l[241],
     pgate_l[238], pgate_l[239], pgate_l[236], pgate_l[237],
     pgate_l[234], pgate_l[235], pgate_l[232], pgate_l[233],
     pgate_l[230], pgate_l[231], pgate_l[228], pgate_l[229],
     pgate_l[226], pgate_l[227], pgate_l[224], pgate_l[225],
     pgate_l[222], pgate_l[223], pgate_l[220], pgate_l[221],
     pgate_l[218], pgate_l[219], pgate_l[216], pgate_l[217],
     pgate_l[214], pgate_l[215], pgate_l[212], pgate_l[213],
     pgate_l[210], pgate_l[211], pgate_l[208], pgate_l[209],
     pgate_l[206], pgate_l[207], pgate_l[204], pgate_l[205],
     pgate_l[202], pgate_l[203], pgate_l[200], pgate_l[201],
     pgate_l[198], pgate_l[199], pgate_l[196], pgate_l[197],
     pgate_l[194], pgate_l[195], pgate_l[192], pgate_l[193],
     pgate_l[190], pgate_l[191], pgate_l[188], pgate_l[189],
     pgate_l[186], pgate_l[187], pgate_l[184], pgate_l[185],
     pgate_l[182], pgate_l[183], pgate_l[180], pgate_l[181],
     pgate_l[178], pgate_l[179], pgate_l[176], pgate_l[177]}),
     .sdo(net1336));
bram_hbuffer_2xbank I20 ( .bm_wdummymux_en_o(net1658),
     .bm_sweb_i(bm_sweb_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_init_i(bm_init_i), .bm_banksel_o(net1671[0:3]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_o(net1651),
     .bm_sreb_o(net1652), .bm_sclk_o(net1653), .bm_sa_o(net1654[0:7]),
     .bm_init_o(net1655), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclkrw_o(net1664), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sdo_o(bm_sdo_o[3:0]), .bm_sdi_o(net1666[0:3]),
     .bm_rcapmux_en_o(net1657), .bm_banksel_i(bm_banksel_i[3:0]),
     .bm_sdo_i(net1667[0:3]));
bram_hbuffer_dff_2xbank I24 ( .bm_sweb_i(net1651), .bm_sreb_i(net1652),
     .bm_sclk_i(net1653), .bm_sa_i(net1654[0:7]), .bm_init_i(net1655),
     .bm_banksel_o(bm_bank30_banksel_o[3:0]),
     .bm_rcapmux_en_i(net1657), .bm_wdummymux_en_i(net1658),
     .bm_sweb_o(net1674), .bm_sreb_o(net1675),
     .bm_sclk_o(bm_bank30_sclk_o[1:0]), .bm_sa_o(net1678[0:7]),
     .bm_init_o(net1679), .bm_sclkrw_i(net1664), .bm_sclkrw_o(net1690),
     .bm_sdi_i(net1666[0:3]), .bm_sdo_o(net1667[0:3]),
     .bm_sdi_o(bm_bank30_sdi_o[3:0]), .bm_rcapmux_en_o(net1681),
     .bm_wdummymux_en_o(net1682), .bm_banksel_i(net1671[0:3]),
     .bm_sdo_i(bm_bank30_sdo_i[3:0]));
bram_hbuffer_1xbank I17 ( .bm_wdummymux_en_o(net1704),
     .bm_sweb_i(net1674), .bm_sreb_i(net1675),
     .bm_sdi_i(bm_bank30_sdi_o[1:0]), .bm_sclk_i(bm_bank30_sclk_o[0]),
     .bm_sa_i(net1678[0:7]), .bm_init_i(net1679),
     .bm_banksel_o(net1715[0:1]), .bm_rcapmux_en_i(net1681),
     .bm_wdummymux_en_i(net1682), .bm_sweb_o(net1696),
     .bm_sreb_o(net1697), .bm_sdi_o(net1698[0:1]), .bm_sclk_o(net1699),
     .bm_sa_o(net1700[0:7]), .bm_init_o(net1701),
     .bm_rcapmux_en_o(net1703), .bm_sclkrw_i(net1690),
     .bm_sclkrw_o(net1712), .bm_sdo_i(net1716[0:1]),
     .bm_banksel_i(bm_bank30_banksel_o[1:0]),
     .bm_sdo_o(bm_bank30_sdo_i[1:0]));
bram_hbuffer_1xbank I2 ( .bm_wdummymux_en_o(net1291),
     .bm_sweb_i(net1696), .bm_sreb_i(net1697), .bm_sdi_i(net1698[0:1]),
     .bm_sclk_i(net1699), .bm_sa_i(net1700[0:7]), .bm_init_i(net1701),
     .bm_banksel_o(bm_bank10_banksel_o[1:0]),
     .bm_rcapmux_en_i(net1703), .bm_wdummymux_en_i(net1704),
     .bm_sweb_o(net1720), .bm_sreb_o(net1293), .bm_sdi_o(net1289[0:1]),
     .bm_sclk_o(net1295), .bm_sa_o(net1296[0:7]), .bm_init_o(net1297),
     .bm_rcapmux_en_o(net1290), .bm_sclkrw_i(net1712),
     .bm_sclkrw_o(net1719), .bm_sdo_i(net1721[0:1]),
     .bm_banksel_i(net1715[0:1]), .bm_sdo_o(net1716[0:1]));
bram_bank_logic_bot I10 ( .bm_sdo_i(net1379[0:1]), .bm_sclk_i(net1295),
     .bm_sclkrw_i(net1719), .bm_sweb_i(net1720),
     .bm_sdo_o(net1721[0:1]), .bm_sweb_o(net1292[0:1]),
     .bm_sclkrw_o(net1294[0:1]),
     .bm_banksel_i(bm_bank10_banksel_o[1:0]));
bram_bank_logic_bot I21 ( .bm_sdo_i(net866[0:1]),
     .bm_sclk_i(bm_bank30_sclk_o[1]), .bm_sclkrw_i(net1690),
     .bm_sweb_i(net1674), .bm_sdo_o(bm_bank30_sdo_i[3:2]),
     .bm_sweb_o(net867[0:1]), .bm_sclkrw_o(net869[0:1]),
     .bm_banksel_i(bm_bank30_banksel_o[3:2]));
cramrow174bl4 I74 ( .vdd_cntl_l(vdd_cntl_l[351:178]),
     .vdd_cntl_r(vdd_cntl_r[351:178]), .reset_r(reset_b_r[351:178]),
     .pgate_r(pgate_r[351:178]), .wl_l(wl_l[351:178]),
     .reset_l(reset_b_l[351:178]), .pgate_l(pgate_l[351:178]),
     .wl_r(wl_r[351:178]), .bl(bl_top[657:654]));
cramrow174bl4 I75 ( .vdd_cntl_l(vdd_cntl_l[173:0]),
     .vdd_cntl_r(vdd_cntl_r[173:0]), .reset_r(reset_b_r[173:0]),
     .pgate_r(pgate_r[173:0]), .wl_l(wl_l[173:0]),
     .reset_l(reset_b_l[173:0]), .pgate_l(pgate_l[173:0]),
     .wl_r(wl_r[173:0]), .bl(bl_bot[657:654]));
clk_mux2to1x4 I_glb_ck_tree_0 ( .vdd_cntl_l({vdd_cntl_l[176],
     vdd_cntl_l[177]}), .wl_l({wl_l[176], wl_l[177]}),
     .reset_l({reset_b_l[176], reset_b_l[177]}),
     .pgate_l({pgate_l[176], pgate_l[177]}), .pgate_r({pgate_r[176],
     pgate_r[177]}), .wl_r({wl_r[176], wl_r[177]}),
     .reset_r({reset_b_r[176], reset_b_r[177]}),
     .vdd_cntl_r({vdd_cntl_r[176], vdd_cntl_r[177]}),
     .bl(bl_top[657:654]), .prog(prog), .min3({padin_163,
     fabric_out_93}), .min2({padin_30, fabric_out_226}),
     .min1({padin_94, fabric_out_30}), .min0({padin_223,
     fabric_out_163}), .gnet(glb_net[5:2]));
clk_mux2to1x4 I_glb_ck_tree_1 ( .vdd_cntl_l({vdd_cntl_l[174],
     vdd_cntl_l[175]}), .wl_l({wl_l[174], wl_l[175]}),
     .reset_l({reset_b_l[174], reset_b_l[175]}),
     .pgate_l({pgate_l[174], pgate_l[175]}), .pgate_r({pgate_r[174],
     pgate_r[175]}), .wl_r({wl_r[174], wl_r[175]}),
     .reset_r({reset_b_r[174], reset_b_r[175]}),
     .vdd_cntl_r({vdd_cntl_r[174], vdd_cntl_r[175]}),
     .bl(bl_bot[657:654]), .prog(prog), .min3({padin_226,
     fabric_out_162}), .min2({padin_93, fabric_out_34}),
     .min1({padin_34, fabric_out_223}), .min0({padin_162,
     fabric_out_94}), .gnet({glb_net[7], glb_net[6], glb_net[1],
     glb_net[0]}));

endmodule
// Library - io, Cell - PVSSRSSTL, View - schematic
// LAST TIME SAVED: Sep  4 18:59:25 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVSSRSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDDSSTLE, View - schematic
// LAST TIME SAVED: Jul 28 17:16:16 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVDDSSTLE (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVSSSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:17:35 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVSSSSTL ( VSSC );
input  VSSC;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDDSSTLD, View - schematic
// LAST TIME SAVED: Jul 28 17:15:51 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVDDSSTLD ( VDDD, VDDSSTLD );
input  VDDD, VDDSSTLD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDDPSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:15:34 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVDDPSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVSSPSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:17:20 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVSSPSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVREFSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:16:31 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVREFSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVSSSSTLD, View - schematic
// LAST TIME SAVED: Jul 28 17:17:58 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVSSSSTLD ( VSSD );
input  VSSD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVD25POCSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:14:18 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PVD25POCSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_lshv_6v_hold, View - schematic
// LAST TIME SAVED: Dec 20 11:32:52 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_lshv_6v_hold ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M7 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(GND_), .G(vddp_tieh), .S(net132));
nch_25  M15 ( .D(net132), .B(GND_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(GND_), .G(vddp_tieh), .S(net140));
nch_25  M14 ( .D(net140), .B(GND_), .G(sel_25), .S(gnd_));

endmodule
// Library - leafcell, Cell - tiehi, View - schematic
// LAST TIME SAVED: Jul  8 16:18:10 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module tiehi ( tiehi );
output  tiehi;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(net4), .B(gnd_), .G(net4), .S(gnd_));
pch_hvt  M0 ( .D(tiehi), .B(vdd_), .G(net4), .S(vdd_));

endmodule
// Library - io, Cell - PMEMIO, View - schematic
// LAST TIME SAVED: Aug 18 15:53:39 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PMEMIO ( C, NET107, PAD, VREF, A2, A6, DS, I, LVCMOS, OEN, PWD,
     S0, S1 );
output  C;

inout  NET107, PAD, VREF;

input  A2, A6, DS, I, LVCMOS, OEN, PWD, S0, S1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PMEMIO_pair, View - schematic
// LAST TIME SAVED: Aug 18 15:54:04 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module PMEMIO_pair ( c_n, c_p, PAD_n, PAD_p, VREFSSTL,
     .cdsNet0(cbit[14]), .cdsNet0(cbit[13]), .cdsNet0(cbit[12]),
     .cdsNet0(cbit[11]), .cdsNet0(cbit[10]), .cdsNet0(cbit[9]),
     .cdsNet0(cbit[8]), .cdsNet0(cbit[7]), .cdsNet0(cbit[6]),
     .cdsNet0(cbit[5]), .cdsNet0(cbit[4]), .cdsNet0(cbit[3]),
     .cdsNet0(cbit[2]), .cdsNet0(cbit[1]), .cdsNet0(cbit[0]), i_n, i_p,
     oen_n, oen_p );
output  c_n, c_p;

inout  PAD_n, PAD_p, VREFSSTL;

input  i_n, i_p, oen_n, oen_p;

input [0:14]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PMEMIO I50 ( .PAD(PAD_p), .VREF(input_), .NET107(net43), .A6(cbit[8]),
     .A2(cbit[9]), .DS(cbit[10]), .LVCMOS(cbit[11]), .S1(cbit[12]),
     .S0(cbit[13]), .PWD(cbit[14]), .C(c_p), .OEN(oen_p), .I(i_p));
PMEMIO I54 ( .PAD(PAD_n), .VREF(VREFSSTL), .NET107(net107),
     .A6(cbit[0]), .A2(cbit[1]), .DS(cbit[2]), .LVCMOS(cbit[3]),
     .S1(cbit[4]), .S0(cbit[5]), .PWD(cbit[6]), .C(c_n), .OEN(oen_n),
     .I(i_n));
LVDS_con I52 ( .VREF(VREFSSTL), .input_(input_), .cbit_7(cbit[7]),
     .Top_Pad_input(net107));

endmodule
// Library - io, Cell - LB_io, View - schematic
// LAST TIME SAVED: Aug 14 15:23:43 2007
// NETLIST TIME: Nov 14 16:12:05 2008
`timescale 1ns / 1ns 

module LB_io ( in, Pad, VREFSSTL, cbit, oen, out );

inout  VREFSSTL;


output [0:19]  in;

inout [0:19]  Pad;

input [0:19]  out;
input [0:19]  oen;
input [0:149]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PMEMIO_pair I60 ( in[8], in[9], Pad[8], Pad[9], VREFSSTL, cbit[60],
     cbit[61], cbit[62], cbit[63], cbit[64], cbit[65], cbit[66],
     cbit[67], cbit[68], cbit[69], cbit[70], cbit[71], cbit[72],
     cbit[73], cbit[74], out[8], out[9], oen[8], oen[9]);
PMEMIO_pair I61 ( in[10], in[11], Pad[10], Pad[11], VREFSSTL, cbit[75],
     cbit[76], cbit[77], cbit[78], cbit[79], cbit[80], cbit[81],
     cbit[82], cbit[83], cbit[84], cbit[85], cbit[86], cbit[87],
     cbit[88], cbit[89], out[10], out[11], oen[10], oen[11]);
PMEMIO_pair I62 ( in[12], in[13], Pad[12], Pad[13], VREFSSTL, cbit[90],
     cbit[91], cbit[92], cbit[93], cbit[94], cbit[95], cbit[96],
     cbit[97], cbit[98], cbit[99], cbit[100], cbit[101], cbit[102],
     cbit[103], cbit[104], out[12], out[13], oen[12], oen[13]);
PMEMIO_pair I63 ( in[14], in[15], Pad[14], Pad[15], VREFSSTL,
     cbit[105], cbit[106], cbit[107], cbit[108], cbit[109], cbit[110],
     cbit[111], cbit[112], cbit[113], cbit[114], cbit[115], cbit[116],
     cbit[117], cbit[118], cbit[119], out[14], out[15], oen[14],
     oen[15]);
PMEMIO_pair I64 ( in[16], in[17], Pad[16], Pad[17], VREFSSTL,
     cbit[120], cbit[121], cbit[122], cbit[123], cbit[124], cbit[125],
     cbit[126], cbit[127], cbit[128], cbit[129], cbit[130], cbit[131],
     cbit[132], cbit[133], cbit[134], out[16], out[17], oen[16],
     oen[17]);
PMEMIO_pair I65 ( in[18], in[19], Pad[18], Pad[19], VREFSSTL,
     cbit[135], cbit[136], cbit[137], cbit[138], cbit[139], cbit[140],
     cbit[141], cbit[142], cbit[143], cbit[144], cbit[145], cbit[146],
     cbit[147], cbit[148], cbit[149], out[18], out[19], oen[18],
     oen[19]);
PMEMIO_pair I56 ( in[0], in[1], Pad[0], Pad[1], VREFSSTL, cbit[0],
     cbit[1], cbit[2], cbit[3], cbit[4], cbit[5], cbit[6], cbit[7],
     cbit[8], cbit[9], cbit[10], cbit[11], cbit[12], cbit[13],
     cbit[14], out[0], out[1], oen[0], oen[1]);
PMEMIO_pair I57 ( in[2], in[3], Pad[2], Pad[3], VREFSSTL, cbit[15],
     cbit[16], cbit[17], cbit[18], cbit[19], cbit[20], cbit[21],
     cbit[22], cbit[23], cbit[24], cbit[25], cbit[26], cbit[27],
     cbit[28], cbit[29], out[2], out[3], oen[2], oen[3]);
PMEMIO_pair I58 ( in[4], in[5], Pad[4], Pad[5], VREFSSTL, cbit[30],
     cbit[31], cbit[32], cbit[33], cbit[34], cbit[35], cbit[36],
     cbit[37], cbit[38], cbit[39], cbit[40], cbit[41], cbit[42],
     cbit[43], cbit[44], out[4], out[5], oen[4], oen[5]);
PMEMIO_pair I59 ( in[6], in[7], Pad[6], Pad[7], VREFSSTL, cbit[45],
     cbit[46], cbit[47], cbit[48], cbit[49], cbit[50], cbit[51],
     cbit[52], cbit[53], cbit[54], cbit[55], cbit[56], cbit[57],
     cbit[58], cbit[59], out[6], out[7], oen[6], oen[7]);

endmodule
// Library - io, Cell - LT_io, View - schematic
// LAST TIME SAVED: Aug 15 10:58:19 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module LT_io ( in, Pad, VREFSSTL, cbit, oen, out );

inout  VREFSSTL;


output [0:19]  in;

inout [0:19]  Pad;

input [0:149]  cbit;
input [0:19]  oen;
input [0:19]  out;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PMEMIO_pair I60 ( in[8], in[9], Pad[8], Pad[9], VREFSSTL, cbit[60],
     cbit[61], cbit[62], cbit[63], cbit[64], cbit[65], cbit[66],
     cbit[67], cbit[68], cbit[69], cbit[70], cbit[71], cbit[72],
     cbit[73], cbit[74], out[8], out[9], oen[8], oen[9]);
PMEMIO_pair I61 ( in[10], in[11], Pad[10], Pad[11], VREFSSTL, cbit[75],
     cbit[76], cbit[77], cbit[78], cbit[79], cbit[80], cbit[81],
     cbit[82], cbit[83], cbit[84], cbit[85], cbit[86], cbit[87],
     cbit[88], cbit[89], out[10], out[11], oen[10], oen[11]);
PMEMIO_pair I62 ( in[12], in[13], Pad[12], Pad[13], VREFSSTL, cbit[90],
     cbit[91], cbit[92], cbit[93], cbit[94], cbit[95], cbit[96],
     cbit[97], cbit[98], cbit[99], cbit[100], cbit[101], cbit[102],
     cbit[103], cbit[104], out[12], out[13], oen[12], oen[13]);
PMEMIO_pair I63 ( in[14], in[15], Pad[14], Pad[15], VREFSSTL,
     cbit[105], cbit[106], cbit[107], cbit[108], cbit[109], cbit[110],
     cbit[111], cbit[112], cbit[113], cbit[114], cbit[115], cbit[116],
     cbit[117], cbit[118], cbit[119], out[14], out[15], oen[14],
     oen[15]);
PMEMIO_pair I64 ( in[16], in[17], Pad[16], Pad[17], VREFSSTL,
     cbit[120], cbit[121], cbit[122], cbit[123], cbit[124], cbit[125],
     cbit[126], cbit[127], cbit[128], cbit[129], cbit[130], cbit[131],
     cbit[132], cbit[133], cbit[134], out[16], out[17], oen[16],
     oen[17]);
PMEMIO_pair I65 ( in[18], in[19], Pad[18], Pad[19], VREFSSTL,
     cbit[135], cbit[136], cbit[137], cbit[138], cbit[139], cbit[140],
     cbit[141], cbit[142], cbit[143], cbit[144], cbit[145], cbit[146],
     cbit[147], cbit[148], cbit[149], out[18], out[19], oen[18],
     oen[19]);
PMEMIO_pair I56 ( in[0], in[1], Pad[0], Pad[1], VREFSSTL, cbit[0],
     cbit[1], cbit[2], cbit[3], cbit[4], cbit[5], cbit[6], cbit[7],
     cbit[8], cbit[9], cbit[10], cbit[11], cbit[12], cbit[13],
     cbit[14], out[0], out[1], oen[0], oen[1]);
PMEMIO_pair I57 ( in[2], in[3], Pad[2], Pad[3], VREFSSTL, cbit[15],
     cbit[16], cbit[17], cbit[18], cbit[19], cbit[20], cbit[21],
     cbit[22], cbit[23], cbit[24], cbit[25], cbit[26], cbit[27],
     cbit[28], cbit[29], out[2], out[3], oen[2], oen[3]);
PMEMIO_pair I58 ( in[4], in[5], Pad[4], Pad[5], VREFSSTL, cbit[30],
     cbit[31], cbit[32], cbit[33], cbit[34], cbit[35], cbit[36],
     cbit[37], cbit[38], cbit[39], cbit[40], cbit[41], cbit[42],
     cbit[43], cbit[44], out[4], out[5], oen[4], oen[5]);
PMEMIO_pair I59 ( in[6], in[7], Pad[6], Pad[7], VREFSSTL, cbit[45],
     cbit[46], cbit[47], cbit[48], cbit[49], cbit[50], cbit[51],
     cbit[52], cbit[53], cbit[54], cbit[55], cbit[56], cbit[57],
     cbit[58], cbit[59], out[6], out[7], oen[6], oen[7]);

endmodule
// Library - io, Cell - IO_LFTCELL, View - schematic
// LAST TIME SAVED: Sep  4 21:02:48 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module IO_LFTCELL ( in, Pad, VREFSSTL, cbit, oen, out );

inout  VREFSSTL;


output [0:39]  in;

inout [0:39]  Pad;

input [0:39]  oen;
input [299:0]  cbit;
input [0:39]  out;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net34;

wire  [0:1]  net037;

wire  [0:1]  net33;



PVSSRSSTL I42 ( );
PVDDSSTLE I40 ( );
PVSSSSTL I39 ( .VSSC(net032));
PVDDSSTLD I38_1_ ( .VDDSSTLD(net33[0]), .VDDD(net34[0]));
PVDDSSTLD I38_0_ ( .VDDSSTLD(net33[1]), .VDDD(net34[1]));
PVDDPSSTL I37_6_ ( );
PVDDPSSTL I37_5_ ( );
PVDDPSSTL I37_4_ ( );
PVDDPSSTL I37_3_ ( );
PVDDPSSTL I37_2_ ( );
PVDDPSSTL I37_1_ ( );
PVDDPSSTL I37_0_ ( );
PVSSPSSTL I36_7_ ( );
PVSSPSSTL I36_6_ ( );
PVSSPSSTL I36_5_ ( );
PVSSPSSTL I36_4_ ( );
PVSSPSSTL I36_3_ ( );
PVSSPSSTL I36_2_ ( );
PVSSPSSTL I36_1_ ( );
PVSSPSSTL I36_0_ ( );
PVREFSSTL I35 ( );
PVSSSSTLD I33_1_ ( .VSSD(net037[0]));
PVSSSSTLD I33_0_ ( .VSSD(net037[1]));
PVD25POCSSTL I32 ( );
LB_io I31 ( .cbit({cbit[150], cbit[151], cbit[152], cbit[153],
     cbit[154], cbit[155], cbit[156], cbit[157], cbit[158], cbit[159],
     cbit[160], cbit[161], cbit[162], cbit[163], cbit[164], cbit[165],
     cbit[166], cbit[167], cbit[168], cbit[169], cbit[170], cbit[171],
     cbit[172], cbit[173], cbit[174], cbit[175], cbit[176], cbit[177],
     cbit[178], cbit[179], cbit[180], cbit[181], cbit[182], cbit[183],
     cbit[184], cbit[185], cbit[186], cbit[187], cbit[188], cbit[189],
     cbit[190], cbit[191], cbit[192], cbit[193], cbit[194], cbit[195],
     cbit[196], cbit[197], cbit[198], cbit[199], cbit[200], cbit[201],
     cbit[202], cbit[203], cbit[204], cbit[205], cbit[206], cbit[207],
     cbit[208], cbit[209], cbit[210], cbit[211], cbit[212], cbit[213],
     cbit[214], cbit[215], cbit[216], cbit[217], cbit[218], cbit[219],
     cbit[220], cbit[221], cbit[222], cbit[223], cbit[224], cbit[225],
     cbit[226], cbit[227], cbit[228], cbit[229], cbit[230], cbit[231],
     cbit[232], cbit[233], cbit[234], cbit[235], cbit[236], cbit[237],
     cbit[238], cbit[239], cbit[240], cbit[241], cbit[242], cbit[243],
     cbit[244], cbit[245], cbit[246], cbit[247], cbit[248], cbit[249],
     cbit[250], cbit[251], cbit[252], cbit[253], cbit[254], cbit[255],
     cbit[256], cbit[257], cbit[258], cbit[259], cbit[260], cbit[261],
     cbit[262], cbit[263], cbit[264], cbit[265], cbit[266], cbit[267],
     cbit[268], cbit[269], cbit[270], cbit[271], cbit[272], cbit[273],
     cbit[274], cbit[275], cbit[276], cbit[277], cbit[278], cbit[279],
     cbit[280], cbit[281], cbit[282], cbit[283], cbit[284], cbit[285],
     cbit[286], cbit[287], cbit[288], cbit[289], cbit[290], cbit[291],
     cbit[292], cbit[293], cbit[294], cbit[295], cbit[296], cbit[297],
     cbit[298], cbit[299]}), .VREFSSTL(VREFSSTL), .Pad(Pad[20:39]),
     .out(out[20:39]), .oen(oen[20:39]), .in(in[20:39]));
LT_io I30 ( .cbit({cbit[0], cbit[1], cbit[2], cbit[3], cbit[4],
     cbit[5], cbit[6], cbit[7], cbit[8], cbit[9], cbit[10], cbit[11],
     cbit[12], cbit[13], cbit[14], cbit[15], cbit[16], cbit[17],
     cbit[18], cbit[19], cbit[20], cbit[21], cbit[22], cbit[23],
     cbit[24], cbit[25], cbit[26], cbit[27], cbit[28], cbit[29],
     cbit[30], cbit[31], cbit[32], cbit[33], cbit[34], cbit[35],
     cbit[36], cbit[37], cbit[38], cbit[39], cbit[40], cbit[41],
     cbit[42], cbit[43], cbit[44], cbit[45], cbit[46], cbit[47],
     cbit[48], cbit[49], cbit[50], cbit[51], cbit[52], cbit[53],
     cbit[54], cbit[55], cbit[56], cbit[57], cbit[58], cbit[59],
     cbit[60], cbit[61], cbit[62], cbit[63], cbit[64], cbit[65],
     cbit[66], cbit[67], cbit[68], cbit[69], cbit[70], cbit[71],
     cbit[72], cbit[73], cbit[74], cbit[75], cbit[76], cbit[77],
     cbit[78], cbit[79], cbit[80], cbit[81], cbit[82], cbit[83],
     cbit[84], cbit[85], cbit[86], cbit[87], cbit[88], cbit[89],
     cbit[90], cbit[91], cbit[92], cbit[93], cbit[94], cbit[95],
     cbit[96], cbit[97], cbit[98], cbit[99], cbit[100], cbit[101],
     cbit[102], cbit[103], cbit[104], cbit[105], cbit[106], cbit[107],
     cbit[108], cbit[109], cbit[110], cbit[111], cbit[112], cbit[113],
     cbit[114], cbit[115], cbit[116], cbit[117], cbit[118], cbit[119],
     cbit[120], cbit[121], cbit[122], cbit[123], cbit[124], cbit[125],
     cbit[126], cbit[127], cbit[128], cbit[129], cbit[130], cbit[131],
     cbit[132], cbit[133], cbit[134], cbit[135], cbit[136], cbit[137],
     cbit[138], cbit[139], cbit[140], cbit[141], cbit[142], cbit[143],
     cbit[144], cbit[145], cbit[146], cbit[147], cbit[148],
     cbit[149]}), .VREFSSTL(VREFSSTL), .Pad(Pad[0:19]),
     .out(out[0:19]), .oen(oen[0:19]), .in(in[0:19]));

endmodule
// Library - io, Cell - PVSS3DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:17:04 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PVSS3DGZ ( VSS );
input  VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD1DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:14:35 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PVDD1DGZ ( VDD );
input  VDD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD2POC, View - schematic
// LAST TIME SAVED: Jul 28 17:15:17 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PVDD2POC ( VDDPST );
input  VDDPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDD2DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:14:57 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PVDD2DGZ ( VDDPST );
input  VDDPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PDT08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 15:32:26 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PDT08DGZ ( PAD, I, OEN );
inout  PAD;

input  I, OEN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_hv_inv, View - schematic
// LAST TIME SAVED: Jan 21 18:15:24 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_hv_inv ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
pch_25  M39 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - io, Cell - PDIDGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:24:26 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PDIDGZ ( C, PAD );
output  C;

input  PAD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PDUW08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 17:52:32 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PDUW08DGZ ( C, PAD, I, OEN, REN );
output  C;

inout  PAD;

input  I, OEN, REN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - RB_io, View - schematic
// LAST TIME SAVED: Sep  5 14:12:55 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module RB_io ( Tdo, c, Pad, I, OEN, REN, TRSTb, Tck, Tdi, Tms );
output  Tdo;


input  TRSTb, Tck, Tdi, Tms;

output [0:23]  c;

inout [0:19]  Pad;

input [0:19]  REN;
input [0:20]  OEN;
input [0:20]  I;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDT08DGZ I23 ( .PAD(Tdo), .OEN(OEN[0]), .I(I[0]));
PDIDGZ I21 ( .C(c[3]), .PAD(TRSTb));
PDIDGZ I22 ( .C(c[2]), .PAD(Tck));
PDIDGZ I58 ( .C(c[0]), .PAD(Tdi));
PDIDGZ I57 ( .C(c[1]), .PAD(Tms));
PDUW08DGZ I49 ( .PAD(Pad[13]), .C(c[17]), .OEN(OEN[14]), .I(I[14]),
     .REN(REN[13]));
PDUW08DGZ I48 ( .PAD(Pad[14]), .C(c[18]), .OEN(OEN[15]), .I(I[15]),
     .REN(REN[14]));
PDUW08DGZ I36 ( .PAD(Pad[15]), .C(c[19]), .OEN(OEN[16]), .I(I[16]),
     .REN(REN[15]));
PDUW08DGZ I37 ( .PAD(Pad[16]), .C(c[20]), .OEN(OEN[17]), .I(I[17]),
     .REN(REN[16]));
PDUW08DGZ I38 ( .PAD(Pad[17]), .C(c[21]), .OEN(OEN[18]), .I(I[18]),
     .REN(REN[17]));
PDUW08DGZ I39 ( .PAD(Pad[18]), .C(c[22]), .OEN(OEN[19]), .I(I[19]),
     .REN(REN[18]));
PDUW08DGZ I40 ( .PAD(Pad[19]), .C(c[23]), .OEN(OEN[20]), .I(I[20]),
     .REN(REN[19]));
PDUW08DGZ I50 ( .PAD(Pad[12]), .C(c[16]), .OEN(OEN[13]), .I(I[13]),
     .REN(REN[12]));
PDUW08DGZ I44 ( .PAD(Pad[7]), .C(c[11]), .OEN(OEN[8]), .I(I[8]),
     .REN(REN[7]));
PDUW08DGZ I15 ( .PAD(Pad[4]), .C(c[8]), .OEN(OEN[5]), .I(I[5]),
     .REN(REN[4]));
PDUW08DGZ I53 ( .PAD(Pad[2]), .C(c[6]), .OEN(OEN[3]), .I(I[3]),
     .REN(REN[2]));
PDUW08DGZ I54 ( .PAD(Pad[1]), .C(c[5]), .OEN(OEN[2]), .I(I[2]),
     .REN(REN[1]));
PDUW08DGZ I55 ( .PAD(Pad[6]), .C(c[10]), .OEN(OEN[7]), .I(I[7]),
     .REN(REN[6]));
PDUW08DGZ I56 ( .PAD(Pad[0]), .C(c[4]), .OEN(OEN[1]), .I(I[1]),
     .REN(REN[0]));
PDUW08DGZ I51 ( .PAD(Pad[11]), .C(c[15]), .OEN(OEN[12]), .I(I[12]),
     .REN(REN[11]));
PDUW08DGZ I32 ( .PAD(Pad[10]), .C(c[14]), .OEN(OEN[11]), .I(I[11]),
     .REN(REN[10]));
PDUW08DGZ I31 ( .PAD(Pad[9]), .C(c[13]), .OEN(OEN[10]), .I(I[10]),
     .REN(REN[9]));
PDUW08DGZ I52 ( .PAD(Pad[3]), .C(c[7]), .OEN(OEN[4]), .I(I[4]),
     .REN(REN[3]));
PDUW08DGZ I43 ( .PAD(Pad[8]), .C(c[12]), .OEN(OEN[9]), .I(I[9]),
     .REN(REN[8]));
PDUW08DGZ I27 ( .PAD(Pad[5]), .C(c[9]), .OEN(OEN[6]), .I(I[6]),
     .REN(REN[5]));

endmodule
// Library - io, Cell - RT_io, View - schematic
// LAST TIME SAVED: Aug 14 15:21:15 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module RT_io ( c, Pad, I, OEN, REN );



output [0:19]  c;

inout [0:19]  Pad;

input [0:19]  REN;
input [0:19]  I;
input [0:19]  OEN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDUW08DGZ I51 ( .PAD(Pad[19]), .C(c[19]), .OEN(OEN[19]), .I(I[19]),
     .REN(REN[19]));
PDUW08DGZ I32 ( .PAD(Pad[0]), .C(c[0]), .OEN(OEN[0]), .I(I[0]),
     .REN(REN[0]));
PDUW08DGZ I33 ( .PAD(Pad[1]), .C(c[1]), .OEN(OEN[1]), .I(I[1]),
     .REN(REN[1]));
PDUW08DGZ I34 ( .PAD(Pad[2]), .C(c[2]), .OEN(OEN[2]), .I(I[2]),
     .REN(REN[2]));
PDUW08DGZ I35 ( .PAD(Pad[3]), .C(c[3]), .OEN(OEN[3]), .I(I[3]),
     .REN(REN[3]));
PDUW08DGZ I36 ( .PAD(Pad[4]), .C(c[4]), .OEN(OEN[4]), .I(I[4]),
     .REN(REN[4]));
PDUW08DGZ I37 ( .PAD(Pad[5]), .C(c[5]), .OEN(OEN[5]), .I(I[5]),
     .REN(REN[5]));
PDUW08DGZ I38 ( .PAD(Pad[6]), .C(c[6]), .OEN(OEN[6]), .I(I[6]),
     .REN(REN[6]));
PDUW08DGZ I39 ( .PAD(Pad[7]), .C(c[7]), .OEN(OEN[7]), .I(I[7]),
     .REN(REN[7]));
PDUW08DGZ I40 ( .PAD(Pad[8]), .C(c[8]), .OEN(OEN[8]), .I(I[8]),
     .REN(REN[8]));
PDUW08DGZ I41 ( .PAD(Pad[9]), .C(c[9]), .OEN(OEN[9]), .I(I[9]),
     .REN(REN[9]));
PDUW08DGZ I42 ( .PAD(Pad[10]), .C(c[10]), .OEN(OEN[10]), .I(I[10]),
     .REN(REN[10]));
PDUW08DGZ I43 ( .PAD(Pad[11]), .C(c[11]), .OEN(OEN[11]), .I(I[11]),
     .REN(REN[11]));
PDUW08DGZ I44 ( .PAD(Pad[12]), .C(c[12]), .OEN(OEN[12]), .I(I[12]),
     .REN(REN[12]));
PDUW08DGZ I45 ( .PAD(Pad[13]), .C(c[13]), .OEN(OEN[13]), .I(I[13]),
     .REN(REN[13]));
PDUW08DGZ I46 ( .PAD(Pad[14]), .C(c[14]), .OEN(OEN[14]), .I(I[14]),
     .REN(REN[14]));
PDUW08DGZ I47 ( .PAD(Pad[15]), .C(c[15]), .OEN(OEN[15]), .I(I[15]),
     .REN(REN[15]));
PDUW08DGZ I48 ( .PAD(Pad[16]), .C(c[16]), .OEN(OEN[16]), .I(I[16]),
     .REN(REN[16]));
PDUW08DGZ I49 ( .PAD(Pad[17]), .C(c[17]), .OEN(OEN[17]), .I(I[17]),
     .REN(REN[17]));
PDUW08DGZ I50 ( .PAD(Pad[18]), .C(c[18]), .OEN(OEN[18]), .I(I[18]),
     .REN(REN[18]));

endmodule
// Library - io, Cell - IO_RGTCELL, View - schematic
// LAST TIME SAVED: Apr 15 11:04:39 2008
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module IO_RGTCELL ( Tdo, in, Pad, REN, TRSTb, Tck, Tdi, Tms, oen, out
     );
output  Tdo;


input  TRSTb, Tck, Tdi, Tms;

output [0:43]  in;

inout [0:39]  Pad;

input [0:40]  oen;
input [0:40]  out;
input [0:39]  REN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:4]  net39;

wire  [0:3]  net37;

wire  [0:6]  net36;



PVSS3DGZ I37_6_ ( .VSS(net36[0]));
PVSS3DGZ I37_5_ ( .VSS(net36[1]));
PVSS3DGZ I37_4_ ( .VSS(net36[2]));
PVSS3DGZ I37_3_ ( .VSS(net36[3]));
PVSS3DGZ I37_2_ ( .VSS(net36[4]));
PVSS3DGZ I37_1_ ( .VSS(net36[5]));
PVSS3DGZ I37_0_ ( .VSS(net36[6]));
PVDD1DGZ I36_3_ ( .VDD(net37[0]));
PVDD1DGZ I36_2_ ( .VDD(net37[1]));
PVDD1DGZ I36_1_ ( .VDD(net37[2]));
PVDD1DGZ I36_0_ ( .VDD(net37[3]));
PVDD2POC I38 ( .VDDPST(vddp_));
PVDD2POC I35 ( .VDDPST(net38));
PVDD2DGZ I34_4_ ( .VDDPST(net39[0]));
PVDD2DGZ I34_3_ ( .VDDPST(net39[1]));
PVDD2DGZ I34_2_ ( .VDDPST(net39[2]));
PVDD2DGZ I34_1_ ( .VDDPST(net39[3]));
PVDD2DGZ I34_0_ ( .VDDPST(net39[4]));
RB_io I26 ( .OEN(oen[0:20]), .Tdi(Tdi), .REN(REN[0:19]), .I(out[0:20]),
     .c(in[0:23]), .Tdo(Tdo), .Pad(Pad[0:19]), .Tck(Tck), .Tms(Tms),
     .TRSTb(TRSTb));
RT_io I27 ( .I(out[21:40]), .c(in[24:43]), .REN(REN[20:39]),
     .OEN(oen[21:40]), .Pad(Pad[20:39]));

endmodule
// Library - ROCK, Cell - vpp_clamp_finger, View - schematic
// LAST TIME SAVED: Jul 30 12:32:02 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module vpp_clamp_finger ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .B(VSS), .D(net12), .G(VSS), .S(VSS));
nch_25  m1 ( .B(VSS), .D(VPP), .G(VDDIO), .S(net12));

endmodule
// Library - ROCK, Cell - vpp_clamp, View - schematic
// LAST TIME SAVED: Jul 30 12:44:43 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module vpp_clamp ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vpp_clamp_finger I3 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I1 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I2 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I5 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I6 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I7 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I8 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I9 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I4 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));

endmodule
// Library - io, Cell - TL_io, View - schematic
// LAST TIME SAVED: Aug 14 15:21:33 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module TL_io ( in, Pad, I, OEN, REN );



output [0:23]  in;

inout [0:23]  Pad;

input [0:23]  OEN;
input [0:23]  I;
input [0:23]  REN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDUW08DGZ I27 ( .PAD(Pad[20]), .C(in[20]), .REN(REN[20]), .I(I[20]),
     .OEN(OEN[20]));
PDUW08DGZ I52 ( .PAD(Pad[21]), .C(in[21]), .OEN(OEN[21]), .I(I[21]),
     .REN(REN[21]));
PDUW08DGZ I53 ( .PAD(Pad[22]), .C(in[22]), .OEN(OEN[22]), .I(I[22]),
     .REN(REN[22]));
PDUW08DGZ I54 ( .PAD(Pad[23]), .C(in[23]), .OEN(OEN[23]), .I(I[23]),
     .REN(REN[23]));
PDUW08DGZ I41 ( .PAD(Pad[10]), .C(in[10]), .OEN(OEN[10]), .I(I[10]),
     .REN(REN[10]));
PDUW08DGZ I38 ( .PAD(Pad[13]), .C(in[13]), .OEN(OEN[13]), .I(I[13]),
     .REN(REN[13]));
PDUW08DGZ I46 ( .PAD(Pad[5]), .C(in[5]), .OEN(OEN[5]), .I(I[5]),
     .REN(REN[5]));
PDUW08DGZ I45 ( .PAD(Pad[6]), .C(in[6]), .OEN(OEN[6]), .I(I[6]),
     .REN(REN[6]));
PDUW08DGZ I49 ( .PAD(Pad[2]), .C(in[2]), .OEN(OEN[2]), .I(I[2]),
     .REN(REN[2]));
PDUW08DGZ I48 ( .PAD(Pad[3]), .C(in[3]), .OEN(OEN[3]), .I(I[3]),
     .REN(REN[3]));
PDUW08DGZ I33 ( .PAD(Pad[17]), .C(in[17]), .OEN(OEN[17]), .I(I[17]),
     .REN(REN[17]));
PDUW08DGZ I50 ( .PAD(Pad[1]), .C(in[1]), .OEN(OEN[1]), .I(I[1]),
     .REN(REN[1]));
PDUW08DGZ I34 ( .PAD(Pad[18]), .C(in[18]), .OEN(OEN[18]), .I(I[18]),
     .REN(REN[18]));
PDUW08DGZ I36 ( .PAD(Pad[15]), .C(in[15]), .OEN(OEN[15]), .I(I[15]),
     .REN(REN[15]));
PDUW08DGZ I42 ( .PAD(Pad[9]), .C(in[9]), .OEN(OEN[9]), .I(I[9]),
     .REN(REN[9]));
PDUW08DGZ I39 ( .PAD(Pad[12]), .C(in[12]), .OEN(OEN[12]), .I(I[12]),
     .REN(REN[12]));
PDUW08DGZ I44 ( .PAD(Pad[7]), .C(in[7]), .OEN(OEN[7]), .I(I[7]),
     .REN(REN[7]));
PDUW08DGZ I35 ( .PAD(Pad[19]), .C(in[19]), .OEN(OEN[19]), .I(I[19]),
     .REN(REN[19]));
PDUW08DGZ I32 ( .PAD(Pad[16]), .C(in[16]), .OEN(OEN[16]), .I(I[16]),
     .REN(REN[16]));
PDUW08DGZ I37 ( .PAD(Pad[14]), .C(in[14]), .OEN(OEN[14]), .I(I[14]),
     .REN(REN[14]));
PDUW08DGZ I40 ( .PAD(Pad[11]), .C(in[11]), .OEN(OEN[11]), .I(I[11]),
     .REN(REN[11]));
PDUW08DGZ I43 ( .PAD(Pad[8]), .C(in[8]), .OEN(OEN[8]), .I(I[8]),
     .REN(REN[8]));
PDUW08DGZ I47 ( .PAD(Pad[4]), .C(in[4]), .OEN(OEN[4]), .I(I[4]),
     .REN(REN[4]));
PDUW08DGZ I51 ( .PAD(Pad[0]), .C(in[0]), .OEN(OEN[0]), .I(I[0]),
     .REN(REN[0]));

endmodule
// Library - io, Cell - TR_io, View - schematic
// LAST TIME SAVED: Aug 14 15:21:47 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module TR_io ( in, Pad, I, OEN, REN );



output [0:23]  in;

inout [0:23]  Pad;

input [0:23]  REN;
input [0:23]  OEN;
input [0:23]  I;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDUW08DGZ I52 ( .PAD(Pad[23]), .C(in[23]), .OEN(OEN[23]), .I(I[23]),
     .REN(REN[23]));
PDUW08DGZ I54 ( .PAD(Pad[21]), .C(in[21]), .OEN(OEN[21]), .I(I[21]),
     .REN(REN[21]));
PDUW08DGZ I53 ( .PAD(Pad[22]), .C(in[22]), .OEN(OEN[22]), .I(I[22]),
     .REN(REN[22]));
PDUW08DGZ I55 ( .PAD(Pad[20]), .C(in[20]), .OEN(OEN[20]), .I(I[20]),
     .REN(REN[20]));
PDUW08DGZ I41 ( .PAD(Pad[10]), .C(in[10]), .OEN(OEN[10]), .I(I[10]),
     .REN(REN[10]));
PDUW08DGZ I38 ( .PAD(Pad[13]), .C(in[13]), .OEN(OEN[13]), .I(I[13]),
     .REN(REN[13]));
PDUW08DGZ I46 ( .PAD(Pad[5]), .C(in[5]), .OEN(OEN[5]), .I(I[5]),
     .REN(REN[5]));
PDUW08DGZ I45 ( .PAD(Pad[6]), .C(in[6]), .OEN(OEN[6]), .I(I[6]),
     .REN(REN[6]));
PDUW08DGZ I49 ( .PAD(Pad[2]), .C(in[2]), .OEN(OEN[2]), .I(I[2]),
     .REN(REN[2]));
PDUW08DGZ I48 ( .PAD(Pad[3]), .C(in[3]), .OEN(OEN[3]), .I(I[3]),
     .REN(REN[3]));
PDUW08DGZ I33 ( .PAD(Pad[17]), .C(in[17]), .OEN(OEN[17]), .I(I[17]),
     .REN(REN[17]));
PDUW08DGZ I50 ( .PAD(Pad[1]), .C(in[1]), .OEN(OEN[1]), .I(I[1]),
     .REN(REN[1]));
PDUW08DGZ I34 ( .PAD(Pad[18]), .C(in[18]), .OEN(OEN[18]), .I(I[18]),
     .REN(REN[18]));
PDUW08DGZ I36 ( .PAD(Pad[15]), .C(in[15]), .OEN(OEN[15]), .I(I[15]),
     .REN(REN[15]));
PDUW08DGZ I42 ( .PAD(Pad[9]), .C(in[9]), .OEN(OEN[9]), .I(I[9]),
     .REN(REN[9]));
PDUW08DGZ I39 ( .PAD(Pad[12]), .C(in[12]), .OEN(OEN[12]), .I(I[12]),
     .REN(REN[12]));
PDUW08DGZ I44 ( .PAD(Pad[7]), .C(in[7]), .OEN(OEN[7]), .I(I[7]),
     .REN(REN[7]));
PDUW08DGZ I35 ( .PAD(Pad[19]), .C(in[19]), .OEN(OEN[19]), .I(I[19]),
     .REN(REN[19]));
PDUW08DGZ I32 ( .PAD(Pad[16]), .C(in[16]), .OEN(OEN[16]), .I(I[16]),
     .REN(REN[16]));
PDUW08DGZ I37 ( .PAD(Pad[14]), .C(in[14]), .OEN(OEN[14]), .I(I[14]),
     .REN(REN[14]));
PDUW08DGZ I40 ( .PAD(Pad[11]), .C(in[11]), .OEN(OEN[11]), .I(I[11]),
     .REN(REN[11]));
PDUW08DGZ I43 ( .PAD(Pad[8]), .C(in[8]), .OEN(OEN[8]), .I(I[8]),
     .REN(REN[8]));
PDUW08DGZ I47 ( .PAD(Pad[4]), .C(in[4]), .OEN(OEN[4]), .I(I[4]),
     .REN(REN[4]));
PDUW08DGZ I51 ( .PAD(Pad[0]), .C(in[0]), .OEN(OEN[0]), .I(I[0]),
     .REN(REN[0]));

endmodule
// Library - io, Cell - IO_TOPCELL, View - schematic
// LAST TIME SAVED: Apr  7 16:35:38 2008
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module IO_TOPCELL ( in, Pad, vpp, vppin, REN, oen, out );

inout  vpp, vppin;


output [0:47]  in;

inout [0:47]  Pad;

input [0:47]  oen;
input [0:47]  out;
input [47:0]  REN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  net045;

wire  [0:3]  net44;

wire  [0:6]  net046;



rppolywo_m  R8 ( .MINUS(vpp), .PLUS(vppin), .BULK(GND_));
vddp_tiehigh I42 ( .vddp_tieh(net040));
vpp_clamp I41 ( .VSS(gnd_), .VDDIO(net040), .VPP(vpp));
TL_io I31 ( .in(in[24:47]), .I(out[24:47]), .REN({REN[24], REN[25],
     REN[26], REN[27], REN[28], REN[29], REN[30], REN[31], REN[32],
     REN[33], REN[34], REN[35], REN[36], REN[37], REN[38], REN[39],
     REN[40], REN[41], REN[42], REN[43], REN[44], REN[45], REN[46],
     REN[47]}), .Pad(Pad[24:47]), .OEN(oen[24:47]));
TR_io I30 ( .in(in[0:23]), .I(out[0:23]), .REN({REN[0], REN[1], REN[2],
     REN[3], REN[4], REN[5], REN[6], REN[7], REN[8], REN[9], REN[10],
     REN[11], REN[12], REN[13], REN[14], REN[15], REN[16], REN[17],
     REN[18], REN[19], REN[20], REN[21], REN[22], REN[23]}),
     .Pad(Pad[0:23]), .OEN(oen[0:23]));
PVDD2POC I35 ( .VDDPST(net43));
PVDD1DGZ I34_0_ ( .VDD(net44[0]));
PVDD1DGZ I34_1_ ( .VDD(net44[1]));
PVDD1DGZ I34_2_ ( .VDD(net44[2]));
PVDD1DGZ I34_3_ ( .VDD(net44[3]));
PVDD2DGZ I33_2_ ( .VDDPST(net045[0]));
PVDD2DGZ I33_1_ ( .VDDPST(net045[1]));
PVDD2DGZ I33_0_ ( .VDDPST(net045[2]));
PVSS3DGZ I32_6_ ( .VSS(net046[0]));
PVSS3DGZ I32_5_ ( .VSS(net046[1]));
PVSS3DGZ I32_4_ ( .VSS(net046[2]));
PVSS3DGZ I32_3_ ( .VSS(net046[3]));
PVSS3DGZ I32_2_ ( .VSS(net046[4]));
PVSS3DGZ I32_1_ ( .VSS(net046[5]));
PVSS3DGZ I32_0_ ( .VSS(net046[6]));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv, View - schematic
// LAST TIME SAVED: Jan  8 14:11:13 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_hv_ls_inv ( in_hv, out_b_hv, sel_25, sel_b_25, vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_lshv_6v_hold Ishv_6v_hold ( .vddp_tieh(vddp_tieh), .out_b_hv(net61),
     .in_hv(in_hv), .sel_b_25(sel_b_25), .sel_25(sel_25),
     .out_hv(sel_hv));
ml_hv_inv Ihv_inv ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));

endmodule
// Library - io, Cell - PDU08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 17:45:09 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module PDU08DGZ ( C, PAD, I, OEN );
output  C;

inout  PAD;

input  I, OEN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - BR_io, View - schematic
// LAST TIME SAVED: Aug 14 15:22:24 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module BR_io ( c, ctst_b_int, Pad, done, I, OEN, REN, ctst_b );
output  ctst_b_int;

inout  done;

input  ctst_b;

output [0:24]  c;

inout [0:23]  Pad;

input [0:23]  REN;
input [0:24]  OEN;
input [0:24]  I;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDIDGZ I55 ( .C(ctst_b_int), .PAD(ctst_b));
PDU08DGZ I26 ( .C(c[20]), .OEN(OEN[20]), .PAD(done), .I(gnd_));
PDUW08DGZ I27 ( .PAD(Pad[20]), .C(c[21]), .REN(REN[20]), .I(I[21]),
     .OEN(OEN[21]));
PDUW08DGZ I52 ( .PAD(Pad[21]), .C(c[22]), .OEN(OEN[22]), .I(I[22]),
     .REN(REN[21]));
PDUW08DGZ I53 ( .PAD(Pad[22]), .C(c[23]), .OEN(OEN[23]), .I(I[23]),
     .REN(REN[22]));
PDUW08DGZ I54 ( .PAD(Pad[23]), .C(c[24]), .OEN(OEN[24]), .I(I[24]),
     .REN(REN[23]));
PDUW08DGZ I41 ( .PAD(Pad[10]), .C(c[10]), .OEN(OEN[10]), .I(I[10]),
     .REN(REN[10]));
PDUW08DGZ I38 ( .PAD(Pad[13]), .C(c[13]), .OEN(OEN[13]), .I(I[13]),
     .REN(REN[13]));
PDUW08DGZ I46 ( .PAD(Pad[5]), .C(c[5]), .OEN(OEN[5]), .I(I[5]),
     .REN(REN[5]));
PDUW08DGZ I45 ( .PAD(Pad[6]), .C(c[6]), .OEN(OEN[6]), .I(I[6]),
     .REN(REN[6]));
PDUW08DGZ I49 ( .PAD(Pad[2]), .C(c[2]), .OEN(OEN[2]), .I(I[2]),
     .REN(REN[2]));
PDUW08DGZ I48 ( .PAD(Pad[3]), .C(c[3]), .OEN(OEN[3]), .I(I[3]),
     .REN(REN[3]));
PDUW08DGZ I33 ( .PAD(Pad[17]), .C(c[17]), .OEN(OEN[17]), .I(I[17]),
     .REN(REN[17]));
PDUW08DGZ I50 ( .PAD(Pad[1]), .C(c[1]), .OEN(OEN[1]), .I(I[1]),
     .REN(REN[1]));
PDUW08DGZ I34 ( .PAD(Pad[18]), .C(c[18]), .OEN(OEN[18]), .I(I[18]),
     .REN(REN[18]));
PDUW08DGZ I36 ( .PAD(Pad[15]), .C(c[15]), .OEN(OEN[15]), .I(I[15]),
     .REN(REN[15]));
PDUW08DGZ I42 ( .PAD(Pad[9]), .C(c[9]), .OEN(OEN[9]), .I(I[9]),
     .REN(REN[9]));
PDUW08DGZ I39 ( .PAD(Pad[12]), .C(c[12]), .OEN(OEN[12]), .I(I[12]),
     .REN(REN[12]));
PDUW08DGZ I44 ( .PAD(Pad[7]), .C(c[7]), .OEN(OEN[7]), .I(I[7]),
     .REN(REN[7]));
PDUW08DGZ I35 ( .PAD(Pad[19]), .C(c[19]), .OEN(OEN[19]), .I(I[19]),
     .REN(REN[19]));
PDUW08DGZ I32 ( .PAD(Pad[16]), .C(c[16]), .OEN(OEN[16]), .I(I[16]),
     .REN(REN[16]));
PDUW08DGZ I37 ( .PAD(Pad[14]), .C(c[14]), .OEN(OEN[14]), .I(I[14]),
     .REN(REN[14]));
PDUW08DGZ I40 ( .PAD(Pad[11]), .C(c[11]), .OEN(OEN[11]), .I(I[11]),
     .REN(REN[11]));
PDUW08DGZ I43 ( .PAD(Pad[8]), .C(c[8]), .OEN(OEN[8]), .I(I[8]),
     .REN(REN[8]));
PDUW08DGZ I47 ( .PAD(Pad[4]), .C(c[4]), .OEN(OEN[4]), .I(I[4]),
     .REN(REN[4]));
PDUW08DGZ I51 ( .PAD(Pad[0]), .C(c[0]), .OEN(OEN[0]), .I(I[0]),
     .REN(REN[0]));

endmodule
// Library - io, Cell - BL_io, View - schematic
// LAST TIME SAVED: Aug 14 15:22:13 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module BL_io ( c, Pad, I, OEN, REN );



output [0:23]  c;

inout [0:23]  Pad;

input [0:23]  REN;
input [0:23]  OEN;
input [0:23]  I;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDUW08DGZ I52 ( .PAD(Pad[23]), .C(c[23]), .OEN(OEN[23]), .I(I[23]),
     .REN(REN[23]));
PDUW08DGZ I54 ( .PAD(Pad[21]), .C(c[21]), .OEN(OEN[21]), .I(I[21]),
     .REN(REN[21]));
PDUW08DGZ I53 ( .PAD(Pad[22]), .C(c[22]), .OEN(OEN[22]), .I(I[22]),
     .REN(REN[22]));
PDUW08DGZ I55 ( .PAD(Pad[20]), .C(c[20]), .OEN(OEN[20]), .I(I[20]),
     .REN(REN[20]));
PDUW08DGZ I41 ( .PAD(Pad[10]), .C(c[10]), .OEN(OEN[10]), .I(I[10]),
     .REN(REN[10]));
PDUW08DGZ I38 ( .PAD(Pad[13]), .C(c[13]), .OEN(OEN[13]), .I(I[13]),
     .REN(REN[13]));
PDUW08DGZ I46 ( .PAD(Pad[5]), .C(c[5]), .OEN(OEN[5]), .I(I[5]),
     .REN(REN[5]));
PDUW08DGZ I45 ( .PAD(Pad[6]), .C(c[6]), .OEN(OEN[6]), .I(I[6]),
     .REN(REN[6]));
PDUW08DGZ I49 ( .PAD(Pad[2]), .C(c[2]), .OEN(OEN[2]), .I(I[2]),
     .REN(REN[2]));
PDUW08DGZ I48 ( .PAD(Pad[3]), .C(c[3]), .OEN(OEN[3]), .I(I[3]),
     .REN(REN[3]));
PDUW08DGZ I33 ( .PAD(Pad[17]), .C(c[17]), .OEN(OEN[17]), .I(I[17]),
     .REN(REN[17]));
PDUW08DGZ I50 ( .PAD(Pad[1]), .C(c[1]), .OEN(OEN[1]), .I(I[1]),
     .REN(REN[1]));
PDUW08DGZ I34 ( .PAD(Pad[18]), .C(c[18]), .OEN(OEN[18]), .I(I[18]),
     .REN(REN[18]));
PDUW08DGZ I36 ( .PAD(Pad[15]), .C(c[15]), .OEN(OEN[15]), .I(I[15]),
     .REN(REN[15]));
PDUW08DGZ I42 ( .PAD(Pad[9]), .C(c[9]), .OEN(OEN[9]), .I(I[9]),
     .REN(REN[9]));
PDUW08DGZ I39 ( .PAD(Pad[12]), .C(c[12]), .OEN(OEN[12]), .I(I[12]),
     .REN(REN[12]));
PDUW08DGZ I44 ( .PAD(Pad[7]), .C(c[7]), .OEN(OEN[7]), .I(I[7]),
     .REN(REN[7]));
PDUW08DGZ I35 ( .PAD(Pad[19]), .C(c[19]), .OEN(OEN[19]), .I(I[19]),
     .REN(REN[19]));
PDUW08DGZ I32 ( .PAD(Pad[16]), .C(c[16]), .OEN(OEN[16]), .I(I[16]),
     .REN(REN[16]));
PDUW08DGZ I37 ( .PAD(Pad[14]), .C(c[14]), .OEN(OEN[14]), .I(I[14]),
     .REN(REN[14]));
PDUW08DGZ I40 ( .PAD(Pad[11]), .C(c[11]), .OEN(OEN[11]), .I(I[11]),
     .REN(REN[11]));
PDUW08DGZ I43 ( .PAD(Pad[8]), .C(c[8]), .OEN(OEN[8]), .I(I[8]),
     .REN(REN[8]));
PDUW08DGZ I47 ( .PAD(Pad[4]), .C(c[4]), .OEN(OEN[4]), .I(I[4]),
     .REN(REN[4]));
PDUW08DGZ I51 ( .PAD(Pad[0]), .C(c[0]), .OEN(OEN[0]), .I(I[0]),
     .REN(REN[0]));

endmodule
// Library - io, Cell - IO_BOTCELL, View - schematic
// LAST TIME SAVED: Aug 14 14:21:13 2007
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module IO_BOTCELL ( ctst_b_int, in, Pad, done, REN, ctst_b, oen, out );
output  ctst_b_int;

inout  done;

input  ctst_b;

output [0:48]  in;

inout [0:47]  Pad;

input [0:48]  oen;
input [0:47]  REN;
input [0:48]  out;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net043;

wire  [0:1]  net044;

wire  [0:2]  net42;

wire  [0:5]  net45;



PVDD1DGZ Ivdd1_2_ ( .VDD(net42[0]));
PVDD1DGZ Ivdd1_1_ ( .VDD(net42[1]));
PVDD1DGZ Ivdd1_0_ ( .VDD(net42[2]));
PVDD2DGZ I35_1_ ( .VDDPST(net043[0]));
PVDD2DGZ I35_0_ ( .VDDPST(net043[1]));
PVDD2POC I36_1_ ( .VDDPST(net044[0]));
PVDD2POC I36_0_ ( .VDDPST(net044[1]));
PVSS3DGZ I37_5_ ( .VSS(net45[0]));
PVSS3DGZ I37_4_ ( .VSS(net45[1]));
PVSS3DGZ I37_3_ ( .VSS(net45[2]));
PVSS3DGZ I37_2_ ( .VSS(net45[3]));
PVSS3DGZ I37_1_ ( .VSS(net45[4]));
PVSS3DGZ I37_0_ ( .VSS(net45[5]));
BR_io Ibr_io ( .Pad(Pad[24:47]), .c(in[24:48]), .I(out[24:48]),
     .ctst_b_int(ctst_b_int), .ctst_b(ctst_b), .done(done),
     .REN(REN[24:47]), .OEN(oen[24:48]));
BL_io Ibl_io ( .I(out[0:23]), .REN(REN[0:23]), .c(in[0:23]),
     .Pad(Pad[0:23]), .OEN(oen[0:23]));

endmodule
// Library - ice4chip, Cell - chip_ice4f, View - schematic
// LAST TIME SAVED: Oct  7 18:00:24 2008
// NETLIST TIME: Nov 14 16:12:06 2008
`timescale 1ns / 1ns 

module chip_ice4f ( tdo, cdone, uio_bbank, uio_lbank, uio_rbank,
     uio_tbank, vpp, VREFSSTL, creset_b, tck, tdi, tms, trstb );

output  tdo;

inout  cdone, vpp;

input  VREFSSTL, creset_b, tck, tdi, tms, trstb;

inout [39:0]  uio_lbank;
inout [0:47]  uio_bbank;
inout [47:0]  uio_tbank;
inout [0:39]  uio_rbank;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  cm_banksel_blbld1;

wire  [47:0]  oen_tbank;

wire  [1:1]  cm_banksel_bltld3;

wire  [47:0]  out_tbank;

wire  [3:0]  bm_sdo_o;

wire  [39:0]  out_lbank;

wire  [1:0]  cm_sdi_u1d;

wire  [1:0]  cm_banksel;

wire  [351:0]  wl_l;

wire  [3:3]  cm_banksel_bltrd1;

wire  [39:0]  oen_lbank;

wire  [39:0]  in_rbank;

wire  [39:0]  out_rbank;

wire  [39:0]  oeb_rbank;

wire  [3:0]  bm_banksel_i;

wire  [351:0]  pgate_l;

wire  [351:0]  vdd_cntl_l;

wire  [7:0]  bm_sa_i;

wire  [479:0]  cf_rbank;

wire  [1:0]  cm_sdi_u1;

wire  [1:0]  monitor_celld2;

wire  [1311:0]  bl_bot;

wire  [3:0]  bm_sdi_i;

wire  [42:47]  spi_ss_in_bbankd;

wire  [351:0]  vdd_cntl_r;

wire  [351:0]  reset_l;

wire  [1:0]  cm_sdi_u1d3;

wire  [1311:0]  bl_top;

wire  [1:0]  cm_sdo_u1;

wire  [39:0]  spi_ss_in_r;

wire  [1:0]  cm_sdo_u3;

wire  [1:0]  cm_sdi_u3d2;

wire  [575:0]  cf_tbank;

wire  [7:1]  psdo;

wire  [1:0]  cm_sdi_u2d;

wire  [1:0]  cm_sdo_u2d1;

wire  [47:24]  spi_ss_in_bbank;

wire  [1:0]  cm_sdo_u1d3;

wire  [2:2]  cm_banksel_blbrd;

wire  [575:0]  cf_bbank;

wire  [1:0]  monitor_celld4;

wire  [1:0]  cm_sdi_u0;

wire  [351:0]  pgate_r;

wire  [47:0]  in_bbank;

wire  [1:0]  cm_sdo_u1d1;

wire  [1:0]  cm_sdo_u0d1;

wire  [39:0]  in_lbank;

wire  [0:19]  net419;

wire  [47:0]  out_bbank;

wire  [47:0]  oen_bbank;

wire  [1:1]  cm_banksel_blbld;

wire  [0:3]  last_rsr;

wire  [47:0]  in_tbank;

wire  [351:0]  wl_r;

wire  [0:479]  cf_lbank;

wire  [351:0]  reset_b_r;



CHIP_route_right_ice4f_guc Ismc_chip_rout_right (
     .nvcm_spi_sdo(nvcm_spi_sdo),
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_relextspi(nvcm_relextspi), .nvcm_rdy(nvcm_rdy),
     .nvcm_boot(nvcm_boot), .bp0(bp0), .smc_load_nvcm_bstream(net082),
     .nvcm_spi_sdi(net081), .nvcm_spi_ss_b(net080), .rst_b(net083),
     .ceb0(ceb), .spi_ss_in_r(spi_ss_in_r[7:1]),
     .smc_write0(smc_write), .cm_banksel_bldld(cm_banksel[1:0]),
     .cm_banksel_bltrd1_3_(cm_banksel_bltrd1[3]),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd[2]), .last_rsr({last_rsr[3],
     last_rsr[2]}), .spi_ss_in_bbank({spi_ss_in_bbankd[47],
     spi_ss_in_bbankd[46], spi_ss_in_bbankd[45], spi_ss_in_bbankd[43],
     spi_ss_in_bbankd[42]}), .cf_r({cf_rbank[479], cf_rbank[40]}),
     .core_por_b_rowu2(core_por_b_rowu2), .core_por_b0(core_por_b0),
     .row_test0(row_test0), .smc_row_inc(smc_row_inc),
     .cram_pgateoff(cram_pgateoff), .core_por_bb(core_por_bb),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .smc_rsr_rst(smc_rsr_rst), .j_rst_b(j_rst_b),
     .smc_wdis_dclk_bltrd1(smc_wdis_dclk_bltrd1),
     .cram_prec_blbrd(cram_prec_blbrd),
     .cram_pullup_b_blbrd(cram_pullup_b_blbrd),
     .cram_write_blbrd(cram_write_blbrd),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .cm_clk_blbrd(cm_clk_blbrd),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .smc_wdis_dclk(smc_wdis_dclk), .smc_clk_out(smc_clk_out),
     .en_8bconfig_b(en_8bconfig_b), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel), .cram_write(cram_write),
     .cram_prec(cram_prec), .cram_pullup_b(cram_pullup_b),
     .last_rsr3(last_rsr3), .core_por_b_rowu3(core_por_b_rowu3),
     .pgate_r(pgate_r[351:0]), .reset_b_r(reset_b_r[351:0]),
     .vdd_cntl_r(vdd_cntl_r[351:0]), .wl_r(wl_r[351:0]),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .cm_sdo_u3(cm_sdo_u3[1:0]), .fabric_out_126(fabric_out_126),
     .fabric_out_122(fabric_out_122), .vddio_rightbank(vddp_),
     .trst_pad(trst_pad), .tms_pad(tms_pad), .tdi_pad(tdi_pad),
     .tck_pad(tck_pad), .monitor_celld4(monitor_celld4[1:0]),
     .fromsdo(fromsdo), .fabric_out_136(fabric_out_136),
     .crst_filterout(crst_filterout), .cm_sdo_u2d1(cm_sdo_u2d1[1:0]),
     .cm_sdo_u1d3(cm_sdo_u1d3[1:0]), .cm_sdo_u0d1(cm_sdo_u0d1[1:0]),
     .cdone_in(cdone_in), .bm_sdo_o(bm_sdo_o[3:0]), .update0(update0),
     .totdopad(totdopad), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .spi_clk_out(spi_clk_out), .shift0(shift0),
     .sdo_enable(sdo_enable), .psdo(psdo[7:1]), .mode0(mode0),
     .md_spi_b(md_spi_b),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .j_tdi(j_tdi), .j_tck(j_tck), .hiz_b0(hiz_b0), .gsr(gsr),
     .gint_hz(gint_hz), .end_of_startup(end_of_startup),
     .en_8bcibfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel1_bltrd1(data_muxsel1_bltrd1),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1), .core_por_b1(core_por_b1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .cm_clk_bltrd1(cm_clk_bltrd1), .cdone_out(cdone_out),
     .bs_en0(bs_en0), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sweb_i(bm_sweb_i), .bm_sreb_i(bm_sreb_i),
     .bm_sdi_i(bm_sdi_i[3:0]), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bm_banksel_i(bm_banksel_i[3:0]),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b));
sg_bufx10 I215 ( .in(spi_clk_out), .out(spi_clk_out2fsm));
nvcm_ml_block Invcm_fsm ( .smc_load_nvcm_bstream(net082),
     .nvcm_relextspi(nvcm_relextspi), .spi_ss_b(net080),
     .spi_sdi(net081), .rst_b(net083), .nvcm_ce_b(end_of_startup),
     .icef_member_sel({tiegnd, tievdd}), .clk(spi_clk_out2fsm),
     .spi_sdo_oe_b(nvcm_spi_sdo_oe_b), .spi_sdo(nvcm_spi_sdo),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .fsm_tm_margin0_read(net093), .fsm_recall(net094), .bp0(bp0),
     .vpp(vppin));
CHIP_route_left Ichip_route_left ( cm_banksel_bltld3[1], cm_clk_bltld3,
     cm_sdi_u1d3[1:0], cm_sdo_u1d1[1:0], core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_b_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, {last_rsr[1], last_rsr[0]},
     monitor_celld2[1:0], pgate_l[351:0], reset_l[351:0],
     smc_wdis_dclk_bltld3r, vdd_cntl_l[351:0], wl_l[351:0],
     cf_lbank[300], cf_lbank[479], cm_banksel_blbld1[0],
     cm_banksel_blbld[1], cm_clk_blbld, cm_sdi_u1d[1:0],
     cm_sdo_u1[1:0], core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0);
CHIP_route_bot Ichip_route_bot (
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .vddio_spi(vddio_spi), .vddio_botbank(vddio_bottombank),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd[2]),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1[0]),
     .cm_banksel_blbld_1_(cm_banksel_blbld[1]), .j_rst_b(j_rst_b),
     .spi_ss_in_bbankd({spi_ss_in_bbankd[47], spi_ss_in_bbankd[46],
     spi_ss_in_bbankd[45], spi_ss_in_bbankd[43],
     spi_ss_in_bbankd[42]}), .spi_ss_in_bbank({spi_ss_in_bbank[47],
     spi_ss_in_bbank[46], spi_ss_in_bbank[45], spi_ss_in_bbank[43],
     spi_ss_in_bbank[42]}), .cm_banksel(cm_banksel[1:0]),
     .monitor_celld2(monitor_celld2[1:0]),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .cram_write_blbld(cram_write_blbld),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld), .cm_clk_blbld(cm_clk_blbld),
     .cram_pullup_b(cram_pullup_b), .cram_write(cram_write),
     .cm_sdi_u2d(cm_sdi_u2d[1:0]), .smc_clk_out(smc_clk_out),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .cm_clk_blbrd(cm_clk_blbrd), .cram_write_blbrd(cram_write_blbrd),
     .cram_pullup_b_blbrd(cram_pullup_b_blbrd),
     .cram_prec_blbrd(cram_prec_blbrd), .bl_bot(bl_bot[1311:0]),
     .smc_write(smc_write), .smc_wdis_dclk(smc_wdis_dclk),
     .smc_rsr_rst(smc_rsr_rst), .smc_row_inc(smc_row_inc),
     .row_test0(row_test0), .last_rsr1(last_rsr0), .j_tck(j_tck),
     .en_8bconfig_b(en_8bconfig_b), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel), .creset_b_int(creset_b_int),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .cram_prec(cram_prec),
     .cram_pgateoff(cram_pgateoff), .core_por_rowu0(core_por_b_rowu0),
     .core_por_bb(core_por_bb), .core_por_b_rowu2(core_por_b_rowu2),
     .core_por_b0(core_por_b0), .cm_sdo_u1d1(cm_sdo_u1d1[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .tck_padl0(tck_padl0), .smc_writel0(smc_writel0),
     .smc_rsr_rstl0(smc_rsr_rstl0), .smc_row_incl0(smc_row_incl0),
     .row_testl1(row_testl1), .monitor_celld4(monitor_celld4[1:0]),
     .last_rsr3(last_rsr3), .j_rst_bl0(j_rst_bl0),
     .crst_filterout(crst_filterout), .cram_wl_enl0(cram_wl_enl0),
     .cram_vddoffl0(cram_vddoffl0), .cram_rstl0(cram_rstl0),
     .cram_pgateoffl0(cram_pgateoffl0), .core_por_bbl0(core_por_bbl0),
     .core_por_b2(core_por_b2), .cm_sdo_u2d1(cm_sdo_u2d1[1:0]),
     .cm_sdo_u1d3(cm_sdo_u1d3[1:0]), .cm_sdo_u0d1(cm_sdo_u0d1[1:0]),
     .cm_sdi_u1d(cm_sdi_u1d[1:0]));
CHIP_route_top Ichip_route_top (
     .data_muxsel1_bltrd1(data_muxsel1_bltrd1),
     .bl_top(bl_top[1311:0]),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3r),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltld3),
     .data_muxsel1_bltld3(data_muxsel1_bltld3),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_b_bltld3),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1),
     .core_por_b_rowu3(core_por_b_rowu3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .cm_prec_bltld3(cram_prec_bltld3), .cm_clk_bltrd1(cm_clk_bltrd1),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cm_banksel_bltrd1(cm_banksel_bltrd1[3]),
     .cm_banksel_bltld3(cm_banksel_bltld3[1]),
     .cm_sdo_u3(cm_sdo_u3[1:0]), .cm_sdo_u1(cm_sdo_u1[1:0]));
PRCUTSSTLSTDR I40cutr ( .VSS(gnd_), .VSSPST(gnd_));
PRCUTSSTLSTDL I40cutl ( .VSS(gnd_), .VSSPST(gnd_));
tielo4x I459 ( .tielo(tiegnd));
tiehi4x I458 ( .tiehi(tievdd));
QUAD_x4 I445 ( .ceb(ceb), .tiegnd(tiegnd), .tievdd(tievdd),
     .fabric_out_126(fabric_out_126), .fabric_out_136(fabric_out_136),
     .fabric_out_122(fabric_out_122), .spi_ss_in_lft_b(net419[0:19]),
     .spiout_lft_b({tiegnd, tiegnd, last_rsr[1], tiegnd, last_rsr[0],
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .spioeb_lft_b({tievdd, tievdd, tiegnd, tievdd, tiegnd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .bm_banksel_i(bm_banksel_i[3:0]), .spiout_b({spi_ss_out_b,
     spi_clk_out, tiegnd, spi_sdo, tiegnd, tiegnd, psdo[7:2], tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd}), .cdone_in_bot_r({end_of_startup,
     end_of_startup, end_of_startup, en_8bconfig_b, en_8bconfig_b,
     en_8bconfig_b, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .spi_ss_in_b(spi_ss_in_bbank[47:24]), .spioeb_b({md_spi_b,
     md_spi_b, tievdd, spi_sdo_oe_b, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .spiout_r({tiegnd, tiegnd, last_rsr[3], tiegnd, last_rsr[2],
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, psdo[1]}),
     .end_of_startup_t({tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd}), .padin_t(in_tbank[47:0]),
     .padin_l(in_lbank[39:0]), .vdd_cntl_l({vdd_cntl_l[176],
     vdd_cntl_l[177], vdd_cntl_l[178], vdd_cntl_l[179],
     vdd_cntl_l[180], vdd_cntl_l[181], vdd_cntl_l[182],
     vdd_cntl_l[183], vdd_cntl_l[184], vdd_cntl_l[185],
     vdd_cntl_l[186], vdd_cntl_l[187], vdd_cntl_l[188],
     vdd_cntl_l[189], vdd_cntl_l[190], vdd_cntl_l[191],
     vdd_cntl_l[192], vdd_cntl_l[193], vdd_cntl_l[194],
     vdd_cntl_l[195], vdd_cntl_l[196], vdd_cntl_l[197],
     vdd_cntl_l[198], vdd_cntl_l[199], vdd_cntl_l[200],
     vdd_cntl_l[201], vdd_cntl_l[202], vdd_cntl_l[203],
     vdd_cntl_l[204], vdd_cntl_l[205], vdd_cntl_l[206],
     vdd_cntl_l[207], vdd_cntl_l[208], vdd_cntl_l[209],
     vdd_cntl_l[210], vdd_cntl_l[211], vdd_cntl_l[212],
     vdd_cntl_l[213], vdd_cntl_l[214], vdd_cntl_l[215],
     vdd_cntl_l[216], vdd_cntl_l[217], vdd_cntl_l[218],
     vdd_cntl_l[219], vdd_cntl_l[220], vdd_cntl_l[221],
     vdd_cntl_l[222], vdd_cntl_l[223], vdd_cntl_l[224],
     vdd_cntl_l[225], vdd_cntl_l[226], vdd_cntl_l[227],
     vdd_cntl_l[228], vdd_cntl_l[229], vdd_cntl_l[230],
     vdd_cntl_l[231], vdd_cntl_l[232], vdd_cntl_l[233],
     vdd_cntl_l[234], vdd_cntl_l[235], vdd_cntl_l[236],
     vdd_cntl_l[237], vdd_cntl_l[238], vdd_cntl_l[239],
     vdd_cntl_l[240], vdd_cntl_l[241], vdd_cntl_l[242],
     vdd_cntl_l[243], vdd_cntl_l[244], vdd_cntl_l[245],
     vdd_cntl_l[246], vdd_cntl_l[247], vdd_cntl_l[248],
     vdd_cntl_l[249], vdd_cntl_l[250], vdd_cntl_l[251],
     vdd_cntl_l[252], vdd_cntl_l[253], vdd_cntl_l[254],
     vdd_cntl_l[255], vdd_cntl_l[256], vdd_cntl_l[257],
     vdd_cntl_l[258], vdd_cntl_l[259], vdd_cntl_l[260],
     vdd_cntl_l[261], vdd_cntl_l[262], vdd_cntl_l[263],
     vdd_cntl_l[264], vdd_cntl_l[265], vdd_cntl_l[266],
     vdd_cntl_l[267], vdd_cntl_l[268], vdd_cntl_l[269],
     vdd_cntl_l[270], vdd_cntl_l[271], vdd_cntl_l[272],
     vdd_cntl_l[273], vdd_cntl_l[274], vdd_cntl_l[275],
     vdd_cntl_l[276], vdd_cntl_l[277], vdd_cntl_l[278],
     vdd_cntl_l[279], vdd_cntl_l[280], vdd_cntl_l[281],
     vdd_cntl_l[282], vdd_cntl_l[283], vdd_cntl_l[284],
     vdd_cntl_l[285], vdd_cntl_l[286], vdd_cntl_l[287],
     vdd_cntl_l[288], vdd_cntl_l[289], vdd_cntl_l[290],
     vdd_cntl_l[291], vdd_cntl_l[292], vdd_cntl_l[293],
     vdd_cntl_l[294], vdd_cntl_l[295], vdd_cntl_l[296],
     vdd_cntl_l[297], vdd_cntl_l[298], vdd_cntl_l[299],
     vdd_cntl_l[300], vdd_cntl_l[301], vdd_cntl_l[302],
     vdd_cntl_l[303], vdd_cntl_l[304], vdd_cntl_l[305],
     vdd_cntl_l[306], vdd_cntl_l[307], vdd_cntl_l[308],
     vdd_cntl_l[309], vdd_cntl_l[310], vdd_cntl_l[311],
     vdd_cntl_l[312], vdd_cntl_l[313], vdd_cntl_l[314],
     vdd_cntl_l[315], vdd_cntl_l[316], vdd_cntl_l[317],
     vdd_cntl_l[318], vdd_cntl_l[319], vdd_cntl_l[320],
     vdd_cntl_l[321], vdd_cntl_l[322], vdd_cntl_l[323],
     vdd_cntl_l[324], vdd_cntl_l[325], vdd_cntl_l[326],
     vdd_cntl_l[327], vdd_cntl_l[328], vdd_cntl_l[329],
     vdd_cntl_l[330], vdd_cntl_l[331], vdd_cntl_l[332],
     vdd_cntl_l[333], vdd_cntl_l[334], vdd_cntl_l[335],
     vdd_cntl_l[336], vdd_cntl_l[337], vdd_cntl_l[338],
     vdd_cntl_l[339], vdd_cntl_l[340], vdd_cntl_l[341],
     vdd_cntl_l[342], vdd_cntl_l[343], vdd_cntl_l[344],
     vdd_cntl_l[345], vdd_cntl_l[346], vdd_cntl_l[347],
     vdd_cntl_l[348], vdd_cntl_l[349], vdd_cntl_l[350],
     vdd_cntl_l[351], vdd_cntl_l[175], vdd_cntl_l[174],
     vdd_cntl_l[173], vdd_cntl_l[172], vdd_cntl_l[171],
     vdd_cntl_l[170], vdd_cntl_l[169], vdd_cntl_l[168],
     vdd_cntl_l[167], vdd_cntl_l[166], vdd_cntl_l[165],
     vdd_cntl_l[164], vdd_cntl_l[163], vdd_cntl_l[162],
     vdd_cntl_l[161], vdd_cntl_l[160], vdd_cntl_l[159],
     vdd_cntl_l[158], vdd_cntl_l[157], vdd_cntl_l[156],
     vdd_cntl_l[155], vdd_cntl_l[154], vdd_cntl_l[153],
     vdd_cntl_l[152], vdd_cntl_l[151], vdd_cntl_l[150],
     vdd_cntl_l[149], vdd_cntl_l[148], vdd_cntl_l[147],
     vdd_cntl_l[146], vdd_cntl_l[145], vdd_cntl_l[144],
     vdd_cntl_l[143], vdd_cntl_l[142], vdd_cntl_l[141],
     vdd_cntl_l[140], vdd_cntl_l[139], vdd_cntl_l[138],
     vdd_cntl_l[137], vdd_cntl_l[136], vdd_cntl_l[135],
     vdd_cntl_l[134], vdd_cntl_l[133], vdd_cntl_l[132],
     vdd_cntl_l[131], vdd_cntl_l[130], vdd_cntl_l[129],
     vdd_cntl_l[128], vdd_cntl_l[127], vdd_cntl_l[126],
     vdd_cntl_l[125], vdd_cntl_l[124], vdd_cntl_l[123],
     vdd_cntl_l[122], vdd_cntl_l[121], vdd_cntl_l[120],
     vdd_cntl_l[119], vdd_cntl_l[118], vdd_cntl_l[117],
     vdd_cntl_l[116], vdd_cntl_l[115], vdd_cntl_l[114],
     vdd_cntl_l[113], vdd_cntl_l[112], vdd_cntl_l[111],
     vdd_cntl_l[110], vdd_cntl_l[109], vdd_cntl_l[108],
     vdd_cntl_l[107], vdd_cntl_l[106], vdd_cntl_l[105],
     vdd_cntl_l[104], vdd_cntl_l[103], vdd_cntl_l[102],
     vdd_cntl_l[101], vdd_cntl_l[100], vdd_cntl_l[99], vdd_cntl_l[98],
     vdd_cntl_l[97], vdd_cntl_l[96], vdd_cntl_l[95], vdd_cntl_l[94],
     vdd_cntl_l[93], vdd_cntl_l[92], vdd_cntl_l[91], vdd_cntl_l[90],
     vdd_cntl_l[89], vdd_cntl_l[88], vdd_cntl_l[87], vdd_cntl_l[86],
     vdd_cntl_l[85], vdd_cntl_l[84], vdd_cntl_l[83], vdd_cntl_l[82],
     vdd_cntl_l[81], vdd_cntl_l[80], vdd_cntl_l[79], vdd_cntl_l[78],
     vdd_cntl_l[77], vdd_cntl_l[76], vdd_cntl_l[75], vdd_cntl_l[74],
     vdd_cntl_l[73], vdd_cntl_l[72], vdd_cntl_l[71], vdd_cntl_l[70],
     vdd_cntl_l[69], vdd_cntl_l[68], vdd_cntl_l[67], vdd_cntl_l[66],
     vdd_cntl_l[65], vdd_cntl_l[64], vdd_cntl_l[63], vdd_cntl_l[62],
     vdd_cntl_l[61], vdd_cntl_l[60], vdd_cntl_l[59], vdd_cntl_l[58],
     vdd_cntl_l[57], vdd_cntl_l[56], vdd_cntl_l[55], vdd_cntl_l[54],
     vdd_cntl_l[53], vdd_cntl_l[52], vdd_cntl_l[51], vdd_cntl_l[50],
     vdd_cntl_l[49], vdd_cntl_l[48], vdd_cntl_l[47], vdd_cntl_l[46],
     vdd_cntl_l[45], vdd_cntl_l[44], vdd_cntl_l[43], vdd_cntl_l[42],
     vdd_cntl_l[41], vdd_cntl_l[40], vdd_cntl_l[39], vdd_cntl_l[38],
     vdd_cntl_l[37], vdd_cntl_l[36], vdd_cntl_l[35], vdd_cntl_l[34],
     vdd_cntl_l[33], vdd_cntl_l[32], vdd_cntl_l[31], vdd_cntl_l[30],
     vdd_cntl_l[29], vdd_cntl_l[28], vdd_cntl_l[27], vdd_cntl_l[26],
     vdd_cntl_l[25], vdd_cntl_l[24], vdd_cntl_l[23], vdd_cntl_l[22],
     vdd_cntl_l[21], vdd_cntl_l[20], vdd_cntl_l[19], vdd_cntl_l[18],
     vdd_cntl_l[17], vdd_cntl_l[16], vdd_cntl_l[15], vdd_cntl_l[14],
     vdd_cntl_l[13], vdd_cntl_l[12], vdd_cntl_l[11], vdd_cntl_l[10],
     vdd_cntl_l[9], vdd_cntl_l[8], vdd_cntl_l[7], vdd_cntl_l[6],
     vdd_cntl_l[5], vdd_cntl_l[4], vdd_cntl_l[3], vdd_cntl_l[2],
     vdd_cntl_l[1], vdd_cntl_l[0]}), .wl_l({wl_l[176], wl_l[177],
     wl_l[178], wl_l[179], wl_l[180], wl_l[181], wl_l[182], wl_l[183],
     wl_l[184], wl_l[185], wl_l[186], wl_l[187], wl_l[188], wl_l[189],
     wl_l[190], wl_l[191], wl_l[192], wl_l[193], wl_l[194], wl_l[195],
     wl_l[196], wl_l[197], wl_l[198], wl_l[199], wl_l[200], wl_l[201],
     wl_l[202], wl_l[203], wl_l[204], wl_l[205], wl_l[206], wl_l[207],
     wl_l[208], wl_l[209], wl_l[210], wl_l[211], wl_l[212], wl_l[213],
     wl_l[214], wl_l[215], wl_l[216], wl_l[217], wl_l[218], wl_l[219],
     wl_l[220], wl_l[221], wl_l[222], wl_l[223], wl_l[224], wl_l[225],
     wl_l[226], wl_l[227], wl_l[228], wl_l[229], wl_l[230], wl_l[231],
     wl_l[232], wl_l[233], wl_l[234], wl_l[235], wl_l[236], wl_l[237],
     wl_l[238], wl_l[239], wl_l[240], wl_l[241], wl_l[242], wl_l[243],
     wl_l[244], wl_l[245], wl_l[246], wl_l[247], wl_l[248], wl_l[249],
     wl_l[250], wl_l[251], wl_l[252], wl_l[253], wl_l[254], wl_l[255],
     wl_l[256], wl_l[257], wl_l[258], wl_l[259], wl_l[260], wl_l[261],
     wl_l[262], wl_l[263], wl_l[264], wl_l[265], wl_l[266], wl_l[267],
     wl_l[268], wl_l[269], wl_l[270], wl_l[271], wl_l[272], wl_l[273],
     wl_l[274], wl_l[275], wl_l[276], wl_l[277], wl_l[278], wl_l[279],
     wl_l[280], wl_l[281], wl_l[282], wl_l[283], wl_l[284], wl_l[285],
     wl_l[286], wl_l[287], wl_l[288], wl_l[289], wl_l[290], wl_l[291],
     wl_l[292], wl_l[293], wl_l[294], wl_l[295], wl_l[296], wl_l[297],
     wl_l[298], wl_l[299], wl_l[300], wl_l[301], wl_l[302], wl_l[303],
     wl_l[304], wl_l[305], wl_l[306], wl_l[307], wl_l[308], wl_l[309],
     wl_l[310], wl_l[311], wl_l[312], wl_l[313], wl_l[314], wl_l[315],
     wl_l[316], wl_l[317], wl_l[318], wl_l[319], wl_l[320], wl_l[321],
     wl_l[322], wl_l[323], wl_l[324], wl_l[325], wl_l[326], wl_l[327],
     wl_l[328], wl_l[329], wl_l[330], wl_l[331], wl_l[332], wl_l[333],
     wl_l[334], wl_l[335], wl_l[336], wl_l[337], wl_l[338], wl_l[339],
     wl_l[340], wl_l[341], wl_l[342], wl_l[343], wl_l[344], wl_l[345],
     wl_l[346], wl_l[347], wl_l[348], wl_l[349], wl_l[350], wl_l[351],
     wl_l[175], wl_l[174], wl_l[173], wl_l[172], wl_l[171], wl_l[170],
     wl_l[169], wl_l[168], wl_l[167], wl_l[166], wl_l[165], wl_l[164],
     wl_l[163], wl_l[162], wl_l[161], wl_l[160], wl_l[159], wl_l[158],
     wl_l[157], wl_l[156], wl_l[155], wl_l[154], wl_l[153], wl_l[152],
     wl_l[151], wl_l[150], wl_l[149], wl_l[148], wl_l[147], wl_l[146],
     wl_l[145], wl_l[144], wl_l[143], wl_l[142], wl_l[141], wl_l[140],
     wl_l[139], wl_l[138], wl_l[137], wl_l[136], wl_l[135], wl_l[134],
     wl_l[133], wl_l[132], wl_l[131], wl_l[130], wl_l[129], wl_l[128],
     wl_l[127], wl_l[126], wl_l[125], wl_l[124], wl_l[123], wl_l[122],
     wl_l[121], wl_l[120], wl_l[119], wl_l[118], wl_l[117], wl_l[116],
     wl_l[115], wl_l[114], wl_l[113], wl_l[112], wl_l[111], wl_l[110],
     wl_l[109], wl_l[108], wl_l[107], wl_l[106], wl_l[105], wl_l[104],
     wl_l[103], wl_l[102], wl_l[101], wl_l[100], wl_l[99], wl_l[98],
     wl_l[97], wl_l[96], wl_l[95], wl_l[94], wl_l[93], wl_l[92],
     wl_l[91], wl_l[90], wl_l[89], wl_l[88], wl_l[87], wl_l[86],
     wl_l[85], wl_l[84], wl_l[83], wl_l[82], wl_l[81], wl_l[80],
     wl_l[79], wl_l[78], wl_l[77], wl_l[76], wl_l[75], wl_l[74],
     wl_l[73], wl_l[72], wl_l[71], wl_l[70], wl_l[69], wl_l[68],
     wl_l[67], wl_l[66], wl_l[65], wl_l[64], wl_l[63], wl_l[62],
     wl_l[61], wl_l[60], wl_l[59], wl_l[58], wl_l[57], wl_l[56],
     wl_l[55], wl_l[54], wl_l[53], wl_l[52], wl_l[51], wl_l[50],
     wl_l[49], wl_l[48], wl_l[47], wl_l[46], wl_l[45], wl_l[44],
     wl_l[43], wl_l[42], wl_l[41], wl_l[40], wl_l[39], wl_l[38],
     wl_l[37], wl_l[36], wl_l[35], wl_l[34], wl_l[33], wl_l[32],
     wl_l[31], wl_l[30], wl_l[29], wl_l[28], wl_l[27], wl_l[26],
     wl_l[25], wl_l[24], wl_l[23], wl_l[22], wl_l[21], wl_l[20],
     wl_l[19], wl_l[18], wl_l[17], wl_l[16], wl_l[15], wl_l[14],
     wl_l[13], wl_l[12], wl_l[11], wl_l[10], wl_l[9], wl_l[8], wl_l[7],
     wl_l[6], wl_l[5], wl_l[4], wl_l[3], wl_l[2], wl_l[1], wl_l[0]}),
     .pado_l(out_lbank[39:0]), .update(update0), .tclk(j_tck),
     .shift(shift0), .padeb_l(oen_lbank[39:0]), .sdi_pad(j_tdi),
     .cf_l({cf_lbank[263], cf_lbank[262], cf_lbank[261], cf_lbank[260],
     cf_lbank[259], cf_lbank[258], cf_lbank[257], cf_lbank[256],
     cf_lbank[255], cf_lbank[254], cf_lbank[253], cf_lbank[252],
     cf_lbank[251], cf_lbank[250], cf_lbank[249], cf_lbank[248],
     cf_lbank[247], cf_lbank[246], cf_lbank[245], cf_lbank[244],
     cf_lbank[243], cf_lbank[242], cf_lbank[241], cf_lbank[240],
     cf_lbank[287], cf_lbank[286], cf_lbank[285], cf_lbank[284],
     cf_lbank[283], cf_lbank[282], cf_lbank[281], cf_lbank[280],
     cf_lbank[279], cf_lbank[278], cf_lbank[277], cf_lbank[276],
     cf_lbank[275], cf_lbank[274], cf_lbank[273], cf_lbank[272],
     cf_lbank[271], cf_lbank[270], cf_lbank[269], cf_lbank[268],
     cf_lbank[267], cf_lbank[266], cf_lbank[265], cf_lbank[264],
     cf_lbank[311], cf_lbank[310], cf_lbank[309], cf_lbank[308],
     cf_lbank[307], cf_lbank[306], cf_lbank[305], cf_lbank[304],
     cf_lbank[303], cf_lbank[302], cf_lbank[301], cf_lbank[300],
     cf_lbank[299], cf_lbank[298], cf_lbank[297], cf_lbank[296],
     cf_lbank[295], cf_lbank[294], cf_lbank[293], cf_lbank[292],
     cf_lbank[291], cf_lbank[290], cf_lbank[289], cf_lbank[288],
     cf_lbank[335], cf_lbank[334], cf_lbank[333], cf_lbank[332],
     cf_lbank[331], cf_lbank[330], cf_lbank[329], cf_lbank[328],
     cf_lbank[327], cf_lbank[326], cf_lbank[325], cf_lbank[324],
     cf_lbank[323], cf_lbank[322], cf_lbank[321], cf_lbank[320],
     cf_lbank[319], cf_lbank[318], cf_lbank[317], cf_lbank[316],
     cf_lbank[315], cf_lbank[314], cf_lbank[313], cf_lbank[312],
     cf_lbank[359], cf_lbank[358], cf_lbank[357], cf_lbank[356],
     cf_lbank[355], cf_lbank[354], cf_lbank[353], cf_lbank[352],
     cf_lbank[351], cf_lbank[350], cf_lbank[349], cf_lbank[348],
     cf_lbank[347], cf_lbank[346], cf_lbank[345], cf_lbank[344],
     cf_lbank[343], cf_lbank[342], cf_lbank[341], cf_lbank[340],
     cf_lbank[339], cf_lbank[338], cf_lbank[337], cf_lbank[336],
     cf_lbank[383], cf_lbank[382], cf_lbank[381], cf_lbank[380],
     cf_lbank[379], cf_lbank[378], cf_lbank[377], cf_lbank[376],
     cf_lbank[375], cf_lbank[374], cf_lbank[373], cf_lbank[372],
     cf_lbank[371], cf_lbank[370], cf_lbank[369], cf_lbank[368],
     cf_lbank[367], cf_lbank[366], cf_lbank[365], cf_lbank[364],
     cf_lbank[363], cf_lbank[362], cf_lbank[361], cf_lbank[360],
     cf_lbank[407], cf_lbank[406], cf_lbank[405], cf_lbank[404],
     cf_lbank[403], cf_lbank[402], cf_lbank[401], cf_lbank[400],
     cf_lbank[399], cf_lbank[398], cf_lbank[397], cf_lbank[396],
     cf_lbank[395], cf_lbank[394], cf_lbank[393], cf_lbank[392],
     cf_lbank[391], cf_lbank[390], cf_lbank[389], cf_lbank[388],
     cf_lbank[387], cf_lbank[386], cf_lbank[385], cf_lbank[384],
     cf_lbank[431], cf_lbank[430], cf_lbank[429], cf_lbank[428],
     cf_lbank[427], cf_lbank[426], cf_lbank[425], cf_lbank[424],
     cf_lbank[423], cf_lbank[422], cf_lbank[421], cf_lbank[420],
     cf_lbank[419], cf_lbank[418], cf_lbank[417], cf_lbank[416],
     cf_lbank[415], cf_lbank[414], cf_lbank[413], cf_lbank[412],
     cf_lbank[411], cf_lbank[410], cf_lbank[409], cf_lbank[408],
     cf_lbank[455], cf_lbank[454], cf_lbank[453], cf_lbank[452],
     cf_lbank[451], cf_lbank[450], cf_lbank[449], cf_lbank[448],
     cf_lbank[447], cf_lbank[446], cf_lbank[445], cf_lbank[444],
     cf_lbank[443], cf_lbank[442], cf_lbank[441], cf_lbank[440],
     cf_lbank[439], cf_lbank[438], cf_lbank[437], cf_lbank[436],
     cf_lbank[435], cf_lbank[434], cf_lbank[433], cf_lbank[432],
     cf_lbank[479], cf_lbank[478], cf_lbank[477], cf_lbank[476],
     cf_lbank[475], cf_lbank[474], cf_lbank[473], cf_lbank[472],
     cf_lbank[471], cf_lbank[470], cf_lbank[469], cf_lbank[468],
     cf_lbank[467], cf_lbank[466], cf_lbank[465], cf_lbank[464],
     cf_lbank[463], cf_lbank[462], cf_lbank[461], cf_lbank[460],
     cf_lbank[459], cf_lbank[458], cf_lbank[457], cf_lbank[456],
     cf_lbank[239], cf_lbank[238], cf_lbank[237], cf_lbank[236],
     cf_lbank[235], cf_lbank[234], cf_lbank[233], cf_lbank[232],
     cf_lbank[231], cf_lbank[230], cf_lbank[229], cf_lbank[228],
     cf_lbank[227], cf_lbank[226], cf_lbank[225], cf_lbank[224],
     cf_lbank[223], cf_lbank[222], cf_lbank[221], cf_lbank[220],
     cf_lbank[219], cf_lbank[218], cf_lbank[217], cf_lbank[216],
     cf_lbank[215], cf_lbank[214], cf_lbank[213], cf_lbank[212],
     cf_lbank[211], cf_lbank[210], cf_lbank[209], cf_lbank[208],
     cf_lbank[207], cf_lbank[206], cf_lbank[205], cf_lbank[204],
     cf_lbank[203], cf_lbank[202], cf_lbank[201], cf_lbank[200],
     cf_lbank[199], cf_lbank[198], cf_lbank[197], cf_lbank[196],
     cf_lbank[195], cf_lbank[194], cf_lbank[193], cf_lbank[192],
     cf_lbank[191], cf_lbank[190], cf_lbank[189], cf_lbank[188],
     cf_lbank[187], cf_lbank[186], cf_lbank[185], cf_lbank[184],
     cf_lbank[183], cf_lbank[182], cf_lbank[181], cf_lbank[180],
     cf_lbank[179], cf_lbank[178], cf_lbank[177], cf_lbank[176],
     cf_lbank[175], cf_lbank[174], cf_lbank[173], cf_lbank[172],
     cf_lbank[171], cf_lbank[170], cf_lbank[169], cf_lbank[168],
     cf_lbank[167], cf_lbank[166], cf_lbank[165], cf_lbank[164],
     cf_lbank[163], cf_lbank[162], cf_lbank[161], cf_lbank[160],
     cf_lbank[159], cf_lbank[158], cf_lbank[157], cf_lbank[156],
     cf_lbank[155], cf_lbank[154], cf_lbank[153], cf_lbank[152],
     cf_lbank[151], cf_lbank[150], cf_lbank[149], cf_lbank[148],
     cf_lbank[147], cf_lbank[146], cf_lbank[145], cf_lbank[144],
     cf_lbank[143], cf_lbank[142], cf_lbank[141], cf_lbank[140],
     cf_lbank[139], cf_lbank[138], cf_lbank[137], cf_lbank[136],
     cf_lbank[135], cf_lbank[134], cf_lbank[133], cf_lbank[132],
     cf_lbank[131], cf_lbank[130], cf_lbank[129], cf_lbank[128],
     cf_lbank[127], cf_lbank[126], cf_lbank[125], cf_lbank[124],
     cf_lbank[123], cf_lbank[122], cf_lbank[121], cf_lbank[120],
     cf_lbank[119], cf_lbank[118], cf_lbank[117], cf_lbank[116],
     cf_lbank[115], cf_lbank[114], cf_lbank[113], cf_lbank[112],
     cf_lbank[111], cf_lbank[110], cf_lbank[109], cf_lbank[108],
     cf_lbank[107], cf_lbank[106], cf_lbank[105], cf_lbank[104],
     cf_lbank[103], cf_lbank[102], cf_lbank[101], cf_lbank[100],
     cf_lbank[99], cf_lbank[98], cf_lbank[97], cf_lbank[96],
     cf_lbank[95], cf_lbank[94], cf_lbank[93], cf_lbank[92],
     cf_lbank[91], cf_lbank[90], cf_lbank[89], cf_lbank[88],
     cf_lbank[87], cf_lbank[86], cf_lbank[85], cf_lbank[84],
     cf_lbank[83], cf_lbank[82], cf_lbank[81], cf_lbank[80],
     cf_lbank[79], cf_lbank[78], cf_lbank[77], cf_lbank[76],
     cf_lbank[75], cf_lbank[74], cf_lbank[73], cf_lbank[72],
     cf_lbank[71], cf_lbank[70], cf_lbank[69], cf_lbank[68],
     cf_lbank[67], cf_lbank[66], cf_lbank[65], cf_lbank[64],
     cf_lbank[63], cf_lbank[62], cf_lbank[61], cf_lbank[60],
     cf_lbank[59], cf_lbank[58], cf_lbank[57], cf_lbank[56],
     cf_lbank[55], cf_lbank[54], cf_lbank[53], cf_lbank[52],
     cf_lbank[51], cf_lbank[50], cf_lbank[49], cf_lbank[48],
     cf_lbank[47], cf_lbank[46], cf_lbank[45], cf_lbank[44],
     cf_lbank[43], cf_lbank[42], cf_lbank[41], cf_lbank[40],
     cf_lbank[39], cf_lbank[38], cf_lbank[37], cf_lbank[36],
     cf_lbank[35], cf_lbank[34], cf_lbank[33], cf_lbank[32],
     cf_lbank[31], cf_lbank[30], cf_lbank[29], cf_lbank[28],
     cf_lbank[27], cf_lbank[26], cf_lbank[25], cf_lbank[24],
     cf_lbank[23], cf_lbank[22], cf_lbank[21], cf_lbank[20],
     cf_lbank[19], cf_lbank[18], cf_lbank[17], cf_lbank[16],
     cf_lbank[15], cf_lbank[14], cf_lbank[13], cf_lbank[12],
     cf_lbank[11], cf_lbank[10], cf_lbank[9], cf_lbank[8], cf_lbank[7],
     cf_lbank[6], cf_lbank[5], cf_lbank[4], cf_lbank[3], cf_lbank[2],
     cf_lbank[1], cf_lbank[0]}), .reset_b_l({reset_l[176],
     reset_l[177], reset_l[178], reset_l[179], reset_l[180],
     reset_l[181], reset_l[182], reset_l[183], reset_l[184],
     reset_l[185], reset_l[186], reset_l[187], reset_l[188],
     reset_l[189], reset_l[190], reset_l[191], reset_l[192],
     reset_l[193], reset_l[194], reset_l[195], reset_l[196],
     reset_l[197], reset_l[198], reset_l[199], reset_l[200],
     reset_l[201], reset_l[202], reset_l[203], reset_l[204],
     reset_l[205], reset_l[206], reset_l[207], reset_l[208],
     reset_l[209], reset_l[210], reset_l[211], reset_l[212],
     reset_l[213], reset_l[214], reset_l[215], reset_l[216],
     reset_l[217], reset_l[218], reset_l[219], reset_l[220],
     reset_l[221], reset_l[222], reset_l[223], reset_l[224],
     reset_l[225], reset_l[226], reset_l[227], reset_l[228],
     reset_l[229], reset_l[230], reset_l[231], reset_l[232],
     reset_l[233], reset_l[234], reset_l[235], reset_l[236],
     reset_l[237], reset_l[238], reset_l[239], reset_l[240],
     reset_l[241], reset_l[242], reset_l[243], reset_l[244],
     reset_l[245], reset_l[246], reset_l[247], reset_l[248],
     reset_l[249], reset_l[250], reset_l[251], reset_l[252],
     reset_l[253], reset_l[254], reset_l[255], reset_l[256],
     reset_l[257], reset_l[258], reset_l[259], reset_l[260],
     reset_l[261], reset_l[262], reset_l[263], reset_l[264],
     reset_l[265], reset_l[266], reset_l[267], reset_l[268],
     reset_l[269], reset_l[270], reset_l[271], reset_l[272],
     reset_l[273], reset_l[274], reset_l[275], reset_l[276],
     reset_l[277], reset_l[278], reset_l[279], reset_l[280],
     reset_l[281], reset_l[282], reset_l[283], reset_l[284],
     reset_l[285], reset_l[286], reset_l[287], reset_l[288],
     reset_l[289], reset_l[290], reset_l[291], reset_l[292],
     reset_l[293], reset_l[294], reset_l[295], reset_l[296],
     reset_l[297], reset_l[298], reset_l[299], reset_l[300],
     reset_l[301], reset_l[302], reset_l[303], reset_l[304],
     reset_l[305], reset_l[306], reset_l[307], reset_l[308],
     reset_l[309], reset_l[310], reset_l[311], reset_l[312],
     reset_l[313], reset_l[314], reset_l[315], reset_l[316],
     reset_l[317], reset_l[318], reset_l[319], reset_l[320],
     reset_l[321], reset_l[322], reset_l[323], reset_l[324],
     reset_l[325], reset_l[326], reset_l[327], reset_l[328],
     reset_l[329], reset_l[330], reset_l[331], reset_l[332],
     reset_l[333], reset_l[334], reset_l[335], reset_l[336],
     reset_l[337], reset_l[338], reset_l[339], reset_l[340],
     reset_l[341], reset_l[342], reset_l[343], reset_l[344],
     reset_l[345], reset_l[346], reset_l[347], reset_l[348],
     reset_l[349], reset_l[350], reset_l[351], reset_l[175],
     reset_l[174], reset_l[173], reset_l[172], reset_l[171],
     reset_l[170], reset_l[169], reset_l[168], reset_l[167],
     reset_l[166], reset_l[165], reset_l[164], reset_l[163],
     reset_l[162], reset_l[161], reset_l[160], reset_l[159],
     reset_l[158], reset_l[157], reset_l[156], reset_l[155],
     reset_l[154], reset_l[153], reset_l[152], reset_l[151],
     reset_l[150], reset_l[149], reset_l[148], reset_l[147],
     reset_l[146], reset_l[145], reset_l[144], reset_l[143],
     reset_l[142], reset_l[141], reset_l[140], reset_l[139],
     reset_l[138], reset_l[137], reset_l[136], reset_l[135],
     reset_l[134], reset_l[133], reset_l[132], reset_l[131],
     reset_l[130], reset_l[129], reset_l[128], reset_l[127],
     reset_l[126], reset_l[125], reset_l[124], reset_l[123],
     reset_l[122], reset_l[121], reset_l[120], reset_l[119],
     reset_l[118], reset_l[117], reset_l[116], reset_l[115],
     reset_l[114], reset_l[113], reset_l[112], reset_l[111],
     reset_l[110], reset_l[109], reset_l[108], reset_l[107],
     reset_l[106], reset_l[105], reset_l[104], reset_l[103],
     reset_l[102], reset_l[101], reset_l[100], reset_l[99],
     reset_l[98], reset_l[97], reset_l[96], reset_l[95], reset_l[94],
     reset_l[93], reset_l[92], reset_l[91], reset_l[90], reset_l[89],
     reset_l[88], reset_l[87], reset_l[86], reset_l[85], reset_l[84],
     reset_l[83], reset_l[82], reset_l[81], reset_l[80], reset_l[79],
     reset_l[78], reset_l[77], reset_l[76], reset_l[75], reset_l[74],
     reset_l[73], reset_l[72], reset_l[71], reset_l[70], reset_l[69],
     reset_l[68], reset_l[67], reset_l[66], reset_l[65], reset_l[64],
     reset_l[63], reset_l[62], reset_l[61], reset_l[60], reset_l[59],
     reset_l[58], reset_l[57], reset_l[56], reset_l[55], reset_l[54],
     reset_l[53], reset_l[52], reset_l[51], reset_l[50], reset_l[49],
     reset_l[48], reset_l[47], reset_l[46], reset_l[45], reset_l[44],
     reset_l[43], reset_l[42], reset_l[41], reset_l[40], reset_l[39],
     reset_l[38], reset_l[37], reset_l[36], reset_l[35], reset_l[34],
     reset_l[33], reset_l[32], reset_l[31], reset_l[30], reset_l[29],
     reset_l[28], reset_l[27], reset_l[26], reset_l[25], reset_l[24],
     reset_l[23], reset_l[22], reset_l[21], reset_l[20], reset_l[19],
     reset_l[18], reset_l[17], reset_l[16], reset_l[15], reset_l[14],
     reset_l[13], reset_l[12], reset_l[11], reset_l[10], reset_l[9],
     reset_l[8], reset_l[7], reset_l[6], reset_l[5], reset_l[4],
     reset_l[3], reset_l[2], reset_l[1], reset_l[0]}), .r(gsr),
     .purst(gsr), .prog(gint_hz), .pgate_l({pgate_l[176], pgate_l[177],
     pgate_l[178], pgate_l[179], pgate_l[180], pgate_l[181],
     pgate_l[182], pgate_l[183], pgate_l[184], pgate_l[185],
     pgate_l[186], pgate_l[187], pgate_l[188], pgate_l[189],
     pgate_l[190], pgate_l[191], pgate_l[192], pgate_l[193],
     pgate_l[194], pgate_l[195], pgate_l[196], pgate_l[197],
     pgate_l[198], pgate_l[199], pgate_l[200], pgate_l[201],
     pgate_l[202], pgate_l[203], pgate_l[204], pgate_l[205],
     pgate_l[206], pgate_l[207], pgate_l[208], pgate_l[209],
     pgate_l[210], pgate_l[211], pgate_l[212], pgate_l[213],
     pgate_l[214], pgate_l[215], pgate_l[216], pgate_l[217],
     pgate_l[218], pgate_l[219], pgate_l[220], pgate_l[221],
     pgate_l[222], pgate_l[223], pgate_l[224], pgate_l[225],
     pgate_l[226], pgate_l[227], pgate_l[228], pgate_l[229],
     pgate_l[230], pgate_l[231], pgate_l[232], pgate_l[233],
     pgate_l[234], pgate_l[235], pgate_l[236], pgate_l[237],
     pgate_l[238], pgate_l[239], pgate_l[240], pgate_l[241],
     pgate_l[242], pgate_l[243], pgate_l[244], pgate_l[245],
     pgate_l[246], pgate_l[247], pgate_l[248], pgate_l[249],
     pgate_l[250], pgate_l[251], pgate_l[252], pgate_l[253],
     pgate_l[254], pgate_l[255], pgate_l[256], pgate_l[257],
     pgate_l[258], pgate_l[259], pgate_l[260], pgate_l[261],
     pgate_l[262], pgate_l[263], pgate_l[264], pgate_l[265],
     pgate_l[266], pgate_l[267], pgate_l[268], pgate_l[269],
     pgate_l[270], pgate_l[271], pgate_l[272], pgate_l[273],
     pgate_l[274], pgate_l[275], pgate_l[276], pgate_l[277],
     pgate_l[278], pgate_l[279], pgate_l[280], pgate_l[281],
     pgate_l[282], pgate_l[283], pgate_l[284], pgate_l[285],
     pgate_l[286], pgate_l[287], pgate_l[288], pgate_l[289],
     pgate_l[290], pgate_l[291], pgate_l[292], pgate_l[293],
     pgate_l[294], pgate_l[295], pgate_l[296], pgate_l[297],
     pgate_l[298], pgate_l[299], pgate_l[300], pgate_l[301],
     pgate_l[302], pgate_l[303], pgate_l[304], pgate_l[305],
     pgate_l[306], pgate_l[307], pgate_l[308], pgate_l[309],
     pgate_l[310], pgate_l[311], pgate_l[312], pgate_l[313],
     pgate_l[314], pgate_l[315], pgate_l[316], pgate_l[317],
     pgate_l[318], pgate_l[319], pgate_l[320], pgate_l[321],
     pgate_l[322], pgate_l[323], pgate_l[324], pgate_l[325],
     pgate_l[326], pgate_l[327], pgate_l[328], pgate_l[329],
     pgate_l[330], pgate_l[331], pgate_l[332], pgate_l[333],
     pgate_l[334], pgate_l[335], pgate_l[336], pgate_l[337],
     pgate_l[338], pgate_l[339], pgate_l[340], pgate_l[341],
     pgate_l[342], pgate_l[343], pgate_l[344], pgate_l[345],
     pgate_l[346], pgate_l[347], pgate_l[348], pgate_l[349],
     pgate_l[350], pgate_l[351], pgate_l[175], pgate_l[174],
     pgate_l[173], pgate_l[172], pgate_l[171], pgate_l[170],
     pgate_l[169], pgate_l[168], pgate_l[167], pgate_l[166],
     pgate_l[165], pgate_l[164], pgate_l[163], pgate_l[162],
     pgate_l[161], pgate_l[160], pgate_l[159], pgate_l[158],
     pgate_l[157], pgate_l[156], pgate_l[155], pgate_l[154],
     pgate_l[153], pgate_l[152], pgate_l[151], pgate_l[150],
     pgate_l[149], pgate_l[148], pgate_l[147], pgate_l[146],
     pgate_l[145], pgate_l[144], pgate_l[143], pgate_l[142],
     pgate_l[141], pgate_l[140], pgate_l[139], pgate_l[138],
     pgate_l[137], pgate_l[136], pgate_l[135], pgate_l[134],
     pgate_l[133], pgate_l[132], pgate_l[131], pgate_l[130],
     pgate_l[129], pgate_l[128], pgate_l[127], pgate_l[126],
     pgate_l[125], pgate_l[124], pgate_l[123], pgate_l[122],
     pgate_l[121], pgate_l[120], pgate_l[119], pgate_l[118],
     pgate_l[117], pgate_l[116], pgate_l[115], pgate_l[114],
     pgate_l[113], pgate_l[112], pgate_l[111], pgate_l[110],
     pgate_l[109], pgate_l[108], pgate_l[107], pgate_l[106],
     pgate_l[105], pgate_l[104], pgate_l[103], pgate_l[102],
     pgate_l[101], pgate_l[100], pgate_l[99], pgate_l[98], pgate_l[97],
     pgate_l[96], pgate_l[95], pgate_l[94], pgate_l[93], pgate_l[92],
     pgate_l[91], pgate_l[90], pgate_l[89], pgate_l[88], pgate_l[87],
     pgate_l[86], pgate_l[85], pgate_l[84], pgate_l[83], pgate_l[82],
     pgate_l[81], pgate_l[80], pgate_l[79], pgate_l[78], pgate_l[77],
     pgate_l[76], pgate_l[75], pgate_l[74], pgate_l[73], pgate_l[72],
     pgate_l[71], pgate_l[70], pgate_l[69], pgate_l[68], pgate_l[67],
     pgate_l[66], pgate_l[65], pgate_l[64], pgate_l[63], pgate_l[62],
     pgate_l[61], pgate_l[60], pgate_l[59], pgate_l[58], pgate_l[57],
     pgate_l[56], pgate_l[55], pgate_l[54], pgate_l[53], pgate_l[52],
     pgate_l[51], pgate_l[50], pgate_l[49], pgate_l[48], pgate_l[47],
     pgate_l[46], pgate_l[45], pgate_l[44], pgate_l[43], pgate_l[42],
     pgate_l[41], pgate_l[40], pgate_l[39], pgate_l[38], pgate_l[37],
     pgate_l[36], pgate_l[35], pgate_l[34], pgate_l[33], pgate_l[32],
     pgate_l[31], pgate_l[30], pgate_l[29], pgate_l[28], pgate_l[27],
     pgate_l[26], pgate_l[25], pgate_l[24], pgate_l[23], pgate_l[22],
     pgate_l[21], pgate_l[20], pgate_l[19], pgate_l[18], pgate_l[17],
     pgate_l[16], pgate_l[15], pgate_l[14], pgate_l[13], pgate_l[12],
     pgate_l[11], pgate_l[10], pgate_l[9], pgate_l[8], pgate_l[7],
     pgate_l[6], pgate_l[5], pgate_l[4], pgate_l[3], pgate_l[2],
     pgate_l[1], pgate_l[0]}), .mode(mode0), .hiz_b(hiz_b0),
     .end_of_startup_l({tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu0_b, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd}), .bs_en(bs_en0),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .spi_ss_in_r(spi_ss_in_r[39:0]),
     .sdo_pad(fromsdo), .pado_r(out_rbank[39:0]),
     .cf_r(cf_rbank[479:0]), .bm_sdo_o(bm_sdo_o[3:0]),
     .wl_r({wl_r[176], wl_r[177], wl_r[178], wl_r[179], wl_r[180],
     wl_r[181], wl_r[182], wl_r[183], wl_r[184], wl_r[185], wl_r[186],
     wl_r[187], wl_r[188], wl_r[189], wl_r[190], wl_r[191], wl_r[192],
     wl_r[193], wl_r[194], wl_r[195], wl_r[196], wl_r[197], wl_r[198],
     wl_r[199], wl_r[200], wl_r[201], wl_r[202], wl_r[203], wl_r[204],
     wl_r[205], wl_r[206], wl_r[207], wl_r[208], wl_r[209], wl_r[210],
     wl_r[211], wl_r[212], wl_r[213], wl_r[214], wl_r[215], wl_r[216],
     wl_r[217], wl_r[218], wl_r[219], wl_r[220], wl_r[221], wl_r[222],
     wl_r[223], wl_r[224], wl_r[225], wl_r[226], wl_r[227], wl_r[228],
     wl_r[229], wl_r[230], wl_r[231], wl_r[232], wl_r[233], wl_r[234],
     wl_r[235], wl_r[236], wl_r[237], wl_r[238], wl_r[239], wl_r[240],
     wl_r[241], wl_r[242], wl_r[243], wl_r[244], wl_r[245], wl_r[246],
     wl_r[247], wl_r[248], wl_r[249], wl_r[250], wl_r[251], wl_r[252],
     wl_r[253], wl_r[254], wl_r[255], wl_r[256], wl_r[257], wl_r[258],
     wl_r[259], wl_r[260], wl_r[261], wl_r[262], wl_r[263], wl_r[264],
     wl_r[265], wl_r[266], wl_r[267], wl_r[268], wl_r[269], wl_r[270],
     wl_r[271], wl_r[272], wl_r[273], wl_r[274], wl_r[275], wl_r[276],
     wl_r[277], wl_r[278], wl_r[279], wl_r[280], wl_r[281], wl_r[282],
     wl_r[283], wl_r[284], wl_r[285], wl_r[286], wl_r[287], wl_r[288],
     wl_r[289], wl_r[290], wl_r[291], wl_r[292], wl_r[293], wl_r[294],
     wl_r[295], wl_r[296], wl_r[297], wl_r[298], wl_r[299], wl_r[300],
     wl_r[301], wl_r[302], wl_r[303], wl_r[304], wl_r[305], wl_r[306],
     wl_r[307], wl_r[308], wl_r[309], wl_r[310], wl_r[311], wl_r[312],
     wl_r[313], wl_r[314], wl_r[315], wl_r[316], wl_r[317], wl_r[318],
     wl_r[319], wl_r[320], wl_r[321], wl_r[322], wl_r[323], wl_r[324],
     wl_r[325], wl_r[326], wl_r[327], wl_r[328], wl_r[329], wl_r[330],
     wl_r[331], wl_r[332], wl_r[333], wl_r[334], wl_r[335], wl_r[336],
     wl_r[337], wl_r[338], wl_r[339], wl_r[340], wl_r[341], wl_r[342],
     wl_r[343], wl_r[344], wl_r[345], wl_r[346], wl_r[347], wl_r[348],
     wl_r[349], wl_r[350], wl_r[351], wl_r[175], wl_r[174], wl_r[173],
     wl_r[172], wl_r[171], wl_r[170], wl_r[169], wl_r[168], wl_r[167],
     wl_r[166], wl_r[165], wl_r[164], wl_r[163], wl_r[162], wl_r[161],
     wl_r[160], wl_r[159], wl_r[158], wl_r[157], wl_r[156], wl_r[155],
     wl_r[154], wl_r[153], wl_r[152], wl_r[151], wl_r[150], wl_r[149],
     wl_r[148], wl_r[147], wl_r[146], wl_r[145], wl_r[144], wl_r[143],
     wl_r[142], wl_r[141], wl_r[140], wl_r[139], wl_r[138], wl_r[137],
     wl_r[136], wl_r[135], wl_r[134], wl_r[133], wl_r[132], wl_r[131],
     wl_r[130], wl_r[129], wl_r[128], wl_r[127], wl_r[126], wl_r[125],
     wl_r[124], wl_r[123], wl_r[122], wl_r[121], wl_r[120], wl_r[119],
     wl_r[118], wl_r[117], wl_r[116], wl_r[115], wl_r[114], wl_r[113],
     wl_r[112], wl_r[111], wl_r[110], wl_r[109], wl_r[108], wl_r[107],
     wl_r[106], wl_r[105], wl_r[104], wl_r[103], wl_r[102], wl_r[101],
     wl_r[100], wl_r[99], wl_r[98], wl_r[97], wl_r[96], wl_r[95],
     wl_r[94], wl_r[93], wl_r[92], wl_r[91], wl_r[90], wl_r[89],
     wl_r[88], wl_r[87], wl_r[86], wl_r[85], wl_r[84], wl_r[83],
     wl_r[82], wl_r[81], wl_r[80], wl_r[79], wl_r[78], wl_r[77],
     wl_r[76], wl_r[75], wl_r[74], wl_r[73], wl_r[72], wl_r[71],
     wl_r[70], wl_r[69], wl_r[68], wl_r[67], wl_r[66], wl_r[65],
     wl_r[64], wl_r[63], wl_r[62], wl_r[61], wl_r[60], wl_r[59],
     wl_r[58], wl_r[57], wl_r[56], wl_r[55], wl_r[54], wl_r[53],
     wl_r[52], wl_r[51], wl_r[50], wl_r[49], wl_r[48], wl_r[47],
     wl_r[46], wl_r[45], wl_r[44], wl_r[43], wl_r[42], wl_r[41],
     wl_r[40], wl_r[39], wl_r[38], wl_r[37], wl_r[36], wl_r[35],
     wl_r[34], wl_r[33], wl_r[32], wl_r[31], wl_r[30], wl_r[29],
     wl_r[28], wl_r[27], wl_r[26], wl_r[25], wl_r[24], wl_r[23],
     wl_r[22], wl_r[21], wl_r[20], wl_r[19], wl_r[18], wl_r[17],
     wl_r[16], wl_r[15], wl_r[14], wl_r[13], wl_r[12], wl_r[11],
     wl_r[10], wl_r[9], wl_r[8], wl_r[7], wl_r[6], wl_r[5], wl_r[4],
     wl_r[3], wl_r[2], wl_r[1], wl_r[0]}),
     .vdd_cntl_r({vdd_cntl_r[176], vdd_cntl_r[177], vdd_cntl_r[178],
     vdd_cntl_r[179], vdd_cntl_r[180], vdd_cntl_r[181],
     vdd_cntl_r[182], vdd_cntl_r[183], vdd_cntl_r[184],
     vdd_cntl_r[185], vdd_cntl_r[186], vdd_cntl_r[187],
     vdd_cntl_r[188], vdd_cntl_r[189], vdd_cntl_r[190],
     vdd_cntl_r[191], vdd_cntl_r[192], vdd_cntl_r[193],
     vdd_cntl_r[194], vdd_cntl_r[195], vdd_cntl_r[196],
     vdd_cntl_r[197], vdd_cntl_r[198], vdd_cntl_r[199],
     vdd_cntl_r[200], vdd_cntl_r[201], vdd_cntl_r[202],
     vdd_cntl_r[203], vdd_cntl_r[204], vdd_cntl_r[205],
     vdd_cntl_r[206], vdd_cntl_r[207], vdd_cntl_r[208],
     vdd_cntl_r[209], vdd_cntl_r[210], vdd_cntl_r[211],
     vdd_cntl_r[212], vdd_cntl_r[213], vdd_cntl_r[214],
     vdd_cntl_r[215], vdd_cntl_r[216], vdd_cntl_r[217],
     vdd_cntl_r[218], vdd_cntl_r[219], vdd_cntl_r[220],
     vdd_cntl_r[221], vdd_cntl_r[222], vdd_cntl_r[223],
     vdd_cntl_r[224], vdd_cntl_r[225], vdd_cntl_r[226],
     vdd_cntl_r[227], vdd_cntl_r[228], vdd_cntl_r[229],
     vdd_cntl_r[230], vdd_cntl_r[231], vdd_cntl_r[232],
     vdd_cntl_r[233], vdd_cntl_r[234], vdd_cntl_r[235],
     vdd_cntl_r[236], vdd_cntl_r[237], vdd_cntl_r[238],
     vdd_cntl_r[239], vdd_cntl_r[240], vdd_cntl_r[241],
     vdd_cntl_r[242], vdd_cntl_r[243], vdd_cntl_r[244],
     vdd_cntl_r[245], vdd_cntl_r[246], vdd_cntl_r[247],
     vdd_cntl_r[248], vdd_cntl_r[249], vdd_cntl_r[250],
     vdd_cntl_r[251], vdd_cntl_r[252], vdd_cntl_r[253],
     vdd_cntl_r[254], vdd_cntl_r[255], vdd_cntl_r[256],
     vdd_cntl_r[257], vdd_cntl_r[258], vdd_cntl_r[259],
     vdd_cntl_r[260], vdd_cntl_r[261], vdd_cntl_r[262],
     vdd_cntl_r[263], vdd_cntl_r[264], vdd_cntl_r[265],
     vdd_cntl_r[266], vdd_cntl_r[267], vdd_cntl_r[268],
     vdd_cntl_r[269], vdd_cntl_r[270], vdd_cntl_r[271],
     vdd_cntl_r[272], vdd_cntl_r[273], vdd_cntl_r[274],
     vdd_cntl_r[275], vdd_cntl_r[276], vdd_cntl_r[277],
     vdd_cntl_r[278], vdd_cntl_r[279], vdd_cntl_r[280],
     vdd_cntl_r[281], vdd_cntl_r[282], vdd_cntl_r[283],
     vdd_cntl_r[284], vdd_cntl_r[285], vdd_cntl_r[286],
     vdd_cntl_r[287], vdd_cntl_r[288], vdd_cntl_r[289],
     vdd_cntl_r[290], vdd_cntl_r[291], vdd_cntl_r[292],
     vdd_cntl_r[293], vdd_cntl_r[294], vdd_cntl_r[295],
     vdd_cntl_r[296], vdd_cntl_r[297], vdd_cntl_r[298],
     vdd_cntl_r[299], vdd_cntl_r[300], vdd_cntl_r[301],
     vdd_cntl_r[302], vdd_cntl_r[303], vdd_cntl_r[304],
     vdd_cntl_r[305], vdd_cntl_r[306], vdd_cntl_r[307],
     vdd_cntl_r[308], vdd_cntl_r[309], vdd_cntl_r[310],
     vdd_cntl_r[311], vdd_cntl_r[312], vdd_cntl_r[313],
     vdd_cntl_r[314], vdd_cntl_r[315], vdd_cntl_r[316],
     vdd_cntl_r[317], vdd_cntl_r[318], vdd_cntl_r[319],
     vdd_cntl_r[320], vdd_cntl_r[321], vdd_cntl_r[322],
     vdd_cntl_r[323], vdd_cntl_r[324], vdd_cntl_r[325],
     vdd_cntl_r[326], vdd_cntl_r[327], vdd_cntl_r[328],
     vdd_cntl_r[329], vdd_cntl_r[330], vdd_cntl_r[331],
     vdd_cntl_r[332], vdd_cntl_r[333], vdd_cntl_r[334],
     vdd_cntl_r[335], vdd_cntl_r[336], vdd_cntl_r[337],
     vdd_cntl_r[338], vdd_cntl_r[339], vdd_cntl_r[340],
     vdd_cntl_r[341], vdd_cntl_r[342], vdd_cntl_r[343],
     vdd_cntl_r[344], vdd_cntl_r[345], vdd_cntl_r[346],
     vdd_cntl_r[347], vdd_cntl_r[348], vdd_cntl_r[349],
     vdd_cntl_r[350], vdd_cntl_r[351], vdd_cntl_r[175],
     vdd_cntl_r[174], vdd_cntl_r[173], vdd_cntl_r[172],
     vdd_cntl_r[171], vdd_cntl_r[170], vdd_cntl_r[169],
     vdd_cntl_r[168], vdd_cntl_r[167], vdd_cntl_r[166],
     vdd_cntl_r[165], vdd_cntl_r[164], vdd_cntl_r[163],
     vdd_cntl_r[162], vdd_cntl_r[161], vdd_cntl_r[160],
     vdd_cntl_r[159], vdd_cntl_r[158], vdd_cntl_r[157],
     vdd_cntl_r[156], vdd_cntl_r[155], vdd_cntl_r[154],
     vdd_cntl_r[153], vdd_cntl_r[152], vdd_cntl_r[151],
     vdd_cntl_r[150], vdd_cntl_r[149], vdd_cntl_r[148],
     vdd_cntl_r[147], vdd_cntl_r[146], vdd_cntl_r[145],
     vdd_cntl_r[144], vdd_cntl_r[143], vdd_cntl_r[142],
     vdd_cntl_r[141], vdd_cntl_r[140], vdd_cntl_r[139],
     vdd_cntl_r[138], vdd_cntl_r[137], vdd_cntl_r[136],
     vdd_cntl_r[135], vdd_cntl_r[134], vdd_cntl_r[133],
     vdd_cntl_r[132], vdd_cntl_r[131], vdd_cntl_r[130],
     vdd_cntl_r[129], vdd_cntl_r[128], vdd_cntl_r[127],
     vdd_cntl_r[126], vdd_cntl_r[125], vdd_cntl_r[124],
     vdd_cntl_r[123], vdd_cntl_r[122], vdd_cntl_r[121],
     vdd_cntl_r[120], vdd_cntl_r[119], vdd_cntl_r[118],
     vdd_cntl_r[117], vdd_cntl_r[116], vdd_cntl_r[115],
     vdd_cntl_r[114], vdd_cntl_r[113], vdd_cntl_r[112],
     vdd_cntl_r[111], vdd_cntl_r[110], vdd_cntl_r[109],
     vdd_cntl_r[108], vdd_cntl_r[107], vdd_cntl_r[106],
     vdd_cntl_r[105], vdd_cntl_r[104], vdd_cntl_r[103],
     vdd_cntl_r[102], vdd_cntl_r[101], vdd_cntl_r[100], vdd_cntl_r[99],
     vdd_cntl_r[98], vdd_cntl_r[97], vdd_cntl_r[96], vdd_cntl_r[95],
     vdd_cntl_r[94], vdd_cntl_r[93], vdd_cntl_r[92], vdd_cntl_r[91],
     vdd_cntl_r[90], vdd_cntl_r[89], vdd_cntl_r[88], vdd_cntl_r[87],
     vdd_cntl_r[86], vdd_cntl_r[85], vdd_cntl_r[84], vdd_cntl_r[83],
     vdd_cntl_r[82], vdd_cntl_r[81], vdd_cntl_r[80], vdd_cntl_r[79],
     vdd_cntl_r[78], vdd_cntl_r[77], vdd_cntl_r[76], vdd_cntl_r[75],
     vdd_cntl_r[74], vdd_cntl_r[73], vdd_cntl_r[72], vdd_cntl_r[71],
     vdd_cntl_r[70], vdd_cntl_r[69], vdd_cntl_r[68], vdd_cntl_r[67],
     vdd_cntl_r[66], vdd_cntl_r[65], vdd_cntl_r[64], vdd_cntl_r[63],
     vdd_cntl_r[62], vdd_cntl_r[61], vdd_cntl_r[60], vdd_cntl_r[59],
     vdd_cntl_r[58], vdd_cntl_r[57], vdd_cntl_r[56], vdd_cntl_r[55],
     vdd_cntl_r[54], vdd_cntl_r[53], vdd_cntl_r[52], vdd_cntl_r[51],
     vdd_cntl_r[50], vdd_cntl_r[49], vdd_cntl_r[48], vdd_cntl_r[47],
     vdd_cntl_r[46], vdd_cntl_r[45], vdd_cntl_r[44], vdd_cntl_r[43],
     vdd_cntl_r[42], vdd_cntl_r[41], vdd_cntl_r[40], vdd_cntl_r[39],
     vdd_cntl_r[38], vdd_cntl_r[37], vdd_cntl_r[36], vdd_cntl_r[35],
     vdd_cntl_r[34], vdd_cntl_r[33], vdd_cntl_r[32], vdd_cntl_r[31],
     vdd_cntl_r[30], vdd_cntl_r[29], vdd_cntl_r[28], vdd_cntl_r[27],
     vdd_cntl_r[26], vdd_cntl_r[25], vdd_cntl_r[24], vdd_cntl_r[23],
     vdd_cntl_r[22], vdd_cntl_r[21], vdd_cntl_r[20], vdd_cntl_r[19],
     vdd_cntl_r[18], vdd_cntl_r[17], vdd_cntl_r[16], vdd_cntl_r[15],
     vdd_cntl_r[14], vdd_cntl_r[13], vdd_cntl_r[12], vdd_cntl_r[11],
     vdd_cntl_r[10], vdd_cntl_r[9], vdd_cntl_r[8], vdd_cntl_r[7],
     vdd_cntl_r[6], vdd_cntl_r[5], vdd_cntl_r[4], vdd_cntl_r[3],
     vdd_cntl_r[2], vdd_cntl_r[1], vdd_cntl_r[0]}),
     .reset_b_r({reset_b_r[176], reset_b_r[177], reset_b_r[178],
     reset_b_r[179], reset_b_r[180], reset_b_r[181], reset_b_r[182],
     reset_b_r[183], reset_b_r[184], reset_b_r[185], reset_b_r[186],
     reset_b_r[187], reset_b_r[188], reset_b_r[189], reset_b_r[190],
     reset_b_r[191], reset_b_r[192], reset_b_r[193], reset_b_r[194],
     reset_b_r[195], reset_b_r[196], reset_b_r[197], reset_b_r[198],
     reset_b_r[199], reset_b_r[200], reset_b_r[201], reset_b_r[202],
     reset_b_r[203], reset_b_r[204], reset_b_r[205], reset_b_r[206],
     reset_b_r[207], reset_b_r[208], reset_b_r[209], reset_b_r[210],
     reset_b_r[211], reset_b_r[212], reset_b_r[213], reset_b_r[214],
     reset_b_r[215], reset_b_r[216], reset_b_r[217], reset_b_r[218],
     reset_b_r[219], reset_b_r[220], reset_b_r[221], reset_b_r[222],
     reset_b_r[223], reset_b_r[224], reset_b_r[225], reset_b_r[226],
     reset_b_r[227], reset_b_r[228], reset_b_r[229], reset_b_r[230],
     reset_b_r[231], reset_b_r[232], reset_b_r[233], reset_b_r[234],
     reset_b_r[235], reset_b_r[236], reset_b_r[237], reset_b_r[238],
     reset_b_r[239], reset_b_r[240], reset_b_r[241], reset_b_r[242],
     reset_b_r[243], reset_b_r[244], reset_b_r[245], reset_b_r[246],
     reset_b_r[247], reset_b_r[248], reset_b_r[249], reset_b_r[250],
     reset_b_r[251], reset_b_r[252], reset_b_r[253], reset_b_r[254],
     reset_b_r[255], reset_b_r[256], reset_b_r[257], reset_b_r[258],
     reset_b_r[259], reset_b_r[260], reset_b_r[261], reset_b_r[262],
     reset_b_r[263], reset_b_r[264], reset_b_r[265], reset_b_r[266],
     reset_b_r[267], reset_b_r[268], reset_b_r[269], reset_b_r[270],
     reset_b_r[271], reset_b_r[272], reset_b_r[273], reset_b_r[274],
     reset_b_r[275], reset_b_r[276], reset_b_r[277], reset_b_r[278],
     reset_b_r[279], reset_b_r[280], reset_b_r[281], reset_b_r[282],
     reset_b_r[283], reset_b_r[284], reset_b_r[285], reset_b_r[286],
     reset_b_r[287], reset_b_r[288], reset_b_r[289], reset_b_r[290],
     reset_b_r[291], reset_b_r[292], reset_b_r[293], reset_b_r[294],
     reset_b_r[295], reset_b_r[296], reset_b_r[297], reset_b_r[298],
     reset_b_r[299], reset_b_r[300], reset_b_r[301], reset_b_r[302],
     reset_b_r[303], reset_b_r[304], reset_b_r[305], reset_b_r[306],
     reset_b_r[307], reset_b_r[308], reset_b_r[309], reset_b_r[310],
     reset_b_r[311], reset_b_r[312], reset_b_r[313], reset_b_r[314],
     reset_b_r[315], reset_b_r[316], reset_b_r[317], reset_b_r[318],
     reset_b_r[319], reset_b_r[320], reset_b_r[321], reset_b_r[322],
     reset_b_r[323], reset_b_r[324], reset_b_r[325], reset_b_r[326],
     reset_b_r[327], reset_b_r[328], reset_b_r[329], reset_b_r[330],
     reset_b_r[331], reset_b_r[332], reset_b_r[333], reset_b_r[334],
     reset_b_r[335], reset_b_r[336], reset_b_r[337], reset_b_r[338],
     reset_b_r[339], reset_b_r[340], reset_b_r[341], reset_b_r[342],
     reset_b_r[343], reset_b_r[344], reset_b_r[345], reset_b_r[346],
     reset_b_r[347], reset_b_r[348], reset_b_r[349], reset_b_r[350],
     reset_b_r[351], reset_b_r[175], reset_b_r[174], reset_b_r[173],
     reset_b_r[172], reset_b_r[171], reset_b_r[170], reset_b_r[169],
     reset_b_r[168], reset_b_r[167], reset_b_r[166], reset_b_r[165],
     reset_b_r[164], reset_b_r[163], reset_b_r[162], reset_b_r[161],
     reset_b_r[160], reset_b_r[159], reset_b_r[158], reset_b_r[157],
     reset_b_r[156], reset_b_r[155], reset_b_r[154], reset_b_r[153],
     reset_b_r[152], reset_b_r[151], reset_b_r[150], reset_b_r[149],
     reset_b_r[148], reset_b_r[147], reset_b_r[146], reset_b_r[145],
     reset_b_r[144], reset_b_r[143], reset_b_r[142], reset_b_r[141],
     reset_b_r[140], reset_b_r[139], reset_b_r[138], reset_b_r[137],
     reset_b_r[136], reset_b_r[135], reset_b_r[134], reset_b_r[133],
     reset_b_r[132], reset_b_r[131], reset_b_r[130], reset_b_r[129],
     reset_b_r[128], reset_b_r[127], reset_b_r[126], reset_b_r[125],
     reset_b_r[124], reset_b_r[123], reset_b_r[122], reset_b_r[121],
     reset_b_r[120], reset_b_r[119], reset_b_r[118], reset_b_r[117],
     reset_b_r[116], reset_b_r[115], reset_b_r[114], reset_b_r[113],
     reset_b_r[112], reset_b_r[111], reset_b_r[110], reset_b_r[109],
     reset_b_r[108], reset_b_r[107], reset_b_r[106], reset_b_r[105],
     reset_b_r[104], reset_b_r[103], reset_b_r[102], reset_b_r[101],
     reset_b_r[100], reset_b_r[99], reset_b_r[98], reset_b_r[97],
     reset_b_r[96], reset_b_r[95], reset_b_r[94], reset_b_r[93],
     reset_b_r[92], reset_b_r[91], reset_b_r[90], reset_b_r[89],
     reset_b_r[88], reset_b_r[87], reset_b_r[86], reset_b_r[85],
     reset_b_r[84], reset_b_r[83], reset_b_r[82], reset_b_r[81],
     reset_b_r[80], reset_b_r[79], reset_b_r[78], reset_b_r[77],
     reset_b_r[76], reset_b_r[75], reset_b_r[74], reset_b_r[73],
     reset_b_r[72], reset_b_r[71], reset_b_r[70], reset_b_r[69],
     reset_b_r[68], reset_b_r[67], reset_b_r[66], reset_b_r[65],
     reset_b_r[64], reset_b_r[63], reset_b_r[62], reset_b_r[61],
     reset_b_r[60], reset_b_r[59], reset_b_r[58], reset_b_r[57],
     reset_b_r[56], reset_b_r[55], reset_b_r[54], reset_b_r[53],
     reset_b_r[52], reset_b_r[51], reset_b_r[50], reset_b_r[49],
     reset_b_r[48], reset_b_r[47], reset_b_r[46], reset_b_r[45],
     reset_b_r[44], reset_b_r[43], reset_b_r[42], reset_b_r[41],
     reset_b_r[40], reset_b_r[39], reset_b_r[38], reset_b_r[37],
     reset_b_r[36], reset_b_r[35], reset_b_r[34], reset_b_r[33],
     reset_b_r[32], reset_b_r[31], reset_b_r[30], reset_b_r[29],
     reset_b_r[28], reset_b_r[27], reset_b_r[26], reset_b_r[25],
     reset_b_r[24], reset_b_r[23], reset_b_r[22], reset_b_r[21],
     reset_b_r[20], reset_b_r[19], reset_b_r[18], reset_b_r[17],
     reset_b_r[16], reset_b_r[15], reset_b_r[14], reset_b_r[13],
     reset_b_r[12], reset_b_r[11], reset_b_r[10], reset_b_r[9],
     reset_b_r[8], reset_b_r[7], reset_b_r[6], reset_b_r[5],
     reset_b_r[4], reset_b_r[3], reset_b_r[2], reset_b_r[1],
     reset_b_r[0]}), .pgate_r({pgate_r[176], pgate_r[177],
     pgate_r[178], pgate_r[179], pgate_r[180], pgate_r[181],
     pgate_r[182], pgate_r[183], pgate_r[184], pgate_r[185],
     pgate_r[186], pgate_r[187], pgate_r[188], pgate_r[189],
     pgate_r[190], pgate_r[191], pgate_r[192], pgate_r[193],
     pgate_r[194], pgate_r[195], pgate_r[196], pgate_r[197],
     pgate_r[198], pgate_r[199], pgate_r[200], pgate_r[201],
     pgate_r[202], pgate_r[203], pgate_r[204], pgate_r[205],
     pgate_r[206], pgate_r[207], pgate_r[208], pgate_r[209],
     pgate_r[210], pgate_r[211], pgate_r[212], pgate_r[213],
     pgate_r[214], pgate_r[215], pgate_r[216], pgate_r[217],
     pgate_r[218], pgate_r[219], pgate_r[220], pgate_r[221],
     pgate_r[222], pgate_r[223], pgate_r[224], pgate_r[225],
     pgate_r[226], pgate_r[227], pgate_r[228], pgate_r[229],
     pgate_r[230], pgate_r[231], pgate_r[232], pgate_r[233],
     pgate_r[234], pgate_r[235], pgate_r[236], pgate_r[237],
     pgate_r[238], pgate_r[239], pgate_r[240], pgate_r[241],
     pgate_r[242], pgate_r[243], pgate_r[244], pgate_r[245],
     pgate_r[246], pgate_r[247], pgate_r[248], pgate_r[249],
     pgate_r[250], pgate_r[251], pgate_r[252], pgate_r[253],
     pgate_r[254], pgate_r[255], pgate_r[256], pgate_r[257],
     pgate_r[258], pgate_r[259], pgate_r[260], pgate_r[261],
     pgate_r[262], pgate_r[263], pgate_r[264], pgate_r[265],
     pgate_r[266], pgate_r[267], pgate_r[268], pgate_r[269],
     pgate_r[270], pgate_r[271], pgate_r[272], pgate_r[273],
     pgate_r[274], pgate_r[275], pgate_r[276], pgate_r[277],
     pgate_r[278], pgate_r[279], pgate_r[280], pgate_r[281],
     pgate_r[282], pgate_r[283], pgate_r[284], pgate_r[285],
     pgate_r[286], pgate_r[287], pgate_r[288], pgate_r[289],
     pgate_r[290], pgate_r[291], pgate_r[292], pgate_r[293],
     pgate_r[294], pgate_r[295], pgate_r[296], pgate_r[297],
     pgate_r[298], pgate_r[299], pgate_r[300], pgate_r[301],
     pgate_r[302], pgate_r[303], pgate_r[304], pgate_r[305],
     pgate_r[306], pgate_r[307], pgate_r[308], pgate_r[309],
     pgate_r[310], pgate_r[311], pgate_r[312], pgate_r[313],
     pgate_r[314], pgate_r[315], pgate_r[316], pgate_r[317],
     pgate_r[318], pgate_r[319], pgate_r[320], pgate_r[321],
     pgate_r[322], pgate_r[323], pgate_r[324], pgate_r[325],
     pgate_r[326], pgate_r[327], pgate_r[328], pgate_r[329],
     pgate_r[330], pgate_r[331], pgate_r[332], pgate_r[333],
     pgate_r[334], pgate_r[335], pgate_r[336], pgate_r[337],
     pgate_r[338], pgate_r[339], pgate_r[340], pgate_r[341],
     pgate_r[342], pgate_r[343], pgate_r[344], pgate_r[345],
     pgate_r[346], pgate_r[347], pgate_r[348], pgate_r[349],
     pgate_r[350], pgate_r[351], pgate_r[175], pgate_r[174],
     pgate_r[173], pgate_r[172], pgate_r[171], pgate_r[170],
     pgate_r[169], pgate_r[168], pgate_r[167], pgate_r[166],
     pgate_r[165], pgate_r[164], pgate_r[163], pgate_r[162],
     pgate_r[161], pgate_r[160], pgate_r[159], pgate_r[158],
     pgate_r[157], pgate_r[156], pgate_r[155], pgate_r[154],
     pgate_r[153], pgate_r[152], pgate_r[151], pgate_r[150],
     pgate_r[149], pgate_r[148], pgate_r[147], pgate_r[146],
     pgate_r[145], pgate_r[144], pgate_r[143], pgate_r[142],
     pgate_r[141], pgate_r[140], pgate_r[139], pgate_r[138],
     pgate_r[137], pgate_r[136], pgate_r[135], pgate_r[134],
     pgate_r[133], pgate_r[132], pgate_r[131], pgate_r[130],
     pgate_r[129], pgate_r[128], pgate_r[127], pgate_r[126],
     pgate_r[125], pgate_r[124], pgate_r[123], pgate_r[122],
     pgate_r[121], pgate_r[120], pgate_r[119], pgate_r[118],
     pgate_r[117], pgate_r[116], pgate_r[115], pgate_r[114],
     pgate_r[113], pgate_r[112], pgate_r[111], pgate_r[110],
     pgate_r[109], pgate_r[108], pgate_r[107], pgate_r[106],
     pgate_r[105], pgate_r[104], pgate_r[103], pgate_r[102],
     pgate_r[101], pgate_r[100], pgate_r[99], pgate_r[98], pgate_r[97],
     pgate_r[96], pgate_r[95], pgate_r[94], pgate_r[93], pgate_r[92],
     pgate_r[91], pgate_r[90], pgate_r[89], pgate_r[88], pgate_r[87],
     pgate_r[86], pgate_r[85], pgate_r[84], pgate_r[83], pgate_r[82],
     pgate_r[81], pgate_r[80], pgate_r[79], pgate_r[78], pgate_r[77],
     pgate_r[76], pgate_r[75], pgate_r[74], pgate_r[73], pgate_r[72],
     pgate_r[71], pgate_r[70], pgate_r[69], pgate_r[68], pgate_r[67],
     pgate_r[66], pgate_r[65], pgate_r[64], pgate_r[63], pgate_r[62],
     pgate_r[61], pgate_r[60], pgate_r[59], pgate_r[58], pgate_r[57],
     pgate_r[56], pgate_r[55], pgate_r[54], pgate_r[53], pgate_r[52],
     pgate_r[51], pgate_r[50], pgate_r[49], pgate_r[48], pgate_r[47],
     pgate_r[46], pgate_r[45], pgate_r[44], pgate_r[43], pgate_r[42],
     pgate_r[41], pgate_r[40], pgate_r[39], pgate_r[38], pgate_r[37],
     pgate_r[36], pgate_r[35], pgate_r[34], pgate_r[33], pgate_r[32],
     pgate_r[31], pgate_r[30], pgate_r[29], pgate_r[28], pgate_r[27],
     pgate_r[26], pgate_r[25], pgate_r[24], pgate_r[23], pgate_r[22],
     pgate_r[21], pgate_r[20], pgate_r[19], pgate_r[18], pgate_r[17],
     pgate_r[16], pgate_r[15], pgate_r[14], pgate_r[13], pgate_r[12],
     pgate_r[11], pgate_r[10], pgate_r[9], pgate_r[8], pgate_r[7],
     pgate_r[6], pgate_r[5], pgate_r[4], pgate_r[3], pgate_r[2],
     pgate_r[1], pgate_r[0]}), .end_of_startup_r({tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, jtag_rowtest_mode_rowu3_b, jtag_rowtest_mode_rowu2_b,
     tievdd, tievdd, tievdd, en_8bconfig_b, en_8bconfig_b,
     en_8bconfig_b, en_8bconfig_b}), .padeb_r(oeb_rbank[39:0]),
     .padin_r(in_rbank[39:0]), .bl_top(bl_top[1311:0]),
     .pado_t(out_tbank[47:0]), .padeb_t(oen_tbank[47:0]),
     .cf_t(cf_tbank[575:0]), .bl_bot(bl_bot[1311:0]),
     .pado_b(out_bbank[47:0]), .cf_b(cf_bbank[575:0]),
     .padeb_b(oen_bbank[47:0]), .padin_b(in_bbank[47:0]));
IO_LFTCELL Iio_lftcell ( .cbit({cf_lbank[0], cf_lbank[1], cf_lbank[2],
     cf_lbank[3], cf_lbank[4], cf_lbank[5], cf_lbank[6], cf_lbank[7],
     cf_lbank[8], cf_lbank[9], cf_lbank[10], cf_lbank[11],
     cf_lbank[12], cf_lbank[13], cf_lbank[14], cf_lbank[24],
     cf_lbank[25], cf_lbank[26], cf_lbank[27], cf_lbank[28],
     cf_lbank[29], cf_lbank[30], cf_lbank[31], cf_lbank[32],
     cf_lbank[33], cf_lbank[34], cf_lbank[35], cf_lbank[36],
     cf_lbank[37], cf_lbank[38], cf_lbank[48], cf_lbank[49],
     cf_lbank[50], cf_lbank[51], cf_lbank[52], cf_lbank[53],
     cf_lbank[54], cf_lbank[55], cf_lbank[56], cf_lbank[57],
     cf_lbank[58], cf_lbank[59], cf_lbank[60], cf_lbank[61],
     cf_lbank[62], cf_lbank[72], cf_lbank[73], cf_lbank[74],
     cf_lbank[75], cf_lbank[76], cf_lbank[77], cf_lbank[78],
     cf_lbank[79], cf_lbank[80], cf_lbank[81], cf_lbank[82],
     cf_lbank[83], cf_lbank[84], cf_lbank[85], cf_lbank[86],
     cf_lbank[96], cf_lbank[97], cf_lbank[98], cf_lbank[99],
     cf_lbank[100], cf_lbank[101], cf_lbank[102], cf_lbank[103],
     cf_lbank[104], cf_lbank[105], cf_lbank[106], cf_lbank[107],
     cf_lbank[108], cf_lbank[109], cf_lbank[110], cf_lbank[120],
     cf_lbank[121], cf_lbank[122], cf_lbank[123], cf_lbank[124],
     cf_lbank[125], cf_lbank[126], cf_lbank[127], cf_lbank[128],
     cf_lbank[129], cf_lbank[130], cf_lbank[131], cf_lbank[132],
     cf_lbank[133], cf_lbank[134], cf_lbank[144], cf_lbank[145],
     cf_lbank[146], cf_lbank[147], cf_lbank[148], cf_lbank[149],
     cf_lbank[150], cf_lbank[151], cf_lbank[152], cf_lbank[153],
     cf_lbank[154], cf_lbank[155], cf_lbank[156], cf_lbank[157],
     cf_lbank[158], cf_lbank[168], cf_lbank[169], cf_lbank[170],
     cf_lbank[171], cf_lbank[172], cf_lbank[173], cf_lbank[174],
     cf_lbank[175], cf_lbank[176], cf_lbank[177], cf_lbank[178],
     cf_lbank[179], cf_lbank[180], cf_lbank[181], cf_lbank[182],
     cf_lbank[192], cf_lbank[193], cf_lbank[194], cf_lbank[195],
     cf_lbank[196], cf_lbank[197], cf_lbank[198], cf_lbank[199],
     cf_lbank[200], cf_lbank[201], cf_lbank[202], cf_lbank[203],
     cf_lbank[204], cf_lbank[205], cf_lbank[206], cf_lbank[216],
     cf_lbank[217], cf_lbank[218], cf_lbank[219], cf_lbank[220],
     cf_lbank[221], cf_lbank[222], cf_lbank[223], cf_lbank[224],
     cf_lbank[225], cf_lbank[226], cf_lbank[227], cf_lbank[228],
     cf_lbank[229], cf_lbank[230], cf_lbank[240], cf_lbank[241],
     cf_lbank[242], cf_lbank[243], cf_lbank[244], cf_lbank[245],
     cf_lbank[246], cf_lbank[247], cf_lbank[248], cf_lbank[249],
     cf_lbank[250], cf_lbank[251], cf_lbank[252], cf_lbank[253],
     cf_lbank[254], cf_lbank[264], cf_lbank[265], cf_lbank[266],
     cf_lbank[267], cf_lbank[268], cf_lbank[269], cf_lbank[270],
     cf_lbank[271], cf_lbank[272], cf_lbank[273], cf_lbank[274],
     cf_lbank[275], cf_lbank[276], cf_lbank[277], cf_lbank[278],
     cf_lbank[288], cf_lbank[289], cf_lbank[290], cf_lbank[291],
     cf_lbank[292], cf_lbank[293], cf_lbank[294], cf_lbank[295],
     cf_lbank[296], cf_lbank[297], cf_lbank[298], cf_lbank[299],
     cf_lbank[300], cf_lbank[301], cf_lbank[302], cf_lbank[312],
     cf_lbank[313], cf_lbank[314], cf_lbank[315], cf_lbank[316],
     cf_lbank[317], cf_lbank[318], cf_lbank[319], cf_lbank[320],
     cf_lbank[321], cf_lbank[322], cf_lbank[323], cf_lbank[324],
     cf_lbank[325], cf_lbank[326], cf_lbank[336], cf_lbank[337],
     cf_lbank[338], cf_lbank[339], cf_lbank[340], cf_lbank[341],
     cf_lbank[342], cf_lbank[343], cf_lbank[344], cf_lbank[345],
     cf_lbank[346], cf_lbank[347], cf_lbank[348], cf_lbank[349],
     cf_lbank[350], cf_lbank[360], cf_lbank[361], cf_lbank[362],
     cf_lbank[363], cf_lbank[364], cf_lbank[365], cf_lbank[366],
     cf_lbank[367], cf_lbank[368], cf_lbank[369], cf_lbank[370],
     cf_lbank[371], cf_lbank[372], cf_lbank[373], cf_lbank[374],
     cf_lbank[384], cf_lbank[385], cf_lbank[386], cf_lbank[387],
     cf_lbank[388], cf_lbank[389], cf_lbank[390], cf_lbank[391],
     cf_lbank[392], cf_lbank[393], cf_lbank[394], cf_lbank[395],
     cf_lbank[396], cf_lbank[397], cf_lbank[398], cf_lbank[408],
     cf_lbank[409], cf_lbank[410], cf_lbank[411], cf_lbank[412],
     cf_lbank[413], cf_lbank[414], cf_lbank[415], cf_lbank[416],
     cf_lbank[417], cf_lbank[418], cf_lbank[419], cf_lbank[420],
     cf_lbank[421], cf_lbank[422], cf_lbank[432], cf_lbank[433],
     cf_lbank[434], cf_lbank[435], cf_lbank[436], cf_lbank[437],
     cf_lbank[438], cf_lbank[439], cf_lbank[440], cf_lbank[441],
     cf_lbank[442], cf_lbank[443], cf_lbank[444], cf_lbank[445],
     cf_lbank[446], cf_lbank[456], cf_lbank[457], cf_lbank[458],
     cf_lbank[459], cf_lbank[460], cf_lbank[461], cf_lbank[462],
     cf_lbank[463], cf_lbank[464], cf_lbank[465], cf_lbank[466],
     cf_lbank[467], cf_lbank[468], cf_lbank[469], cf_lbank[470]}),
     .out(out_lbank[39:0]), .oen(oen_lbank[39:0]), .in(in_lbank[39:0]),
     .VREFSSTL(VREFSSTL), .Pad(uio_lbank[39:0]));
IO_RGTCELL Iright_bank ( .REN({cf_rbank[0], cf_rbank[10], cf_rbank[24],
     cf_rbank[34], cf_rbank[48], cf_rbank[58], cf_rbank[72],
     cf_rbank[82], cf_rbank[96], cf_rbank[106], cf_rbank[120],
     cf_rbank[130], cf_rbank[144], cf_rbank[154], cf_rbank[168],
     cf_rbank[178], cf_rbank[192], cf_rbank[202], cf_rbank[216],
     cf_rbank[226], cf_rbank[240], cf_rbank[250], cf_rbank[264],
     cf_rbank[274], cf_rbank[288], cf_rbank[298], cf_rbank[312],
     cf_rbank[322], cf_rbank[336], cf_rbank[346], cf_rbank[360],
     cf_rbank[370], cf_rbank[384], cf_rbank[394], cf_rbank[408],
     cf_rbank[418], cf_rbank[432], cf_rbank[442], cf_rbank[456],
     cf_rbank[466]}), .Pad(uio_rbank[0:39]), .out({totdopad,
     out_rbank[0], out_rbank[1], out_rbank[2], out_rbank[3],
     out_rbank[4], out_rbank[5], out_rbank[6], out_rbank[7],
     out_rbank[8], out_rbank[9], out_rbank[10], out_rbank[11],
     out_rbank[12], out_rbank[13], out_rbank[14], out_rbank[15],
     out_rbank[16], out_rbank[17], out_rbank[18], out_rbank[19],
     out_rbank[20], out_rbank[21], out_rbank[22], out_rbank[23],
     out_rbank[24], out_rbank[25], out_rbank[26], out_rbank[27],
     out_rbank[28], out_rbank[29], out_rbank[30], out_rbank[31],
     out_rbank[32], out_rbank[33], out_rbank[34], out_rbank[35],
     out_rbank[36], out_rbank[37], out_rbank[38], out_rbank[39]}),
     .in({tdi_pad, tms_pad, tck_pad, trst_pad, in_rbank[0],
     in_rbank[1], in_rbank[2], in_rbank[3], in_rbank[4], in_rbank[5],
     in_rbank[6], in_rbank[7], in_rbank[8], in_rbank[9], in_rbank[10],
     in_rbank[11], in_rbank[12], in_rbank[13], in_rbank[14],
     in_rbank[15], in_rbank[16], in_rbank[17], in_rbank[18],
     in_rbank[19], in_rbank[20], in_rbank[21], in_rbank[22],
     in_rbank[23], in_rbank[24], in_rbank[25], in_rbank[26],
     in_rbank[27], in_rbank[28], in_rbank[29], in_rbank[30],
     in_rbank[31], in_rbank[32], in_rbank[33], in_rbank[34],
     in_rbank[35], in_rbank[36], in_rbank[37], in_rbank[38],
     in_rbank[39]}), .Tdo(tdo), .TRSTb(trstb), .Tdi(tdi), .Tms(tms),
     .Tck(tck), .oen({sdo_enable, oeb_rbank[0], oeb_rbank[1],
     oeb_rbank[2], oeb_rbank[3], oeb_rbank[4], oeb_rbank[5],
     oeb_rbank[6], oeb_rbank[7], oeb_rbank[8], oeb_rbank[9],
     oeb_rbank[10], oeb_rbank[11], oeb_rbank[12], oeb_rbank[13],
     oeb_rbank[14], oeb_rbank[15], oeb_rbank[16], oeb_rbank[17],
     oeb_rbank[18], oeb_rbank[19], oeb_rbank[20], oeb_rbank[21],
     oeb_rbank[22], oeb_rbank[23], oeb_rbank[24], oeb_rbank[25],
     oeb_rbank[26], oeb_rbank[27], oeb_rbank[28], oeb_rbank[29],
     oeb_rbank[30], oeb_rbank[31], oeb_rbank[32], oeb_rbank[33],
     oeb_rbank[34], oeb_rbank[35], oeb_rbank[36], oeb_rbank[37],
     oeb_rbank[38], oeb_rbank[39]}));
IO_TOPCELL Iio_topcell ( .vppin(vppin), .vpp(vpp), .REN({cf_tbank[0],
     cf_tbank[10], cf_tbank[24], cf_tbank[34], cf_tbank[48],
     cf_tbank[58], cf_tbank[72], cf_tbank[82], cf_tbank[96],
     cf_tbank[106], cf_tbank[120], cf_tbank[130], cf_tbank[144],
     cf_tbank[154], cf_tbank[168], cf_tbank[178], cf_tbank[192],
     cf_tbank[202], cf_tbank[216], cf_tbank[226], cf_tbank[240],
     cf_tbank[250], cf_tbank[264], cf_tbank[274], cf_tbank[288],
     cf_tbank[298], cf_tbank[312], cf_tbank[322], cf_tbank[336],
     cf_tbank[346], cf_tbank[360], cf_tbank[370], cf_tbank[384],
     cf_tbank[394], cf_tbank[408], cf_tbank[418], cf_tbank[432],
     cf_tbank[442], cf_tbank[456], cf_tbank[466], cf_tbank[480],
     cf_tbank[490], cf_tbank[504], cf_tbank[514], cf_tbank[528],
     cf_tbank[538], cf_tbank[552], cf_tbank[562]}),
     .Pad(uio_tbank[47:0]), .out(out_tbank[47:0]),
     .oen(oen_tbank[47:0]), .in(in_tbank[47:0]));
IO_BOTCELL Iio_botcell ( .done(cdone), .ctst_b(creset_b),
     .REN({cf_bbank[0], cf_bbank[10], cf_bbank[24], cf_bbank[34],
     cf_bbank[48], cf_bbank[58], cf_bbank[72], cf_bbank[82],
     cf_bbank[96], cf_bbank[106], cf_bbank[120], cf_bbank[130],
     cf_bbank[144], cf_bbank[154], cf_bbank[168], cf_bbank[178],
     cf_bbank[192], cf_bbank[202], cf_bbank[216], cf_bbank[226],
     cf_bbank[240], cf_bbank[250], cf_bbank[264], cf_bbank[274],
     cf_bbank[288], cf_bbank[298], cf_bbank[312], cf_bbank[322],
     cf_bbank[336], cf_bbank[346], cf_bbank[360], cf_bbank[370],
     cf_bbank[384], cf_bbank[394], cf_bbank[408], cf_bbank[418],
     cf_bbank[432], cf_bbank[442], cf_bbank[456], cf_bbank[466],
     cf_bbank[480], cf_bbank[490], cf_bbank[504], cf_bbank[514],
     cf_bbank[528], cf_bbank[538], cf_bbank[552], cf_bbank[562]}),
     .Pad(uio_bbank[0:47]), .in({in_bbank[0], in_bbank[1], in_bbank[2],
     in_bbank[3], in_bbank[4], in_bbank[5], in_bbank[6], in_bbank[7],
     in_bbank[8], in_bbank[9], in_bbank[10], in_bbank[11],
     in_bbank[12], in_bbank[13], in_bbank[14], in_bbank[15],
     in_bbank[16], in_bbank[17], in_bbank[18], in_bbank[19],
     in_bbank[20], in_bbank[21], in_bbank[22], in_bbank[23],
     in_bbank[24], in_bbank[25], in_bbank[26], in_bbank[27],
     in_bbank[28], in_bbank[29], in_bbank[30], in_bbank[31],
     in_bbank[32], in_bbank[33], in_bbank[34], in_bbank[35],
     in_bbank[36], in_bbank[37], in_bbank[38], in_bbank[39],
     in_bbank[40], in_bbank[41], in_bbank[42], in_bbank[43], cdone_in,
     in_bbank[44], in_bbank[45], in_bbank[46], in_bbank[47]}),
     .ctst_b_int(creset_b_int), .oen({oen_bbank[0], oen_bbank[1],
     oen_bbank[2], oen_bbank[3], oen_bbank[4], oen_bbank[5],
     oen_bbank[6], oen_bbank[7], oen_bbank[8], oen_bbank[9],
     oen_bbank[10], oen_bbank[11], oen_bbank[12], oen_bbank[13],
     oen_bbank[14], oen_bbank[15], oen_bbank[16], oen_bbank[17],
     oen_bbank[18], oen_bbank[19], oen_bbank[20], oen_bbank[21],
     oen_bbank[22], oen_bbank[23], oen_bbank[24], oen_bbank[25],
     oen_bbank[26], oen_bbank[27], oen_bbank[28], oen_bbank[29],
     oen_bbank[30], oen_bbank[31], oen_bbank[32], oen_bbank[33],
     oen_bbank[34], oen_bbank[35], oen_bbank[36], oen_bbank[37],
     oen_bbank[38], oen_bbank[39], oen_bbank[40], oen_bbank[41],
     oen_bbank[42], oen_bbank[43], cdone_out, oen_bbank[44],
     oen_bbank[45], oen_bbank[46], oen_bbank[47]}), .out({out_bbank[0],
     out_bbank[1], out_bbank[2], out_bbank[3], out_bbank[4],
     out_bbank[5], out_bbank[6], out_bbank[7], out_bbank[8],
     out_bbank[9], out_bbank[10], out_bbank[11], out_bbank[12],
     out_bbank[13], out_bbank[14], out_bbank[15], out_bbank[16],
     out_bbank[17], out_bbank[18], out_bbank[19], out_bbank[20],
     out_bbank[21], out_bbank[22], out_bbank[23], out_bbank[24],
     out_bbank[25], out_bbank[26], out_bbank[27], out_bbank[28],
     out_bbank[29], out_bbank[30], out_bbank[31], out_bbank[32],
     out_bbank[33], out_bbank[34], out_bbank[35], out_bbank[36],
     out_bbank[37], out_bbank[38], out_bbank[39], out_bbank[40],
     out_bbank[41], out_bbank[42], out_bbank[43], tievdd,
     out_bbank[44], out_bbank[45], out_bbank[46], out_bbank[47]}));

endmodule
// Library - tsmcN65lo, Cell - nand3_25, View - schematic
// LAST TIME SAVED: Mar 29 20:19:50 2006
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module nand3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(net21), .B(Gb), .G(C), .S(G));
nch_25  M2 ( .D(net25), .B(Gb), .G(B), .S(net21));
nch_25  NM1 ( .D(Y), .B(Gb), .G(A), .S(net25));
pch_25  PM1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M1 ( .D(Y), .B(Pb), .G(C), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(P));

endmodule
// Library - tsmcN65lo, Cell - nor3_25, View - schematic
// LAST TIME SAVED: Mar 29 20:26:16 2006
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module nor3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M2 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  M3 ( .D(Y), .B(Gb), .G(C), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  M1 ( .D(Y), .B(Pb), .G(C), .S(net16));
pch_25  PM1 ( .D(net12), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(net16), .B(Pb), .G(B), .S(net12));

endmodule
// Library - NVCM, Cell - ml_ls_vdd2vdd25, View - schematic
// LAST TIME SAVED: Apr  4 14:26:57 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
pch_25  M13 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
pch_25  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));
pch_25  M6 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
nch_25  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
nch_25  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));

endmodule
// Library - tsmcN65lo, Cell - inv_25, View - schematic
// LAST TIME SAVED: Mar 29 20:14:12 2006
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module inv_25 ( OUT, G, Gb, IN, P, Pb );
output  OUT;

input  G, Gb, IN, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  NM1 ( .D(OUT), .B(Gb), .G(IN), .S(G));
pch_25  PM1 ( .D(OUT), .B(Pb), .G(IN), .S(P));

endmodule
// Library - sbtlibn65lp, Cell - vddp_tiehigh, View - schematic
// LAST TIME SAVED: May  8 16:23:22 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module vddp_tiehigh ( vddp_tieh );
inout  vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M8 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net9), .S(vddp_));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tielow, View - schematic
// LAST TIME SAVED: May  8 16:23:59 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module vdd_tielow ( gnd_tiel );
inout  gnd_tiel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(gnd_tiel), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(net9), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_chip_spare, View - schematic
// LAST TIME SAVED: Sep 11 18:02:11 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_chip_spare (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(net96), .B(net85), .G(net286), .S(net85));
pch_25  M5 ( .D(net85), .B(net123), .G(net114), .S(net123));
pch_25  M3 ( .D(net108), .B(net89), .G(net316), .S(net89));
pch_25  M2 ( .D(net89), .B(net126), .G(net119), .S(net126));
nch_25  M7 ( .D(net100), .B(GND_), .G(net286), .S(gnd_));
nch_25  M1 ( .D(net96), .B(GND_), .G(net121), .S(net100));
nch_25  M6 ( .D(net104), .B(GND_), .G(net316), .S(gnd_));
nch_25  M4 ( .D(net108), .B(GND_), .G(net121), .S(net104));
ml_hv_ls_inv I132 ( .sel_b_25(net316), .sel_25(net405),
     .out_b_hv(net119), .in_hv(net126), .vddp_tieh(net121));
ml_hv_ls_inv Iml_hv_ls_inv_vppt ( .sel_b_25(net286), .sel_25(net404),
     .out_b_hv(net114), .in_hv(net123), .vddp_tieh(net121));
rppolywo_m  R8 ( .MINUS(vddp_), .PLUS(net123), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(vddp_), .PLUS(net126), .BULK(gnd_));
nand3_25 I257 ( .B(net0373), .A(net0373), .Y(net0397), .C(net0373),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I256 ( .B(net0381), .A(net0381), .Y(net0373), .C(net0381),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I255 ( .B(net215), .A(net215), .Y(net0381), .C(net215),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I248 ( .B(net0397), .A(net0397), .Y(net0405), .C(net0397),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I247 ( .B(net0405), .A(net0405), .Y(net0413), .C(net0405),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I245 ( .B(net0413), .A(net0413), .Y(net0421), .C(net0413),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I244 ( .B(net0421), .A(net0421), .Y(net0453), .C(net0421),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I231 ( .B(net0453), .A(net0453), .Y(net0445), .C(net0453),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I233 ( .B(net0437), .A(net0437), .Y(net0429), .C(net0437),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I234 ( .B(net0429), .A(net0429), .Y(net0595), .C(net0429),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I232 ( .B(net0445), .A(net0445), .Y(net0437), .C(net0445),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nor3_25 I215 ( .B(net0460), .A(net0460), .C(net0460), .Y(net0594),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I214 ( .B(net0468), .A(net0468), .C(net0468), .Y(net0460),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I212 ( .B(net0476), .A(net0476), .C(net0476), .Y(net0468),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I211 ( .B(net160), .A(net160), .C(net160), .Y(net0492),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I209 ( .B(net0500), .A(net0500), .C(net0500), .Y(net0476),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I42 ( .B(net191), .A(net191), .C(net191), .Y(net160), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I78 ( .B(net199), .A(net199), .C(net199), .Y(net191), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I83 ( .B(net207), .A(net207), .C(net207), .Y(net199), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I84 ( .B(net215), .A(net215), .C(net215), .Y(net207), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I210 ( .B(net0492), .A(net0492), .C(net0492), .Y(net0500),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
inv_hvt I120 ( .A(net253), .Y(net249));
inv_hvt I119 ( .A(net231), .Y(net253));
inv_hvt I118 ( .A(net231), .Y(net258));
inv_hvt I117 ( .A(net258), .Y(net254));
inv_hvt I319 ( .A(net263), .Y(net259));
inv_hvt I323 ( .A(net231), .Y(net263));
inv_hvt I57 ( .A(net231), .Y(net268));
inv_hvt I58 ( .A(net268), .Y(net264));
ml_ls_vdd2vdd25 I122 ( .in(net249), .sup(vddp_), .out_vddio_b(net291),
     .out_vddio(net252), .in_b(net253));
ml_ls_vdd2vdd25 I121 ( .in(net254), .sup(vddp_), .out_vddio_b(net297),
     .out_vddio(net257), .in_b(net258));
ml_ls_vdd2vdd25 I335 ( .in(net259), .sup(vddp_), .out_vddio_b(net303),
     .out_vddio(net262), .in_b(net263));
ml_ls_vdd2vdd25 I56 ( .in(net264), .sup(vddp_), .out_vddio_b(net309),
     .out_vddio(net267), .in_b(net268));
inv_25 I126 ( .IN(net291), .OUT(net271), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I125 ( .IN(net297), .OUT(net272), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I139 ( .IN(net405), .OUT(net316), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(net404), .OUT(net286), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I384 ( .IN(net303), .OUT(net274), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I54 ( .IN(net309), .OUT(net273), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nand3_hvt I185 ( .Y(net0665), .B(net0661), .C(net0661), .A(net0661));
nand3_hvt I186 ( .Y(net0661), .B(net0657), .C(net0657), .A(net0657));
nand3_hvt I187 ( .Y(net0657), .B(net0653), .C(net0653), .A(net0653));
nand3_hvt I188 ( .Y(net0653), .B(net0649), .C(net0649), .A(net0649));
nand3_hvt I183 ( .Y(net0649), .B(net281), .C(net281), .A(net281));
nand3_hvt I246 ( .Y(net328), .B(net324), .C(net324), .A(net324));
nand3_hvt I61 ( .Y(net332), .B(net328), .C(net328), .A(net328));
nand3_hvt I62 ( .Y(net336), .B(net332), .C(net332), .A(net332));
nand3_hvt I63 ( .Y(net340), .B(net336), .C(net336), .A(net336));
nand3_hvt I64 ( .Y(net360), .B(net340), .C(net340), .A(net340));
nand3_hvt I104 ( .Y(net281), .B(net344), .C(net344), .A(net344));
nand3_hvt I105 ( .Y(net344), .B(net348), .C(net348), .A(net348));
nand3_hvt I106 ( .Y(net348), .B(net352), .C(net352), .A(net352));
nand3_hvt I107 ( .Y(net352), .B(net356), .C(net356), .A(net356));
nand3_hvt I108 ( .Y(net356), .B(net360), .C(net360), .A(net360));
nand3_hvt I184 ( .Y(net0596), .B(net0665), .C(net0665), .A(net0665));
nor3_hvt I177 ( .B(net0732), .Y(net0728), .A(net0732), .C(net0732));
nor3_hvt I178 ( .B(net0728), .Y(net0724), .A(net0728), .C(net0728));
nor3_hvt I179 ( .B(net0724), .Y(net0720), .A(net0724), .C(net0724));
nor3_hvt I180 ( .B(net0720), .Y(net0716), .A(net0720), .C(net0720));
nor3_hvt I181 ( .B(net0716), .Y(net0712), .A(net0716), .C(net0716));
nor3_hvt I182 ( .B(net0712), .Y(net0597), .A(net0712), .C(net0712));
nor3_hvt I65 ( .B(net363), .Y(net383), .A(net363), .C(net363));
nor3_hvt I70 ( .B(net367), .Y(net363), .A(net367), .C(net367));
nor3_hvt I71 ( .B(net371), .Y(net367), .A(net371), .C(net371));
nor3_hvt I72 ( .B(net375), .Y(net371), .A(net375), .C(net375));
nor3_hvt I73 ( .B(net379), .Y(net375), .A(net379), .C(net379));
nor3_hvt I99 ( .B(net383), .Y(net387), .A(net383), .C(net383));
nor3_hvt I100 ( .B(net387), .Y(net391), .A(net387), .C(net387));
nor3_hvt I101 ( .B(net391), .Y(net395), .A(net391), .C(net391));
nor3_hvt I102 ( .B(net395), .Y(net399), .A(net395), .C(net395));
nor3_hvt I103 ( .B(net399), .Y(net0732), .A(net399), .C(net399));
vddp_tiehigh I140 ( .vddp_tieh(net121));
vdd_tielow I154 ( .gnd_tiel(net405));
vdd_tielow I155 ( .gnd_tiel(net404));
vdd_tielow I153 ( .gnd_tiel(net231));
vdd_tielow I146 ( .gnd_tiel(net215));
vdd_tielow I145 ( .gnd_tiel(net324));
vdd_tielow I144 ( .gnd_tiel(net379));

endmodule
// Library - NVCM, Cell - ml_chip_buf, View - schematic
// LAST TIME SAVED: Feb 26 16:35:06 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_chip_buf ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(in), .Y(net120));
inv_hvt I45 ( .A(net120), .Y(out));

endmodule
// Library - misc, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jun  5 11:34:46 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - NVCM, Cell - ml_chip_buf_top, View - schematic
// LAST TIME SAVED: Apr 21 14:59:16 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_chip_buf_top ( fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_trim_vbg_buf, fsm_vpgmwl_buf,
     fsm_wgnden_buf, fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmvfy, fsm_trim_vbg, fsm_vpgmwl, fsm_wgnden );
output  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_wgnden_buf;

input  fsm_lshven, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmvfy,
     fsm_wgnden;

output [2:0]  fsm_vpgmwl_buf;
output [3:0]  fsm_trim_vbg_buf;

input [3:0]  fsm_trim_vbg;
input [2:0]  fsm_vpgmwl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_chip_buf I50_2_ ( .in(fsm_vpgmwl[2]), .out(fsm_vpgmwl_buf[2]));
ml_chip_buf I50_1_ ( .in(fsm_vpgmwl[1]), .out(fsm_vpgmwl_buf[1]));
ml_chip_buf I50_0_ ( .in(fsm_vpgmwl[0]), .out(fsm_vpgmwl_buf[0]));
ml_chip_buf I56 ( .in(fsm_wgnden), .out(fsm_wgnden_buf));
ml_chip_buf I49_3_ ( .in(fsm_trim_vbg[3]), .out(fsm_trim_vbg_buf[3]));
ml_chip_buf I49_2_ ( .in(fsm_trim_vbg[2]), .out(fsm_trim_vbg_buf[2]));
ml_chip_buf I49_1_ ( .in(fsm_trim_vbg[1]), .out(fsm_trim_vbg_buf[1]));
ml_chip_buf I49_0_ ( .in(fsm_trim_vbg[0]), .out(fsm_trim_vbg_buf[0]));
ml_chip_buf I51 ( .in(fsm_lshven), .out(fsm_lshven_buf));
ml_chip_buf I53 ( .in(fsm_nvcmen), .out(fsm_nvcmen_buf));
ml_chip_buf I54 ( .in(fsm_pgmdisc), .out(fsm_pgmdisc_buf));
ml_chip_buf I57 ( .in(fsm_pgmvfy), .out(fsm_pgmvfy_buf));
ml_chip_buf I55 ( .in(fsm_pgm), .out(fsm_pgm_buf));

endmodule
// Library - NVCM, Cell - ml_hv_invx3, View - schematic
// LAST TIME SAVED: Jan 25 09:27:09 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv_invx3 ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_switch, View - schematic
// LAST TIME SAVED: Feb  1 16:53:01 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_lshv_6v_switch ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M11 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv_hotsw, View - schematic
// LAST TIME SAVED: Jan 24 11:18:40 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3 Ihv_invx3 ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));
ml_lshv_6v_switch Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM, Cell - ml_hv2vddp_sw, View - schematic
// LAST TIME SAVED: May  1 11:01:33 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv2vddp_sw ( out_hv, hv2vddp, vddp_tieh );
inout  out_hv;

input  hv2vddp, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(sw_vddp_b),
     .sel_25(net035), .out_b_hv(sw_vpp_b), .in_hv(out_hv),
     .vddp_tieh(vddp_tieh));
pch_25  M1 ( .D(net27), .B(out_hv), .G(sw_vpp_b), .S(out_hv));
pch_25  M0 ( .D(net27), .B(vddp_), .G(sw_vddp_b), .S(vddp_));
inv_25 I62 ( .IN(net37), .OUT(sw_vddp_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I71 ( .IN(net060), .OUT(net035), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net060),
     .out_vddio(net37), .in_b(net46));
inv_hvt I65 ( .A(hv2vddp), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));

endmodule
// Library - NVCM, Cell - ml_vpp_ref_sw, View - schematic
// LAST TIME SAVED: Mar 21 16:41:35 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpp_ref_sw ( in, out, sel_b_25 );
inout  in, out;

input  sel_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I281 ( .IN(sel_b_25), .OUT(net122), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M12 ( .D(out), .B(GND_), .G(net122), .S(in));
pch_25  M14 ( .D(in), .B(vddp_), .G(sel_b_25), .S(out));

endmodule
// Library - NVCM, Cell - ml_vpp_ref, View - schematic
// LAST TIME SAVED: Apr  7 18:49:59 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpp_ref ( vref_25, bgr, pumpen_25, vppwl_25 );
inout  vref_25;

input  bgr, pumpen_25;

input [2:0]  vppwl_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_b_25;

wire  [7:0]  red_dec_25;



nch_na25  M0 ( .D(net179), .B(GND_), .G(ctrl_gate_25),
     .S(bgr_mirror_25));
nand3_25 I44_7_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[7]),
     .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_6_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[6]),
     .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_5_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[5]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_4_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[4]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_3_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[3]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_2_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[2]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_1_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[1]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_0_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[0]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
ml_vpp_ref_sw I281 ( .in(net92), .out(vref_25),
     .sel_b_25(red_dec_25[6]));
ml_vpp_ref_sw I287 ( .in(net95), .out(vref_25),
     .sel_b_25(red_dec_25[4]));
ml_vpp_ref_sw I283 ( .in(net98), .out(vref_25),
     .sel_b_25(red_dec_25[7]));
ml_vpp_ref_sw I290 ( .in(net0100), .out(vref_25),
     .sel_b_25(red_dec_25[0]));
ml_vpp_ref_sw I288 ( .in(net104), .out(vref_25),
     .sel_b_25(red_dec_25[3]));
ml_vpp_ref_sw I284 ( .in(net139), .out(vref_25),
     .sel_b_25(red_dec_25[5]));
ml_vpp_ref_sw I291 ( .in(net110), .out(vref_25),
     .sel_b_25(red_dec_25[1]));
ml_vpp_ref_sw I292 ( .in(net113), .out(vref_25),
     .sel_b_25(red_dec_25[2]));
nmoscap_25  C3 ( .MINUS(net0129), .PLUS(net0113));
nmoscap_25  C2 ( .MINUS(gnd_), .PLUS(ctrl_gate_25));
inv_25 I38 ( .IN(pumpen_25), .OUT(vppref_en_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_2_ ( .IN(vppwl_25[2]), .OUT(vppwl_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_1_ ( .IN(vppwl_25[1]), .OUT(vppwl_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_0_ ( .IN(vppwl_25[0]), .OUT(vppwl_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
rppolywo_m  R11 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R13 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R14 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R15 ( .MINUS(net104), .PLUS(net95), .BULK(GND_));
rppolywo_m  R16 ( .MINUS(net104), .PLUS(net95), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net95), .PLUS(net139), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net95), .PLUS(net139), .BULK(GND_));
rppolywo_m  R19 ( .MINUS(net139), .PLUS(net92), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(net139), .PLUS(net92), .BULK(GND_));
rppolywo_m  R21 ( .MINUS(net92), .PLUS(net98), .BULK(GND_));
rppolywo_m  R22 ( .MINUS(net92), .PLUS(net98), .BULK(GND_));
rppolywo_m  R25 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R24 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(net0100), .BULK(GND_));
rppolywo_m  R5 ( .MINUS(net0100), .PLUS(net110), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net0100), .PLUS(net110), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(bgr_mirror_25), .PLUS(net0129), .BULK(GND_));
nch_25  M10 ( .D(net163), .B(GND_), .G(bgr), .S(gnd_));
nch_25  M14 ( .D(net0113), .B(GND_), .G(vppref_en_b_25), .S(gnd_));
nch_25  M15 ( .D(ctrl_gate_25), .B(GND_), .G(vppref_en_b_25),
     .S(gnd_));
nch_25  M8 ( .D(ctrl_gate_25), .B(GND_), .G(bgr_mirror_25),
     .S(net163));
nch_25  M13 ( .D(net0113), .B(GND_), .G(bgr), .S(net163));
pch_25  M18 ( .D(net179), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
pch_25  M5 ( .D(ctrl_gate_25), .B(vddp_), .G(net0113), .S(net175));
pch_25  M6 ( .D(net0113), .B(vddp_), .G(net0113), .S(net175));
pch_25  M7 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Aug  3 14:03:13 2007
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module sbtlibn65lp_ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - NVCM, Cell - ml_vpp_ctrl, View - schematic
// LAST TIME SAVED: Apr 30 14:24:32 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpp_ctrl ( pumpen_25, vpint_en, vpp_2_vdd, vppdisc_25,
     vppwl_25, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_vpgmwl_buf, fsm_wgnden );
output  pumpen_25, vpint_en, vpp_2_vdd, vppdisc_25;

input  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint, fsm_wgnden;

output [2:0]  vppwl_25;

input [2:0]  fsm_vpgmwl_buf;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  net068;

wire  [0:2]  net038;

wire  [0:2]  net082;

wire  [0:2]  net092;



nand4_hvt I75 ( .D(fsm_pgm_buf), .C(fsm_lshven_buf), .A(net0127),
     .Y(net046), .B(net0127));
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(net0122));
nor2_hvt I111 ( .A(vpp_pumpen_b), .B(net080), .Y(net0133));
nor2_hvt I87 ( .A(vpp_pumpen), .Y(net036), .B(fsm_pgmdisc_buf));
sbtlibn65lp_ml_dff_schematic I77 ( .CLK(net084), .QN(vpp_pumpen_b),
     .R(pgm_dis), .D(vdd_tieh), .Q(vpp_pumpen));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
nand3_hvt I79 ( .C(net086), .A(fsm_pgm_buf), .Y(pgm_dis),
     .B(fsm_nvcmen_buf));
nand2_hvt I104 ( .A(fsm_tm_xforce), .Y(net049), .B(fsm_tm_xvppint));
inv_25 I95_2_ ( .IN(net068[0]), .OUT(vppwl_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_1_ ( .IN(net068[1]), .OUT(vppwl_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_0_ ( .IN(net068[2]), .OUT(vppwl_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I81 ( .IN(net073), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(net088), .OUT(vppdisc_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I96_2_ ( .in(net082[0]), .sup(vddp_),
     .out_vddio_b(net068[0]), .out_vddio(net038[0]), .in_b(net092[0]));
ml_ls_vdd2vdd25 I96_1_ ( .in(net082[1]), .sup(vddp_),
     .out_vddio_b(net068[1]), .out_vddio(net038[1]), .in_b(net092[1]));
ml_ls_vdd2vdd25 I96_0_ ( .in(net082[2]), .sup(vddp_),
     .out_vddio_b(net068[2]), .out_vddio(net038[2]), .in_b(net092[2]));
ml_ls_vdd2vdd25 I84 ( .in(net0133), .sup(vddp_), .out_vddio_b(net073),
     .out_vddio(net074), .in_b(net0134));
ml_ls_vdd2vdd25 I173 ( .in(fsm_pgmdisc_buf), .sup(vddp_),
     .out_vddio_b(net088), .out_vddio(net048), .in_b(net0106));
inv_hvt I107 ( .A(net0122), .Y(net0124));
inv_hvt I109 ( .A(fsm_pgmvfy_buf), .Y(net0127));
inv_hvt I131 ( .A(net049), .Y(net080));
inv_hvt I110_2_ ( .A(net092[0]), .Y(net082[0]));
inv_hvt I110_1_ ( .A(net092[1]), .Y(net082[1]));
inv_hvt I110_0_ ( .A(net092[2]), .Y(net082[2]));
inv_hvt I76 ( .A(net046), .Y(net084));
inv_hvt I108 ( .A(fsm_pgmdisc_buf), .Y(net0122));
inv_hvt I78 ( .A(net0124), .Y(net086));
inv_hvt I113 ( .A(vpp_pumpen_b), .Y(vpint_en));
inv_hvt I91 ( .A(net036), .Y(net089));
inv_hvt I90 ( .A(net089), .Y(vpp_2_vdd));
inv_hvt I98_2_ ( .A(fsm_vpgmwl_buf[2]), .Y(net092[0]));
inv_hvt I98_1_ ( .A(fsm_vpgmwl_buf[1]), .Y(net092[1]));
inv_hvt I98_0_ ( .A(fsm_vpgmwl_buf[0]), .Y(net092[2]));
inv_hvt I112 ( .A(net0133), .Y(net0134));
inv_hvt I101 ( .A(fsm_pgmdisc_buf), .Y(net0106));

endmodule
// Library - NVCM, Cell - ml_vpp_reg, View - schematic
// LAST TIME SAVED: May  3 15:48:51 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpp_reg ( slow_25, bgr, pbias_25, pump_in, vpp_int,
     pumpen_25, vppdisc_25, vref_25 );
output  slow_25;

inout  bgr, pbias_25, pump_in, vpp_int;

input  pumpen_25, vppdisc_25, vref_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I261 ( .vddp_tieh(net0208));
nch_na25  M11 ( .D(net0199), .B(GND_), .G(vppdisc_25), .S(VDD_));
nch_na25  M22 ( .D(vpp_int), .B(GND_), .G(pump_gate), .S(pump_in));
nch_na25  M1 ( .D(GND_), .B(GND_), .G(pump_gate), .S(GND_));
nch_na25  M10 ( .D(net0203), .B(GND_), .G(net0208), .S(net0199));
nch_na25  M5 ( .D(pump_opamp_out), .B(GND_), .G(vpp_int),
     .S(pump_opamp_out));
inv_25 I211 ( .IN(en_buf_b_25), .OUT(en_buf_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I212 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
pch_25  M31 ( .D(net0203), .B(net0165), .G(dis_pgate_25), .S(net0165));
pch_25  M0 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
pch_25  M9 ( .D(net0166), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
pch_25  M14 ( .D(pump_opamp_out), .B(net125), .G(vref_25), .S(net125));
pch_25  M18 ( .D(net122), .B(vpp_int), .G(net122), .S(vpp_int));
pch_25  M13 ( .D(net124), .B(net125), .G(vdiv), .S(net125));
pch_25  M32 ( .D(dis_pgate_25), .B(vddp_), .G(dis_pgate_25),
     .S(vddp_));
pch_25  M33 ( .D(dis_pgate_25), .B(vddp_), .G(vppdisc_25), .S(vddp_));
pch_25  M12 ( .D(net125), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M19 ( .D(net134), .B(net122), .G(net134), .S(net122));
pch_25  M21 ( .D(net138), .B(net134), .G(net138), .S(net134));
pch_25  M23 ( .D(net142), .B(net138), .G(net142), .S(net138));
pch_25  M24 ( .D(vdiv), .B(net142), .G(vdiv), .S(net142));
pch_25  M25 ( .D(net0224), .B(vdiv), .G(net0224), .S(vdiv));
pch_25  M4_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
pch_25  M4_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
nch_25  M40 ( .D(dis_pgate_25), .B(GND_), .G(vppdisc_25), .S(gnd_));
nch_25  M8 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
nch_25  M16 ( .D(net124), .B(GND_), .G(net124), .S(net155));
nch_25  M17 ( .D(net155), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M6 ( .D(vpp_int), .B(GND_), .G(en_buf_25), .S(net168));
nch_25  M20 ( .D(slow_25), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M7 ( .D(net168), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M41 ( .D(net0224), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M15 ( .D(pump_opamp_out), .B(GND_), .G(net124), .S(net155));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net0250));
rppolywo_m  R5 ( .MINUS(net0165), .PLUS(vpp_int), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(pump_gate), .PLUS(pump_in), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net0247), .PLUS(net0250), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net0247), .BULK(GND_));

endmodule
// Library - misc, Cell - ml_mux3_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:41 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_mux3_hvt ( out, in0, in1, in2, sel );
output  out;

input  in0, in1, in2;

input [3:0]  sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I25 ( .A(sel[2]), .Y(net26));
inv_hvt I24 ( .A(sel[1]), .Y(net28));
inv_hvt I21 ( .A(sel[0]), .Y(net30));
txgate_hvt I23 ( .in(in1), .out(out), .pp(net28), .nn(sel[1]));
txgate_hvt I20 ( .in(in0), .out(out), .pp(net30), .nn(sel[0]));
txgate_hvt I26 ( .in(in2), .out(out), .pp(net26), .nn(sel[2]));
nch_hvt  MN19 ( .D(out), .B(gnd_), .G(sel[3]), .S(gnd_));

endmodule
// Library - tsmcN65lo, Cell - nand2_25, View - schematic
// LAST TIME SAVED: Mar 29 20:17:19 2006
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module nand2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(net16), .B(Gb), .G(B), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(A), .S(net16));
pch_25  M2 ( .D(Y), .B(Pb), .G(B), .S(P));
pch_25  PM1 ( .D(Y), .B(Pb), .G(A), .S(P));

endmodule
// Library - NVCM, Cell - ml_vpp_vco, View - schematic
// LAST TIME SAVED: Apr  8 16:31:55 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpp_vco ( clk_25_0, pbias_25, slow_25, en_25, freq_25 );
output  clk_25_0;

inout  pbias_25, slow_25;

input  en_25;

input [1:0]  freq_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:1]  freq_b_25;



nch_na25  M4 ( .D(GND_), .B(GND_), .G(net173), .S(GND_));
nch_na25  M15 ( .D(GND_), .B(GND_), .G(net185), .S(GND_));
nch_na25  M16 ( .D(GND_), .B(GND_), .G(net193), .S(GND_));
nch_na25  M2 ( .D(GND_), .B(GND_), .G(net189), .S(GND_));
nch_25  M5 ( .D(net173), .B(GND_), .G(net185), .S(net177));
nch_25  M6 ( .D(net177), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M13 ( .D(net181), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M14 ( .D(net185), .B(GND_), .G(net193), .S(net181));
nch_25  M8 ( .D(net189), .B(GND_), .G(net173), .S(net201));
nch_25  M17 ( .D(net193), .B(GND_), .G(net195), .S(net197));
nch_25  M18 ( .D(net197), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M1 ( .D(net201), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M23 ( .D(pbias_osc_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M24 ( .D(slow_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M25 ( .D(nbias_osc_25), .B(GND_), .G(en_25), .S(slow_25));
pch_25  M7 ( .D(net173), .B(vddp_), .G(net185), .S(net236));
pch_25  M10 ( .D(net236), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M9 ( .D(net248), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M3 ( .D(net189), .B(vddp_), .G(net173), .S(net248));
pch_25  M11 ( .D(net256), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M12 ( .D(net185), .B(vddp_), .G(net193), .S(net256));
pch_25  M19 ( .D(net193), .B(vddp_), .G(net195), .S(net260));
pch_25  M20 ( .D(net260), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M22 ( .D(pbias_osc_25), .B(vddp_), .G(en_b_25), .S(net228));
pch_25  M26_1_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M26_0_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_1_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_0_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M28 ( .D(net212), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M29 ( .D(nbias_osc_25), .B(vddp_), .G(freq_25[0]), .S(net212));
pch_25  M30 ( .D(nbias_osc_25), .B(vddp_), .G(freq_b_25[1]),
     .S(net208));
pch_25  M21 ( .D(net228), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
nand2_25 I96 ( .G(GND_), .Pb(vddp_), .A(net189), .Y(net195), .P(vddp_),
     .B(en_25), .Gb(GND_));
inv_25 I201 ( .IN(net195), .OUT(clk_25_0), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I188 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I199 ( .IN(freq_25[1]), .OUT(freq_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));

endmodule
// Library - NVCM, Cell - ml_vpp_pump, View - schematic
// LAST TIME SAVED: Apr  7 18:25:20 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpp_pump ( pump_in, clkin_25, en_25 );
inout  pump_in;

input  clkin_25, en_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));
nmoscap_25  C1 ( .MINUS(clk_b_25), .PLUS(s_3));
pch_25  M0 ( .D(net23), .B(vddp_), .G(net64), .S(vddp_));
inv_25 I194 ( .IN(clkin_25), .OUT(net70), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(en_25), .OUT(net64), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I210 ( .IN(net28), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I219 ( .IN(net40), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I220 ( .IN(net34), .OUT(net46), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I221 ( .IN(net46), .OUT(net40), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I224 ( .IN(clkin_25), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I209 ( .IN(net70), .OUT(net28), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
nch_na25  M10 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
nch_na25  M11 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
nch_na25  M12 ( .D(s_2), .B(GND_), .G(s_2), .S(s_3));
nch_na25  M22 ( .D(net23), .B(GND_), .G(net23), .S(s_0));
nch_na25  M1 ( .D(s_3), .B(GND_), .G(s_3), .S(pump_in));

endmodule
// Library - NVCM, Cell - ml_vpp_pumpx3, View - schematic
// LAST TIME SAVED: Apr  8 17:28:05 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpp_pumpx3 ( pump_in, clkin_0_25, pumpen_25 );
inout  pump_in;

input  clkin_0_25, pumpen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I195 ( .IN(clkin_0_25), .OUT(net13), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I84 ( .IN(net13), .OUT(net024), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
ml_vpp_pump Ivpp_pump_0 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(clkin_0_25));
ml_vpp_pump I79 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net024));
ml_vpp_pump Ivpp_pump_1 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net13));

endmodule
// Library - NVCM, Cell - ml_vppint_top, View - schematic
// LAST TIME SAVED: May  1 11:06:26 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vppint_top ( vpint_en, vpp_int, bgr, fsm_lshven_buf,
     fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf, fsm_pgmvfy_buf,
     fsm_tm_xforce, fsm_tm_xvppint, fsm_vpgmwl_buf, fsm_wgnden_buf );
output  vpint_en;

inout  vpp_int;

input  bgr, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_wgnden_buf;

input [2:0]  fsm_vpgmwl_buf;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_25;

wire  [1:0]  freq_25;



ml_hv2vddp_sw Ivpxa_2vddp_sw ( .hv2vddp(vpp_2_vdd),
     .vddp_tieh(vddp_tieh), .out_hv(vpp_int));
inv_25 I38 ( .IN(vddp_tieh), .OUT(freq_25[1]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I86 ( .IN(vddp_tieh), .OUT(freq_25[0]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
ml_vpp_ref Ivpp_ref ( .vref_25(vref_25), .vppwl_25(vppwl_25[2:0]),
     .pumpen_25(pumpen_25), .bgr(bgr));
ml_vpp_ctrl Ivpp_ctrl ( .vpint_en(vpint_en),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .vppdisc_25(vppdisc_25), .fsm_wgnden(fsm_wgnden_buf),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf), .vppwl_25(vppwl_25[2:0]),
     .vpp_2_vdd(vpp_2_vdd), .pumpen_25(pumpen_25));
ml_vpp_reg Ivpp_reg ( .bgr(bgr), .slow_25(slow_25),
     .pbias_25(pbias_25), .vref_25(vref_25), .vppdisc_25(vppdisc_25),
     .pumpen_25(pumpen_25), .pump_in(pump_in), .vpp_int(vpp_int));
ml_vpp_vco Ivpp_vco ( .pbias_25(pbias_25), .slow_25(slow_25),
     .freq_25(freq_25[1:0]), .en_25(pumpen_25), .clk_25_0(clkin_0_25));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));
nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpp_int));
ml_vpp_pumpx3 Ivpp_pumpx3 ( .pump_in(pump_in), .pumpen_25(pumpen_25),
     .clkin_0_25(clkin_0_25));

endmodule
// Library - NVCM, Cell - UBGR_2511_065_FLAT, View - schematic
// LAST TIME SAVED: Apr  1 15:53:36 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module UBGR_2511_065_FLAT ( VREF, PDN, T0, T1, T2, T3, TEN, VDD25, VSS
     );
output  VREF;

input  PDN, T0, T1, T2, T3, TEN, VDD25, VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_bgr_top, View - schematic
// LAST TIME SAVED: Apr  7 14:19:14 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_bgr_top ( bgr_int, fsm_nvcmen_buf, fsm_trim_vbg_buf );
inout  bgr_int;

input  fsm_nvcmen_buf;

input [3:0]  fsm_trim_vbg_buf;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  bgr_trim_25;

wire  [0:3]  net48;

wire  [0:3]  net53;

wire  [0:3]  net44;



inv_25 I38 ( .IN(net58), .OUT(PDN), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
vddp_tiehigh I85 ( .vddp_tieh(TEN));
UBGR_2511_065_FLAT Ibgr ( .TEN(TEN), .VSS(gnd_), .VDD25(vddp_),
     .VREF(bgr_int), .T3(bgr_trim_25[3]), .T2(bgr_trim_25[2]),
     .T1(bgr_trim_25[1]), .T0(bgr_trim_25[0]), .PDN(PDN));
inv_hvt I88_3_ ( .A(fsm_trim_vbg_buf[3]), .Y(net48[0]));
inv_hvt I88_2_ ( .A(fsm_trim_vbg_buf[2]), .Y(net48[1]));
inv_hvt I88_1_ ( .A(fsm_trim_vbg_buf[1]), .Y(net48[2]));
inv_hvt I88_0_ ( .A(fsm_trim_vbg_buf[0]), .Y(net48[3]));
inv_hvt I319 ( .A(net50), .Y(net46));
inv_hvt I87_3_ ( .A(net48[0]), .Y(net44[0]));
inv_hvt I87_2_ ( .A(net48[1]), .Y(net44[1]));
inv_hvt I87_1_ ( .A(net48[2]), .Y(net44[2]));
inv_hvt I87_0_ ( .A(net48[3]), .Y(net44[3]));
inv_hvt I323 ( .A(fsm_nvcmen_buf), .Y(net50));
ml_ls_vdd2vdd25 I80_3_ ( .in(net44[0]), .sup(vddp_),
     .out_vddio_b(net53[0]), .out_vddio(bgr_trim_25[3]),
     .in_b(net48[0]));
ml_ls_vdd2vdd25 I80_2_ ( .in(net44[1]), .sup(vddp_),
     .out_vddio_b(net53[1]), .out_vddio(bgr_trim_25[2]),
     .in_b(net48[1]));
ml_ls_vdd2vdd25 I80_1_ ( .in(net44[2]), .sup(vddp_),
     .out_vddio_b(net53[2]), .out_vddio(bgr_trim_25[1]),
     .in_b(net48[2]));
ml_ls_vdd2vdd25 I80_0_ ( .in(net44[3]), .sup(vddp_),
     .out_vddio_b(net53[3]), .out_vddio(bgr_trim_25[0]),
     .in_b(net48[3]));
ml_ls_vdd2vdd25 I335 ( .in(net46), .sup(vddp_), .out_vddio_b(net58),
     .out_vddio(bgr_en_25), .in_b(net50));

endmodule
// Library - NVCM, Cell - ml_pump_vpxa_3.3v, View - schematic
// LAST TIME SAVED: Nov 14 11:45:03 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_pump_vpxa_3_3v ( out, clkin_25, en );
inout  out;

input  clkin_25, en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M10 ( .B(GND_), .D(s_0), .G(s_0), .S(s_1));
nch_na25  M11 ( .B(GND_), .D(s_1), .G(s_1), .S(s_2));
nch_na25  M12 ( .B(GND_), .D(s_2), .G(s_2), .S(out));
nch_na25  M22 ( .B(GND_), .D(net0115), .G(net0115), .S(s_0));
inv_25 I194 ( .IN(clkin_25), .OUT(net064), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(en), .OUT(net042), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I210 ( .IN(net076), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I219 ( .IN(net040), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I220 ( .IN(net034), .OUT(net046), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I221 ( .IN(net046), .OUT(net040), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I224 ( .IN(clkin_25), .OUT(net034), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I209 ( .IN(net064), .OUT(net076), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
pch_25  M0 ( .D(net0115), .B(vddp_), .G(net042), .S(vddp_));
nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));

endmodule
// Library - tsmcN65lo, Cell - nor2_25, View - schematic
// LAST TIME SAVED: Mar 29 20:24:25 2006
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module nor2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  PM1 ( .D(net15), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(net15));

endmodule
// Library - sbtlibn65lp, Cell - ml_dlatch_25, View - schematic
// LAST TIME SAVED: Feb 21 13:49:32 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_dlatch_25 ( Q_25, D_25, EN_25, R_25 );
output  Q_25;

input  D_25, EN_25, R_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M9 ( .D(net31), .B(vddp_), .G(EN_25), .S(vddp_));
pch_25  M7 ( .D(net39), .B(vddp_), .G(EN_B_25), .S(vddp_));
pch_25  M3 ( .D(net52), .B(vddp_), .G(D_25), .S(net39));
pch_25  M4 ( .D(net52), .B(vddp_), .G(Q_25), .S(net31));
nch_25  M8 ( .D(net52), .B(GND_), .G(D_25), .S(net48));
nch_25  M1 ( .D(net48), .B(GND_), .G(EN_25), .S(GND_));
nch_25  M5 ( .D(net40), .B(GND_), .G(EN_B_25), .S(GND_));
nch_25  M6 ( .D(net52), .B(GND_), .G(Q_25), .S(net40));
inv_25 I156 ( .IN(EN_25), .OUT(EN_B_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nor2_25 I161 ( .A(net52), .Y(Q_25), .Gb(GND_), .G(GND_), .Pb(vddp_),
     .P(vddp_), .B(R_25));

endmodule
// Library - misc, Cell - ml_osc_stage, View - schematic
// LAST TIME SAVED: Sep  8 19:15:04 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_osc_stage ( out, clkin, oscen_b, pbias, sel_trim );
output  out;

input  clkin, oscen_b, pbias;

input [3:0]  sel_trim;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_mux3_hvt Iml_mux3_hvt_bot ( .in1(loadbot_1), .in0(loadbot_0),
     .out(in_bot), .sel(sel_trim[3:0]), .in2(loadbot_2));
nor2_hvt I228 ( .A(clkin), .B(oscen_b), .Y(net403));
inv_hvt I229 ( .A(net403), .Y(net419));
nch_hvt  MN41 ( .D(loadbot_0), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN39 ( .D(loadbot_2), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN29 ( .D(out), .B(gnd_), .G(in_bot), .S(gnd_));
nch_hvt  MN42 ( .D(loadbot_1), .B(gnd_), .G(net419), .S(gnd_));
pch_hvt  M82 ( .D(vdd_), .B(vdd_), .G(loadbot_1), .S(vdd_));
pch_hvt  M83 ( .D(vdd_), .B(vdd_), .G(loadbot_0), .S(vdd_));
pch_hvt  M85 ( .D(vdd_), .B(vdd_), .G(loadbot_2), .S(vdd_));
pch_hvt  M84 ( .D(vdd_), .B(vdd_), .G(loadbot_1), .S(vdd_));
pch_hvt  M81 ( .D(vdd_), .B(vdd_), .G(loadbot_2), .S(vdd_));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(loadbot_0), .S(vdd_));
pch_hvt  MP73 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net456));
pch_hvt  MP30 ( .D(net452), .B(vdd_), .G(oscen_b), .S(vdd_));
pch_hvt  MP72 ( .D(net456), .B(vdd_), .G(sel_trim[2]), .S(net452));
pch_hvt  MP33 ( .D(out), .B(vdd_), .G(in_bot), .S(vdd_));
pch_hvt  MP74 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net452));

endmodule
// Library - NVCM, Cell - ml_pump_clk_reg, View - schematic
// LAST TIME SAVED: Feb 13 16:09:37 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_pump_clk_reg ( clk_out_25, clk_in_25, pump_chrg_25,
     pump_on_25 );
output  clk_out_25;

input  clk_in_25, pump_chrg_25, pump_on_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



exor2_25 I85 ( .A(clk_in_25), .Y(net020), .B(clk_out_25));
nand2_25 I78 ( .G(GND_), .Pb(vddp_), .A(pump_chrg_25), .Y(clk_freeze),
     .P(vddp_), .B(pump_on_25), .Gb(GND_));
inv_25 I72 ( .IN(net020), .OUT(clk_equal), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(vddp_tieh), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
vddp_tiehigh I117 ( .vddp_tieh(vddp_tieh));
ml_dlatch_25 I63 ( .D_25(clk_in_25), .EN_25(clk_go), .R_25(net34),
     .Q_25(clk_out_25));
ml_dlatch_25 I64 ( .D_25(vddp_tieh), .EN_25(clk_equal),
     .R_25(clk_freeze), .Q_25(clk_go));

endmodule
// Library - NVCM, Cell - ml_pump_vpxa_x2, View - schematic
// LAST TIME SAVED: Nov 14 11:48:00 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_pump_vpxa_x2 ( vpxa_int, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, pumpen, pumpen_25, vpxa_clk_25, vpxa_clk_b_25 );
inout  vpxa_int;

input  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25, pumpen,
     pumpen_25, vpxa_clk_25, vpxa_clk_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_pump_vpxa_3_3v Ivpxa_pump_0 ( .en(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_0_25));
ml_pump_vpxa_3_3v Ivpxa_pump_2 ( .en(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_2_25));
ml_pump_vpxa_3_3v Ivpxa_pump_1 ( .en(pumpen_25), .clkin_25(clkin_1_25),
     .out(vpxa_int));
ml_pump_clk_reg Iclk_reg_0 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_0_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_0_25));
ml_pump_clk_reg Iclk_reg_2 ( .clk_in_25(vpxa_clk_b_25),
     .pump_chrg_25(pump_chrg_2_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_2_25));
ml_pump_clk_reg Iclk_reg_1 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_1_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_1_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_osc, View - schematic
// LAST TIME SAVED: Mar 14 15:11:03 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpxa_osc ( vpxa_clk_25, bgr, freq_25, pumpen_25 );
output  vpxa_clk_25;

inout  bgr;

input  pumpen_25;

input [1:0]  freq_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  freq_buf_b_25;



inv_25 I38 ( .IN(pumpen_25), .OUT(pbiasen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I195 ( .IN(freq_25[0]), .OUT(freq_buf_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
pch_25  M9 ( .D(net64), .B(vddp_), .G(pbiasen_b_25), .S(vddp_));
pch_25  M4_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
pch_25  M4_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
pch_25  M0 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
nch_25  M8 ( .D(pbias_25), .B(GND_), .G(pbiasen_b_25), .S(gnd_));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net74));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net83), .PLUS(net74), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net83), .BULK(GND_));
ml_vpp_vco Ivpx_vpp_vco ( .pbias_25(pbias_25), .slow_25(net86),
     .freq_25({freq_25[1], freq_buf_b_25[0]}), .en_25(pumpen_25),
     .clk_25_0(vpxa_clk_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_ctrl, View - schematic
// LAST TIME SAVED: Oct 28 15:47:22 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpxa_ctrl ( pumpen, pumpen_25, vpxa_2_vdd, fsm_pumpen,
     fsm_tm_xforce, fsm_tm_xvpxaint );
output  pumpen, pumpen_25, vpxa_2_vdd;

input  fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I73 ( .A(fsm_tm_xvpxaint), .B(fsm_tm_xforce), .Y(net042));
inv_25 I38 ( .IN(net045), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I173 ( .in(net049), .sup(vddp_), .out_vddio_b(net045),
     .out_vddio(net046), .in_b(net075));
nor2_hvt I72 ( .A(vpxa_off), .B(net065), .Y(net049));
nor2_hvt I69 ( .A(vpxa_2_vdd), .B(vpxa_2_vdd), .Y(net043));
inv_hvt I75 ( .A(net049), .Y(net056));
inv_hvt I76 ( .A(net056), .Y(pumpen));
inv_hvt I110 ( .A(net049), .Y(net075));
inv_hvt I74 ( .A(net042), .Y(net065));
inv_hvt I131 ( .A(fsm_pumpen), .Y(vpxa_2_vdd));
inv_hvt I70 ( .A(net043), .Y(vpxa_off));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff_25, View - schematic
// LAST TIME SAVED: Feb 11 11:37:05 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_dff_25 ( Q_25, Q_B_25, CLK_25, D_25, R_25 );
output  Q_25, Q_B_25;

input  CLK_25, D_25, R_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I87 ( .IN(net044), .OUT(net038), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I72 ( .IN(CLK_25), .OUT(net044), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I90 ( .IN(Q_25), .OUT(Q_B_25), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
ml_dlatch_25 Ilatch2 ( .D_25(net053), .EN_25(net038), .R_25(R_25),
     .Q_25(Q_25));
ml_dlatch_25 Ilatch1 ( .Q_25(net053), .EN_25(net044), .D_25(D_25),
     .R_25(R_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_n, View - schematic
// LAST TIME SAVED: Feb  5 15:08:44 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp_n ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M0 ( .D(out_div), .B(vddp_), .G(out_ref), .S(vddp_));
pch_25  M4 ( .D(out_ref), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M5 ( .D(out_div), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M7 ( .D(out_ref), .B(vddp_), .G(out_ref), .S(vddp_));
nch_25  M1 ( .D(out_div), .B(GND_), .G(in_div), .S(net049));
nch_25  M2 ( .D(out_ref), .B(GND_), .G(in_ref), .S(net049));
nch_25  M6_1_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_top_n, View - schematic
// LAST TIME SAVED: Feb 21 13:55:00 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp_top_n ( pump_chrg_25, in_div, in_ref, sa_bias,
     saen_25 );
output  pump_chrg_25;

input  in_div, in_ref, sa_bias, saen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_25 I103 ( .G(gnd_), .Pb(vddp_), .A(saen_25), .Y(chrg_b_25),
     .P(vddp_), .B(net27), .Gb(gnd_));
nch_25  M6_1_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
inv_25 I102 ( .IN(chrg_b_25), .OUT(pump_chrg_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I104 ( .IN(out_div2), .OUT(net27), .P(vddp_), .Pb(vddp_),
     .G(net087), .Gb(gnd_));
ml_core_sa_comp_n Icore_sa_comp_n0 ( .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp_n Iml_core_sa_comp_n1 ( .out_div(out_div2),
     .out_ref(out_ref2), .in_div(in_div2), .in_ref(in_ref2),
     .sa_bias(sa_bias), .saen_25(saen_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_reg, View - schematic
// LAST TIME SAVED: May  3 13:50:36 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpxa_reg ( freq_25, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, vpxa_int, bgr, fsm_vrdwl, pumpen, vpxa_clk_25 );
output  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25;

inout  vpxa_int;

input  bgr, pumpen, vpxa_clk_25;

output [1:0]  freq_25;

input [2:0]  fsm_vrdwl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  freq_in_25;

wire  [0:2]  vrdwl_vpxa;

wire  [0:2]  vrdwl_b_vpxa;



nand2_25 I145 ( .G(GND_), .Pb(vddp_), .A(net0171), .Y(freq_in_25[0]),
     .P(vddp_), .B(net0179), .Gb(GND_));
nand2_25 I158 ( .G(GND_), .Pb(vddp_), .A(net0179), .Y(freq_in_25[1]),
     .P(vddp_), .B(net0163), .Gb(GND_));
nand3_25 I44 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0179),
     .C(pump_chrg_0_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I149 ( .B(pump_chrg_1_b_25), .A(pump_chrg_2_25), .Y(net0171),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I159 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0163),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
ml_dff_25 I125 ( .Q_B_25(net0187), .R_25(saen_b_25),
     .D_25(freq_in_25[1]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[1]));
ml_dff_25 I126 ( .Q_B_25(net0192), .R_25(saen_b_25),
     .D_25(freq_in_25[0]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[0]));
inv_hvt I85 ( .A(net171), .Y(net175));
inv_hvt I183 ( .A(fsm_vrdwl[2]), .Y(net171));
inv_hvt I83 ( .A(pumpen), .Y(net143));
inv_hvt I82 ( .A(net143), .Y(net145));
inv_hvt I184 ( .A(fsm_vrdwl[1]), .Y(net176));
inv_hvt I187 ( .A(fsm_vrdwl[0]), .Y(net181));
inv_hvt I186 ( .A(net181), .Y(net185));
inv_hvt I185 ( .A(net176), .Y(net180));
inv_25 I155 ( .IN(pump_chrg_0_25), .OUT(pump_chrg_0_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
inv_25 I63 ( .IN(net169), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(net168), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I154 ( .IN(pump_chrg_1_25), .OUT(pump_chrg_1_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_ls_vdd2vdd25 I191 ( .in(saen_25), .sup(vpxa_int),
     .out_vddio_b(saen_b_vpxa), .out_vddio(net0210), .in_b(saen_b_25));
ml_ls_vdd2vdd25 I335 ( .in(net145), .sup(vddp_), .out_vddio_b(net168),
     .out_vddio(net169), .in_b(net143));
ml_ls_vdd2vdd25 I87 ( .in(net171), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[2]), .out_vddio(vrdwl_b_vpxa[2]),
     .in_b(net175));
ml_ls_vdd2vdd25 I98 ( .in(net176), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[1]), .out_vddio(vrdwl_b_vpxa[1]),
     .in_b(net180));
ml_ls_vdd2vdd25 I99 ( .in(net181), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[0]), .out_vddio(vrdwl_b_vpxa[0]),
     .in_b(net185));
ml_core_sa_comp_top_n Icore_sa_comp_top_n2 (
     .pump_chrg_25(pump_chrg_2_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_2));
ml_core_sa_comp_top_n core_sa_comp_top_n0 (
     .pump_chrg_25(pump_chrg_0_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_0));
ml_core_sa_comp_top_n Icore_sa_comp_top_n1 (
     .pump_chrg_25(pump_chrg_1_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_1));
rppolywo_m  R29 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R28 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R27 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(in_div_0), .PLUS(net202), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net232), .PLUS(net223), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(net270), .PLUS(net226), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net226), .PLUS(net229), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(sa_bias), .PLUS(net232), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net202), .PLUS(net237), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(net237), .PLUS(net270), .BULK(GND_));
rppolywo_m  R30 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(gnd_), .PLUS(in_div_2), .BULK(GND_));
rppolywo_m  R31 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
pch_25  M3 ( .D(net229), .B(vpxa_int), .G(saen_b_vpxa), .S(vpxa_int));
pch_25  M11_1_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M11_0_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M15 ( .D(net237), .B(vpxa_int), .G(vrdwl_vpxa[0]), .S(net270));
pch_25  M37 ( .D(net226), .B(vpxa_int), .G(vrdwl_vpxa[2]), .S(net229));
pch_25  M1 ( .D(net223), .B(vddp_), .G(saen_b_25), .S(vddp_));
pch_25  M14 ( .D(net270), .B(vpxa_int), .G(vrdwl_vpxa[1]), .S(net226));
pch_25  M8_1_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
pch_25  M8_0_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
nch_25  M2 ( .D(sa_bias), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M32 ( .D(net229), .B(GND_), .G(vrdwl_b_vpxa[2]), .S(net226));
nch_25  M0_3_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_2_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_1_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_0_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M9 ( .D(net270), .B(GND_), .G(vrdwl_b_vpxa[0]), .S(net237));
nch_25  M7 ( .D(net226), .B(GND_), .G(vrdwl_b_vpxa[1]), .S(net270));

endmodule
// Library - NVCM, Cell - ml_hv2vdd_sw, View - schematic
// LAST TIME SAVED: Apr  8 14:27:39 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv2vdd_sw ( out_hv, hv2vdd, vddp_tieh );
inout  out_hv;

input  hv2vdd, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M1 ( .D(net27), .B(GND_), .G(vddp_tieh), .S(out_hv));
nch_na25  M2 ( .D(vdd_), .B(GND_), .G(hv2vdd_25), .S(net27));
inv_25 I62 ( .IN(net40), .OUT(hv2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net40),
     .out_vddio(net37), .in_b(net46));
inv_hvt I65 ( .A(hv2vdd), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));

endmodule
// Library - NVCM, Cell - ml_vpxa_top, View - schematic
// LAST TIME SAVED: Sep  4 16:21:42 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_vpxa_top ( vpxa_int, bgr, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint, fsm_vrdwl );
inout  vpxa_int;

input  bgr, fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;

input [2:0]  fsm_vrdwl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  freq_25;



nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpxa_int));
ml_pump_vpxa_x2 Ipump_vpxa_x3 ( .pumpen(pumpen),
     .vpxa_clk_b_25(vpxa_clk_b_25), .vpxa_clk_25(vpxa_clk_25),
     .pumpen_25(pumpen_25), .pump_chrg_2_25(pump_chrg_2_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_0_25(pump_chrg_0_25),
     .vpxa_int(vpxa_int));
inv_25 I73 ( .IN(vpxa_clk_25), .OUT(vpxa_clk_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_vpxa_osc Ivpxa_osc ( .freq_25(freq_25[1:0]), .bgr(bgr),
     .pumpen_25(pumpen_25), .vpxa_clk_25(vpxa_clk_25));
ml_vpxa_ctrl Ivpxa_ctrl ( .fsm_pumpen(fsm_pumpen), .pumpen(pumpen),
     .pumpen_25(pumpen_25), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .vpxa_2_vdd(vpxa_2_vdd));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));
ml_vpxa_reg Ivpxa_reg ( .pump_chrg_0_25(pump_chrg_0_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_2_25(pump_chrg_2_25),
     .freq_25(freq_25[1:0]), .vpxa_clk_25(vpxa_clk_25),
     .pumpen(pumpen), .fsm_vrdwl(fsm_vrdwl[2:0]), .bgr(bgr),
     .vpxa_int(vpxa_int));
ml_hv2vdd_sw Ivpxa_2vdd_sw ( .vddp_tieh(vddp_tieh),
     .hv2vdd(vpxa_2_vdd), .out_hv(vpxa_int));

endmodule
// Library - misc, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:59 2007
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_mux2_hvt ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - NVCM, Cell - ml_hv_invx3_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:19:36 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv_invx3_enhance ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh
     );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_switch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 14:46:53 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_lshv_6v_switch_enhance ( out_b_hv, out_hv, in_hv, sel_25,
     sel_b_25, vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M11 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv_hotsw_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:16:13 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw_enhance ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3_enhance Ihv_invx3 ( .vddp_tieh(vddp_tieh),
     .out_b_hv(out_b_hv), .sel_25(sel_25), .in_hv(in_hv),
     .sel_hv(sel_hv));
ml_lshv_6v_switch_enhance Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM, Cell - ml_hv_hotswitch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:15:29 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv_hotswitch_enhance ( hv_in_hv, hv_out_hv, selhv_25,
     vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M7 ( .D(net12), .B(GND_), .G(selhv_25), .S(net15));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
pch_25  M0 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_pump_a_clkdly, View - schematic
// LAST TIME SAVED: Feb 11 09:24:13 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_pump_a_clkdly ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(net66), .S(vdd_));
pch_hvt  M0 ( .D(vdd_), .B(vdd_), .G(net62), .S(vdd_));
inv_hvt I206 ( .A(in), .Y(net66));
inv_hvt I204 ( .A(net64), .Y(net62));
inv_hvt I205 ( .A(net66), .Y(net64));
inv_hvt I207 ( .A(net70), .Y(out));
inv_hvt I208 ( .A(net62), .Y(net70));

endmodule
// Library - NVCM, Cell - ml_hvmux_top_ctrl, View - schematic
// LAST TIME SAVED: May  2 18:30:47 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hvmux_top_ctrl ( bgrext_en, bgrint_en, en_vblinhi,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp, fsm_lshven,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint, fsm_wgnden,
     fsm_wpen, tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );
output  bgrext_en, bgrint_en, en_vblinhi, ngate_vddp, ngate_vpxa,
     sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint,
     vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint, vpxaint_ext,
     vtmode, ysup25_2vdd, ysup25_2vddp;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_testdec,
     tm_wleqbl, vpint_en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



mux2_hvt I260 ( .in1(fsm_wgnden), .in0(fsm_wpen), .out(net0217),
     .sel(pgmpulse_b));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
anor21_hvt I245 ( .A(net0189), .B(net0193), .Y(vppint_ext),
     .C(net0188));
anor21_hvt I109 ( .A(net0201), .B(net0199), .Y(vpxa_ext), .C(net0188));
nand3_hvt I248 ( .Y(net0189), .B(vpint_en), .C(fsm_tm_xvppint),
     .A(fsm_tm_xforce));
nand3_hvt I246 ( .Y(net0201), .B(vddp_rd_b), .C(fsm_tm_xvpxa),
     .A(fsm_tm_xforce));
nand3_hvt I247 ( .Y(net0193), .B(pmprd), .C(pmprd),
     .A(fsm_tm_xvppint));
nand3_hvt I35 ( .C(fsm_lshven), .A(fsm_pgm), .Y(pgmpulse_b),
     .B(net0327));
nand3_hvt I205 ( .Y(net0213), .B(net0321), .C(pgmpulse_b),
     .A(net0321));
nand3_hvt I240 ( .C(pmprd), .A(fsm_tm_xvpxa), .Y(net0199), .B(pmprd));
nor2_hvt I213 ( .A(net0324), .B(fsm_nvcmen_b), .Y(net0251));
nor2_hvt I224 ( .A(vddp_rd_b), .B(net0258), .Y(vpxa_vppd));
nor2_hvt I214 ( .A(net0251), .B(net0266), .Y(sbhvsup_vppint));
nor2_hvt I215 ( .A(net0264), .B(net0311), .Y(sbhvsup_vddp));
nor2_hvt I183 ( .A(net87), .B(net73), .Y(ysup25_2vddp));
nor2_hvt I14 ( .A(net75), .B(net93), .Y(ysup25_2vdd));
nor2_hvt I207 ( .A(net0325), .B(net0260), .Y(sb25sup_vddp));
nor2_hvt I206 ( .A(net0268), .B(net0213), .Y(sb25sup_vpxa));
nor2_hvt I185 ( .A(gnd_tiel), .B(gnd_tiel), .Y(net0240));
nor2_hvt I223 ( .B(net0240), .Y(vddp_rd), .A(net0349));
nor2_hvt I195 ( .A(net0272), .B(rd_vddp), .Y(ngate_vpxa));
nor2_hvt I196 ( .A(net0331), .B(net0270), .Y(ngate_vddp));
nor2_hvt I225 ( .A(net0256), .B(vddp_rd), .Y(vpxa_vpxaint));
ml_pump_a_clkdly I219 ( .in(ysup25_2vddp_b), .out(net75));
ml_pump_a_clkdly I227 ( .in(net0297), .out(net0256));
ml_pump_a_clkdly I226 ( .in(net0319), .out(net0258));
ml_pump_a_clkdly I209 ( .in(net0323), .out(net0260));
ml_pump_a_clkdly I184 ( .in(ysup25_2vdd_b), .out(net73));
ml_pump_a_clkdly I217 ( .in(net0313), .out(net0264));
ml_pump_a_clkdly I216 ( .in(net0309), .out(net0266));
ml_pump_a_clkdly I208 ( .in(net0329), .out(net0268));
ml_pump_a_clkdly I198 ( .in(net0339), .out(net0270));
ml_pump_a_clkdly I197 ( .in(net0335), .out(net0272));
nand2_hvt I254 ( .A(bgrext_en), .Y(bgrint_en), .B(fsm_tm_xforce));
nand2_hvt I104 ( .A(fsm_nvcmen), .Y(net77), .B(tm_wleqbl));
nand2_hvt I179 ( .A(fsm_nvcmen), .Y(net80), .B(net0217));
nand2_hvt I252 ( .A(fsm_nvcmen_buf), .Y(net0277), .B(fsm_tm_xvbg));
nand2_hvt I234 ( .A(fsm_pumpen), .Y(net0286), .B(fsm_tm_xvpxaint));
inv_hvt I259 ( .A(pgmpulse_b), .Y(net0324));
inv_hvt I229 ( .A(vpxa_vppd), .Y(net0297));
inv_hvt I250 ( .A(fsm_pumpen), .Y(net0188));
inv_hvt I182 ( .A(ysup25_2vdd), .Y(ysup25_2vdd_b));
inv_hvt I230 ( .A(vddp_rd), .Y(vddp_rd_b));
inv_hvt I249 ( .A(pgmpulse_b), .Y(pgmpulse));
inv_hvt I131 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I178 ( .A(net77), .Y(vtmode));
inv_hvt I180 ( .A(net80), .Y(net93));
inv_hvt I253 ( .A(net0277), .Y(bgrext_en));
inv_hvt I218 ( .A(sbhvsup_vddp), .Y(net0309));
inv_hvt I221 ( .A(net0251), .Y(net0311));
inv_hvt I220 ( .A(sbhvsup_vppint), .Y(net0313));
inv_hvt I134 ( .A(net93), .Y(net87));
inv_hvt I181 ( .A(ysup25_2vddp), .Y(ysup25_2vddp_b));
inv_hvt I228 ( .A(vpxa_vpxaint), .Y(net0319));
inv_hvt I204 ( .A(rd_vddp), .Y(net0321));
inv_hvt I212 ( .A(sb25sup_vpxa), .Y(net0323));
inv_hvt I210 ( .A(net0213), .Y(net0325));
inv_hvt I202 ( .A(fsm_pgmvfy), .Y(net0327));
inv_hvt I211 ( .A(sb25sup_vddp), .Y(net0329));
inv_hvt I199 ( .A(rd_vddp), .Y(net0331));
inv_hvt I236 ( .A(fsm_tm_xforce), .Y(pmprd));
inv_hvt I200 ( .A(ngate_vddp), .Y(net0335));
inv_hvt I235 ( .A(net0286), .Y(vpxaint_ext));
inv_hvt I201 ( .A(ngate_vpxa), .Y(net0339));
inv_hvt I233 ( .A(fsm_nvcmen_b), .Y(fsm_nvcmen_buf));
nor3_hvt I105 ( .B(tm_testdec), .Y(en_vblinhi), .A(fsm_nvcmen_b),
     .C(tm_allbl_l));
nor3_hvt I186 ( .C(fsm_rd), .A(fsm_tm_rd_mode), .B(fsm_pgmvfy),
     .Y(net0349));
nor3_hvt I187 ( .B(net0240), .Y(rd_vddp), .A(net0349),
     .C(fsm_nvcmen_b));

endmodule
// Library - NVCM, Cell - ml_hvmux_ls25, View - schematic
// LAST TIME SAVED: Feb 15 14:23:11 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hvmux_ls25 ( bgrext_en_25, bgrint_en_25, ngate_vddp_25,
     ngate_vpxa_25, sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25, bgrext_en, bgrint_en,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp );
output  bgrext_en_25, bgrint_en_25, ngate_vddp_25, ngate_vpxa_25,
     sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25;

input  bgrext_en, bgrint_en, ngate_vddp, ngate_vpxa, sb25sup_vddp,
     sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint, vppint_ext, vpxa_ext,
     vpxa_vppd, vpxa_vpxaint, vpxaint_ext, vtmode, ysup25_2vdd,
     ysup25_2vddp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I317 ( .A(net054), .Y(net052));
inv_hvt I314 ( .A(vpxa_vppd), .Y(net054));
inv_hvt I327 ( .A(net066), .Y(net056));
inv_hvt I329 ( .A(bgrint_en), .Y(net058));
inv_hvt I321 ( .A(vpxaint_ext), .Y(net060));
inv_hvt I320 ( .A(net060), .Y(net062));
inv_hvt I325 ( .A(net082), .Y(net064));
inv_hvt I326 ( .A(vppint_ext), .Y(net066));
inv_hvt I312 ( .A(bgrext_en), .Y(net068));
inv_hvt I313 ( .A(net068), .Y(net070));
inv_hvt I328 ( .A(net058), .Y(net0487));
inv_hvt I239 ( .A(sb25sup_vpxa), .Y(net0486));
inv_hvt I319 ( .A(net0112), .Y(net0488));
inv_hvt I240 ( .A(net0486), .Y(net080));
inv_hvt I324 ( .A(vpxa_ext), .Y(net082));
inv_hvt I206 ( .A(vtmode), .Y(net084));
inv_hvt I213 ( .A(ysup25_2vdd), .Y(net086));
inv_hvt I214 ( .A(net086), .Y(net088));
inv_hvt I205 ( .A(net084), .Y(net090));
inv_hvt I216 ( .A(net088), .Y(net092));
inv_hvt I110 ( .A(net072), .Y(net074));
inv_hvt I227 ( .A(net098), .Y(net096));
inv_hvt I228 ( .A(ngate_vddp), .Y(net098));
inv_hvt I217 ( .A(net092), .Y(ysup25_2vdd_buf));
inv_hvt I190 ( .A(ysup25_2vddp), .Y(net072));
inv_hvt I219 ( .A(ngate_vpxa), .Y(net0104));
inv_hvt I220 ( .A(net0104), .Y(net0106));
inv_hvt I232 ( .A(sb25sup_vddp), .Y(net0108));
inv_hvt I231 ( .A(net0108), .Y(net0110));
inv_hvt I323 ( .A(vpxa_vpxaint), .Y(net0112));
inv_hvt I256 ( .A(net0116), .Y(net0114));
inv_hvt I257 ( .A(sbhvsup_vddp), .Y(net0116));
inv_hvt I258 ( .A(net0120), .Y(net0118));
inv_hvt I259 ( .A(sbhvsup_vppint), .Y(net0120));
ml_ls_vdd2vdd25 I336 ( .in(net064), .sup(vddp_), .out_vddio_b(net0123),
     .out_vddio(net0207), .in_b(net082));
ml_ls_vdd2vdd25 I337 ( .in(net056), .sup(vddp_), .out_vddio_b(net0128),
     .out_vddio(net0208), .in_b(net066));
ml_ls_vdd2vdd25 I338 ( .in(net052), .sup(vddp_), .out_vddio_b(net0133),
     .out_vddio(net0211), .in_b(net054));
ml_ls_vdd2vdd25 I339 ( .in(net0487), .sup(vddp_),
     .out_vddio_b(net0138), .out_vddio(net0209), .in_b(net058));
ml_ls_vdd2vdd25 I332 ( .in(net070), .sup(vddp_), .out_vddio_b(net0148),
     .out_vddio(net0149), .in_b(net068));
ml_ls_vdd2vdd25 I238 ( .in(net080), .sup(vddp_), .out_vddio_b(net0153),
     .out_vddio(net0154), .in_b(net0486));
ml_ls_vdd2vdd25 I334 ( .in(net062), .sup(vddp_), .out_vddio_b(net0158),
     .out_vddio(net0214), .in_b(net060));
ml_ls_vdd2vdd25 I335 ( .in(net0488), .sup(vddp_),
     .out_vddio_b(net0163), .out_vddio(net0206), .in_b(net0112));
ml_ls_vdd2vdd25 I212 ( .in(net088), .sup(vddp_), .out_vddio_b(net0168),
     .out_vddio(net0169), .in_b(net086));
ml_ls_vdd2vdd25 I226 ( .in(net096), .sup(vddp_), .out_vddio_b(net0173),
     .out_vddio(net0174), .in_b(net098));
ml_ls_vdd2vdd25 I203 ( .in(net072), .sup(vddp_), .out_vddio_b(net077),
     .out_vddio(net078), .in_b(net074));
ml_ls_vdd2vdd25 I221 ( .in(net0106), .sup(vddp_),
     .out_vddio_b(net0183), .out_vddio(net0184), .in_b(net0104));
ml_ls_vdd2vdd25 I233 ( .in(net0110), .sup(vddp_),
     .out_vddio_b(net0188), .out_vddio(net0219), .in_b(net0108));
ml_ls_vdd2vdd25 I207 ( .in(net090), .sup(vddp_), .out_vddio_b(net0193),
     .out_vddio(net0194), .in_b(net084));
ml_ls_vdd2vdd25 I260 ( .in(net0114), .sup(vddp_),
     .out_vddio_b(net0198), .out_vddio(net0220), .in_b(net0116));
ml_ls_vdd2vdd25 I261 ( .in(net0118), .sup(vddp_),
     .out_vddio_b(net0203), .out_vddio(net0204), .in_b(net0120));
inv_25 I390 ( .IN(net0148), .OUT(bgrext_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I384 ( .IN(net0163), .OUT(vpxa_vpxaint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I386 ( .IN(net0133), .OUT(vpxa_vppd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I388 ( .IN(net0123), .OUT(vpxa_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I376 ( .IN(net0168), .OUT(ysup25_2vdd_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I387 ( .IN(net0158), .OUT(vpxaint_ext_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I389 ( .IN(net0128), .OUT(vppint_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I362 ( .IN(net077), .OUT(ysup25_2vddp_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I383 ( .IN(net0203), .OUT(sbhvsup_vppint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I379 ( .IN(net0183), .OUT(ngate_vpxa_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I377 ( .IN(net0193), .OUT(vtmode_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I378 ( .IN(net0173), .OUT(ngate_vddp_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I381 ( .IN(net0153), .OUT(sb25sup_vpxa_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I382 ( .IN(net0198), .OUT(sbhvsup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I380 ( .IN(net0188), .OUT(sb25sup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I391 ( .IN(net0138), .OUT(bgrint_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_bgrxcvr, View - schematic
// LAST TIME SAVED: Apr  8 10:30:41 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hvmux_bgrxcvr ( bgr, bgr_int, bgrint_en_25, vpp,
     bgrext_en_25, vddp_tieh );
inout  bgr, bgr_int, bgrint_en_25, vpp;

input  bgrext_en_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M0 ( .D(bgr), .B(GND_), .G(bgrint_en_25), .S(bgr_int));
nch_25  M2 ( .D(vpp), .B(GND_), .G(vddp_tieh), .S(net53));
nch_25  M3 ( .D(net53), .B(GND_), .G(bgrext_en_25), .S(bgr));

endmodule
// Library - NVCM, Cell - ml_hv_hotswitch, View - schematic
// LAST TIME SAVED: Jan 25 09:27:57 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hv_hotswitch ( hv_in_hv, hv_out_hv, selhv_25, vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M7 ( .D(net12), .B(GND_), .G(selhv_25), .S(net15));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
pch_25  M0 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_hotswitch, View - schematic
// LAST TIME SAVED: Jan 26 19:35:53 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch ( hvin_a_hv, hvin_b_hv, out_hv, sel_hv_a_25,
     sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - misc, Cell - ml_osc_logic, View - schematic
// LAST TIME SAVED: Aug 28 14:12:11 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_osc_logic ( sel_trim, clkin, smc_osc_fsel, smc_oscen );

input  clkin, smc_oscen;

output [3:0]  sel_trim;

input [1:0]  smc_osc_fsel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:2]  in_sel;



tiehi I281 ( .tiehi(net058));
ml_dff I174 ( .R(reset_ff), .D(net050), .CLK(clkin_buf_b), .QN(net150),
     .Q(net172));
ml_dff I238 ( .R(reset_ff), .D(net050), .CLK(clkin_buf), .QN(net154),
     .Q(net177));
ml_dff I244 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf),
     .QN(net155), .Q(net182));
ml_dff I245 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf_b),
     .QN(net153), .Q(net187));
ml_dff I242 ( .R(reset_ff), .D(net048), .CLK(clkin_buf_b), .QN(net191),
     .Q(net192));
ml_dff I243 ( .R(reset_ff), .D(net048), .CLK(clkin_buf), .QN(net152),
     .Q(net197));
ml_mux2_hvt I279 ( .in1(net182), .in0(net187), .out(sel_trim[0]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I277 ( .in1(net057), .in0(net061), .out(sel_trim[2]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I278 ( .in1(net052), .in0(net054), .out(sel_trim[1]),
     .sel(clkin_buf_delay));
nor2_hvt I256 ( .A(smc_osc_fsel[1]), .B(smc_osc_fsel[0]),
     .Y(in_sel[2]));
inv_hvt I263 ( .A(clkin_buf), .Y(net065));
inv_hvt I252 ( .A(smc_oscen), .Y(reset_ff));
inv_hvt I264 ( .A(net065), .Y(net063));
inv_hvt I253 ( .A(clkin_buf_b), .Y(clkin_buf));
inv_hvt I254 ( .A(clkin), .Y(clkin_buf_b));
inv_hvt I255 ( .A(smc_osc_fsel[1]), .Y(in_sel[1]));
inv_hvt I266 ( .A(net063), .Y(net059));
inv_hvt I265 ( .A(net059), .Y(net0143));
inv_hvt I274 ( .A(net177), .Y(net057));
inv_hvt I273 ( .A(net172), .Y(net061));
inv_hvt I275 ( .A(net192), .Y(net054));
inv_hvt I276 ( .A(net197), .Y(net052));
inv_hvt I261 ( .A(in_sel[2]), .Y(net050));
inv_hvt I267 ( .A(net0143), .Y(net0144));
inv_hvt I262 ( .A(in_sel[1]), .Y(net048));
inv_hvt I268 ( .A(net0144), .Y(net0145));
inv_hvt I269 ( .A(net0142), .Y(clkin_buf_delay));
inv_hvt I270 ( .A(net0145), .Y(net0142));
inv_hvt I176 ( .A(net058), .Y(sel_trim[3]));

endmodule
// Library - NVCM, Cell - ml_ysup_25_switch, View - schematic
// LAST TIME SAVED: Apr  8 10:33:54 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_ysup_25_switch ( vdd, vddp, ysup_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25 );
inout  vdd, vddp, ysup_25;

input  ysup25_2vdd_25, ysup25_2vdd_buf, ysup25_2vddp_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd), .B(GND_), .G(ysup25_2vdd_25), .S(ysup_25));
pch_25  M5 ( .D(net73), .B(vddp), .G(ysup25_2vddp_b_25), .S(vddp));
pch_25  M0 ( .D(ysup_25), .B(ysup_25), .G(ysup25_2vdd_buf), .S(net73));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_vblinhi, View - schematic
// LAST TIME SAVED: Feb  1 08:51:27 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_vblinhi ( vblinhi, vpxa, en_vblinhi, vtmode,
     vtmode_25 );
inout  vblinhi, vpxa;

input  en_vblinhi, vtmode, vtmode_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I191 ( .A(en_vblinhi), .B(vtmode_buf), .Y(ngate_inhi_lv));
nand2_hvt I104 ( .A(net063), .Y(pgate_inhi_lv), .B(en_vblinhi));
inv_hvt I110 ( .A(net063), .Y(vtmode_buf));
inv_hvt I190 ( .A(vtmode), .Y(net063));
nch_25  M9 ( .D(net062), .B(GND_), .G(net062), .S(vblinhi));
nch_25  M8 ( .D(vpxa), .B(GND_), .G(vtmode_25), .S(net062));
pch_hvt  M7_1_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_0_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
nch_hvt  M0_1_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_0_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_top, View - schematic
// LAST TIME SAVED: May  2 18:49:30 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hvmux_top ( bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi, vpp, vpp_int, vpxa, vpxa_int, ysup_25, fsm_lshven,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint, fsm_wgnden,
     fsm_wpen, tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );
inout  bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi, vpp,
     vpp_int, vpxa, vpxa_int, ysup_25;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_testdec,
     tm_wleqbl, vpint_en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ixcvr_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(vppint_ext_25), .hv_in_hv(vpp_int), .hv_out_hv(vpp));
ml_hvmux_top_ctrl Ihvmux_top_ctrl ( .vpint_en(vpint_en),
     .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl),
     .tm_testdec(tm_testdec), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvpxa(fsm_tm_xvpxa), .fsm_tm_xvppint(fsm_tm_xvppint),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .ysup25_2vddp(ysup25_2vddp), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vppint(sbhvsup_vppint), .sbhvsup_vddp(sbhvsup_vddp),
     .sb25sup_vpxa(sb25sup_vpxa), .sb25sup_vddp(sb25sup_vddp),
     .ngate_vpxa(ngate_vpxa), .ngate_vddp(ngate_vddp),
     .en_vblinhi(en_vblinhi), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en));
ml_hvmux_ls25 Ihvmux_ls25 ( .ysup25_2vddp(ysup25_2vddp),
     .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vppint_25(sbhvsup_vppint_25), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en), .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vtmode_25(vtmode_25),
     .vpxaint_ext_25(vpxaint_ext_25),
     .vpxa_vpxaint_25(vpxa_vpxaint_25), .vpxa_vppd_25(vpxa_vppd_25),
     .vpxa_ext_25(net164), .vppint_ext_25(vppint_ext_25),
     .sbhvsup_vddp_25(sbhvsup_vddp_25),
     .sb25sup_vpxa_25(sb25sup_vpxa_25),
     .sb25sup_vddp_25(sb25sup_vddp_25), .ngate_vpxa_25(ngate_vpxa_25),
     .ngate_vddp_25(ngate_vddp_25), .bgrint_en_25(bgrint_en_25),
     .bgrext_en_25(bgrext_en_25));
ml_hvmux_bgrxcvr Ixcvr_bgr ( .vddp_tieh(vddp_tieh),
     .bgrext_en_25(bgrext_en_25), .vpp(vpp),
     .bgrint_en_25(bgrint_en_25), .bgr_int(bgr_int), .bgr(bgr));
ml_hv_hotswitch Ixcvr_vpxa_int ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa_int), .hv_out_hv(vpp));
ml_hv_hotswitch Ixcvr_vpxa ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa), .hv_out_hv(vpp));
ml_hvmux_hotswitch Isw_sbhvsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(sbhvsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sb25sup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sb25sup_vpxa_25), .sel_hv_a_25(sb25sup_vddp_25),
     .out_hv(sb25sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_ngate ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(ngate_vpxa_25), .sel_hv_a_25(ngate_vddp_25),
     .out_hv(ngate_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_1_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vpxa_int), .hvin_a_hv(vpxa_int));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_0_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vpxa_int), .hvin_a_hv(vpxa_int));
ml_ysup_25_switch Isw_ysup25_1_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ysup_25_switch Isw_ysup25_0_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
vddp_tiehigh I188_9_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_8_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_0_ ( .vddp_tieh(vddp_tieh));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_1_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_0_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));

endmodule
// Library - NVCM, Cell - ml_hvmux_hotswitch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:28:27 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch_enhance ( hvin_a_hv, hvin_b_hv, out_hv,
     sel_hv_a_25, sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch_enhance Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - sbtlibn65lp, Cell - oai22x2_hvt, View - schematic
// LAST TIME SAVED: Jan 24 13:53:38 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module oai22x2_hvt ( Y, A0, A1, B0, B1 );
output  Y;

input  A0, A1, B0, B1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(Y), .B(GND_), .G(A0), .S(net024));
nch_hvt  M8 ( .D(Y), .B(GND_), .G(A1), .S(net024));
nch_hvt  M10 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M4 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - sbtlibn65lp, Cell - anor31_hvt, View - schematic
// LAST TIME SAVED: Feb 13 14:15:10 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module anor31_hvt ( Y, A, B, C, D );
output  Y;

input  A, B, C, D;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(Y), .B(gnd_), .G(A), .S(net23));
nch_hvt  M8 ( .D(net030), .B(gnd_), .G(C), .S(gnd_));
nch_hvt  M6 ( .D(net23), .B(gnd_), .G(B), .S(net030));
nch_hvt  M7 ( .D(Y), .B(gnd_), .G(D), .S(gnd_));
pch_hvt  M5 ( .D(Y), .B(vdd_), .G(D), .S(net35));
pch_hvt  M4 ( .D(net35), .B(vdd_), .G(A), .S(vdd_));
pch_hvt  M3 ( .D(net35), .B(vdd_), .G(B), .S(vdd_));
pch_hvt  M2 ( .D(net35), .B(vdd_), .G(C), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_logic, View - schematic
// LAST TIME SAVED: May  9 14:35:36 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_logic ( gnv, gred, gwl_misc, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, s, sa_trim, saen, testdec_en_b, testdec_even_b,
     testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd, fsm_coladd, fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_trow, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_dma, tm_testdec, tm_testdec_wr );
output  gwl_misc, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, saen, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [1:0]  gred;
output [3:0]  s;
output [2:0]  sa_trim;
output [5:0]  gnv;

input [2:0]  fsm_trim_rrefpgm;
input [0:0]  fsm_coladd;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_b;

wire  [5:0]  gnv_b;

wire  [1:0]  xadd_b;

wire  [1:0]  gred_b;

wire  [1:0]  xadd;

wire  [0:2]  net390;

wire  [2:0]  sa_trim_b;

wire  [0:1]  net386;



vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
anor21_hvt I109_1_ ( .A(net386[0]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I109_0_ ( .A(net386[1]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
oai22x2_hvt I93 ( .A1(fsm_rd), .Y(net196), .A0(fsm_pgmvfy),
     .B0(gnd_tiel), .B1(gnd_tiel));
ml_pump_a_clkdly I230 ( .in(net0231), .out(net0232));
ml_pump_a_clkdly I208 ( .in(net200), .out(net201));
ml_pump_a_clkdly I202 ( .in(net202), .out(net203));
ml_pump_a_clkdly I198 ( .in(net204), .out(net205));
ml_pump_a_clkdly I207 ( .in(net206), .out(net207));
nor4_hvt I175 ( .D(fsm_tm_allwl_h), .B(fsm_pgmvfy), .Y(net211),
     .A(fsm_pgmvfy), .C(fsm_rd));
nor4_hvt I176 ( .D(testdec_wp), .B(fsm_nvcmen_b), .Y(net216),
     .A(fsm_wren_b), .C(net331));
nor4_hvt I218 ( .D(net282), .B(fsm_tm_allbl_l), .Y(net0258),
     .A(fsm_tm_allbl_l), .C(fsm_nvcmen_b));
nor4_hvt I191 ( .B(pgm_hvpulse), .Y(wrsup_2vdd_int), .D(fsm_nvcmen_b),
     .A(pgm_hvpulse), .C(testdec_wr));
nor4_hvt I171 ( .D(fsm_wpen_b), .B(fsm_nvcmen_b), .Y(net226),
     .A(testdec_wr), .C(fsm_tm_allwl_l));
nor2_hvt I233 ( .A(fsm_pgm), .B(fsm_pgmvfy), .Y(net0176));
nor2_hvt I228 ( .A(fsm_pgmdisc), .B(fsm_pgmhv), .Y(net0231));
nor2_hvt I231 ( .A(net0258), .B(tm_testdec), .Y(pgminhi_dmmy_b));
nor2_hvt I165 ( .B(fsm_nv_sisi_ui), .Y(x1_desel_b),
     .A(fsm_nv_rri_trim));
nor2_hvt I186 ( .A(fsm_pgmvfy), .B(fsm_pgm_b), .Y(stress2));
nor2_hvt I216 ( .A(fsm_nvcmen_b), .B(tm_dma), .Y(saen));
nor2_hvt I203 ( .A(net203), .B(net351), .Y(gwlbsup_vpxa));
nor2_hvt I209 ( .A(net207), .B(net246), .Y(gwphv_vppint));
nor2_hvt I214 ( .A(net0232), .B(fsm_nvcmen_b), .Y(net246));
nor2_hvt I210 ( .A(net359), .B(net201), .Y(gwphv_vddp));
nor2_hvt I226 ( .A(net0288), .B(net0390), .Y(gwlb_en));
nor2_hvt I201 ( .A(net196), .B(net205), .Y(gwlbsup_vddp));
nor3_hvt I182 ( .B(fsm_tm_allwl_l), .Y(net330), .A(fsm_tm_allwl_l),
     .C(fsm_tm_allwl_l));
nor3_hvt I105 ( .B(fsm_tm_allwl_h), .Y(net0288), .A(fsm_tm_allwl_h),
     .C(fsm_tm_allwl_h));
nor3_hvt I162 ( .Y(net0274), .B(fsm_tm_trow), .C(fsm_nv_sisi_ui),
     .A(fsm_nv_rri_trim));
anor31_hvt I121_3_ ( .A(net365), .D(net345), .B(xadd[1]), .Y(s_b[3]),
     .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net365), .D(net345), .B(xadd[1]), .Y(s_b[2]),
     .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net365), .D(net345), .B(xadd_b[1]), .Y(s_b[1]),
     .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net365), .D(net345), .B(xadd_b[1]), .Y(s_b[0]),
     .C(xadd_b[0]));
nand3_hvt I167 ( .B(fsm_nvcmen), .Y(gwlb_dis), .A(net0332),
     .C(testwr_wpgnd_b));
nand3_hvt I184 ( .Y(net274), .B(fsm_tm_allwl_h), .C(fsm_tm_allwl_h),
     .A(stress2));
nand3_hvt I125 ( .C(fsm_ymuxdis), .A(tm_testdec), .Y(testdec_prec_b),
     .B(fsm_rd));
nand3_hvt I195 ( .Y(net282), .B(net341), .C(fsm_lshven), .A(fsm_pgm));
nand3_hvt I154 ( .Y(net286), .B(fsm_pgm), .C(fsm_tm_allwl_h),
     .A(fsm_wren));
nand3_hvt I122 ( .A(fsm_nvcmen), .C(net307), .Y(net292),
     .B(tm_allwl_l_b));
nand2_hvt I170 ( .A(tm_testdec_wr), .Y(testwr_wpgnd_b),
     .B(tm_testdec));
nand2_hvt I188 ( .A(testdec_en), .Y(testdec_odd_b), .B(fsm_coladd[0]));
nand2_hvt I189 ( .A(net355), .Y(testdec_even_b), .B(testdec_en));
nand2_hvt I155 ( .A(net377), .Y(net307), .B(tm_testdec));
nand2_hvt I89 ( .A(fsm_rd), .Y(testdec_en_b), .B(tm_testdec));
inv_hvt I232 ( .A(net0176), .Y(net0365));
inv_hvt I174 ( .A(net211), .Y(wp_frcen));
inv_hvt I163 ( .A(net0274), .Y(gwl_misc));
inv_hvt I187 ( .A(fsm_pgm), .Y(fsm_pgm_b));
inv_hvt I131 ( .A(testdec_en_b), .Y(testdec_en));
inv_hvt I178 ( .A(net307), .Y(testdec_wp));
inv_hvt I196 ( .A(net282), .Y(pgm_hvpulse));
inv_hvt I185 ( .A(net274), .Y(wr_frcen));
inv_hvt I206 ( .A(gwlbsup_vpxa), .Y(net204));
inv_hvt I177 ( .A(net216), .Y(wr_dis));
inv_hvt I183 ( .A(net330), .Y(net331));
inv_hvt I192 ( .A(wrsup_2vdd_int), .Y(net333));
inv_hvt I179 ( .A(fsm_wpen), .Y(fsm_wpen_b));
inv_hvt I194 ( .A(testwr_wpgnd_b), .Y(testdec_wr));
inv_hvt I212 ( .A(gwphv_vddp), .Y(net206));
inv_hvt I197 ( .A(fsm_pgmvfy), .Y(net341));
inv_hvt I205 ( .A(gwlbsup_vddp), .Y(net202));
inv_hvt I152 ( .A(net286), .Y(net345));
inv_hvt I120_5_ ( .A(gnv_b[5]), .Y(gnv[5]));
inv_hvt I120_4_ ( .A(gnv_b[4]), .Y(gnv[4]));
inv_hvt I120_3_ ( .A(gnv_b[3]), .Y(gnv[3]));
inv_hvt I120_2_ ( .A(gnv_b[2]), .Y(gnv[2]));
inv_hvt I120_1_ ( .A(gnv_b[1]), .Y(gnv[1]));
inv_hvt I120_0_ ( .A(gnv_b[0]), .Y(gnv[0]));
inv_hvt I172 ( .A(net226), .Y(wp_dis));
inv_hvt I204 ( .A(net196), .Y(net351));
inv_hvt I160_1_ ( .A(gred_b[1]), .Y(gred[1]));
inv_hvt I160_0_ ( .A(gred_b[0]), .Y(gred[0]));
inv_hvt I190 ( .A(fsm_coladd[0]), .Y(net355));
inv_hvt I150_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I150_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I215 ( .A(net246), .Y(net359));
inv_hvt I225 ( .A(pgm_hvpulse), .Y(net0390));
inv_hvt I213 ( .A(gwphv_vppint), .Y(net200));
inv_hvt I161_1_ ( .A(fsm_rowadd[3]), .Y(gred_b[1]));
inv_hvt I161_0_ ( .A(fsm_rowadd[2]), .Y(gred_b[0]));
inv_hvt I151 ( .A(net292), .Y(net365));
inv_hvt I119_5_ ( .A(fsm_rowadd[7]), .Y(gnv_b[5]));
inv_hvt I119_4_ ( .A(fsm_rowadd[6]), .Y(gnv_b[4]));
inv_hvt I119_3_ ( .A(fsm_rowadd[5]), .Y(gnv_b[3]));
inv_hvt I119_2_ ( .A(fsm_rowadd[4]), .Y(gnv_b[2]));
inv_hvt I119_1_ ( .A(fsm_rowadd[3]), .Y(gnv_b[1]));
inv_hvt I119_0_ ( .A(fsm_rowadd[2]), .Y(gnv_b[0]));
inv_hvt I157 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I153 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I193 ( .A(net333), .Y(wrsup_2vdd));
inv_hvt I181 ( .A(fsm_wren), .Y(fsm_wren_b));
inv_hvt I156 ( .A(tm_testdec_wr), .Y(net377));
inv_hvt I147_3_ ( .A(s_b[3]), .Y(s[3]));
inv_hvt I147_2_ ( .A(s_b[2]), .Y(s[2]));
inv_hvt I147_1_ ( .A(s_b[1]), .Y(s[1]));
inv_hvt I147_0_ ( .A(s_b[0]), .Y(s[0]));
inv_hvt I25_2_ ( .A(sa_trim_b[2]), .Y(sa_trim[2]));
inv_hvt I25_1_ ( .A(sa_trim_b[1]), .Y(sa_trim[1]));
inv_hvt I25_0_ ( .A(sa_trim_b[0]), .Y(sa_trim[0]));
inv_hvt I24_2_ ( .A(net390[0]), .Y(sa_trim_b[2]));
inv_hvt I24_1_ ( .A(net390[1]), .Y(sa_trim_b[1]));
inv_hvt I24_0_ ( .A(net390[2]), .Y(sa_trim_b[0]));
mux2_hvt I180_1_ ( .in1(fsm_rowadd[1]), .in0(fsm_rowadd[1]),
     .out(net386[0]), .sel(fsm_nv_rrow));
mux2_hvt I180_0_ ( .in1(fsm_rowadd[0]), .in0(fsm_rowadd[0]),
     .out(net386[1]), .sel(fsm_nv_rrow));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net390[0]), .sel(net0365));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net390[1]), .sel(net0365));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net390[2]), .sel(net0365));
mux2_hvt I221 ( .in1(fsm_wpen), .in0(fsm_wgnden), .out(net0332),
     .sel(pgm_hvpulse));

endmodule
// Library - NVCM, Cell - ml_gwlwr_bldrv, View - schematic
// LAST TIME SAVED: Apr  9 11:04:12 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwlwr_bldrv ( bgr, bl_pgm_glb, bl_frc_gnd, fsm_din, fsm_pgm,
     fsm_pgmien, fsm_trim_ipp, tm_dma );
inout  bgr, bl_pgm_glb;

input  bl_frc_gnd, fsm_din, fsm_pgm, fsm_pgmien, tm_dma;

input [3:0]  fsm_trim_ipp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net0152;

wire  [0:3]  net0172;

wire  [0:3]  net0156;

wire  [0:7]  net0115;

wire  [0:1]  net0180;

wire  [0:1]  net0160;



nand2_hvt I71 ( .B(fsm_din), .A(fsm_pgmien), .Y(fsm_pgmien_b_buf));
nor2_hvt I121 ( .A(net086), .B(fsm_pgmien_b_buf), .Y(pgm_trim0_en));
nor2_hvt I114 ( .B(tm_dma), .Y(net0116), .A(tm_dma));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
nor4_hvt I105 ( .D(fsm_trim_ipp[0]), .B(fsm_trim_ipp[2]), .Y(net086),
     .A(fsm_trim_ipp[3]), .C(fsm_trim_ipp[1]));
nch_hvt  M36 ( .D(net0173), .B(GND_), .G(pgm_trim0_en), .S(net0107));
nch_hvt  M37 ( .D(net0107), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M31_7_ ( .D(net0115[0]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[0]));
nch_hvt  M31_6_ ( .D(net0115[1]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[1]));
nch_hvt  M31_5_ ( .D(net0115[2]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[2]));
nch_hvt  M31_4_ ( .D(net0115[3]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[3]));
nch_hvt  M31_3_ ( .D(net0115[4]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[4]));
nch_hvt  M31_2_ ( .D(net0115[5]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[5]));
nch_hvt  M31_1_ ( .D(net0115[6]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[6]));
nch_hvt  M31_0_ ( .D(net0115[7]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[7]));
nch_hvt  M19 ( .D(net0135), .B(GND_), .G(fsm_trim_ipp[0]),
     .S(net0131));
nch_hvt  M38_7_ ( .D(net0152[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_6_ ( .D(net0152[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_5_ ( .D(net0152[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_4_ ( .D(net0152[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_3_ ( .D(net0152[4]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_2_ ( .D(net0152[5]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_1_ ( .D(net0152[6]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_0_ ( .D(net0152[7]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_3_ ( .D(net0156[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_2_ ( .D(net0156[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_1_ ( .D(net0156[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_0_ ( .D(net0156[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_1_ ( .D(net0160[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_0_ ( .D(net0160[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M26 ( .D(net0131), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M33 ( .D(bl_pgm_glb), .B(GND_), .G(net0187), .S(gnd_));
nch_hvt  M30_3_ ( .D(net0172[0]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[0]));
nch_hvt  M30_2_ ( .D(net0172[1]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[1]));
nch_hvt  M30_1_ ( .D(net0172[2]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[2]));
nch_hvt  M30_0_ ( .D(net0172[3]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[3]));
nch_hvt  M34 ( .D(net089), .B(GND_), .G(pgm_trim0_en), .S(gnd_));
nch_hvt  M27_1_ ( .D(net0180[0]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[0]));
nch_hvt  M27_0_ ( .D(net0180[1]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[1]));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net0114), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net0114), .PLUS(net0141), .BULK(GND_));
inv_hvt I115 ( .A(net0116), .Y(net0187));
inv_hvt I58 ( .A(pgmen_b), .Y(pgmen));
inv_hvt I131 ( .A(fsm_pgm), .Y(pgmen_b));
inv_hvt I72 ( .A(fsm_pgmien_b_buf), .Y(fsm_pgmien_buf));
ml_ls_vdd2vdd25 I56 ( .in(pgmen), .sup(vddp_),
     .out_vddio_b(pgmen_b_25), .out_vddio(pgmen_25), .in_b(pgmen_b));
nch_25  M20 ( .D(net0173), .B(GND_), .G(pgm_inhi_bias),
     .S(bl_pgm_glb));
nch_25  M21 ( .D(pgm_inhi_bias), .B(GND_), .G(pgm_inhi_bias),
     .S(gnd_));
nch_25  M12_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[0]));
nch_25  M12_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[1]));
nch_25  M13_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[0]));
nch_25  M13_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[1]));
nch_25  M13_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[2]));
nch_25  M13_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[3]));
nch_25  M6 ( .D(net0164), .B(GND_), .G(net0164), .S(gnd_));
nch_25  M3 ( .D(dec_bias_p), .B(GND_), .G(bgr), .S(net0141));
nch_25  M10 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net089));
nch_25  M18_7_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[0]));
nch_25  M18_6_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[1]));
nch_25  M18_5_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[2]));
nch_25  M18_4_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[3]));
nch_25  M18_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[4]));
nch_25  M18_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[5]));
nch_25  M18_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[6]));
nch_25  M18_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[7]));
nch_25  M9 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net0135));
nch_25  M8 ( .D(net0164), .B(GND_), .G(pgmen_b_25), .S(gnd_));
pch_25  M11 ( .D(pgm_inhi_bias), .B(vddp_), .G(vdd_tieh), .S(net0259));
pch_25  M14_1_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M14_0_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M5 ( .D(net0164), .B(vddp_), .G(dec_bias_p), .S(net0199));
pch_25  M7_1_ ( .D(net0199), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M7_0_ ( .D(net0199), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M4 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p), .S(net0199));

endmodule
// Library - NVCM, Cell - ml_ymux_vblinhi_pgm_drv, View - schematic
// LAST TIME SAVED: Apr  8 10:44:07 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_ymux_vblinhi_pgm_drv ( vblinhi_pgm_25, ysup_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25 );
inout  vblinhi_pgm_25, ysup_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd_), .B(GND_), .G(en_blinhi_pgm_b_ysup_25),
     .S(vblinhi_pgm_25));
pch_25  M5 ( .D(net10), .B(ysup_25), .G(en_blinhi_pgm_b_ysup_25),
     .S(ysup_25));
pch_25  M0 ( .D(net10), .B(vblinhi_pgm_25), .G(en_blinhi_pgm_b),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_wr_sup, View - schematic
// LAST TIME SAVED: Jan 24 10:11:13 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_wr_sup ( wr_sup_25, wrsup_2vdd, wrsup_2vdd_25 );
inout  wr_sup_25;

input  wrsup_2vdd, wrsup_2vdd_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I120 ( .A(net19), .Y(wrsup_vdd_in));
inv_hvt I131 ( .A(wrsup_2vdd), .Y(net19));
inv_25 I119 ( .IN(net20), .OUT(wrsup_vdd_in_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(wrsup_2vdd_25), .OUT(net20), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_2_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_1_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_0_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));

endmodule
// Library - misc, Cell - ml_osc, View - schematic
// LAST TIME SAVED: Aug 28 14:10:03 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_osc ( clk_out, smc_osc_fsel, smc_oscen );
output  clk_out;

input  smc_oscen;

input [1:0]  smc_osc_fsel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sel_trim;



tielo I272 ( .tielo(net0103));
tiehi I219 ( .tiehi(net0106));
ml_osc_stage I254 ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_b_buf), .out(out_bot), .sel_trim(sel_trim[3:0]));
ml_osc_stage I255 ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_buf), .out(out_top), .sel_trim(sel_trim[3:0]));
ml_osc_logic Iosc_logic ( .sel_trim(sel_trim[3:0]),
     .smc_oscen(smc_oscen), .smc_osc_fsel(smc_osc_fsel[1:0]),
     .clkin(clk_out));
ml_dff I174 ( .R(oscen_b), .D(clkby2_b), .CLK(clk_dffin),
     .QN(clkby2_b), .Q(clkby2));
nor3_hvt I256 ( .B(net079), .Y(net075), .A(net079), .C(net079));
nor3_hvt I218 ( .B(net083), .Y(net079), .A(net083), .C(net083));
nor3_hvt I217 ( .B(net0106), .Y(net083), .A(net0106), .C(net0106));
nand3_hvt I224 ( .Y(net088), .B(net0106), .C(net0106), .A(net0106));
nand3_hvt I230 ( .Y(net092), .B(net088), .C(net088), .A(net088));
nand3_hvt I231 ( .Y(net096), .B(net092), .C(net092), .A(net092));
rppolywo_m  R18 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net362), .PLUS(net356), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net356), .PLUS(pbias), .BULK(gnd_));
rppolywo_m  R7 ( .BULK(gnd_), .MINUS(net383), .PLUS(net366));
rppolywo_m  R2 ( .MINUS(net366), .PLUS(net362), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net437), .PLUS(net383), .BULK(gnd_));
nand2_hvt I175 ( .A(out_bot), .Y(clk_dffin), .B(out_top));
inv_hvt I222 ( .A(clkby2), .Y(clkby2_b_buf));
inv_hvt I220 ( .A(clkby2_b), .Y(clkby2_buf));
inv_hvt I176 ( .A(clkby2_b), .Y(clk_out));
inv_hvt I248 ( .A(net0103), .Y(net0226));
inv_hvt I198 ( .A(smc_oscen), .Y(oscen_b));
nch_hvt  M45 ( .D(gnd_), .B(gnd_), .G(gnd_), .S(gnd_));
nch_hvt  MN31 ( .D(net437), .B(gnd_), .G(smc_oscen), .S(gnd_));
nch_hvt  MN44 ( .D(pbias), .B(gnd_), .G(net0103), .S(net371));
pch_hvt  MP77 ( .D(net371), .B(vdd_), .G(net0226), .S(pbias));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(vdd_), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(smc_oscen), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_ls25_1b, View - schematic
// LAST TIME SAVED: Jan 23 16:20:39 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25_1b ( out_25, in );
output  out_25;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I145 ( .A(in), .Y(net45));
inv_25 I153 ( .IN(out_b_25), .OUT(out_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I112 ( .in(in), .sup(vddp_), .out_vddio_b(out_b_25),
     .out_vddio(net025), .in_b(net45));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_ls25, View - schematic
// LAST TIME SAVED: May  1 10:33:06 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25 ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25,
     gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25, s_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wrsup_2vdd_25, fsm_gwlbdis, gnv, gred, gwl_misc, gwl_nvcm,
     gwl_red, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, s, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wrsup_2vdd_25;

input  fsm_gwlbdis, gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, testdec_en_b, testdec_even_b, testdec_odd_b,
     testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen, wrsup_2vdd;

output [5:0]  gnv_b_25;
output [3:0]  s_25;
output [1:0]  gred_25;
output [5:0]  gnv_25;
output [1:0]  gred_b_25;

input [5:0]  gnv;
input [3:0]  s;
input [1:0]  gred;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I_1_ ( .IN(gred_25[1]), .OUT(gred_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I_0_ ( .IN(gred_25[0]), .OUT(gred_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I143 ( .IN(net101), .OUT(fsm_gwlbdis_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_5_ ( .IN(gnv_25[5]), .OUT(gnv_b_25[5]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_4_ ( .IN(gnv_25[4]), .OUT(gnv_b_25[4]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_3_ ( .IN(gnv_25[3]), .OUT(gnv_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_2_ ( .IN(gnv_25[2]), .OUT(gnv_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_1_ ( .IN(gnv_25[1]), .OUT(gnv_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_0_ ( .IN(gnv_25[0]), .OUT(gnv_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_gwlwr_ctrl_ls25_1b I133 ( .in(testdec_en_b),
     .out_25(testdec_en_b_25));
ml_gwlwr_ctrl_ls25_1b I139 ( .in(gwlb_dis), .out_25(gwlb_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_frcen ( .in(wr_frcen),
     .out_25(wr_frcen_25));
ml_gwlwr_ctrl_ls25_1b I144 ( .in(gwlb_en), .out_25(gwlb_en_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vpp ( .in(gwphv_vppint),
     .out_25(gwphv_vppint_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwlb_vddp ( .in(gwlbsup_vddp),
     .out_25(gwlbsup_vddp_25));
ml_gwlwr_ctrl_ls25_1b ls25_gwlb_vpp ( .in(gwlbsup_vpxa),
     .out_25(gwlbsup_vpxa_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_vdd ( .in(wrsup_2vdd),
     .out_25(wrsup_2vdd_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_dis ( .in(wr_dis), .out_25(wr_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vddp ( .in(gwphv_vddp),
     .out_25(gwphv_vddp_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_frcen ( .in(wp_frcen),
     .out_25(wp_frcen_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_dis ( .in(wp_dis), .out_25(wp_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwl_red ( .in(gwl_red),
     .out_25(gwl_red_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_nvcm ( .in(gwl_nvcm),
     .out_25(gwl_nvcm_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_misc ( .in(gwl_misc),
     .out_25(gwl_misc_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_1_ ( .in(gred[1]),
     .out_25(gred_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_0_ ( .in(gred[0]),
     .out_25(gred_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_5_ ( .in(gnv[5]), .out_25(gnv_25[5]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_4_ ( .in(gnv[4]), .out_25(gnv_25[4]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_3_ ( .in(gnv[3]), .out_25(gnv_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_2_ ( .in(gnv[2]), .out_25(gnv_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_1_ ( .in(gnv[1]), .out_25(gnv_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_0_ ( .in(gnv[0]), .out_25(gnv_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_3_ ( .in(s[3]), .out_25(s_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_2_ ( .in(s[2]), .out_25(s_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_1_ ( .in(s[1]), .out_25(s_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_0_ ( .in(s[0]), .out_25(s_25[0]));
ml_gwlwr_ctrl_ls25_1b I134 ( .in(testdec_prec_b),
     .out_25(testdec_prec_b_25));
ml_gwlwr_ctrl_ls25_1b I136 ( .in(pgminhi_dmmy_b),
     .out_25(pgminhi_dmmy_b_25));
ml_gwlwr_ctrl_ls25_1b I140 ( .in(fsm_gwlbdis), .out_25(net101));
ml_gwlwr_ctrl_ls25_1b I137 ( .in(testdec_even_b),
     .out_25(testdec_even_b_25));
ml_gwlwr_ctrl_ls25_1b I138 ( .in(testdec_odd_b),
     .out_25(testdec_odd_b_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_npgate_gen, View - schematic
// LAST TIME SAVED: Sep 15 17:21:19 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_core_sa_npgate_gen ( dec_trim, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, vpxa, fsm_tm_testdec, saen, satrim,
     vddp_tieh );
output  saen_25, saen_b_vpxa;

inout  vpxa;

input  fsm_tm_testdec, saen, vddp_tieh;

output [4:1]  sa_ngate_25;
output [7:0]  dec_trim;
output [4:1]  sa_pgate_vpxa;

input [2:0]  satrim;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  ydec_b;

wire  [2:0]  ydec;

wire  [7:0]  dec_trim_b;

wire  [4:1]  pgate_in;

wire  [4:1]  ngate_in_25_b;

wire  [4:1]  trim;

wire  [4:1]  trim_b;

wire  [0:3]  net53;

wire  [0:3]  net48;

wire  [0:3]  net36;



nor4_hvt I102 ( .D(fsm_tm_testdec), .C(dec_trim[7]), .A(dec_trim[5]),
     .B(dec_trim[6]), .Y(net47));
ml_hv_invx3 I135 ( .sel_hv(net048), .sel_25(net048),
     .vddp_tieh(vddp_tieh), .out_b_hv(saen_b_vpxa), .in_hv(vpxa));
ml_hv_invx3 I130_4_ ( .sel_hv(pgate_in[4]), .sel_25(pgate_in[4]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[4]), .in_hv(vpxa));
ml_hv_invx3 I130_3_ ( .sel_hv(pgate_in[3]), .sel_25(pgate_in[3]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[3]), .in_hv(vpxa));
ml_hv_invx3 I130_2_ ( .sel_hv(pgate_in[2]), .sel_25(pgate_in[2]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[2]), .in_hv(vpxa));
ml_hv_invx3 I130_1_ ( .sel_hv(pgate_in[1]), .sel_25(pgate_in[1]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[1]), .in_hv(vpxa));
inv_25 I149 ( .IN(net052), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I153_4_ ( .IN(ngate_in_25_b[4]), .OUT(sa_ngate_25[4]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_3_ ( .IN(ngate_in_25_b[3]), .OUT(sa_ngate_25[3]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_2_ ( .IN(ngate_in_25_b[2]), .OUT(sa_ngate_25[2]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_1_ ( .IN(ngate_in_25_b[1]), .OUT(sa_ngate_25[1]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_4_ ( .Y(dec_trim_b[4]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_3_ ( .Y(dec_trim_b[3]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_2_ ( .Y(dec_trim_b[2]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nand3_hvt I37_1_ ( .Y(dec_trim_b[1]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_0_ ( .Y(dec_trim_b[0]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nor2_hvt I75_4_ ( .Y(net48[0]), .B(dec_trim[4]), .A(sa_high_res));
nor2_hvt I75_3_ ( .Y(net48[1]), .B(dec_trim[3]), .A(trim[4]));
nor2_hvt I75_2_ ( .Y(net48[2]), .B(dec_trim[2]), .A(trim[3]));
nor2_hvt I75_1_ ( .Y(net48[3]), .B(dec_trim[1]), .A(trim[2]));
inv_hvt I145 ( .A(net076), .Y(net078));
inv_hvt I143 ( .A(net078), .Y(net080));
inv_hvt I146 ( .A(saen), .Y(net076));
inv_hvt I114 ( .A(net47), .Y(sa_high_res));
inv_hvt I38_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I38_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I38_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I38_4_ ( .A(dec_trim_b[4]), .Y(dec_trim[4]));
inv_hvt I38_3_ ( .A(dec_trim_b[3]), .Y(dec_trim[3]));
inv_hvt I38_2_ ( .A(dec_trim_b[2]), .Y(dec_trim[2]));
inv_hvt I38_1_ ( .A(dec_trim_b[1]), .Y(dec_trim[1]));
inv_hvt I38_0_ ( .A(dec_trim_b[0]), .Y(dec_trim[0]));
inv_hvt I40_2_ ( .A(ydec_b[2]), .Y(ydec[2]));
inv_hvt I40_1_ ( .A(ydec_b[1]), .Y(ydec[1]));
inv_hvt I40_0_ ( .A(ydec_b[0]), .Y(ydec[0]));
inv_hvt I76_4_ ( .A(net48[0]), .Y(trim[4]));
inv_hvt I76_3_ ( .A(net48[1]), .Y(trim[3]));
inv_hvt I76_2_ ( .A(net48[2]), .Y(trim[2]));
inv_hvt I76_1_ ( .A(net48[3]), .Y(trim[1]));
inv_hvt I39_2_ ( .A(satrim[2]), .Y(ydec_b[2]));
inv_hvt I39_1_ ( .A(satrim[1]), .Y(ydec_b[1]));
inv_hvt I39_0_ ( .A(satrim[0]), .Y(ydec_b[0]));
inv_hvt I78_4_ ( .A(trim[4]), .Y(trim_b[4]));
inv_hvt I78_3_ ( .A(trim[3]), .Y(trim_b[3]));
inv_hvt I78_2_ ( .A(trim[2]), .Y(trim_b[2]));
inv_hvt I78_1_ ( .A(trim[1]), .Y(trim_b[1]));
ml_ls_vdd2vdd25 I128_4_ ( .in(ngate_in_25_b[4]), .sup(vpxa),
     .out_vddio_b(pgate_in[4]), .out_vddio(net53[0]), .in_b(net36[0]));
ml_ls_vdd2vdd25 I128_3_ ( .in(ngate_in_25_b[3]), .sup(vpxa),
     .out_vddio_b(pgate_in[3]), .out_vddio(net53[1]), .in_b(net36[1]));
ml_ls_vdd2vdd25 I128_2_ ( .in(ngate_in_25_b[2]), .sup(vpxa),
     .out_vddio_b(pgate_in[2]), .out_vddio(net53[2]), .in_b(net36[2]));
ml_ls_vdd2vdd25 I128_1_ ( .in(ngate_in_25_b[1]), .sup(vpxa),
     .out_vddio_b(pgate_in[1]), .out_vddio(net53[3]), .in_b(net36[3]));
ml_ls_vdd2vdd25 I136 ( .in(net053), .sup(vpxa), .out_vddio_b(net047),
     .out_vddio(net048), .in_b(net052));
ml_ls_vdd2vdd25 I137 ( .in(net078), .sup(vddp_), .out_vddio_b(net052),
     .out_vddio(net053), .in_b(net080));
ml_ls_vdd2vdd25 I129_4_ ( .in(trim[4]), .sup(vddp_),
     .out_vddio_b(net36[0]), .out_vddio(ngate_in_25_b[4]),
     .in_b(trim_b[4]));
ml_ls_vdd2vdd25 I129_3_ ( .in(trim[3]), .sup(vddp_),
     .out_vddio_b(net36[1]), .out_vddio(ngate_in_25_b[3]),
     .in_b(trim_b[3]));
ml_ls_vdd2vdd25 I129_2_ ( .in(trim[2]), .sup(vddp_),
     .out_vddio_b(net36[2]), .out_vddio(ngate_in_25_b[2]),
     .in_b(trim_b[2]));
ml_ls_vdd2vdd25 I129_1_ ( .in(trim[1]), .sup(vddp_),
     .out_vddio_b(net36[3]), .out_vddio(ngate_in_25_b[1]),
     .in_b(trim_b[1]));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl, View - schematic
// LAST TIME SAVED: May  1 11:11:08 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25, gred_25,
     gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25,
     gwlb_en_25, pgminhi_dmmy_b_25, s_25, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv,
     vddp_tieh, vpp_int, vpxa, wr_sup_25, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

inout  bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv, vddp_tieh, vpp_int,
     vpxa, wr_sup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [5:0]  gnv_25;
output [5:0]  gnv_b_25;
output [1:0]  gred_25;
output [4:1]  sa_ngate_25;
output [3:0]  s_25;
output [1:0]  gred_b_25;
output [4:1]  sa_pgate_vpxa;

input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
input [0:0]  fsm_coladd;
input [3:0]  fsm_trim_ipp;
input [7:0]  fsm_rowadd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  sa_trim;

wire  [3:0]  s;

wire  [1:0]  gred;

wire  [5:0]  gnv;

wire  [7:0]  dec_trim;



ml_hvmux_hotswitch_enhance Ihvmux_gwpsup_hv ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwphv_vppint_25), .sel_hv_a_25(gwphv_vddp_25),
     .out_hv(gwp_sup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_gwlwr_ctrl_logic Igwlwr_ctrl_logic ( .fsm_pgmdisc(fsm_pgmdisc),
     .gwlb_en(gwlb_en), .tm_testdec_wr(tm_testdec_wr),
     .tm_testdec(tm_testdec), .tm_dma(tm_dma),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_rd(fsm_rd), .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[0]), .wrsup_2vdd(wrsup_2vdd),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .testdec_prec_b(net172),
     .testdec_odd_b(testdec_odd_b), .testdec_even_b(testdec_even_b),
     .testdec_en_b(net175), .saen(saen), .sa_trim(sa_trim[2:0]),
     .s(s[3:0]), .pgminhi_dmmy_b(net179), .gwphv_vppint(gwphv_vppint),
     .gwphv_vddp(gwphv_vddp), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vddp(gwlbsup_vddp), .gwlb_dis(gwlb_dis),
     .gwl_misc(gwl_misc), .gred(gred[1:0]), .gnv(gnv[5:0]));
ml_hvmux_hotswitch Ihvmux_gwlbsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwlbsup_vpxa_25), .sel_hv_a_25(gwlbsup_vddp_25),
     .out_hv(gwl_b_sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_gwlwr_bldrv Igwlwr_bldrv ( .fsm_din(fsm_din), .tm_dma(tm_dma),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .bl_frc_gnd(gnd_), .bgr(bgr),
     .bl_pgm_glb(bl_pgm_glb));
ml_gwlwr_ctrl_wr_sup Igwlwr_ctrl_wr_sup ( .wrsup_2vdd(wrsup_2vdd),
     .wrsup_2vdd_25(wrsup_2vdd_25), .wr_sup_25(wr_sup_25));
ml_gwlwr_ctrl_ls25 Igwlwr_ctrl_ls25 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_en(gwlb_en), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwlb_dis(gwlb_dis), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vpxa_25(gwlbsup_vpxa_25), .wrsup_2vdd_25(wrsup_2vdd_25),
     .wrsup_2vdd(wrsup_2vdd), .testdec_odd_b(testdec_odd_b),
     .testdec_even_b(testdec_even_b),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .testdec_prec_b(net172),
     .testdec_en_b(net175), .pgminhi_dmmy_b(net179),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwphv_vddp(gwphv_vddp),
     .gwlbsup_vddp(gwlbsup_vddp), .gwphv_vppint(gwphv_vppint),
     .gwlbsup_vddp_25(gwlbsup_vddp_25),
     .gwphv_vppint_25(gwphv_vppint_25), .gwphv_vddp_25(gwphv_vddp_25),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .s(s[3:0]), .gwl_red(fsm_nv_rrow),
     .gwl_nvcm(fsm_nv_bstream), .gwl_misc(gwl_misc), .gred(gred[1:0]),
     .gnv(gnv[5:0]), .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]));
vddp_tiehigh Ivddp_tiehigh_15_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_14_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_13_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_12_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_11_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_10_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_9_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_8_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_0_ ( .vddp_tieh(vddp_tieh));
ml_core_sa_npgate_gen Icore_sa_npgate_gen (
     .fsm_tm_testdec(tm_testdec), .satrim(sa_trim[2:0]),
     .vddp_tieh(vddp_tieh), .saen(saen), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .dec_trim(dec_trim[7:0]),
     .vpxa(vpxa));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr, View - schematic
// LAST TIME SAVED: Feb 25 14:20:48 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr ( wr, gwl_wr_25, s_25, wr_sup_25 );
output  wr;

input  gwl_wr_25, s_25, wr_sup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_25 I59 ( .A(gwl_wr_25), .Y(net27), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(s_25));
inv_25 I38 ( .IN(net27), .OUT(wr), .P(wr_sup_25), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr_x4, View - schematic
// LAST TIME SAVED: Jan 21 18:09:38 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x4 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  gwl_wr_25, wr_sup_25;

output [3:0]  wr;

input [3:0]  s_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr Iml_lwldrv_2 ( .gwl_wr_25(gwl_wr_25), .wr(wr[2]),
     .s_25(s_25[2]), .wr_sup_25(wr_sup_25));
ml_rock_lwldrv_wr Iml_lwldrv_1 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[1]), .wr(wr[1]));
ml_rock_lwldrv_wr Iml_lwldrv_3 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3]), .wr(wr[3]));
ml_rock_lwldrv_wr Iml_lwldrv_0 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[0]), .wr(wr[0]));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr_x228, View - schematic
// LAST TIME SAVED: Jan 23 13:37:56 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x228 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  wr_sup_25;

output [227:0]  wr;

input [56:0]  gwl_wr_25;
input [3:0]  s_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_56_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[227:224]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[56]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_55_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[223:220]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[55]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_54_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[219:216]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[54]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_53_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[215:212]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[53]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_52_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[211:208]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[52]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_51_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[207:204]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[51]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_50_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[203:200]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[50]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_49_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[199:196]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[49]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_48_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[195:192]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[48]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_47_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[191:188]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[47]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_46_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[187:184]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[46]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_45_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[183:180]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[45]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_44_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[179:176]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[44]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_43_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[175:172]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[43]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_42_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[171:168]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[42]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_41_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[167:164]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[41]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_40_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[163:160]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[40]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_39_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[159:156]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[39]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_38_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[155:152]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[38]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_37_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[151:148]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[37]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_36_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[147:144]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[36]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_35_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[143:140]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[35]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_34_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[139:136]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[34]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_33_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[135:132]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[33]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_32_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[131:128]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[32]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_31_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[127:124]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[31]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_30_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[123:120]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[30]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_29_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[119:116]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[29]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_28_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[115:112]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[28]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_27_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[111:108]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[27]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_26_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[107:104]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[26]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_25_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[103:100]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[25]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_24_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[99:96]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[24]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_23_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[95:92]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[23]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_22_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[91:88]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[22]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_21_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[87:84]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[21]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_20_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[83:80]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[20]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_19_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[79:76]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[19]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_18_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[75:72]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[18]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_17_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[71:68]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[17]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_16_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[67:64]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[16]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_15_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[63:60]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[15]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_14_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[59:56]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[14]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_13_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[55:52]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[13]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_12_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[51:48]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[12]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_11_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[47:44]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[11]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_10_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[43:40]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[10]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_9_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[39:36]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[9]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_8_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[35:32]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[8]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_7_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[31:28]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[7]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_6_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[27:24]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[6]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_5_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[23:20]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[5]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_4_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[19:16]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[4]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_3_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[15:12]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[3]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_2_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[11:8]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[2]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_1_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[7:4]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[1]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_0_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[3:0]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[0]));

endmodule
// Library - NVCM, Cell - ml_ls_vddp2vpxa, View - schematic
// LAST TIME SAVED: Dec 30 20:36:23 2007
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_ls_vddp2vpxa ( out_33, out_b_33, sup, in_25, in_b_25 );
output  out_33, out_b_33;

inout  sup;

input  in_25, in_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(out_b_33), .B(sup), .G(in_25), .S(net29));
pch_25  M13 ( .D(out_33), .B(sup), .G(in_b_25), .S(net33));
pch_25  M4 ( .D(net29), .B(sup), .G(out_33), .S(sup));
pch_25  M6 ( .D(net33), .B(sup), .G(out_b_33), .S(sup));
nch_25  M9 ( .D(out_33), .B(gnd_), .G(in_b_25), .S(gnd_));
nch_25  M15 ( .D(out_b_33), .B(gnd_), .G(in_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_gwhv, View - schematic
// LAST TIME SAVED: May 16 11:27:16 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_gwhv ( gwp_hv, gwp_sup_hv, gwl_25, gwl_25_b,
     vddp_tieh );
output  gwp_hv;

inout  gwp_sup_hv;

input  gwl_25, gwl_25_b, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M10 ( .D(net0129), .B(gnd_), .G(vddp_tieh), .S(net050));
nch_25  M12 ( .D(gwp_hv), .B(gnd_), .G(vddp_tieh), .S(net034));
nch_25  M11 ( .D(net034), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M13 ( .D(net050), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M14 ( .D(net054), .B(gnd_), .G(vddp_tieh), .S(net058));
nch_25  M15 ( .D(net058), .B(gnd_), .G(gwl_25), .S(gnd_));
pch_25  M6 ( .D(net067), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M16 ( .D(gwp_hv), .B(net067), .G(gwl_25_b), .S(net067));
pch_25  M5 ( .D(net054), .B(net087), .G(gwl_25), .S(net087));
pch_25  M8 ( .D(net087), .B(gwp_sup_hv), .G(net0129), .S(gwp_sup_hv));
pch_25  M9 ( .D(net091), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M7 ( .D(net0129), .B(net091), .G(gwl_25_b), .S(net091));

endmodule
// Library - NVCM, Cell - ml_gwl_drv, View - schematic
// LAST TIME SAVED: Apr 30 15:58:52 2008
// NETLIST TIME: Nov 14 16:11:59 2008
`timescale 1ns / 1ns 

module ml_gwl_drv ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25,
     radd_1_25, radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );
output  gwl_b_25, gwl_wr_25, gwp_hv;

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25, radd_1_25,
     radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_ls_vddp2vpxa I99 ( .in_25(gwlb_25), .sup(gwl_b_sup_25),
     .in_b_25(gwlb_b_25), .out_33(out_33), .out_b_33(net053));
nor3_25 I76 ( .C(net84), .A(net68), .Y(dec_sel_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(net76));
nor2_25 I111 ( .A(net096), .Y(gwlb_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_dis_25));
nor2_25 I79 ( .A(wr_dis_25), .Y(gwl_wr_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(net056));
nor2_25 I117 ( .A(dec_sel_25), .Y(net096), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_en_25));
nor2_25 I82 ( .A(dec_sel_25), .Y(net058), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_frcen_25));
nor2_25 I85 ( .A(net058), .Y(gwl_wp_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_dis_25));
nor2_25 I59 ( .B(dec_sel_25), .A(wr_frcen_25), .Y(net056), .P(vddp_),
     .Pb(vddp_), .Gb(gnd_), .G(gnd_));
ml_rock_lwldrv_gwhv Iml_rock_lwldrv_gwhv ( .gwp_sup_hv(gwp_sup_hv),
     .vddp_tieh(vddp_tieh), .gwp_hv(gwp_hv), .gwl_25(gwl_wp_25),
     .gwl_25_b(gwl_wp_b_25));
nand3_25 I44 ( .B(radd_4_25), .A(radd_5_25), .Y(net76), .C(radd_3_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I47 ( .B(radd_1_25), .A(radd_2_25), .Y(net84), .C(radd_0_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I104 ( .B(gwlgrpsel_25), .A(gwlgrpsel_25), .Y(net68),
     .C(radd_6_25), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
inv_25 I38 ( .IN(gwl_wp_25), .OUT(gwl_wp_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I100 ( .IN(out_33), .OUT(gwl_b_25), .P(gwl_b_sup_25),
     .Pb(gwl_b_sup_25), .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(gwlb_25), .OUT(gwlb_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - misc, Cell - ml_osc_top, View - schematic
// LAST TIME SAVED: Oct 14 15:50:05 2008
// NETLIST TIME: Nov 14 16:11:58 2008
`timescale 1ns / 1ns 

module ml_osc_top ( cnt_podt_out, smc_clk, crst_b, por_b, smc_osc_fsel,
     smc_oscoff_b, smc_podt_off, smc_podt_rst );
output  cnt_podt_out, smc_clk;

input  crst_b, por_b, smc_oscoff_b, smc_podt_off, smc_podt_rst;

input [1:0]  smc_osc_fsel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  q_b;

wire  [10:0]  q;



tiehi I179 ( .tiehi(net076));
nor2_hvt I256 ( .A(rst_osc_b), .B(smc_oscoff_b), .Y(net066));
nor2_hvt I266 ( .A(clk_out), .B(smc_podt_off), .Y(net078));
nor2_hvt I257 ( .A(disable_osc), .B(net066), .Y(smc_oscen));
nor2_hvt I264 ( .A(smc_podt_rst), .B(net090), .Y(net054));
nor2_hvt I252 ( .A(cnt_rst), .B(smc_oscoff_b), .Y(net0124));
nand2_hvt I227 ( .A(smc_off_b), .B(rst_osc_b), .Y(disable_osc));
nand2_hvt I270 ( .A(crst_b), .Y(net064), .B(por_b));
ml_dff I230 ( .R(cnt_rst), .D(net076), .CLK(q_b[10]), .QN(net067),
     .Q(net063));
ml_dff I243 ( .R(rst_off_latch), .D(net0174), .CLK(clk_out_b),
     .QN(smc_off_b), .Q(net0152));
ml_dff I228_10_ ( .R(cnt_rst), .D(q_b[10]), .CLK(q[9]), .QN(q_b[10]),
     .Q(q[10]));
ml_dff I228_9_ ( .R(cnt_rst), .D(q_b[9]), .CLK(q[8]), .QN(q_b[9]),
     .Q(q[9]));
ml_dff I228_8_ ( .R(cnt_rst), .D(q_b[8]), .CLK(q[7]), .QN(q_b[8]),
     .Q(q[8]));
ml_dff I228_7_ ( .R(cnt_rst), .D(q_b[7]), .CLK(q[6]), .QN(q_b[7]),
     .Q(q[7]));
ml_dff I228_6_ ( .R(cnt_rst), .D(q_b[6]), .CLK(q[5]), .QN(q_b[6]),
     .Q(q[6]));
ml_dff I228_5_ ( .R(cnt_rst), .D(q_b[5]), .CLK(q[4]), .QN(q_b[5]),
     .Q(q[5]));
ml_dff I228_4_ ( .R(cnt_rst), .D(q_b[4]), .CLK(q[3]), .QN(q_b[4]),
     .Q(q[4]));
ml_dff I228_3_ ( .R(cnt_rst), .D(q_b[3]), .CLK(q[2]), .QN(q_b[3]),
     .Q(q[3]));
ml_dff I228_2_ ( .R(cnt_rst), .D(q_b[2]), .CLK(q[1]), .QN(q_b[2]),
     .Q(q[2]));
ml_dff I228_1_ ( .R(cnt_rst), .D(q_b[1]), .CLK(q[0]), .QN(q_b[1]),
     .Q(q[1]));
ml_dff I228_0_ ( .R(cnt_rst), .D(q_b[0]), .CLK(clk_in), .QN(q_b[0]),
     .Q(q[0]));
inv_hvt I233 ( .A(clk_out), .Y(clk_out_b));
inv_hvt I271 ( .A(net064), .Y(rst_osc_b));
inv_hvt I267 ( .A(net078), .Y(clk_in));
inv_hvt I262 ( .A(net067), .Y(cnt_podt_out));
inv_hvt I244 ( .A(smc_oscoff_b), .Y(net0174));
inv_hvt I265 ( .A(net054), .Y(cnt_rst));
inv_hvt I229 ( .A(rst_osc_b), .Y(net090));
inv_hvt I253 ( .A(net0124), .Y(rst_off_latch));
inv_hvt I232 ( .A(clk_out_b), .Y(smc_clk));
ml_osc Iml_osc ( .smc_osc_fsel(smc_osc_fsel[1:0]), .clk_out(clk_out),
     .smc_oscen(smc_oscen));

endmodule
