---------------------------------------------------------------------------
---------------------------------------------------------------------------
--
--      KEYBOARD SCANNING SYSTEM MODULE
-- 
--      FOR THE LOW-END CIJ PLATFORM FPGA
--
--      VHDL DESIGN FILE :KBD7.VHD
--
--      by: S. Kozich, M. Stamer
--      VIDEOJET TECHNOLOGIES INC.
--
---------------------------------------------------------------------------
---------------------------------------------------------------------------
--
-------------------------------------------------------------------------------
--
-- Copyright 2002 Videojet Technologies Inc. All Rights Reserved. 
--
-- An unpublished work of Videojet Technologies Inc. The software and 
-- documentation contained herein are copyrighted works which include 
-- confidential information and trade secrets proprietary to Videojet 
-- Technologies Inc. and shall not be copied, duplicated, disclosed or used, 
-- in whole or in part, except pursuant to the License Agreement or as 
-- otherwise expressly approved by Videojet Technologies Inc.
--
-------------------------------------------------------------------------------
--
-- The following entity was generated by the Altera Quartus software.  It 
-- implements a block of embedded RAM with the pescribed proerties.
--
-- Below that is the enitity for the low-end keyboard scanning function.  
-- It consists of several state machines and related logic to continually
-- scan and debounce the keyboard.  When a stable change is detected, an
-- interrupt is generated.  The logic will store all new key stroke coordinate
-- values in a FIFO.  From there, software will read the FIFO contents to
-- determine which keys have changed their up/down status since the last
-- interrupt.
--
-- KBD6.VHD is modified from the previous version used on the low-end prototype.
-- That system used 16 column drivers and 8 row inputs.  This system uses 8
-- column drivers, 8 row inputs plus separate inputs for shift, ALT and CONTROL
-- keys.  The later 3 keys are always driven by a ground.  Their outputs are used
-- as qualifier bits, but are not used for key down/ key up sensing.  An
-- 11 bit value is debounced output.
-- 
-- KBD7.VHD brings in another interrupt signal, kbdio_intr.
--
-------------------------------------------------------------------------------
-- megafunction wizard: %LPM_RAM_DP%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_ram_dp 

-- ============================================================
-- File Name: dpram8x11.vhd
-- Megafunction Name(s):
-- 			lpm_ram_dp
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
-- ************************************************************


--Copyright (C) 1991-2003 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY dpram8x11 IS
	PORT
	(
		clk             : IN STD_LOGIC;
	        data		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wraddress	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		rdaddress	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		wren		: IN STD_LOGIC  := '1';
		rden		: IN STD_LOGIC  := '1';
		q		: OUT STD_LOGIC_VECTOR (10 DOWNTO 0)
	);
END dpram8x11;


ARCHITECTURE SYN OF dpram8x11 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (10 DOWNTO 0);

COMPONENT lpm_ram_dp

    port (
        WrAddress: in  std_logic_vector(3 downto 0); 
        Data: in  std_logic_vector(10 downto 0); 
        WrClock: in  std_logic; 
        WE: in  std_logic; 
        RdAddress: in  std_logic_vector(3 downto 0); 
        Q: out  std_logic_vector(10 downto 0));

END COMPONENT;

signal low :std_logic;

BEGIN
	q    <= sub_wire0(10 DOWNTO 0);

	lpm_ram_dp_component : lpm_ram_dp
	PORT MAP (
        WrAddress   => '0' & wraddress,
        RdAddress   => '0' & rdaddress,
        Data        => data,
        WrClock     => clk,
        WE          => wren,
        Q           => sub_wire0
	);

	low <= '0';

END SYN;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library synplify;
use synplify.attributes.all;

ENTITY kbd7 IS
	port(mclk, Nreset, scan_col_tick, kbd_intr, kbd_intr_flag,
		Nkbd_alt_in, Nkbd_ctrl_in, Nkbd_shift_in : in std_logic;

		kbd_int_trig, key_down_click : out std_logic;

		col : out std_logic_vector(7 downto 0);

		rowin : in std_logic_vector(7 downto 0);

		KBD_reg_read_strobe, KBD_fifo_clr_strobe : in std_logic;

		-- debug outputs

		kbdsig1, kbdsig2, kbdsig3, kbdsig4, kbdsig5, kbdsig6, kbdsig7 : out std_logic;

	    fifo_reg_out : out std_logic_vector(9 downto 0));
END kbd7;

ARCHITECTURE archkbd7 OF kbd7 IS

	attribute syn_hier of archkbd7: architecture is "remove";


	SIGNAL reset, start_scan1, start_scan2, scan_inc, scan_complete,
		col_inc, scanreset, scan_clear, ram1_we_en, ram2_we_en, colgate,
		ram3_we_en, ram_we, ram1_we, ram1_enab, ram2_we, ram2_enab, ram3_we, 
		ram3_enab, scan1_pointer_regen, scan2_pointer_regen, 
		high, low, compare_inc, fifo_inc, ram_match,
		start_compare1, start_compare2, ram_data_latch_en, ram_init, 
		init_inc, init_clr, init_wr_en, init_we, scan1_active, old_noteq_new,
		scan2_active, new_noteq_sec, sec_noteq_old, start_fifo_ld, fifo_ld_active,
		ram_rd, compare_new_regen, compare_noteq, compare_noteq_in, compare_old_regen,
		ram_rd2, compare_old_new, compare_old_new_in, old_latch_regen, new_stable_regen,
		bit_pos_inc, bit_pos_reset, fifowrreq, fifordreq, fifoclr, fifofull, 
		fifoempty, fifo_buffer_overflow, ram_data_latch_bit, ramdata_bit,
	 	set_fifo_buffer_overflow, pos_ctr_reset,
		scan_pointer_update_tick, fifo_pointer_update_tick, ram_read_en, ram_rd_en,
		ram_rd_en2, ram_rd_strobe, Nalt_in, Nctrl_in, Nshift_in,
		Nalt, Nctrl, Nshift, column_0, kbdsig1_del, kbdsig2_del, kbdsig3_del, 
		kbdsig4_del, test_state, mid_column_tick1, mid_column_tick2, test_key,
		kbdsig5_del, kbdsig6_del,kbdsig7_del, strobe_del, test_key_strobe, 
		test_key_down, key_down_click_start, key_down_click_temp : std_logic;

	SIGNAL ramdata, ramdatain, ram_data_latch, combined_row, combined_row_latched,
			ram1data, ram2data, ram3data, ramdatain_latch : std_logic_vector(10 downto 0);
 
	SIGNAL  fifo_data, fifo_qout : std_logic_vector(7 downto 0);
	SIGNAL  rowin_del, row : std_logic_vector(7 downto 0);
	SIGNAL coladdr : std_logic_vector(2 downto 0);
	SIGNAL fifo_pointer, scan_pointer, compare_pointer : std_logic_vector(1 downto 0);
	SIGNAL bitpos : std_logic_vector(3 downto 0);
	SIGNAL keycount : std_logic_vector(4 downto 0);

	SIGNAL pointreg : std_logic_vector(5 downto 0);

-- Examples of Synplicity attributes that help avoid the pointreg state problem.

attribute syn_encoding of pointreg : signal is "safe, onehot";

-- attribute syn_state_machine of pointreg : signal is FALSE;

	constant abc	: std_logic_vector(5 downto 0) := "000110";
	constant acb	: std_logic_vector(5 downto 0) := "001001";
	constant bac	: std_logic_vector(5 downto 0) := "010010";
	constant bca	: std_logic_vector(5 downto 0) := "011000";
	constant cab	: std_logic_vector(5 downto 0) := "100001";
	constant cba	: std_logic_vector(5 downto 0) := "100100";


    
	type fifoload_states is (idle, load_old_pointer, wait1, latch_old_ram, wait_old,
		wait2, wait3, wait4, wait5, wait6, wait7, wait8, wait9, waita, waitb, waitc, load_new_pointer, 
		waitd, waite, waitf, test_new_eq_old, start_bit_chk, reset_bit_ctr, 
		bit_test, test_fifofull, test_flags, write_fifo, fifo_write_wait,
		inc_bit_pos_counter, count_settle2, test_count_complete, 
		 inc_addr, count_settle, test_count_dun, set_kbd_int
		  );
	
	SIGNAL fifoloadstate : fifoload_states;

    type kbdscan_states is(idle, load_scan1_pointer, load_scan2_pointer, 
		scan_init, scan_wait, compare_new1, new_ptr_delay, compare_wait1,
		compare_wait2, compare_wait3, compare_wait4, compare_wait5, compare_new2, compare_new3,
		compare_new4, compare_old1, old_ptr_delay, compare_old_wait1, compare_old_wait2, compare_old_wait3,
		compare_old_wait4, compare_old_wait5, compare_old2, compare_old3, 
		compare_old4, store_wait, store_kbd_wait, store_kbd1, store_kbd2, inc_scan_addr, 
		count_settle, test_scan_done);

    SIGNAL kbdscanstate : kbdscan_states;

 
	type kbdtop_states is(idle, clr_off, init_wait1, init_wait2, write_to_ram, testforend, inc_addr_ctr,
		end_init, scan1, test_start1, test_scan_done1, test_scan1_bit, scan2, test_start2,
		test_scan_done2, test_scan_new_sec, test_scan_sec_old, load_fifo, test_fifo_dun, 
		wait_update, update_ram_pointers);

    SIGNAL kbdtopstate : kbdtop_states;
	
    type fifo_clk_gate_states is(idle, gen_read_clk, wait1);

    SIGNAL fifoclk_gatestate : fifo_clk_gate_states;


COMPONENT dpram8x11 IS
	PORT
	(
		clk         : IN STD_LOGIC;
	        data		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wraddress		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		rdaddress		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		wren		: IN STD_LOGIC  := '1';
		rden		: IN STD_LOGIC  := '1';
		q		: OUT STD_LOGIC_VECTOR (10 DOWNTO 0)
	);
END COMPONENT;


COMPONENT fifo16x8b IS
	PORT
	(
		data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		wrreq		: IN STD_LOGIC ;
		rdreq		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		sclr		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		full		: OUT STD_LOGIC ;
		empty		: OUT STD_LOGIC 
	);
END COMPONENT;

COMPONENT enreg11
	port(d : in std_logic_vector(10 downto 0);
		 en, clk, Nreset : in std_logic;
		 q : out std_logic_vector(10 downto 0));
END COMPONENT;

COMPONENT enreg2
	port(d : in std_logic_vector(1 downto 0);
		 en, clk, Nreset : in std_logic;
		 q : out std_logic_vector(1 downto 0));
END COMPONENT;

COMPONENT pulse_5 
    PORT(mclk, Nreset, clk_tick, pulse_in : in std_logic;
		pulse_out : out std_logic);
END COMPONENT;

attribute altera_implement_in_eab : boolean;
attribute altera_implement_in_eab of ram1, ram2, ram3 : label is true;

attribute altera_implement_in_eab of fifo1: label is true;


BEGIN

---------------------------- Miscellaneous -------------------------------

	reset <= not(Nreset);

	high <= '1';
	low  <= '0';

-- Resync external keyboard input signals to the processor clock.	
	
	row_resync : process (mclk, Nreset)
	BEGIN
	if(Nreset='0') then
	    row <= (others=> '1');
	    rowin_del <= (others=> '1');
		Nalt <= '1';
		Nctrl <= '1';
		Nshift <= '1';
		Nalt_in <= '1';
		Nctrl_in <= '1';
		Nshift_in <= '1';
	elsif(rising_edge(mclk)) then
		rowin_del <= rowin;
		row <= rowin_del;
		Nalt_in <= Nkbd_alt_in;
		Nctrl_in <= Nkbd_ctrl_in;
		Nshift_in <= Nkbd_shift_in;
		Nalt <= Nalt_in;
		Nctrl <= Nctrl_in;
		Nshift <= Nshift_in;
	end if;
	END process row_resync;	  
	
    column_0 <= '0' when (coladdr="000") else '1';

	combined_row(10) <=	Nalt OR column_0;   -- OR needed to get single reading per scan
	combined_row(9) <=	Nctrl OR column_0;  -- since these 3 keys are driven by constant
	combined_row(8) <=	Nshift OR column_0; -- ground.  This avoids getting 8 key actuations
	combined_row(7 downto 0) <=	row;		-- per key operation.


----------------------------Keyboard Top Level State Machine -----------------

	kbdtop: process (mclk, Nreset, KBD_fifo_clr_strobe)
	BEGIN
	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
	    kbdtopstate <= idle;
 
		init_clr <= '1';
		ram_init <= '0';
		start_scan1 <= '0';
		start_scan2 <= '0';
		start_fifo_ld <= '0';
		init_we <= '0';

	elsif(rising_edge(mclk)) then
	
		case kbdtopstate is		
			when idle => ---  Initialize RAM to all '1's
				init_clr <= '1';
				ram_init <= '1';
	    		start_scan1 <= '0';
				start_scan2 <= '0';
				start_fifo_ld <= '0';
				init_we <= '0';
				kbdtopstate <= clr_off;

			when clr_off =>
				init_clr <= '0';
	    		kbdtopstate <= init_wait1;

			when init_wait1 =>
				kbdtopstate <= init_wait2;

			when init_wait2 =>
				kbdtopstate <= write_to_ram;

			when write_to_ram =>
				init_we <= '1';
				kbdtopstate <= testforend;

			when testforend =>
				init_we <= '0';
				if (coladdr = "111") then
					kbdtopstate <= end_init;
					ram_init <= '0';
				else 
					kbdtopstate <= inc_addr_ctr ; -- increment address counter (3 bit)
				end if;
			
			when inc_addr_ctr =>
				kbdtopstate <= init_wait1;

			when end_init =>				-- end ram initialization
				init_clr <= '1';	    -- Clears Address counter for new scan
				kbdtopstate <= scan1;


			--- Start Main State Machine -------------

			when scan1 =>
				init_clr <= '0';								
				start_scan1 <= '1'; 		-- Starts Scan1 - writes data to "New" Ram
				kbdtopstate <= test_start1;

			when test_start1 =>
				if (scan1_active='1') then -- Hand shake with state machine to insure
				start_scan1 <= '0';		   -- start of scan
				kbdtopstate <= test_scan_done1;
				end if;

			when test_scan_done1 =>
				if (scan1_active='0') then
				kbdtopstate <= test_scan1_bit;
				end if;

			when test_scan1_bit =>
				if (old_noteq_new='1') then
				kbdtopstate <= scan2;
				else 
				kbdtopstate <=scan1;
				end if;

			when scan2 =>
				start_scan2 <= '1'; 		-- Starts Scan2 - writes data to "Sec" Ram
				kbdtopstate <= test_start2;

			when test_start2 =>
				if (scan2_active='1') then	-- Hand shake with state machine to insure
				start_scan2 <= '0'; 		-- start of scan
				kbdtopstate <= test_scan_done2;
				end if;

			when test_scan_done2 =>
				if (scan2_active='0') then
				kbdtopstate <= test_scan_new_sec;
				end if;

			when test_scan_new_sec =>
				if (new_noteq_sec='1') then	 -- compare latched row with ram (which ram?)
				kbdtopstate <= test_scan_sec_old;
				else 
				kbdtopstate <=load_fifo;
				end if;					
			
			when test_scan_sec_old =>
				if (sec_noteq_old='1') then	
				kbdtopstate <= scan2;		 -- then scan_pointer_update_tick
				else 
				kbdtopstate <=scan1;
				end if;
			
			when load_fifo =>
				start_fifo_ld <= '1';
				if (fifo_ld_active='1') then
				kbdtopstate <= test_fifo_dun;
				else kbdtopstate <= load_fifo;
				end if;

			when test_fifo_dun =>  -- Wait for FIFO load process to complete.
				start_fifo_ld <= '0';
				if (fifo_ld_active='0') then
				kbdtopstate <= update_ram_pointers;
				else kbdtopstate <= test_fifo_dun;
				end if;

			when update_ram_pointers =>
				kbdtopstate <= wait_update;

			when wait_update =>
				kbdtopstate <= scan1;

			when others =>
					kbdtopstate <= idle;

		end case;
	end if;
	END process kbdtop;

	scan_pointer_update_tick <= '1' 
				when(kbdtopstate=test_scan_sec_old AND sec_noteq_old='1') else '0';
	
	fifo_pointer_update_tick <= '1' 
				when(kbdtopstate=update_ram_pointers) else '0';
	
	init_inc <= '1' when (kbdtopstate = inc_addr_ctr) else '0';
--	init_we <= '1' when (kbdtopstate=write_to_ram) else '0';--- Sets WR active for all 3 RAMs

	-- temporary debug signal outputs
	-- scan1_active_out, scan2_active_out, fifowrreq_out, fifoempty_out

--	scan1_active_out <= scan1_active;
--	scan2_active_out <= scan2_active;
--	fifoempty_out <= fifoempty;
--	new_noteq_sec_out <= new_noteq_sec;
--	compare_old_new_out <= compare_old_new;
-- 	fifo_ld_active_out <= fifo_ld_active;



	tempdebug: process (mclk, Nreset)
	BEGIN
	if(Nreset='0') then
		kbdsig1_del <= '0';
		kbdsig1     <= '0';
		kbdsig2_del <= '0';
		kbdsig2     <= '0';
		kbdsig3_del <= '0';
		kbdsig3     <= '0';
		kbdsig4_del <= '0';
		kbdsig4     <= '0';
		kbdsig5_del <= '0';
		kbdsig5     <= '0';
		kbdsig6_del <= '0';
		kbdsig6     <= '0';
		kbdsig7_del <= '0';
		kbdsig7     <= '0';
	elsif(rising_edge(mclk)) then 
		kbdsig1_del <= fifo_ld_active; 
		kbdsig2_del <= scan2_active; 
		kbdsig3_del <= fifowrreq;
		kbdsig4_del <= pointreg(4); -- fifowrreq;
		kbdsig5_del <= pointreg(5); -- kbd_intr_flag;
		kbdsig6_del <= key_down_click_start;
		kbdsig7_del <= fifoempty;
		
		kbdsig1 <= kbdsig1_del;
		kbdsig2 <= kbdsig2_del;
		kbdsig3 <= kbdsig3_del;
		kbdsig4 <= kbdsig4_del;
		kbdsig5 <= kbdsig5_del;
		kbdsig6 <= kbdsig6_del;
		kbdsig7 <= kbdsig7_del;
		-- ramdata = combined_row_latched
		-- new_stable_regen
--	kbdsig1 <= fifoempty;
--	kbdsig2 <= fifo_ld_active;
--	kbdsig3 <= '0';
--	kbdsig4 <= '0';
	end if;
	END process tempdebug;
	
-- new_noteq_sec	
-- scan_col_tick, key_down_click_start, key_down_click	

------ ram pointers - old_pointer, temp1_pointer, new_pointer

--  Scans Keyboard & Compares each Keyboard Value (11 bits) to 11 bits in RAM.

	kbdscan1: process (mclk, Nreset, KBD_fifo_clr_strobe, start_scan1)
	BEGIN
	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
	    kbdscanstate    <= idle;
		colgate <= '0';
		new_noteq_sec <= '0';
		sec_noteq_old <= '0';
		old_noteq_new <= '0';
		scan1_active <= '0';
		scan2_active <= '0';
		ram_rd_en <= '0';
		ram_rd <= '0';
		ram_we <= '0';
		mid_column_tick1 <= '0';
		mid_column_tick2 <= '0';

		elsif(rising_edge(mclk)) then
		case kbdscanstate is
			when idle =>
				colgate <= '0';
				scan1_active <= '0';
				scan2_active <= '0';
				ram_rd_en <= '0';
				ram_rd <= '0';
				ram_we <= '0';
				mid_column_tick1 <= '0';
				mid_column_tick2 <= '0';

				if(start_scan1='1' AND scan_col_tick='1') then
					colgate <= '1';
					scan1_active <= '1';
    				kbdscanstate  <= load_scan1_pointer;

				elsif(start_scan2='1' AND scan_col_tick='1') then
					colgate <= '1';
					scan2_active <= '1';
					kbdscanstate  <= load_scan2_pointer;

				end if;

            when load_scan1_pointer => -- state decode for pointer select
                kbdscanstate <= scan_init;

            when load_scan2_pointer => -- state decode for pointer select
                kbdscanstate <= scan_init;

			when scan_init =>   -- reset column counter
--				colgate <= '1'; -- moved earlier & then delayed scan for full debounce tick
				new_noteq_sec <= '0';  -- clear here instead of in idle state, since
				sec_noteq_old <= '0';  -- scan needs to end, yet retain values measured.
				old_noteq_new <= '0';
                kbdscanstate <= scan_wait;

 			when scan_wait =>    -- Wait for a period of time, then proceed.
				if(scan_col_tick='1') then  -- The sum of all waits = scan interval
				    mid_column_tick1 <= '1';
                	kbdscanstate <= compare_new1; 
				end if;

			when compare_new1 =>		-- compare_new_regen - in scan 2, 
			    mid_column_tick1 <= '0';   -- sets up compare ptr of ROW to NEW	ram
				kbdscanstate <= new_ptr_delay; -- mid_column_tick1 controls latch of row data

			when new_ptr_delay =>
				kbdscanstate <= compare_wait1;

			when compare_wait1 => 
			 	ram_rd_en <= '1';
				kbdscanstate <= compare_wait2;
			
			when compare_wait2 =>
				ram_rd <= '1';
				kbdscanstate <= compare_wait3;
 
			when compare_wait3 =>
				kbdscanstate <= compare_wait4;

			when compare_wait4 =>
				ram_rd <= '0';
				kbdscanstate <= compare_wait5;

			when compare_wait5 =>
				kbdscanstate <= compare_new2;

			when compare_new2 =>
				kbdscanstate <= compare_new3;

			when compare_new3 =>
				kbdscanstate <= compare_new4;

			when compare_new4 =>
				if compare_noteq = '1' then new_noteq_sec <= '1';  --  Not needed for scan1
				end if;
				ram_rd_en <= '0';
				kbdscanstate <= compare_old1;

			when compare_old1 =>		-- compare_old_regen - sets up compare ptr of ROW to OLD
				kbdscanstate <= old_ptr_delay; 

			when old_ptr_delay =>
				kbdscanstate <= compare_old_wait1;

			when compare_old_wait1 =>
				ram_rd_en <= '1';
				kbdscanstate <= compare_old_wait2;

			when compare_old_wait2 =>
				ram_rd <= '1';
				kbdscanstate <= compare_old_wait3;

			when compare_old_wait3 =>
				kbdscanstate <= compare_old_wait4;

			when compare_old_wait4 =>
				ram_rd <= '0';
				kbdscanstate <= compare_old_wait5;

			when compare_old_wait5 =>
				kbdscanstate <= compare_old2;

			when compare_old2 =>
				kbdscanstate <= compare_old3;

			when compare_old3 =>
				kbdscanstate <= compare_old4;

			when compare_old4 =>
				if compare_noteq = '1' AND scan1_active = '1' then old_noteq_new <= '1'; 
				elsif compare_noteq = '1' AND scan2_active = '1' then sec_noteq_old <= '1'; 
				end if;
				ram_rd <= '0';
				kbdscanstate <= store_wait;

			when store_wait =>
 				ram_rd_en <= '0';
				ram_we <= '1';
				kbdscanstate <= store_kbd1;

			when store_kbd1 =>     -- Generate RAM write pulse to store row value
                kbdscanstate <= store_kbd2;

			when store_kbd2 =>     -- Generate RAM write pulse to store row value
				ram_we <= '0';
                kbdscanstate <= store_kbd_wait;

			when store_kbd_wait =>     -- Generate RAM write pulse to store row value
----				if(scan_col_tick='1') then  -- The sum of all waits = scan interval
----                	kbdscanstate <= inc_scan_addr;
----				end if;
                kbdscanstate <= inc_scan_addr;

			when inc_scan_addr =>    -- Increment column pointer and continue
			    kbdscanstate <= count_settle;

			when count_settle =>    -- Increment column pointer and continue
                kbdscanstate <= test_scan_done;

            when test_scan_done =>	-- test if read of all 8 columns are done 
            	if (coladdr="000") then
                    kbdscanstate <= idle;  -- scan done
				else							
                    kbdscanstate <= scan_wait;
                end if;

			when others =>
					kbdscanstate <= idle;

			end case;
		end if;
		END process kbdscan1;


	scan1_pointer_regen <= '1' when(kbdscanstate=load_scan1_pointer) else '0';
	scan2_pointer_regen <= '1' when(kbdscanstate=load_scan2_pointer) else '0';

	compare_new_regen <= '1' when (kbdscanstate=compare_new1) else '0';
	compare_old_regen <= '1' when (kbdscanstate=compare_old1) else '0';
	scan_clear <= '1' when(kbdscanstate=scan_init) else '0';
--	ram_we <= '1' when(kbdscanstate=store_kbd) else '0';
	scan_inc <= '1' when(kbdscanstate=inc_scan_addr) else '0';

	
---------------------------- SCAN COMPARE LOGIC ----------------------------------

	scanlatch: process (mclk, Nreset, KBD_fifo_clr_strobe)
	BEGIN
	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
		combined_row_latched <= (others =>'1');
	elsif rising_edge(mclk) then
		if(mid_column_tick1='1') then
			combined_row_latched <= combined_row;
		end if;
	end if;
	END process scanlatch;

	compare_noteq_in <= '0' when(ramdata = combined_row_latched) else '1';	

	ramdatain <= "11111111111" when(ram_init='1') else combined_row_latched;

    ramdatainlatch: process (mclk, Nreset, KBD_fifo_clr_strobe)
    BEGIN
	-- process intended to insure against routing delay ambiguities
	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
		ramdatain_latch <= (others => '1');
	elsif rising_edge(mclk) then
		ramdatain_latch <= ramdatain;
    end if;
    END process ramdatainlatch;

		
    scan_cmpr_latch: process (mclk, Nreset, KBD_fifo_clr_strobe, compare_noteq_in)
    BEGIN

	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
		compare_noteq <= '0';
	elsif rising_edge(mclk) then
		compare_noteq <= compare_noteq_in;
    end if;
    END process scan_cmpr_latch;


 ------------------  FIFO LOAD State Machine -------------------------------------------------

	fifoload: process (mclk, Nreset, KBD_fifo_clr_strobe, start_fifo_ld, compare_old_new,
						ram_data_latch_bit, ramdata_bit, fifofull, fifoempty, kbd_intr_flag,
						bitpos, coladdr)
	BEGIN
	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
	    fifoloadstate <= idle;
		bit_pos_reset <= '1';
--		bit_pos_inc <= '0';
		ram_rd_en2 <= '0';
		ram_rd2 <= '0';
		elsif(rising_edge(mclk)) then
		case fifoloadstate is
			when idle =>
				ram_rd_en2 <= '0';
				ram_rd2 <= '0';
				bit_pos_reset <= '1';	-- Clear bit position counter
				if(start_fifo_ld='1') then
    				fifoloadstate  <= load_old_pointer;
				end if;

            when load_old_pointer => -- state decode for pointer select (see State Decode below for output)
				bit_pos_reset <= '0';	--  Enable bit position counter
 				fifoloadstate <= wait1;

             when wait1 => -- Wait for a period of time, then proceed.
				ram_rd_en2<= '1';
				fifoloadstate <= wait5;
 
             when wait5 => -- Wait for a period of time, then proceed.				
				ram_rd2 <= '1';
				fifoloadstate <= wait6;				

            when wait6 => -- Wait for a period of time, then proceed.
				fifoloadstate <= waitb;				
						
            when waitb => -- Wait for a period of time, then proceed.
				ram_rd2 <= '0';
				fifoloadstate <= waitc;				
						
            when waitc => -- Wait for a period of time, then proceed.
				fifoloadstate <= waite;				
						
            when waite => -- Wait for a period of time, then proceed.
				ram_rd_en2<= '0';
				fifoloadstate <= latch_old_ram;				
						
           when latch_old_ram => -- - state decode (see State Decode below for output)
				--				ram_rd_en2<= '0'; -- ram_data_latch_en
            	fifoloadstate <= wait_old;

            when wait_old => -- Wait for a period of time, then proceed.
				fifoloadstate <= load_new_pointer;

         	when load_new_pointer => -- state decode for pointer select (see State Decode below for output)
 				fifoloadstate <= wait2;	 -- new_stable_regen

             when wait2 => -- Wait for a period of time, then proceed.
				ram_rd_en2<= '1';
				fifoloadstate <= wait3;

             when wait3 => -- Wait for a period of time, then proceed.
				ram_rd2 <= '1';
				fifoloadstate <= wait4;
				
            when wait4 => -- Wait for a period of time, then proceed.
				fifoloadstate <= waitf;					

            when waitf => -- Wait for a period of time, then proceed.
			 	ram_rd2 <= '0';
				fifoloadstate <= wait7;					
				
            when wait7 => -- Wait for a period of time, then proceed.
				fifoloadstate <= waita;					
				
            when waita => -- Wait for a period of time, then proceed.
				fifoloadstate <= waitd;					
				
            when waitd => -- Wait for a period of time, then proceed.
				fifoloadstate <= test_new_eq_old;					
				
             when test_new_eq_old =>            
				if compare_old_new = '1' then   -- If new and old byte not eq. then 
				fifoloadstate <= start_bit_chk; -- determine bit position that is different
				else fifoloadstate <= inc_addr;
                end if;

			when start_bit_chk =>
				bit_pos_reset <= '1';  
				fifoloadstate <= reset_bit_ctr;

			when reset_bit_ctr =>
				bit_pos_reset <= '0';
				fifoloadstate <= wait8;

            when wait8 => -- Wait for a period of time, then proceed.
				fifoloadstate <= wait9;					
				
            when wait9 => -- Wait for a period of time, then proceed.
				fifoloadstate <= bit_test;					
				
			when bit_test =>
				if ram_data_latch_bit = ramdata_bit then 
				fifoloadstate <= inc_bit_pos_counter;
				else fifoloadstate <= test_fifofull;
                end if;

			when test_fifofull =>
				if fifofull = '1' then
--				if low = '1' then  -- used for debug only; ignores fifo full condition
				fifoloadstate <= inc_bit_pos_counter;   -- If FIFO full skip write and set Overflow Flag
				else fifoloadstate <= test_flags;
                end if;

			 -- If FIFO empty and Int flag set then assume Processor is completing Kbd Interrupt routine
			 -- and about to exit. Wait for exit (Int Flg cleared) before writing data to avoid possibility
			 -- of writing data to FIFO and not setting Int Flag.
			when test_flags =>
				if (fifoempty = '1' AND kbd_intr='0' AND kbd_intr_flag = '1') then 
				fifoloadstate <= test_flags;
				else fifoloadstate <= write_fifo;
                end if;				

			when write_fifo =>
				fifoloadstate <= fifo_write_wait;

			when fifo_write_wait =>
--				bit_pos_inc <= '1';
				fifoloadstate <= inc_bit_pos_counter; 

			when inc_bit_pos_counter =>              -- Increment bit position counter
--				bit_pos_inc <= '0';
			    fifoloadstate <= count_settle2;

			when count_settle2 =>    -- 
                    fifoloadstate <= test_count_complete;
		
            when test_count_complete =>	-- test if compare of all 11 bits done
            	if (bitpos="0000") then
				    ram_rd_en2 <= '0';
                    fifoloadstate <= inc_addr;  -- End bit pos. test - return to main FIFO Loop
				else							
                    fifoloadstate <= wait8;
                end if;

			when inc_addr =>    -- Increment ram pointer and continue
			    fifoloadstate <= count_settle;

			when count_settle =>    -- Increment ram pointer and continue
                    fifoloadstate <= test_count_dun;
		
            when test_count_dun =>	-- test if compare of all 16 bytes are done 
            	if (coladdr="000") then
                    fifoloadstate <= set_kbd_int;  -- FIFO Load Complete
				else							
                    fifoloadstate <= load_old_pointer;  -- Continue FIFO Laod
                end if;

			when set_kbd_int =>		 -- State Decode. Only set Kbd Int if FIFO not empty & Int Flag not set
                fifoloadstate <= idle;

			when others =>
					fifoloadstate <= idle;

			end case;
		end if;
		END process fifoload;


	fifo_ld_active <= '1' when (fifoloadstate/=idle) else '0';
	fifowrreq <= '1' when (fifoloadstate=write_fifo) else '0';
				 
	set_fifo_buffer_overflow <= '1' when (fifoloadstate=test_fifofull AND fifofull = '1') else '0';
	old_latch_regen <= '1' when(fifoloadstate=load_old_pointer) else '0';
	ram_data_latch_en <= '1' when(fifoloadstate=latch_old_ram) else '0';
	new_stable_regen <= '1' when(fifoloadstate=load_new_pointer) else '0';

	bit_pos_inc <= '1' when(fifoloadstate=inc_bit_pos_counter) else '0';
	fifo_inc <= '1' when(fifoloadstate=inc_addr) else '0';
	kbd_int_trig <= '1' when (fifoloadstate=set_kbd_int AND fifoempty = '0' AND kbd_intr_flag = '0') else '0';
						-- Only set Kbd Int if FIFO not empty & Int Flag not set

	test_state <= '1' when(fifoloadstate=test_new_eq_old) else '0'; -- used for debug

		
  ----------------- Keyboard Beeper --------------------------------------------

    -- The keyboard will beep each time a key down event is detected.  If they are
    -- too close together, the pulse_5 timer  just runs out.  It could be changed
	-- to retriggerable if anybody need this.
		
	key_down_click_start <= '1' when (fifowrreq='1' AND fifo_data(7)='0') else '0';
		
	pulser: pulse_5 
    PORT MAP(mclk, Nreset, scan_col_tick, key_down_click_start, key_down_click_temp);

	key_down_click <= key_down_click_temp;
	
  ------------ Overflow Bit Register--------------------------------------------
  
	overflowreg: process (mclk, Nreset, set_fifo_buffer_overflow, KBD_reg_read_strobe)
	BEGIN
	if(Nreset='0') then     
 		fifo_buffer_overflow <= '0'; 
	elsif(rising_edge(mclk)) then
		if set_fifo_buffer_overflow = '1' then fifo_buffer_overflow <= '1';
		elsif KBD_reg_read_strobe = '1' then fifo_buffer_overflow <= '0';
		end if;
     end if;
    END process overflowreg;
---------------------------------------------------------------------------------




    -----  Data Byte Loaded Into FIFO  ---------------------------------
	fifo_data(2 downto 0) <= coladdr;  --  Keyboard Switch Matrix Column 
	fifo_data(6 downto 3) <= bitpos;   --  Keyboard Switch Matrix Row 

	fifo_data(7) <= ramdata_bit;   	   --  Note: 1 represents switch open
									   --		 0 represents switch closed			

	data_bit_mux: process (mclk, Nreset, bitpos, ramdata)
	BEGIN
	if(Nreset='0') then     
 		ramdata_bit <= '1'; 
	elsif(rising_edge(mclk)) then
				case bitpos is

					when "0000" =>
						ramdata_bit <= ramdata(0);
							
					when "0001" =>
						ramdata_bit <= ramdata(1);	
 
					when "0010" =>
						ramdata_bit <= ramdata(2);	
 
					when "0011" =>
						ramdata_bit <= ramdata(3);	
 
					when "0100" =>
						ramdata_bit <= ramdata(4);	
 
					when "0101" =>
						ramdata_bit <= ramdata(5);	
 
					when "0110" =>
						ramdata_bit <= ramdata(6);	
 
					when "0111" =>
						ramdata_bit <= ramdata(7);	
 
					when "1000" =>
						ramdata_bit <= ramdata(8);	
 
					when "1001" =>
						ramdata_bit <= ramdata(9);	
 
					when "1010" =>
						ramdata_bit <= ramdata(10);	
 
					when others =>
						ramdata_bit <= '1';
							
				end case;
     end if;
    END process data_bit_mux;
	


	ram_latch_bit_mux: process (mclk, Nreset, bitpos, ram_data_latch)
	BEGIN
	if(Nreset='0') then     
 		ram_data_latch_bit <= '1'; 
	elsif(rising_edge(mclk)) then
				case bitpos is

					when "0000" =>
						ram_data_latch_bit <= ram_data_latch(0);
							
					when "0001" =>
						ram_data_latch_bit <= ram_data_latch(1);	
 
					when "0010" =>
						ram_data_latch_bit <= ram_data_latch(2);	
 
					when "0011" =>
						ram_data_latch_bit <= ram_data_latch(3);	
 
					when "0100" =>
						ram_data_latch_bit <= ram_data_latch(4);	
 
					when "0101" =>
						ram_data_latch_bit <= ram_data_latch(5);	
 
					when "0110" =>
						ram_data_latch_bit <= ram_data_latch(6);	
 
					when "0111" =>
						ram_data_latch_bit <= ram_data_latch(7);	
 
					when "1000" =>
						ram_data_latch_bit <= ram_data_latch(8);	
 
					when "1001" =>
						ram_data_latch_bit <= ram_data_latch(9);	
 
					when "1010" =>
						ram_data_latch_bit <= ram_data_latch(10);	
 
					when others =>
						ram_data_latch_bit <= '1';
							
				end case;
     end if;
    END process ram_latch_bit_mux;


------------------- FIFO Compare Logic ------------------------------------

	compare_old_new_in <= '0' when(ramdata = ram_data_latch) else '1';	

    fifo_cmpr_latch: process (mclk, Nreset, KBD_fifo_clr_strobe, compare_old_new_in)
    BEGIN

	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
		compare_old_new <= '0';
	elsif rising_edge(mclk) then
		compare_old_new <= compare_old_new_in; -- a '1' when different; '0'=same 
    end if;									   
    END process fifo_cmpr_latch;


----------------------------------------------------------------------------
	pos_ctr_reset <= bit_pos_reset OR NOT(Nreset);

------------------- Bit Position Counter (4 bit, 0 through 10) ---------------------------

    bitcount: process (mclk, bit_pos_inc, pos_ctr_reset)
    BEGIN

	if(pos_ctr_reset='1') then
        bitpos <= (others=> '0');
	elsif rising_edge(mclk) then
		if(bit_pos_inc='1') then -- count up
			if(bitpos="1010") then
			    bitpos <= "0000";
			else
			    bitpos <= bitpos + 1;
	        end if;
		end if;
    end if;
    END process bitcount;


   scanaddrlatch: process (mclk, Nreset, scan1_pointer_regen, scan2_pointer_regen)
    BEGIN
	if(Nreset='0') then
        scan_pointer <= (others=> '0');
	elsif rising_edge(mclk) then
		if(scan1_pointer_regen='1') then
		    scan_pointer <= pointreg(1 downto 0);
		elsif(scan2_pointer_regen='1') then
		    scan_pointer <= pointreg(3 downto 2);
		elsif(ram_init='1') then
			scan_pointer <= "11"; 
        end if;
    end if;
    END process scanaddrlatch;


    ramwritemux1: process (mclk, Nreset)
    BEGIN
	if(Nreset='0') then
        ram1_we_en <= '0';
        ram2_we_en <= '0';
        ram3_we_en <= '0';
	elsif rising_edge(mclk) then
			case scan_pointer IS

				when "00" =>
					ram1_we_en <= '1';
					ram2_we_en <= '0';
					ram3_we_en <= '0';

				when "01" =>
					ram1_we_en <= '0';
					ram2_we_en <= '1';
					ram3_we_en <= '0';

				when "10" =>
					ram1_we_en <= '0';
					ram2_we_en <= '0';
					ram3_we_en <= '1';

				when "11" =>
					ram1_we_en <= '1';
					ram2_we_en <= '1';
					ram3_we_en <= '1';				

				when others =>
					ram1_we_en <= '0';
					ram2_we_en <= '0';
					ram3_we_en <= '0';

			end case;
    end if;
    END process ramwritemux1;

	ram1_we <= ram1_we_en AND (ram_we OR init_we);
	ram2_we <= ram2_we_en AND (ram_we OR init_we);
	ram3_we <= ram3_we_en AND (ram_we OR init_we);


----------------------- RAM Pointer Registers ------------------------------

------------ Case Statements for Pointer updating --------------------------


-- So far, we did not need this 3 bit decision basis, just the one input condition.

--	input <= new_stable_value & new_old_same & new_sec_same; -- concatinate test bits for
                             		  -- evaluation in case statements.

	-- Note that the format of the pointreg sequence from left to right
	-- is OLD, SEC, NEW.  Each of these pointers consists of a 2 bit value.
	-- This value is encoded into the constants defined above and used here
	-- to simplify the case statement readability.
	-- The symbols a, b and c are abreviations for the 2 bit address pointers,
	-- where:
	--			a = 00
	--			b = 01
	-- 			c = 10

----	constant abc	: std_logic_vector(5 downto 0) := "000110";
----	constant acb	: std_logic_vector(5 downto 0) := "001001";
----	constant bac	: std_logic_vector(5 downto 0) := "010010";
----	constant bca	: std_logic_vector(5 downto 0) := "011000";
----	constant cab	: std_logic_vector(5 downto 0) := "100001";
----	constant cba	: std_logic_vector(5 downto 0) := "100100";


	pointerlogic: process (mclk, Nreset, scan_pointer_update_tick, fifo_pointer_update_tick)
	BEGIN
	if(Nreset='0') then     
 		pointreg <= abc; 
	elsif(rising_edge(mclk)) then
			case pointreg is

				when abc =>
					if(scan_pointer_update_tick='1') then
						pointreg <= acb; -- assumes that NEW and SEC pointer
										 -- always exchange values regardless
										 -- of the compare results (simplest).
 					elsif(fifo_pointer_update_tick='1') then
						pointreg <= bca;
					end if;


				when acb =>
					if(scan_pointer_update_tick='1') then
						pointreg <= abc; -- assumes that NEW and SEC pointer
										 -- always exchange values regardless
										 -- of the compare results (simplest).
 					elsif(fifo_pointer_update_tick='1') then
						pointreg <= cba;
					end if;

				when bac =>
					if(scan_pointer_update_tick='1') then
						pointreg <= bca; -- assumes that NEW and SEC pointer
										 -- always exchange values regardless
										 -- of the compare results (simplest).
 					elsif(fifo_pointer_update_tick='1') then
						pointreg <= acb;
					end if;

				when bca =>
					if(scan_pointer_update_tick='1') then
						pointreg <= bac; -- assumes that NEW and SEC pointer
										 -- always exchange values regardless
										 -- of the compare results (simplest).
 					elsif(fifo_pointer_update_tick='1') then
						pointreg <= cab;
					end if;

				when cab =>
					if(scan_pointer_update_tick='1') then
						pointreg <= cba; -- assumes that NEW and SEC pointer
										 -- always exchange values regardless
										 -- of the compare results (simplest).
 					elsif(fifo_pointer_update_tick='1') then
						pointreg <= abc;
					end if;

				when cba =>
					if(scan_pointer_update_tick='1') then
						pointreg <= cab; -- assumes that NEW and SEC pointer
										 -- always exchange values regardless
										 -- of the compare results (simplest).
 					elsif(fifo_pointer_update_tick='1') then
						pointreg <= bac;
					end if;

				when others =>  -- Default from unknown or illegal cases.
					pointreg <= abc;

			end case;
	end if;
	END process pointerlogic;


------------------------- FIFO Instantiation -------------------------------

	fifo1 : fifo16x8b
	PORT MAP
	(fifo_data, fifowrreq, fifordreq, mclk, KBD_fifo_clr_strobe, fifo_qout, fifofull, fifoempty);

----------------------------------------------------------------------------

------Define 10 bit Output Reg. --------------------------------------------
	fifo_reg_out(7 downto 0) <= fifo_qout;
	fifo_reg_out(8) <= fifoempty;
	fifo_reg_out(9) <=	fifo_buffer_overflow;


------------------  FIFO Clock Gate State Machine --------------------------

	fifo_clk_gate: process (mclk, Nreset, KBD_fifo_clr_strobe, KBD_reg_read_strobe)
	BEGIN
	if(Nreset='0' OR KBD_fifo_clr_strobe = '1') then
	    fifoclk_gatestate <= idle;
		fifordreq <= '0';
	elsif(rising_edge(mclk)) then
		case fifoclk_gatestate is
			when idle =>

				if(KBD_reg_read_strobe='1') then
					fifordreq <= '1';
    				fifoclk_gatestate  <= gen_read_clk;
				end if;

            when gen_read_clk => -- state decode FIFO read pulse (1 clock wide) 
				fifordreq <= '0';
 				fifoclk_gatestate <= wait1;
	
			when wait1 =>    -- Wait unit  KBD_reg_read_strobe inactive	
				if 	(KBD_reg_read_strobe='0') then 
				fifoclk_gatestate <= idle;
				else fifoclk_gatestate <= wait1;
				end if;

			when others =>  -- Default from unknown or illegal cases.
					fifoclk_gatestate <= idle;

			end case;
		end if;
		END process fifo_clk_gate;			 
				 
--	fifordreq <= '1' when (fifoclk_gatestate=gen_read_clk) else '0';	 
				 
	
------------------------- RAM Instantiations -------------------------------

	ram1 : dpram8x11
	PORT MAP
	(mclk, ramdatain_latch, coladdr, coladdr, ram1_we, ram_read_en, ram1data);

	ram2 : dpram8x11
	PORT MAP
	(mclk, ramdatain_latch, coladdr, coladdr, ram2_we, ram_read_en, ram2data);

	ram3 : dpram8x11
	PORT MAP
	(mclk, ramdatain_latch, coladdr, coladdr, ram3_we, ram_read_en, ram3data);


---------------------------- RAM DATA LATCH ---------------------------------

	ramdatalatch : enreg11 port map(
		 ramdata, ram_data_latch_en, mclk, Nreset, ram_data_latch);

    compareaddrlatch: process (mclk, Nreset, compare_old_regen, compare_new_regen,
								old_latch_regen, new_stable_regen)
    BEGIN
	if(Nreset='0') then
        compare_pointer <= (others=> '1');
	elsif rising_edge(mclk) then
		if(compare_old_regen='1' OR old_latch_regen = '1') then
		    compare_pointer <= pointreg(5 downto 4);		-- Point to Old RAM for compare
		elsif(compare_new_regen='1' OR new_stable_regen = '1') then
		    compare_pointer <= pointreg(1 downto 0);		-- Point to New RAM for compare
		elsif(ram_init='1') then
			compare_pointer <= "11";
       end if;
    end if;
    END process compareaddrlatch;


   ramreadmux1: process (mclk, Nreset )
    BEGIN
	if(Nreset='0') then
		ramdata <= (others=> '1');	
	elsif rising_edge(mclk) then
		if(ram_rd_strobe='1') then
			case compare_pointer IS

				when "00" =>
					ramdata <= ram1data;

				when "01" =>
					ramdata <= ram2data;

				when "10" =>
					ramdata <= ram3data;

				when others =>
					ramdata <= (others=> '1');

			end case;
		end if;
    end if;
    END process ramreadmux1;

	ram_read_en <= '1'; -- ram_rd_en OR ram_rd_en2;

	ram_rd_strobe <= ram_rd OR ram_rd2;

--	ramdata_reg : process (mclk, Nreset, ram1_rd_en, ram2_rd_en, ram3_rd_en)
--	BEGIN
--	if(Nreset='0') then
--		ramdata <= (others=> '1');
--	elsif(rising_edge(mclk)) then
--		if(ram_rd_strobe='1') then
--			if(ram1_rd_en='1') then
--				ramdata <= ram1data;
--			elsif(ram2_rd_en='1') then
--				ramdata <= ram2data;
--			elsif(ram3_rd_en='1') then
--				ramdata <= ram3data;
--			else
--				ramdata <= (others=> '1');
--			end if;
--		end if;
--	end if;
--	END process ramdata_reg;


------------------- Keyboard Scan Counter ---------------------------

	col_inc <= scan_inc OR  fifo_inc OR init_inc;

	scanreset <= '1' when (Nreset='0' OR scan_clear='1' OR init_clr='1' OR start_fifo_ld='1') else '0';

    colcount: process (mclk, col_inc, scanreset)
    BEGIN

	if(scanreset='1') then
        coladdr <= (others=> '0');
	elsif rising_edge(mclk) then
		if(col_inc='1') then -- count up
		    coladdr <= coladdr + 1;
        end if;
    end if;
    END process colcount;

-------------------- Column Demux Logic --------------------------

-- Used for simulation runs only.
--    col(0) <='0' 	when (coladdr(3 downto 0)="0000" AND colgate='1') else '1';
--    col(1) <='0' 	when (coladdr(3 downto 0)="0001" AND colgate='1') else '1';
--    col(2) <='0' 	when (coladdr(3 downto 0)="0010" AND colgate='1') else '1';
--    col(3) <='0' 	when (coladdr(3 downto 0)="0011" AND colgate='1') else '1';
--    col(4) <='0' 	when (coladdr(3 downto 0)="0100" AND colgate='1') else '1';
--    col(5) <='0' 	when (coladdr(3 downto 0)="0101" AND colgate='1') else '1';
--    col(6) <='0' 	when (coladdr(3 downto 0)="0110" AND colgate='1') else '1';
--    col(7) <='0' 	when (coladdr(3 downto 0)="0111" AND colgate='1') else '1';

    col(0) <='0' 	when (coladdr="000" AND colgate='1') else 'Z';
    col(1) <='0' 	when (coladdr="001" AND colgate='1') else 'Z';
    col(2) <='0' 	when (coladdr="010" AND colgate='1') else 'Z';
    col(3) <='0' 	when (coladdr="011" AND colgate='1') else 'Z';
    col(4) <='0' 	when (coladdr="100" AND colgate='1') else 'Z';
    col(5) <='0' 	when (coladdr="101" AND colgate='1') else 'Z';
    col(6) <='0' 	when (coladdr="110" AND colgate='1') else 'Z';
    col(7) <='0' 	when (coladdr="111" AND colgate='1') else 'Z';


END archkbd7;
