%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_method=rsa
%%% protect key_block
SsjfE8XxZlfNb/NT05/qnu4Dd+u6OVyWw0B2Y9DjTKWTyzKDCjyYUOuE4EJyX2gPaoluhfHCsKEjAU+8vIGyMkYKyDBe7DIfUTtx9JMw9MyXqx4pYK7d2ScYkuBA6fNfp3sCB3/YJluOHuXEKOFLgfaPmrIR2IMvlAmwQE3KVOj78vPxgAqgtuDZ+q38HnJvZyKmCKoZqpTfhV1EJkf3nZOvkXZ3nGSAmBJp5Mccx0pPMm21KaC5+gdC/CcHte8aK4+NrQZcrNsWSAVYSXsv5Yz8EDV/mjg339V6UMIruoFsOQbuNybaFfjYzrxvRmAVD6HnXETgnvOBXK63WSJ2Hy==
%%% protect author=Lattice Semiconductor Corp.
%%% protect data_method=blowfish
%%% protect data_keyowner=LatticeSemiCorp
%%% protect data_keyname=lte_datapath
%%% protect data_block
tIJeCh/F2NAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsAyrlX0gor6tVKtg7aPDoVB3ByGK/VBOniK3a0yLM5mRQQDm0+FyW5cCrRrGz4N4qPFHzx41G1TX5KcFXXGVwNLFN64LgH5CMAyrlX0gor6tNzUEBQoLQ8H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC4kq3srN7+p8pYtFYwwZhWqsyMGi2gKJIToC639UCAtrpWuXtbdXdq/CTJmvKVExS6nbMVREOZFXX7FJuNkvS4F3yRFNELvN/RfBjge+BTkeL6VzlnGc/+S3a0wy44Ms6JA0MhusifFfriGawGO8GqSUbYzptWFRza6Jxq/NewlqMHl3CYoq3QYm/MXoS8jXO8MRFxW0sPFOLWt2Yt/8Gl8qSTHFiH1kTCqQ+hVhIitbxlBn6uUFJLTfQ5erSelw4OXh7EFjYzOwZtft2qgKkqdvQUyhBqn1GkqbmLtngTq+UAnTvq7uXQisIturjZfZOBNa91oqLi39bpJBPqqb6wdeJayjcn3gyYma9s1iOOrpjAE9+MWUwntRXogseZtwmfwNKRm55vIEtKqHu2CSdDtVYycmWZhaXVxRPQDZoVN04h/FG23lS/anr5lh1ouzFM0Ac+YVBs5zFlXGHWUlNRC17beq/m+CEpnmH7dxq6r+KX0DdpkLh6mJPjRr0jh/uxGa4TM8NBEjJEsgFM1hTLE4wFWY4OAFkxVzPHOsvPGs/9lwpWOYitytNe2hTN8U5JW+oLGHK1SV/4cIAducePjNZbtkU1JgtRYCUJz0CJQrwgDn6YE2issSXVqVgAVEUF1qjFJUHWvH5bq5w1SPcLfX/o+2eMA2lC671jZPPTfIERaBBzAvnjcm2utZi+wc2R+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC1pURxGQczVlcLpMDZXOk/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwt3gjIEtmkGJUn/JVTdmWYH6MQhTMtwAUK7cvUi1o/TGoQ1R4UUhLal0nUbGM+SWQTJ5r1xzfDXClC+R9yUfoJ0Gb8Ye9mOhQPlT58qADgnayba61mL7BzZLgSgz8KdKfq6G1G9T48ue8LT3JSAFfVg2jmz4lCH4bEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsvZXzvFjDk/E8jCmrTA34ECueWGoonK3GY9BCSCKyXy1idipxlUuI0S33hUU5oIdEEWH4+LwrdSY1qeF/3xLYVZd6RBKNM6Eip9JBxvAjUFxuqimyh3chzS/77koXJE7AV+wVeeATG8+xJbku+DGjG1qOiGQvRf+TwELQPrOCdhhVKl4Jhni0OKly64myqQ5ES0xiBngYr5XiBFjJ+vOQ+LCcdI1c8QA76xKl+nv/xy6Sx/H94hLTY1ph9EJwygYpsFvYoh5TYxtaYfRCcMoGK9ovv3izTod5K+W6keJ03eG6rEFd7QSuNKly64myqQ5ES0xiBngYr5XiBFjJ+vOQ+LCcdI1c8QA5kHQ5ddmeoBYwV5wNiRJ/ZDPbkBzQdmF4GMmRgScitOVcQF0znFJaHrmeXx2d9TysWVW0lhSZI/BRw56OPkg/Sr4YFewe2llmZ66FqCFbUCzpEo49KB6oCDhLedypjXa3Wo6IZC9F/5Fldw/XOl282BqbfOJJ3OrAU5cw5MiWQAd13JG6BZzlTZ4itJqwS47yoz5Qt65ma3xO7Gfeo0MjEzI4C2OHqUZL2+riRMkQMuEwe+YWZZrOl46FnwlZdCSgU5cw5MiWQAd13JG6BZzlTZ4itJqwS47yoz5Qt65ma35p2odmtdTjYf5Lu66NXfxHWo6IZC9F/5KMoSqOcxZ4FzHV0f9xyNDjWJsSfx9OMCW3gjXOEok0SYW10OsWEUi9pizNGOcBESL4RbG7OXtJWreh8mIljtYPUQMX56yVAEuysWb8bvfkBGKFCf6+tQ+EGpt84knc6sBTlzDkyJZABwctBB7RV8e/g/0d+fL3g8YRhYKpgEmx9HQ8wFO/M7GW/me1x9h61evPd/Y2AL5TevE/MsZ9IBFfS4GZUdz+Zlq0Lj2lFxsKTbMnQlCZwBr2uOTBnkKfyaMCQeuDZHbLsJu/um9PrknouMa06uX55ehZVbSWFJkj8RiUBsRRrZezjoWfCVl0JKBTlzDkyJZABwctBB7RV8e/g/0d+fL3g8YRhYKpgEmx94KIxjBb7VISt6HyYiWO1g9RAxfnrJUASNXJgNi/c0jgGpt84knc6sBTlzDkyJZAB3XckboFnOVNniK0mrBLjvKjPlC3rmZrfE7sZ96jQyMTMjgLY4epRkvb6uJEyRAy4HPUIn0+NIcPYg8PKAP8lICp/YNXMMo+zDzAyIDd8ANpZoW/GvRb062mLM0Y5wERIVXa5ZfbCiuiHSutWIY+S0iwnHSNXPEAOKqejPHy7NHQd8sYoPw3z5JKHozjh0OSjzlRNGHp1OjPUJ7+7dTW2IAS1GUT/Suh2wJB64Nkdsuwm7+6b0+uSei4xrTq5fnl6FlVtJYUmSPwXkZANSEarGPxVKcyA/TL/1ibEn8fTjAlt4I1zhKJNEuEx/UufzCpLWlEx0cJjq1IS0xiBngYr5X+S7uujV38R1qOiGQvRf+RUtXGBgtkskKGY8Sonln5ecKKzspNYOJFNz7Ynn829T5G7yIHZVSLdxj2xuG2LhpZsFvYoh5TYxlM2bu+WFHT1Vg+UOWjJwK7tugxD2QId+S5ZPPacqIdUrIQIzWFAzziWLd95iKP6KRO8bfwEMJbFLlk89pyoh1Q+b9iDlAwW6GzaUnbp7B7W8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9mAXBJjTEirtO+XpO/51g8HWK8opvpitytZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkxeZMP5Ziang59RsG3YsO+QDpz23nyyck0YNHhdfKXcBbcmCydlEwqDfEUpIDdRqEB8pWXSZSj1O0kfhGIVJ+sqJsEbX0JalsIP99gw1gQgWqDXxlkXGyt+Ze7uy/i2WPQRM5a3QoG6c/gWHRCvm82pAFBpperUxu1eN6cKE8PL2ajkcM0HTJMWiAiNHs4agN/b6uJEyRAy4gMjCLCS/c5twIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk5ObRzSM0cQs8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEdvF3B3A6aoB1e0P0BJnYqhlJH4Ity3OeXLPGMpkOr+nPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx8939jYAvlN5uJENWVgUTMCccP57iyXMCHZIVgGmGPplkLbvqjM5nGQVI8CB0DIrjJ6b+11OiNzEAGkuTHgN5IEc1LYXpf5P82K6hMdSPTRxAFBpperUxu1LGkp384+Kj1i5t3ireDk+Rx6G6Y3CZNbii90ZSwmGhgz5oQLaYuGZrHszq1lh4rjbQpprNa4fn+sSpfp7/8ctLuRgyX6MnyvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk2wB+7h+Ops6cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM4gYI4+CnS6Q87gw/X+LIlG7mKWiqxBZI6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUctajohkL0X/kwj/ltX+8gJ4QhXX1FYfhX2w7svVw9oCOK0RjtJINLBLTVr8ikO3n6QNccOO/XLE6ACDwf94yKK4wynzEPEEV7Q4S3ncqY12tJ6b+11OiNzHGyf/zw7r0uC0j3r0EOM4eEJ23uxQ2QhqNMp6W7hWfPoZDoeS7S0Oc4Lwn2kgjW7dC9k6h5Y71X81lmcYIz62/qPYQEx3C56YYa77f8vmAHaRmk52OiAavoQcjBsP0HrSDKkvY++Zbwb6IhgkZZbtUVEbpeCnAPqBm1/WBNgQD87Hw9Ya4xpPW8Xu6CjZDTW2CUGnKO+XO3RZVbSWFJkj8mRd8k2q1hq06JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcjI9RKJpATlw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/Hv/ScZwIEtcwp2udCckVWEWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMXmTD+WYmp4D+60Wnki7pOv6rlTyE6svQFCuQ94pGXg7qOyDGL4z8pCWjtIDJjfhO9XTEYfeTIji8V8b58GG7aG1QhNxWUqndD+L1J6e9gnwVkL6lrP3Ai82wOMSIWNIEvYcLyVDJh9h68GeGPd97Abo6pi85pwqtNZKzY4pJfX8xBPmd3IyJn0uQRHxqQ8BZFU8UVcBXwAuYiqiWWtCZqQBQaaXq1MbubM/2Rj+cdugBKVBuglOW+ax7M6tZYeK7HVbaI9yUfqqiElkWPOTuY/OZUX9y2RFcgCkD7Ytwz0DbQpprNa4fnZB0OXXZnqAUcHhx5xnkZgnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR97XL1oK/jHfF9J8j7SYid2/ZNayljPTQfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8yL325+3J+sFlVtJYUmSPwUcOejj5IP0q+GBXsHtpZZmeuhaghW1As6RKOPSgeqAjUe9kkxijWfP+uWm9UhzbEfUxVuCXS5Y5cRiFXk5lH5QWLmVx0vBuU3AAYs20Uay36xikhqd3RcZji/ODKCZ180YXyVXWerMNaYfRCcMoGKfID8LDeXPCoZVduYZlaoCgo2jp1ruGht2K6hMdSPTRwZW38nhD0S7p1+11Tf6mJKkNEPMoCb13phZozdt25vcB+pBQUd/IzhcfToHZ5ByWeUPQ5KkdgkjMDBYzeHuk3SM1ILnQKCFfPz3f2NgC+U3rxRLu0XWMpK6BphuFXO8gny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+To4dhv1qMaw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9nzVgO1RRXmAASlbnNB3Y0l8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEf2+riRMkQMuEwe+YWZZrOlkoejOOHQ5KPOVE0YenU6M9Qnv7t1NbYgBLUZRP9K6HbAkHrg2R2y7Cbv7pvT65J6ULPvvK7PC69RpeXrPc92ZGrlJlIW7JGDnMQvunqozFDGPbG4bYuGliVZc0BIPe+mSRsolPlb3m5RpeXrPc92ZEXlAuVY+wJdzh509K8ZDkar73Isr9tVv4YN2vW5rDpG2HUbSjO/lROTsRdHHlLuegKAWAUt8Nn7NWYnM+lVTISe0ux4QFEQFLhO0R4gvDoi4cMmgMS30D0bmKMy8DBAMqjV813ehqxtJeX0C8xw+w81Zicz6VVMhOL580Ku4o0cNyPPFFXDCrVr0IpCVjxOwtfzyeLG5RUgvCjy3WV9golDPcV+8IRxTEydRzqij1whbuUxToA3iR1hdlLCHWbufkvT0GdGV6gL2fWwA4yVPNerUxF/KHyDoOjqSFmk3zYp0fsaZDC8Afknz76s+NvFevXsWtrJKq4Ml72uaVM7kctr4ovML7SUr0od6lH+0tGho+vy87Qhp/sw0mP3skyStAVQO2qyBK5ZZofMwHrUCMVAFBpperUxuwGznUfbr9n6BqGVcD+0rY50cRI00EQFLfgAboRs8l9qWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmspIqjZ4KdmCy6W0OuJKSNlM2bu+WFHT1t6Z8lyqB3GtwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkywnHSNXPEAON8CYNU16QSihmPEqJ5Z+XnCis7KTWDiRTc+2J5/NvU+Ru8iB2VUi3cY9sbhti4aWbBb2KIeU2MZTNm7vlhR09QHYTm0EAuqWOMKA1BJV2ZOK4S462vJR2uEx/UufzCpLv3T+/Q7PTTl782x0Hz5p0SdtPUJet6W/OMKA1BJV2ZPCFVAlm/B5ypzEL7p6qMxQxj2xuG2LhpY+cf6JceQfkH5RcNB0Y414IKLVRP+gR5DFldxS0KnQs564K/wQvn7OKhA+sNVVs3E3I88UVcMKtWvQikJWPE7CA1xw479csToAIPB/3jIorujqSFmk3zYpQcj1oMvj/BObX0PIDZBZLNTEWtiGVkNRHEcuJ+RvSwbcckoVRMuvumRXZEp4UN23tnUuFoUtsdADhU75otEOOxuNFnTiwyZmlArXMaWD0mMw96eqkUwxp5NMii1sPd31YcVURn/Kv+qtX1L25Mc6zZfc7WVs9nmeUQlm3kjqGg3mJGcwwwWk+7QR9MkxrqogmvBLVs07DaKtTcTiRY5uTTjgq5bS0R062Hcxa4XBoETvlas30N2OIbHw9Ya4xpPWCoKkBwTO4RWdlAok5s4rKowe9+D+FNx6MbpURTIzzpZwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk5ObRzSM0cQs8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEdx6zntlvw61+8cZztlcmOkdHESNNBEBS3Oa3aSjowxtvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx8939jYAvlN4PFNV1xWiLU+tgJtISb6v6koejOOHQ5KPOVE0YenU6M1Znz26sJMu7NrBKvbSWGzh1ros83AXh2nYzi4h7qnN8AdhObQQC6pY4woDUElXZk4rhLjra8lHa4TH9S5/MKku/dP79Ds9NOXvzbHQfPmnRJ209Ql63pb84woDUElXZk8IVUCWb8HnKnMQvunqozFDWmH0QnDKBihFlpWoLRMoV5bpT/tkBZNQOA8iS2QMlvf7rFS/YCcMmp09XPYzEI6LPVIHPSNemf9z9wV7kUOSO9bMpVXuOVT9YggAh2zYxKrOm4GNjZXJtIKLVRP+gR5D+E20KsWCsj+p1Yg9VOK0ooXGvPCY6toFYggAh2zYxKrOm4GNjZXJtIKLVRP+gR5DtEgXdQXEbmCNZ2jA6uqcZr4ePFoHgHvgBq8OYNNE4kSHtmpgoIVG9S9ktXJmTRafPyHEDU6aYFCGsk4fQlnIs22RPOjd1Wncw0mP3skyStFRWHJYQ/HeH5v3z4BoloQPZPhptMRKt7jEfL8or/UgqxaL58fFmwD5je6gc3gi9wHMETKfbOj03oe+eSd+ASXXwjJg8usv7SsMiO/n7dyRrLm7LTOpN6IrVezX+/1O8veuXOdiXA4/o4SSlnUTC2Qg42Me5quvq0vXFawSPwn81vmgjkm09k5bCzY5w6IKJWujqSFmk3zYpXJcgOF5iXjhyinP1PwyLrOL580Ku4o0c6PGVuhZTck4MK41UJTu/SpKpq0ectclzEfaEaaVB8n4lUIzcVNuR9/sS+mV6bOK8RN7coAtNOaScofEdYXXbBrJtDR8wyWEqqDXxlkXGyt+dlHXYVfdTkVHM2yVOm3MlBEzlrdCgbpz+BYdEK+bzakf0KAuwLMe8Y9H7UTLSrNo03Omv+l8qHUTe3KALTTmkfDi9IlOSviSfm2aPk+DQ3i5JNQbS9Kln3URzjzJp067j2grARZwQ4hSJrXT7TbAS8jfGqseA0SqXdToO7KQt0kr15D2mwrLWYob7wXVXN80Ql5U7vYUivVSswSnK9VcWVJu9hEbmsEHj5RcgwgjQhTQp5xaLaiGlKA//vtqa/HWRarXObm18SpTM4+MW9kctkuS1mgx2ReqT/su5/Z/5bcLNjnDogolaeMICCqyxpgTOfv8bha5Tti9nAOXMoiDEQvZOoeWO9V8EtZlyUyk3a3EK95r9tEWszlQhkJuH3ClUQvxTMwUD+rbfULmuke0DhGYkdUTkyweoNfGWRcbK33eqkj2k9wy59nPA40Hoxh+bSVormCaLsMkk0V06BxHN1JlOQ1p7hKXOQsr7ApO696g18ZZFxsrfx1W2iPclH6qohJZFjzk7mBD0ExRs9ghb0uwTtBtpz0SwpGBD4G1Yc5fKlaij9lr/Yob7wXVXN82VtLSIlgruvy8QB0k6Z5z9fBOCByfhll3/U30/DvApyDJwqq0pLPf5Lx0KNW8GR0iDomWkfWEta/XsWtrJKq4MWFNijlx/13A/78RUp/uizbl1ldhQw+Y3NEgk0Xpg0PDhhQd5G/Xq5OYiqiWWtCZqlA3m4ke0h7AxDEQ14u2USDQ68/3TNPUeGmM340wuvpGzpuBjY2VybWo5HDNB0yTFAoHnaArgPt00CwarNCE7L2ouaB4FXMSJwZgHw80d0FyWD+M7jr76jvx8qk47WgppoqIdLq2gfy8KY7iD29xKuQRM5a3QoG6cNv1C5IcM115gp3oNnw3RHXDLvEmaOuprPC7n3244wpk20KaazWuH5+JGv3ZDsRT7SnzTo33N4Er7iNLGpBz65fL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk2wB+7h+Ops6cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMjmJGmnDlH5Y2zKMO9BcVGyhjpcragxsOXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZtRAxfnrJUASQjgSq+42WaeK49tLLbRTxCp/YNXMMo+ztCYYJvd31+JpkvUKCEqQl6jPlC3rmZrfE7sZ96jQyMSAogKCi1mhFJ8LjLxV4aFo8nr+ei788bGj6/LztCGn+zawSr20lhs4bGgSEMsSQH9htPbp57vxxZ8LjLxV4aFo8nr+ei788bFoq3EIk8EtRyBkfl83H8VOV/I5oZBSb5slUIzcVNuR93Xr+PkTzya0MHRKiVWorhuZW8Gn8vZC/bE6/8NUMa+/msAgkAG5f2ej6/LztCGn+zDSY/eyTJK0VFYclhD8d4cnejDXJspPjJEN/e+4dvrvRqd42lmOPEPCCD8Qa/jQUObV9EPoBEz3VFYclhD8d4cnejDXJspPjGxjXDZKiHt3VDJ2qFMJOwGawCCQAbl/Z2ircQiTwS1HNp+ipJFgnO/C4OEyxUpTDy8V8b58GG7aakY/FF8AzWiOlDRqsyXhhQa/k5mtKf0tjl6qMQBreSbxDac8D3GtNToxuWMoEH3sPL/sSLuLBfTLApOQol6t3+L580Ku4o0cQ7DbMqsIswCj6/LztCGn+3EK95r9tEWskYxlJQ1vSfSCk1ezLNPwKGDg+W9R36aPqDXxlkXGyt+dlHXYVfdTkf9o8oOEEXMG1GNCSUw7966SqatHnLXJc+iPsIb6KJrZ9xikmyUKNrNJYhE/0QKEvcINnKKON5bzntLseEBREBS63iLFularIZ8A84lnmGTMq6mJ4B7GgmZxisOaoSCGPrEddF643SlECoKkBwTO4RVKNFsMVU+AuxUjqW31aQvzqXz7T3JZ9rjZPhptMRKt7pQ30dN/N5xBCdjN2EKA1FDwlfaMSUKA/M8CDbHYXDumaktTFvAbh44VjKY+ZWouQ9a++NL1ZZOQdQVtBqkwhRajIXoWCtX8ZEaneNpZjjxDZSAvcTbQPR9ghAz2KDowHHrWMIpBrA1QRN7coAtNOaRf6xMSxaklGp+bZo+T4NDe4OfE/m2jeCcKgqQHBM7hFUo0WwxVT4C7Trol1QmPg0Z/F8tPnMoYuK8n4nHtlKBlQ/NL6qMs778MoY/p6Q9WXIM+aEC2mLhmax7M6tZYeK6x8PWGuMaT1gqCpAcEzuEVnZQKJObOKyqMHvfg/hTcekI4EqvuNlmn/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNbwb5RoGmEZTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyHX3S639fwE5uM7mYuvgPmoVq81GdeMIoLWE+J/CFJL46JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUctajohkL0X/kT3Eqg2+sX1fetIEggrRU2NYmxJ/H04wJbeCNc4SiTRJhbXQ6xYRSL2mLM0Y5wERIvhFsbs5e0lbnfJYL4GyuiJrs6rcE5ddzG6h96qoENi0lUIzcVNuR9yBkfl83H8VONL6qjRMpM1v7xMVeykU9PJrs6rcE5ddzG6h96qoENi0ubstM6k3oivawMr5DqsStWWIE7b+X8v6e0ux4QFEQFNdTKUFHOYgB9o/Dy0NcnK4gotVE/6BHkMWV3FLQqdCzKgE7/Wg2oF8lUIzcVNuR9zafoqSRYJzvwuDhMsVKUw/+6xUv2AnDJtOzjAXFxvcUl97XTDoneesqATv9aDagXy5uy0zqTeiKuE7RHiC8OiLhwyaAxLfQPSem/tdTojcxNuF9Szb8bc8e57RD9aSuRb/4fWEjYA+4NVFi3rYRA4AeL+Nz/rOr6LnwzU+G8vcN33gJ70sm/+NqPwv0nP0sPyXl9AvMcPsPg5KHxlT5WSIlUIzcVNuR9zafoqSRYJzvryfice2UoGWnNOR1VEMsPXIn7VbSoM5uR5yUa6qpw2AzUgudAoIV84Q4FE3t1NdWOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHdpsyj1Cur7DQFURKM+r0PEZ8qp5acqR9YioH+dNlQhry/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR/b6uJEyRAy4/XqXE5gXOKv+Cp9jwX0mA9YmxJ/H04wJbeCNc4SiTRJhbXQ6xYRSL2mLM0Y5wERIVXa5ZfbCiui2tqhYUB7+BPq6OCYUYhVgTc+2J5/NvU+/paFmRb2SaWN3V2MCtXJ08xEJr05kfCqh7LJLT39acH5RcNB0Y414Tc+2J5/NvU+SqatHnLXJc8pJ7Grijx5007ZvP/PYbvGhnqiQkZnUWTyAJ9PHzeXvkt8vesj/3ckh7ZqYKCFRvYGffOuD9aSmQcj1oMvj/BPc/cFe5FDkjvWzKVV7jlU/WIIAIds2MSqzpuBjY2VybSCi1UT/oEeQCoKkBwTO4RVDbVXqhBiWBiGsk4fQlnIs22RPOjd1Wncw0mP3skyStFRWHJYQ/HeH5v3z4BoloQPZPhptMRKt7jEfL8or/UgqxaL58fFmwD5je6gc3gi9wHMETKfbOj03oe+eSd+ASXXwjJg8usv7SrQR9MkxrqogivQjeGQ1Z4QmxL5kTsVGAq1NxOJFjm5NOOCrltLRHTqmwc/MfC2LfpQ9DkqR2CSMdY1jTjDML4h3YPzVvainmEx9tPmLwgRlkxABqgeVZ5ry/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiZ0kzHopDoC3Lkwh3dD2oRE8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/Hz3f2NgC+U3l9v0LT2OLyvkoejOOHQ5KPOVE0YenU6M9Qnv7t1NbYgBLUZRP9K6HbAkHrg2R2y7Cbv7pvT65J6ULPvvK7PC69RpeXrPc92ZEXlAuVY+wJdzh509K8ZDkar73Isr9tVv4YN2vW5rDpG2HUbSjO/lRPET/gv9cMW9dB+DvHKS5GYWaFvxr0W9Ot7A827fZ/94YYylKdDZ5Rs2HUbSjO/lROTsRdHHlLuegKAWAUt8Nn7NWYnM+lVTISe0ux4QFEQFLhO0R4gvDoi4cMmgMS30D0bmKMy8DBAMqjV813ehqxtJeX0C8xw+w81Zicz6VVMhOL580Ku4o0cNyPPFFXDCrVr0IpCVjxOwtfzyeLG5RUgvCjy3WV9golDPcV+8IRxTEydRzqij1whbuUxToA3iR1hdlLCHWbufkvT0GdGV6gL2fWwA4yVPNcycLNVmspuhEliET/RAoS9phE0HWhuiJue0ux4QFEQFLreIsW6VqshnwDziWeYZMzZ69vQf60huQ0RUQQFakJD+fu3S3MoLDCtX1L25Mc6zYVTiGXHOnHGAodA/dD5hHsByVASsWw8eNWiqZnaehAmgGwFmQkytbiowJ6U1UDbBc4edPSvGQ5GoZ6okJGZ1Fk7ZOEinR1yI+YiqiWWtCZqRqhT9zYkEL5Gs0INCZgPqpzAiNYJyQuINAsGqzQhOy9qLmgeBVzEie+VqzfQ3Y4h1i5t3ireDk9K9eQ9psKy1iXl9AvMcPsPg5KHxlT5WSIubstM6k3oirhO0R4gvDoi4cMmgMS30D2DPmhAtpi4ZmsezOrWWHiusfD1hrjGk9YyBdfreKUHqvDqITd5qHgol1o8dKovrKRZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk1vBvlGgaYRlOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHKmevqGssw+r2tm9VWt6ZjYcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMsJx0jVzxADujz8jlDsWTRMlMoTQR8oTGHSutWIY+S0sRP+C/1wxb1HLNm3JqNigKr73Isr9tVv0oqZTsfwuk5KykLxLUCU+pQs++8rs8Lr1Gl5es9z3ZkReUC5Vj7Al3OHnT0rxkORqvvciyv21W/hg3a9bmsOkbYdRtKM7+VE8RP+C/1wxb10H4O8cpLkZhZoW/GvRb063sDzbt9n/3hhjKUp0NnlGzYdRtKM7+VE5OxF0ceUu56AoBYBS3w2ftTNm7vlhR09doJHToildnuAT+C4N5bcirsY21T3uRMTTB0SolVqK4bmVvBp/L2Qv2dlHXYVfdTkeOhZ8JWXQkoSCiDkMrkG5MGg46/2mOgtjjgq5bS0R06bUXfYiX6zhTSR+EYhUn6yme31JapRDb5qqmdnk+XrXCgAN3cKhu7CypXQNWliz1950zf1hEgFpZcWonor9aLdBqh3FPNHl8IJb53+keb6tRoq3EIk8EtR1o6zbS+gixVQQ7dOXKu15bYrqEx1I9NHOy6HZ2gx4ddzwINsdhcO6YlBxxtJgi6DUr15D2mwrLWJeX0C8xw+w9/VE+0/jpYRj/Nb4tQS9QVLm7LTOpN6IrHRNnd95WGxPcaLydpsQM04vnzQq7ijRz6dpx44IiSf6Pr8vO0Iaf7cQr3mv20RayRjGUlDW9J9I+p5o2nQMwYmvDvlbHCB5XCzY5w6IKJWujqSFmk3zYpPzs6sp9JqVqAbAWZCTK1uIMoNZA6HRxHrV9S9uTHOs2SSSjLMyW2Zjt9KaKl6V6O1MRa2IZWQ1EcRy4n5G9LBnPKxSUCjyIDYWaM3bdub3AQ/MD4EOyOKzkaVkh5MO7Yzjd1O/hTjTyOToSWgnr1A1f6SWwJmJhB8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxUEbKCKe8/aTtOsxCli+ng8tVBiPHRYISYItlvXDeXPsXGFHZhHbqA3BXOJ7Al3cioSTfRYOQZ8fCazLeXjMuBwTYtOoT7nIVV7QHkSimC8Hitk6rHgYBLJe3Z6TrsGRdHpmvw+nYI9ikRLId1/SlzSAGi83ij4iMpHglQLSQ90MYTs2hyfwtsUdZzrukmRrK+SrE9dUdiwRlFg8z0q1SDnXWCzISwE5ie09MiKx/k4LOOMnhu/92K+vmgpkrEgeQ8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/Hz3f2NgC+U3m15chBRdA8s/FUpzID9Mv/WJsSfx9OMCW3gjXOEok0S4TH9S5/MKktaUTHRwmOrUhLTGIGeBivl+zTNpRthTdAVsrIUVylWzm3gjXOEok0S4vnzQq7ijRxniK0mrBLjvIlZunU3QS6KYWm+lCgt4TCfC4y8VeGhaPJ6/nou/PGxo+vy87Qhp/s2sEq9tJYbOGxoEhDLEkB/YbT26ee78cWfC4y8VeGhaPJ6/nou/PGxo89YgelNuZyIMNoQVj4Gs2HW9k/xEsA/V7jGBFTBKPdxtNQwKIvW4OL580Ku4o0c3JT1QvxKJI84woDUElXZkyVHgMd9t6ID5YWVd4d4l5hoEpoGKVb/tJqOfUlpK0V+4vnzQq7ijRyIHludb1tJ1gNccOO/XLE6ACDwf94yKK5xRf+bc+4/TIFEj6WZn/ACrU3E4kWObk044KuW0tEdOm1F32Il+s4UIe2amCghUb3/mAIK5xKYqUM96lkPB7qLUzMxN3ZVssADXHDjv1yxOgAg8H/eMiiuwnHR8qg4ByusPWg6FSenyE7slFv/HsQ4k7EXRx5S7noMff42vU+310M96lkPB7qLUzMxN3ZVssADXHDjv1yxOgAg8H/eMiiuPChdvtgo24zs6rpTEkAOrMIKQH9xapKWG5ijMvAwQDKo1fNd3oasbSXl9AvMcPsPNWYnM+lVTITi+fNCruKNHDcjzxRVwwq1a9CKQlY8TsLX88nixuUVILwo8t1lfYKJQz3FfvCEcUxMnUc6oo9cIW7lMU6AN4kdYXZSwh1m7n5L09BnRleoC9n1sAOMlTzXuzQXK640z5WSqatHnLXJc0kslYxRg4xuJVCM3FTbkff7EvplemzivETe3KALTTmkWeqvSSURVaDFqLXblKCxf4o9UZjnVVXWCoKkBwTO4RU5182bLPIFv1vno5JkABvrdbUMg2MTlGyengKjTN/dQWi6syZn5bD0lysnx2MJWB56lBe6jEjSCb+loWZFvZJpEM1QdQlGyXaoNfGWRcbK341j2fEH9Oosv8b3F8OzqIrdKnc/75K1rK1fUvbkxzrNkkkoyzMltmZazGgsBo3y6L23f9HiueSykYxlJQ1vSfQD7ww01GJMJlxzvvbPTG8YqDXxlkXGyt8/Ogktwxzt8blUUQ1CB5q7TV2sVx5eG9Qj8PMGgN1syV78Qt31rEhQf7jkko578xx9YwHCJqSKDsLNjnDogolaypi6g8qNJM4i6t4AwQan2sLNjnDogolawnHR8qg4Byt2qGJ/T63OOMxBPmd3IyJnzMkjNxwm/oFIfZMPk8JQzqmp7k7PXJLm2K6hMdSPTRzX2DqWnVX7sU/qWQ5Hv1Gd4lNUvbW+wOrumjuFj/OguLOm4GNjZXJt29vsizn5Nq30Ip8kzGNVVa6YsNpgi+6Rnf4aANrGCDCQ0Q8ygJvXeoyPK02G2zKy8QPM73BnLVOhIrQczov2YiRc92bxqcgZ4Lwn2kgjW7fAWCwd+65pMISBp+5AZSzfS3AJxkqhA/xLlPG6JlS1qEWdCC77flxk05W1Xe7Ip3XWvBynW3Y8Oxhrvt/y+YAd29vsizn5Nq1U9OR63hmifhkAQQQY5wT4dc5GUn5akNxOuiXVCY+DRo+BzrtiRr+8kNEPMoCb13pURul4KcA+oGbX9YE2BAPzvasFSgZCszBdaN+5BSM4t5GMZSUNb0n0dJ/RNhdhV/pLGi5soS1D8WZjTk7CmTdKATIba/4QQIeYu0LpoYV/jgxV4Cag/UNQrNwDQdgHXttOuiXVCY+DRsvIxndlw2/n67Cu6nIIXDbnlTdP1SVD7WircQiTwS1Hb7uKklN0PMxYsKM8Nhsvic85VY7vR1UdEuXr+96W9ByqgmkyYRIDFafSxnyK4ka8Su4PQa3bVmprBIDG5Zi+cJDRDzKAm9d6WGtfBT+QcukQG6+W18Oav/zQP48ppIldgfSTdzgr2TOumLDaYIvukZ3+GgDaxggwkNEPMoCb13rY0WYKPte0DMqYuoPKjSTO0KLXf18FbUXgPnqxhI4HtwaNbUPylerWwTjsYrKP2fWl8/e2DgUY8GSfNthhrTQkSd4c8Yu7QP4RIEOGmj3TD/Pa4x/Ly7vx33L5JCUdUrUUmaMupkARDHMOR5HIz51KtY2ChAhRVj8IV+I0T08S252UddhV91ORiDoBkY+ZqSzqTaFEFAnw5x9zLFcFVb+2wFgsHfuuaTCXEYhV5OZR+b0Q2e188EyvmWa6iigPwWyY4gkNBzSsqWT96yf7j6DAbPYtzNG8cPr0IwMM62rQqhhrvt/y+YAdNAsGqzQhOy+4Nj3gfp+GzbVJaQM6SNVzoA5WSPvdW+2oNfGWRcbK38dVtoj3JR+qG6CItCHO0RREiguf16CD8EMk0TSM9YNtF/bivOH/eXnztYY2GvLYDJzMkw3X8uxoby2ENhBK+YAYR3JLHcsoZuhftE1O0pRzNAsGqzQhOy80WfwostzGmqlcH8CGu5cFYRP8ZSQnUiGQ0Q8ygJvXer23f9HiueSytY2ChAhRVj/o6khZpN82KSZ41Foxsw8WnZR12FX3U5F7miPT05xQ/ag18ZZFxsrfrTIP0x/AMDCDPmhAtpi4ZsmhdMzPTwDOYKd6DZ8N0R34Aq0nlxxOjLSnI9mdW9A2E9aLO1aROYygq7qQppQ+pjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZl0qVcZcc1OySCORHUxrAk6KBMumk01vK8FMGJBTLArALd28KpRgYyHQygPuei+tZLKRdtogVez5+BSRXN0q1v9wlaCEIJsXPISJX44lCihvx0KLunvl9r/4eMBQbspR45fyRLNIwGcde09MiKx/k4IogQlVyKQ3wgIVcrD3junMe09MiKx/k4KWfCqIW9Q3Z8zL57mip0pnxyI1jDuM17KP6fzvgkmmTqREsh3X9KXNelChvXg131VZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQky75E0BqC5xoT3/8LhTT0HO0pJAd2bC8Morj20sttFPEKn9g1cwyj7MPMDIgN3wA2lmhb8a9FvTraYszRjnAREi+EWxuzl7SVud8lgvgbK6ImuzqtwTl13MbqH3qqgQ2LS5uy0zqTeiK6RwhYBBfYwiajn1JaStFfgprFl6y4oojwZ5ff3+sY3+F4bvjTw1YNeuXOdiXA4/oq+9yLK/bVb/7BSLiIsxb60N1XstUC8zIwZ5ff3+sY3///9Fq9m2cXxKMlhs4Fj2GcV5R/T9Pl+jTtm8/89hu8aGeqJCRmdRZV6WfOUHHLPQubstM6k3oith1G0ozv5UTxE/4L/XDFvVplFNjUrP3jbNaS5yFK/KSAs8/nrduZqGR3etd7eKWGS5uy0zqTeiKYH16AdxVud0bmKMy8DBAMqjV813ehqxt+dsmPeGkoTvIPtJ7Q7V2DtTEWtiGVkNRHEcuJ+RvSwZzysUlAo8iA5OxF0ceUu56eNMYVsOex/3CPzgAeAtcvsIKQH9xapKWG5ijMvAwQDKo1fNd3oasbdzvuiD6mPSTlM7FV/qoydnBYUSx7a+c9iCi1UT/oEeQFoahIdILFGvCPzgAeAtcvsIKQH9xapKWG5ijMvAwQDKo1fNd3oasbSXl9AvMcPsPNWYnM+lVTITi+fNCruKNHDcjzxRVwwq1a9CKQlY8TsLX88nixuUVILwo8t1lfYKJQz3FfvCEcUxMnUc6oo9cIW7lMU6AN4kdYXZSwh1m7n5L09BnRleoC9n1sAOMlTzXMnCzVZrKboRJYhE/0QKEvaYRNB1oboibntLseEBREBS63iLFularIZ8A84lnmGTM2evb0H+tIbkNEVEEBWpCQ/n7t0tzKCwwrV9S9uTHOs2FU4hlxzpxxgKHQP3Q+YR7AclQErFsPHjVoqmZ2noQJoBsBZkJMrW4qMCelNVA2wXOHnT0rxkORqGeqJCRmdRZO2ThIp0dciPmIqollrQmakaoU/c2JBC+RrNCDQmYD6qcwIjWCckLiDQLBqs0ITsvai5oHgVcxInvlas30N2OIdYubd4q3g5PRN7coAtNOaRf6xMSxaklGvO1hjYa8tgM4OfE/m2jeCfBlJytqBJLIWRREyO/wGvVn+kA3veXZRXOD6zkVh0pQo8ICLvkw7wFYZeb6Q6Wi8tPNKkcPeR6uag18ZZFxsrfCDFi8Mf5UOeMuPJoWygEHE66JdUJj4NGy8jGd2XDb+eDl8oJk8rmQOECmS4PkR1u4lNUvbW+wOrumjuFj/OguLOm4GNjZXJtx2+/7YFOZyPd+7pXgYUtFBXAm1jHB9QJDAFQSVKp0VEDDmo0qbnltrWNgoQIUVY/ypi6g8qNJM4bxysRTdQaKDa8G1mrpGGUdsK/EIw/FDMXGXv+C8GK148WnUzHK6u6tY2ChAhRVj8dhKXsebYhCfvhfGCISCKWoCVkGWUa/AZ2wr8QjD8UMxcZe/4LwYrXjxadTMcrq7q9qwVKBkKzMPkMAgbd8Bdcws2OcOiCiVpp8nkoyvI3slHM2yVOm3Ml34OYrTLIinG7jev7ZxFV+owE0Pvr7BLriqrQM+5Iw+y9SDXlQX4nbbhIUzjiYs5wljEgz1df4qG1vax5gFRFqGhtqFLJbS9mxXsrV/Uqglz3/YTEDcbPj/jd3N6U8G3M1m5/BXeuazIYa77f8vmAHQqCpAcEzuEVadzH5P/DyrCS67yTOwGGySTRDeAGWcxZ3sbpvd9KN36oNfGWRcbK38dvv+2BTmcjpytwHsV5Z1yuyPGmGhT7Vmt/vre0En4v5ufktSkWo4tdkINk58cbd0r15D2mwrLWf8WT5B6Iqhl+jMPgFUFmaxaGoSHSCxRrPW7loPnU47sASlQboJTlvhLubMjDCne3FpziG0dVJueDKDWQOh0cR7QR9MkxrqogivQjeGQ1Z4RMhkqnWgnKzL4HehfI+P95eRio3fZ/ac4ASlQboJTlvmsezOrWWHiuajkcM0HTJMUCgedoCuA+3fzmVF/ctkRXnZR12FX3U5FmZVD+LBdvK0KuWnwI9ksmewEsd18WgyHy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/Fkb5u9pEAHWTxAPOfM63n+4JpjUSIgOcHBi7fQX9B3GfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxH9vq4kTJEDLhvV9DG8U+Z+diDw8oA/yUgKn9g1cwyj7MPMDIgN3wA2lmhb8a9FvTraYszRjnAREhVdrll9sKK6La2qFhQHv4E+ro4JhRiFWBNz7Ynn829T5Kpq0ectclzWaFvxr0W9Ot7A827fZ/94aTEtCM6JTfemuzqtwTl13MbqH3qqgQ2LSVQjNxU25H3BLUZRP9K6HZGB9L8oDlvzfvExV7KRT08muzqtwTl13MbqH3qqgQ2LSMEdkLgw0dQWZpE83DjuVDWmH0QnDKBihFlpWoLRMoV5bpT/tkBZNSSqatHnLXJc8ucSVbkTUA0J3ow1ybKT4yxQZ6gRrrYU+OhZ8JWXQkoyD7Se0O1dg7UxFrYhlZDURxHLifkb0sGc8rFJQKPIgOTsRdHHlLuegyy8elbgDrZMimRuJCPMe9TMzE3dlWywANccOO/XLE6ACDwf94yKK7o6khZpN82KUHI9aDL4/wTm19DyA2QWSzUxFrYhlZDURxHLifkb0sG3HJKFUTLr7pkV2RKeFDdt7Z1LhaFLbHQA4VO+aLRDjsbjRZ04sMmZpQK1zGlg9JjMPenqpFMMaeTTIotbD3d9WHFVEZ/yr/qO90dSaW1lw3bZE86N3Vad6CFpiqCEM806aIZAGVoM765YOX7gU6yaCto6qRcTrPRohmYNO0SazC0//yLJZNFE39byhFoSVL8edW1WpNGyKaCAIczG/6hgJ1gOr6ApWoLaKtxCJPBLUdj7jimXIKZPAuZhbu0EawqLm7LTOpN6IqRPRnBG0f+2OuXOdiXA4/o4SSlnUTC2QgWCK4BxSW31QM1bFVqXuaXoA7EpVKE/qVK9eQ9psKy1iXl9AvMcPsP7+lZSmsI8XRourMmZ+Ww9LEddF643SlEbYHdoSwozNmn3stXColEBnpz07QGDrdWx2+/7YFOZyNFgBHmCWp1lRXAm1jHB9QJ+0wRCQqLE1zEDX+2RjgsecBYLB37rmkwpP+F8h81xcWJgOL/ulWbggMffkOTIQ1Tc8KnL/Vuix4lUIzcVNuR9x4RxoT/hZ3vkNEPMoCb13pYa18FP5By6aFOWhvQIMdbnm+KT6SkUD1qNyl9rew/ihE7nNp8sszc5iKqJZa0Jmoyt2j8t2e5uQpGpqBkhI+ESXRDKGDxasa1jYKECFFWP+jqSFmk3zYp0fsaZDC8AflInN/tpiHunC/Ey5zgjnpOm+FBP5/V+6sYa77f8vmAHQqCpAcEzuEVSjRbDFVPgLuipIaLgfXlFPWzKVV7jlU/WIIAIds2MSqzpuBjY2VybWo5HDNB0yTFBEzlrdCgbpw2/ULkhwzXXmCneg2fDdEdcMu8SZo66ms8LuffbjjCmTbQpprNa4fnVRENgWJj/mAJ7Wsg6VowrO26DEPZAh35/sCusBCkCcidKCAKe7ioPJUzaieDhIg70ruTV91SZC4fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwuJKt7Kze/qfEg2GBGWdp6+ba4tYSGGu76g6WVlzc1l0pOTpOcBgaCoXHACojHgtWWxd7lNh/wwskDvGcVrJOJStW35N7S1tYN/XtlbBqfF9En+237qd7yev+Z0zNMzgG65t1JqDfV34q2zEUq06bqVnBZlDDWPRc0fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv19JhV0Bg8FAX8cYC1vw6ZInrSOdnQKWp0tGcGsxfg0omtQ797AIb1pn5zUaoL+FImERhWsm5kQkFnNNo97vtpDsuOAuWahUAp+b8/epKVm2q5gyM5K/Ntm+rPKsEBPe9BDw5nl0nob9ZJwV5YQzzonSggCnu4qDywUBTkL2d8ouiUB+Pgbq2QWwqNIEAgjQzsSW5LvgxoxhwTBtm/clkkpmH7SyfPW5XKPLOlfCEauVCpCbUnTKAL3fB4M+H++XZqz9ZhWHvovNaYfRCcMoGKrHEBNYVWkOfy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8aYPOpim5d4PnBEjSImSjA2v0M01y2Iovb+WL68jVja08v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEfET/gv9cMW9XNx0AXermK1jiY81PWGBDdTVBqJB8oL4SR64g5RIKvAmo59SWkrRX50fcyomcziLRuofeqqBDYtBLw1PtszppFN5jzmcA/oCD0t08jyjY9hq+9yLK/bVb8XU6Ay9J9uOHAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcrpLydPnYbDpNRZtho2r7ijuy29NHSztQNYWhWcUDcHCHkVZjqqtrl7s4Nv7JQ/3RiXTDn68kBVjWGKdeOXNrhuofeqqBDYtvkUOfzCMW1ngGdmu3V7h+lgELcI2cuHlq+9yLK/bVb8XU6Ay9J9uOMGOdbJ9JQtT0IfOTurgDkODQg7c6oNYCJwwKNE35BB990roM54EK1imaNlzPwo5sDE+uVqwwM28qKgl+Cl8oUobqH3qqgQ2LZibnm2Aoe5zTeY85nAP6AjE/jD0Aosqt790/v0Oz005Vi0YdZUWnCP4ykDFWmiWvVO9d4D4TNSLZe+SbrxqF+p2mh1DDys6gRPtTqKOd5yP6d7Q0qQ2F//7emgPJ/N2ZPh4xY5V2Uraub5YVOrHt7hh5ejBTYOD3dDsO7YCStYgvF5XbSxEKXkbqH3qqgQ2LZgQMrMQdTH1+SgywgfpGdAxVnjt2EkDC3sDzbt9n/3hrB0of9AwQRIqzj6lr8nqicGOdbJ9JQtToAKIHjDKC8IuxinGJGN23/ZSw9kAR1Fo4epBBCThubgnfB1/43zu/PVA1C21mBZ6XmKwwVwQ8HJ4E8aLOHGahWW50JAXJVSX9fCtUq8mxCLsY21T3uRMTSlT50JpQ6IZO03oo5dzY8Lsqu+J2ZpR9fJl5c4BOSEjCH6ltDmp5o31F1pdw6Brx22tQXIXOnN3zRhCO1/voFBYggAh2zYxKiMkpe6qB+YHgvk2ra7jWnjkRIonLHIBpMaBW4VdPXXgv3T+/Q7PTTktLeagn/bBLuUI5d3wGEtsT6hkAxz4gJkcRy4n5G9LBpY57gFx+WW+14kypcIU8Y5+aXlLqSGkYj4dPRBoau9wqXPmbxtDMhHdw0PrZsWx+12bKts26arYo42UxL+43zqBxl0y+KwUu21F32Il+s4UdRi6xiCt9dd+uoW8v7QTlAWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w8oACBRsXpDAAAHguAl8GJ9CdlDjFnY5zlRWHJYQ/HeHYVd/hmcRcoXVgxNv1+NZ8Mo8s6V8IRq5UKkJtSdMoAvd8Hgz4f75dmrP1mFYe+i8GmzRe6RhG4gsAUx65quh4+HDJoDEt9A9HBMG2b9yWSTdBKi0KQJgsSd8HX/jfO789UDULbWYFnpeYrDBXBDwcngTxos4cZqFZbnQkBclVJdewcwKoALhOViCACHbNjEqIySl7qoH5geC+TatruNaeJflwNcfg3u+Ph09EGhq73Cpc+ZvG0MyEd3DQ+tmxbH7XZsq2zbpqtijjZTEv7jfOii+G04JfRlAVFYclhD8d4dhV3+GZxFyhansBGLG4sVHyjyzpXwhGrlQqQm1J0ygC93weDPh/vl2as/WYVh76LwabNF7pGEbiMC7q/CTDcNca9CKQlY8TsL2UsPZAEdRaPxKE4tbCfjG7KrvidmaUfXyZeXOATkhIwh+pbQ5qeaN9RdaXcOga8dtrUFyFzpzdy/b13kGAN8SHEcuJ+RvSwaWOe4BcfllvteJMqXCFPGOruVZFG1win0FlZovy43TGHwWSnEfLS8kUlBsfAG9u8PKAAgUbF6QwAAB4LgJfBif2W3a3wXw4fbC4OEyxUpTDzGkUbScpd8XbpzZDEZfO5bKPLOlfCEaua89lpwFAvlQ/OYyC6BzaD6R+8P9B+Li0pTOxVf6qMnZI4vTKyHBGc+ia3IMTTWunlRWHJYQ/HeHYVd/hmcRcoVcKm1mS6TjY5uh67W335M2+VTcuF60a3lSUGx8Ab27w/MqTOuUQB8jAWDQJ3KBpIOSxWonF3FK3IHGXTL4rBS7bUXfYiX6zhRax+85yFK1KCG+kpyK5fDDm6Hrtbffkzb5VNy4XrRreVJQbHwBvbvD8ypM65RAHyMBYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h2FXf4ZnEXKFILyjQAbRjKXKPLOlfCEaua89lpwFAvlQ/OYyC6BzaD6R+8P9B+Li0pTOxVf6qMnZI4vTKyHBGc/8kzRDBuhudcLg4TLFSlMPMaRRtJyl3xe9mX55Mj8TWu0DWuO35dXhtp4a0882wVTd8Hgz4f75dmrP1mFYe+i8rD1oOhUnp8jqbdmcoQYqPLL7BcGqqvAn4cMmgMS30D0cEwbZv3JZJBLsyBh6i0eBm6HrtbffkzZiSiR2u+FIv/zmMgugc2g+kfvD/Qfi4tKeuCv8EL5+zubV9EPoBEz3VFYclhD8d4dhV3+GZxFyhfofWMA7BUp5Ph09EGhq73Cpc+ZvG0MyEd3DQ+tmxbH7+cAw5ftJgkGj99yOUBIgrBxHLifkb0sGljnuAXH5Zb4CfVy7pt5w0uyq74nZmlH18mXlzgE5ISMIfqW0OanmjfUXWl3DoGvHu7lyLWw/4bda9Sh843vJFuxjbVPe5ExNKVPnQmlDohlPMdwAOegRpO0DWuO35dXhEYNU9Coc9yLK1hAN0qkLhMxbYEEvvZM2QxYn9XKnHX3nkjRpdXAmkuHDJoDEt9A9HBMG2b9yWSQSU16jowa3gZuh67W335M2YkokdrvhSL/85jILoHNoPpH7w/0H4uLSnrgr/BC+fs6IhdTrbbAMB1RWHJYQ/HeHYVd/hmcRcoWBzVKEGOd7EAWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N15P/MTFnKkSFRWHJYQ/HeHYVd/hmcRcoWDTEp1chIgHwWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N3F+qHBRdksN1RWHJYQ/HeHYVd/hmcRcoXVx4fVE8v8xgWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N38ChqcrOjAqlRWHJYQ/HeHYVd/hmcRcoUdLF9iBgfSAwWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N0ovhtOCX0ZQFRWHJYQ/HeHYVd/hmcRcoXVb6LEz/gTpAWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N3u+49+N5j8NVRWHJYQ/HeHYVd/hmcRcoVyxlXOC0CSCQWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N0uiOCvAh4SdFRWHJYQ/HeHYVd/hmcRcoWbCjAfTt0nhgWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N0hpOPYobPKzVRWHJYQ/HeHYVd/hmcRcoW3OkOIJwzyigWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N1hw4ye9aQIFVRWHJYQ/HeHYVd/hmcRcoX56anHvshnkz4dPRBoau9wqXPmbxtDMhHdw0PrZsWx+6W6jAtQ7NSzr5EQVKqlJmfsY21T3uRMTSlT50JpQ6IZN7/isUTshhvtA1rjt+XV4RGDVPQqHPciytYQDdKpC4TMW2BBL72TNm10LBNExmx6QnZQ4xZ2Oc5UVhyWEPx3h2FXf4ZnEXKFQ9W6qBwySEUFlZovy43TGHwWSnEfLS8kUlBsfAG9u8PzKkzrlEAfI/XN0ECXBOZLHEcuJ+RvSwaWOe4BcfllvppGQqsJ6lhA+UqBclH1Zl3GgVuFXT114L90/v0Oz005LS3moJ/2wS4Nj/ycJBqmvjGTzC+tFdi17GNtU97kTE0pU+dCaUOiGVilk/aamdD5J3wdf+N87vz1QNQttZgWel5isMFcEPByeBPGizhxmoWKOIoVfakQ1O95b3xuiqJ14cMmgMS30D0cEwbZv3JZJHDplIOR+P+UyjyzpXwhGrlQqQm1J0ygC93weDPh/vl2as/WYVh76Lw1Zicz6VVMhO77j343mPw1VFYclhD8d4dhV3+GZxFyhW6hQp6saxA9BZWaL8uN0xh8FkpxHy0vJFJQbHwBvbvD8ypM65RAHyMwbMyLOKdd9xxHLifkb0sGljnuAXH5Zb5jntRuL2GVHTM7C1rqEbUDxoFbhV09deC/dP79Ds9NOS0t5qCf9sEuDY/8nCQapr6u0ywU1a9xp+xjbVPe5ExNKVPnQmlDohmlwHaaMzfqAid8HX/jfO789UDULbWYFnpeYrDBXBDwcngTxos4cZqFijiKFX2pENT6uiDHkJbnkeHDJoDEt9A9HBMG2b9yWSRBN5++Ce9cpso8s6V8IRq5UKkJtSdMoAvd8Hgz4f75dmrP1mFYe+i8NWYnM+lVTISKQvleug2OFFRWHJYQ/HeHYVd/hmcRcoWKfKy8M4NGjwWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w/MqTOuUQB8j0kN21EY3p3ocRy4n5G9LBpY57gFx+WW+Y57Ubi9hlR1VHhHX/SSnmMaBW4VdPXXgv3T+/Q7PTTktLeagn/bBLg2P/JwkGqa+03ZTtguYRprsY21T3uRMTSlT50JpQ6IZHAFuQufF58knfB1/43zu/PVA1C21mBZ6XmKwwVwQ8HJ4E8aLOHGahYo4ihV9qRDUjvRVbRyIZJ3hwyaAxLfQPRwTBtm/clkk2CSCFOiBbunKPLOlfCEauVCpCbUnTKAL3fB4M+H++XZqz9ZhWHvovDVmJzPpVUyEIaTj2KGzys1UVhyWEPx3h2FXf4ZnEXKFeRgyryh/lyQFlZovy43TGHwWSnEfLS8kUlBsfAG9u8PzKkzrlEAfI2pYUdsbq6MZHEcuJ+RvSwaWOe4BcfllvvAH9QMRnGQyYeNhmqjn/dnGgVuFXT114L90/v0Oz005LS3moJ/2wS4Nj/ycJBqmvhWvX6YGThMv7GNtU97kTE0pU+dCaUOiGQRCDBBhTdtkJ3wdf+N87vz1QNQttZgWel5isMFcEPByeBPGizhxmoWKOIoVfakQ1IEJ4xPIApjN4cMmgMS30D0cEwbZv3JZJNBJUOSJNtKnyjyzpXwhGrlQqQm1J0ygC93weDPh/vl2as/WYVh76Lw1Zicz6VVMhKuMjhEadZ2SKwToSBd2MuLWo6IZC9F/5AuYOyEp0EiDcFRBBy7QQJjQRGEpx5qru9IsonT1uyPaHZIVgGmGPplkLbvqjM5nGQyr/RDaViH/9vq4kTJEDLgykUV9ihzFkEOuXINAhUEU/xQ8kLqYeSmvaczVN04/GowJz7XvC21mv/O5YA6k/Chr+KVDNFYgINajohkL0X/kQ28OwGFrYstHUBIp6wAdhJsXNgTamt+dq+SjTAfWpdAS0xiBngYr5Z64K/wQvn7O9ovv3izTod7Ew4MATawI+z5RBZzJV+rYoOM0qWobbY9JfV5hnmgGTcIu+AmZSzjIJu/um9PrknouMa06uX55ehZVbSWFJkj8Cl+chz497fKScCX1DB23583NonL3dWzRuvv15QtiSAUcRy4n5G9LBrQ4aS4ILKhEhmTvfwks6l8CLmfIM/UTQK0PJJjKTd001EDF+eslQBKmCq+celbcYEoalaCF9VPhr4ePFoHgHviag7zoWYYl9wlo7SAyY34TT8j3mV/adLlVVHZWTNJI9NwLW+qZfNqtbCnBr9+eQ+dh+kp+lXpT4zuOlTZns5Df7EluS74MaMZwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkw0p9NLVo8qpEzy5fugPzVh8qWiurn64jyeKJKsvCqSZittbmMoORLNZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkxeZMP5ZiangoBU0R0N7y8PNghawJfC4752ZIevvosDue6cqmYFapnOZ66FqCFbUCzpEo49KB6oCNR72STGKNZ8/65ab1SHNsR9TFW4JdLljSFRmxday5j7mIqollrQmahLTGIGeBivl8IMB0jorXOipfPtPcln2uGCneg2fDdEd/z66MD8vr54Q9BMUbPYIWyzSrZCTRoPljB734P4U3Hp0pNR7i8zmhVnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTNyQ3dT7+qhvy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8YG5Ur/Px+18LdRrUx4jyWDA11Kefwq9Itu3ycR4iwxc0/Jjl2gKHf/y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR/b6uJEyRAy4MpFFfYocxZBDrlyDQIVBFP8UPJC6mHkpr2nM1TdOPxqMCc+17wttZr/zuWAOpPwo4USuAIYBNog/65ab1SHNsR9TFW4JdLljSFRmxday5j7mIqollrQmahLTGIGeBivl8IMB0jorXOipfPtPcln2uGCneg2fDdEd/z66MD8vr54Q9BMUbPYIWyzSrZCTRoPljB734P4U3Hp0pNR7i8zmhVnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT5XqQCbH0FUzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR9aGpozh3oald5P/T3smJtqUwzuvBwcZEzR97ojYf/rqG89ZeNx4SsDB1W6jSiFKuqKbTsfrBcDdcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMsJx0jVzxADh2RncgRHF44Ei9MOj2bCw3vt5NFMJVwX+mVkwDpd1m52PfXMMKi7udVdrll9sKK6La2qFhQHv4E+ro4JhRiFWBNz7Ynn829T86uDXg701h016zdY+7gque/dP79Ds9NORxz2aV72P1tf+U4Ljxdhslj7jimXIKZPMRP+C/1wxb1jFTVC1da57Sj6/LztCGn+zawSr20lhs4b4GoSMHqf5g8MB1RyZzk9H5RcNB0Y414Tc+2J5/NvU9S/7I+O20A1eEx/UufzCpLv3T+/Q7PTTnvS0yqfLfA/fHdVw9HuBxh9gcP5UVItPZxmKdMzxK6vdK8WJrcBtKGCo4Eo10lmgSfouWrei5nHgWVmi/LjdMYfBZKcR8tLyRSUGx8Ab27w2zwfmoz/VQbVMz8s7lE/N1Uf6nM7ZL9IQE/guDeW3Iq7GNtU97kTE3SvFia3AbShiuJDlhnagBgbVMhG5GuSU2NJx7w8tHUsEc5WGRlNKj62gvpG5cakkBZ/P03QpcfEy39OmVUNK9WWyf/KMIBsqkHj8SxtqN1mNTSRCRalyta4cMmgMS30D0bmKMy8DBAMqjV813ehqxtKqYdaOM7pm6zLzf7kXdle/7rFS/YCcMmzJVhSlJVabaVONf5mDWVfAS1GUT/Suh2qmA+PLbqdMrSR+EYhUn6ylu8EVTQ6nd0mvv76RJp8q1cXqKMo9pFVgmN2zjTSiaErf+Zxr0GVxzulW6ndXTiulEPp5ISEdMkO9tf7B5akt+yO+C6dwgZCf41lnblFWJq6th7ZrHrv1wyo4ep/ZN/+64xKFFcwID19prjrMmAo7dQ0Eb6lzyhs8OTyNLgcNdkQIaAy+tSTHHkQK/WNyYU+xpjN+NMLr6RHJ7TLaX4iiLHb7/tgU5nI0WAEeYJanWVpzXSFAaeCde4S5g4i6k1L8LNjnDogolaCBIImGH29F0Hj8SxtqN1mKe/e1fD7vJlNcz3Y3VAXWaCKXglvNDwpQ1s8E7IYjG8s6bgY2Nlcm3zEHuynralTQKB52gK4D7dNBl4YnPWAp7dJBylX5VGYgePxLG2o3WY1NJEJFqXK1rm5+S1KRaji12Qg2Tnxxt3UJORqUMJszKkaob/OPpUhWKYlE/Yt7+1lCcmFqKbx7DXM4IM299D551CQG+whAA3PC26ZBtIw7wjdaFtlHxN9BZRTCWZ9HtRws2OcOiCiVohlqoYVn4UaY7j2M5Jh+x9PwGopGN5FQ4E3CZyf4wRpBhSWCXX+Sr1NCCopbgUiKnGLJsafJl7FuuwrupyCFw2Q/i9SenvYJ9k1474miVzp9v+Wb4/9gqpXZCDZOfHG3c3Z/t23jIIOSGItpwm5WaApBalGmZgvwDR5ieZM43Z8VBs5MeygkjUFUjOeyYmrRmB8tYSRba22yGWqhhWfhRpM/CfthWsoLvDUday3LKTASGItpwm5WaABqQi7S79Wz3TWRy6M7nz0w1s8E7IYjG87tPw8w01uGC/StlC46lljpDRDzKAm9d6WGtfBT+QcumhTlob0CDHW/MQe7KetqVNpzTkdVRDLD3Uv7mFxss7EPj+2GZTnoEGodDra8bnlyp0cRI00EQFLUNvDsBha2LLR1ASKesAHYTLVhrhazZewPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk2wB+7h+Ops6cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPk3fhOuSioAbyq8Wm2xhak16Tsf03QXLBjEInwZUrqv+RmWtChEHxJcC1JNnembCXAM0a3l1uLja6oLHpVV8Np8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/Hz3f2NgC+U3u5Xklg/cjEu+E5fChEDzRvrX986XsstBA1kl9fhw5akjAnPte8LbWYdDzAU78zsZV61fZAhUbixwZ5ff3+sY3///9Fq9m2cX0c5WGRlNKj6rjkwZ5Cn8mgZdtSKwYfzVzPM706mht6Qy3DswB+taRyfC4y8VeGhaPJ6/nou/PGxuijQhG1j7mxZoW/GvRb063sDzbt9n/3hVg7HWcWxg4hDdV7LVAvMyMGeX39/rGN/cKiq3FWcSYmVONf5mDWVfAS1GUT/Suh2kd3rXe3ilhk/AaikY3kVDgTcJnJ/jBGkGFJYJdf5KvUgZ4hsPBG1l/1ugukkm/R3qKEn8e9LDB8nfB1/43zu/PVA1C21mBZ6XmKwwVwQ8HJ4E8aLOHGahYo4ihV9qRDUjVvLkc6jddHUxFrYhlZDURxHLifkb0sGc8rFJQKPIgNhV3+GZxFyhRQYjbUyBeePA9+EfURL1ORFy1NiCVwoZF5KT7GfnZ0hAlqEL3jNxSe133Aes06zPeqCaUBDDGzaGFJYJdf5KvU5XbGukr+cOuxjbVPe5ExNMHRKiVWorhuZW8Gn8vZC/Xl1J0pu3JgRIz4gTwMALcgDXHDjv1yxOgAg8H/eMiiuIZaqGFZ+FGlniK0mrBLjvDc94ADxNcvlLxXxvnwYbtpqRj8UXwDNaMxxKz/86jqUS5jc2cXxjiQNC3dqTDDPFNFtrzx2NQD3m6ydiF3BQUIKGnCbdGF8+hhwSrMeIlNeHbyceMIolwf/T6desC057vkjT1RpnTbPPN4pLEffj7/F1ehkOX2pljdn+3beMgg5miSFpFyxOAdRCWbeSOoaDbtwcZyZxxotq7z0WNseUXcT1zWClEYtH2qRdR2rIf5Pnt7wAqyJilkETGOhmusAceVJru0SfqKaEIR3B87jZMXPOVWO70dVHSjgX4SQvpv2GFJYJdf5KvUl0kVd6I9XC+upeoVu8P7o9mM58TmWawAtr5YOpIy1GsdE2d33lYbEx1W2iPclH6oboIi0Ic7RFPoyMQRQMJ3tJYswwyzV738YUlgl1/kq9Tldsa6Sv5w66GJOJWzoaHcDDmo0qbnltuQnfxo58a0Pqkerb9/0PJf5gEIOUMJDT2pZH0Js0UgvFdE6F4ndwAWkaob/OPpUhSwNneBEclq7YdmMIq6KJs1r3cbOwbtgy7EddF643SlEZv/aciMOengXywxn5DqdtsWCeqU8hMhX65c52JcDj+hifLLRb46RFItsnj7/eesYuvr9GEghadTjqS2b4yIpdlRC/FMzBQP6fgnLAPM7YegCL4kAwql+gAMOajSpueW2SvXkPabCstZKPfagA4hoTR+HX+e+EyQb8x1TTbZl0m58l/bcat7/iv0EIgS6cOQBzaFE8TZHJv1m/9pyIw56eA1Cy3rAnd8hsH/3oQTw5E1KPfagA4hoTcKiLnxbeT333HXdzFORfHctr5YOpIy1GkwiNg1tb/y8lTjX+Zg1lXxj7jimXIKZPFRG6XgpwD6gZtf1gTYEA/PHVbaI9yUfqqiElkWPOTuYEtMYgZ4GK+X66zThkS01sfXWaUqncgTFLH70chck88rEw4MATawI+z5RBZzJV+rYzgNfLR1CceqXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiZJfJT2nt/Oy0V4GR+KKys4E2lMnDQinRNiw0JFvUEcZaDQcLL1lV9/N9rtkCuXVOQ4rZgEWPOx111oFCWRqiOJWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMXmTD+WYmp4JCx7LDjAJnDnh1SEIcIwkM9zQjfrwajONWZoiiFN4qH0dLAGo5XTXHsY21T3uRMTWwW9iiHlNjGrD1oOhUnp8jqbdmcoQYqPB8pWXSZSj1OIe2amCghUb1L2S1cmZNFpxm4dksQUX+Wzc2icvd1bNG6+/XlC2JIBRxHLifkb0sGc8rFJQKPIgOTsRdHHlLueui6Xf2SSSRmr4ePFoHgHvgBq8OYNNE4kdJH4RiFSfrKEjZKLX3iONXV3XOfIx3XI2U5KTI6ttYRb580ad4N6sEOXwcdMyM2dhFXqcS8alUjQyqPvE1DdKlbrQ/WgDUlb61fUvbkxzrNkkkoyzMltmZp6IyCaraU/UdkfOMwP5zO8Rp7kdD9W9cQ/MD4EOyOK3rV0TQIge02eG2gKRi7tthAFr9VUDtbw5/zHEc2XEGvStSnt59bBhjUQMX56yVAEqYKr5x6VtxgShqVoIX1U+Gvh48WgeAe+JqDvOhZhiX3CWjtIDJjfhO9XTEYfeTIji8V8b58GG7aywKTkKJerd/dYrG9IrDBnIdMPQli8g1QpbBDjLCMeZRVW3DiKRkzwhA0iiIzyl97gGwFmQkytbiDKDWQOh0cR7Hw9Ya4xpPWVTgwMqe8P9lhZozdt25vcDNSC50CghXz8939jYAvlN4Vdf0sP8GLr/Ryz82RAliHewOuTFQXEC836fokJVW7b9HLht3g0Q+viRBEiIwu/d8K55YaiicrcZj0EJIIrJfLWJ2KnGVS4jRLfeFRTmgh0QRYfj4vCt1JjWp4X/fEthVl3pEEo0zoSKn0kHG8CNQXnAz/tY0NP4c0p6jWOL6R+qToshz/rweqZIKw64sLmaNz7xqqm7aS44an4nrK5j1oJfQStDLFQ01WNbV8zjtZu00HjFkuFs/ULsF05dGSf7A0Pn/VgPsBDy/3hOVKUaEJRnoIJ9g2lpY0Pn/VgPsBD18+HpiKWFvZINmgGWztr9IgiU2dFg3BccQ960qIFlK2Trls1ZJGB1d8EgNGoYoA+k86/2QZrtGw0/wt2HmmrlUrGxeGBUye7EzMVeZioIlterSgAUVblC1zUrhyMHPiGEWJtq0XfVEwOO2pnU0JrydZyQd1HCuO7NO9vZgYpLhuDPbkBzQdmF4C3GyeKu1sA3++zESfaqtLSmbLgxsBVvDnzu2uMSHUtm24UXWZ93SqcltH5Z1YRBNrqwyQz6t696xxATWFVpDn37tbLbwCTCAv3//9gJQ1aB6UrcHEtN1hdptYTo5RyvvWv3HztEjAKsA7RoU50YOI+kjjWGn+pRRbAuMDzpUVy9ajohkL0X/kLQjENVqBRl6yji1SZLbhRg6AfcIZ55g+bBb2KIeU2MbWmH0QnDKBiqxxATWFVpDn0uKnh3OBU5PHTlNvSDCf1IIFAqqIZbzyEHmW84XT8GDia6ZdiOLlNHKfmA/tO6HvkXqa2e0qgYuJZP14xGil+iwnHSNXPEAOxxOjV76ilQDeGhbaHcPyvTNr7qP1MQecrxhl00PxBAr+ryY68bCm3y/UPIBUiTHQhGvSy7s0Z6J9gFA6FCVksETk5O5KbTx7Y2kOcbirTHMiqbC1oZrO/Tmipoug+x8neOP6qAdbkf4a++4I5TsFsDZxlBfyw/CMuYbXdfjgjJ+jnZHlAzqm8mbYOSeSyvPJBHBRNy+iSjfE0DsuyXaXntCftbikVuLR1EDF+eslQBK8PTBk3PdvfN4aFtodw/K9M2vuo/UxB5yvGGXTQ/EECv6vJjrxsKbfA3W/qowsOlW52Cn0JLAPGxgWSxfSmmX+hGFgqmASbH3TxEcWWioEB7BMRycdGw+mu1djm6U5DOY+eVd+Dcwcu2BarwBHj96D4mumXYji5TRyn5gP7Tuh782a0SxqIBG+rOBnT9RdRge/em5oaCkppiWatKptj5ooXCUgcjrg4tegxqG99BVMRcb+/0YvzP1s96NuItgiCOzAWCwd+65pMAo87QNhWHJ8beCNc4SiTRIv/pq+69lgIUIGkWjGk/dNQLw4iiueoOKrx7tK8uVfzeLf2aGIOmIFuRicv7dGsbMggW261MLKN4prYSX/XBo2uPCPwMD3gx6DqdjTzTnd1sbTnRb7om7LdflakqN+CvvWo6IZC9F/5C0IxDVagUZeCJ/eyJoULDX+ryY68bCm39PC1od5iM1b9xRdkFrqZV/GPbG4bYuGlj7RsYEc9qLvREgFhSGKf/yg6MEj4Km9XV8vaYQ+E+yqsfD1hrjGk9ag1uT5qIfGpXK6S8nT52GwYU5I7tctEXGsPWg6FSenyOpt2ZyhBio8wRllQdqKbSSdsiWbLnZgOxyhQeVck280U/PU54Vd/wsaVdzDZB/7WXyvkUO4cdh/AWDQJ3KBpIPFkEyXaEK48BLTGIGeBivlfRcDUIWlX52bKbFVC8Y13XjU82hxwyKEs16wVUTREvHTYmgpGkHqNp0aURK7nY7emCNB/Ui+52gdYCA0bKI1vI7Vcpa3x0Xt9vq4kTJEDLitDbjdUkbb94bFiEQK5urj1ph9EJwygYpSBYRmj2zA6L90/v0Oz005grgujKbUrP8dYCA0bKI1vATf5WfIrTTcwY51sn0lC1Mu2x8fIx2HCGHW9k/xEsA/flgzdT+AQOqnDtGy5QsDkUrrNyOtQq7jrnWI0Litikm4ZCyeZ0RWDmerIhIt8k+Oj+zl3OsGIozoh5KoxCdYwoR1KYRjmxKfeIEWMn685D7TWena3neGC5nroWoIVtQLvhFsbs5e0laneSSYQwnU1Davr2hlLruV+FJpoRBNj49boTyYFjhMlNFPNU9RZoP8y31CPaOtq8ukZDRZFGinJhv78VamsGoVOFeAQZMniyn2UZvXgfthisBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMRP+C/1wxb1FKSRUZJW2f1doPDqTAXZ+Ln9p8BFGkEDYO2fkMaHs6pDRDwuChd04SYu4KqWvjvGBna6Apbqv55x8tfLfHJerR9H39suf2qrm0KHQBZSWjaII3XwmDHYkCHtmpgoIVG91OrVDwu8mOlrRYw+DambdLVa+SA+X+xJG5ijMvAwQDKo1fNd3oasbWsEfBjq7CmJnImtp5chWA73bXmhrVVT3BuYozLwMEAyqNXzXd6GrG1CrpurXlNjtKQLHHvANWXU5H3EcBCUCEiscQE1hVaQ59kuOd+Yq6yoFLMzJpytedSaApkQAR3YQ3O+g8+YjV+OZMAtFuUZoekxLggftS1lBbjEZRpET6MzG5ijMvAwQDKo1fNd3oasbQE9TCAjedSZuu1UUbXXuUVRAMRfiUZYrCCi1UT/oEeQVj74zqI4xqFOxEzEHoOHOtaG+TeZLE8ymlYqV8JzNNQgotVE/6BHkH2Uk6QzKssaGvyf9BN60rEabNF7pGEbiM2LjsOLP3OvmnUzvAfa8R/0EKCRztvjRvA3JkPT22pdBna6Apbqv55x8tfLfHJerR9H39suf2qrD5Cqsc7yA3Bx4q7T19FIoxOl5wm/+vjTDBCw04mzFx4DXHDjv1yxOgAg8H/eMiiukIGZiKmzQHzt1tRQtVbTvj967mUGBG8jk7EXRx5S7noXQb6fB2gviI9onXBLEFsaATdyZWdPOzlVX8TPGNYDIfxlIluSA10xqjGGlBfkgc0LoJ4pAAg2LDQBmQSaJS8irOBnT9RdRgdKMURBn49/9bwYiE/IZiK5yHmsxtb6EWrtCTG6bpheMuLrGZzfM7WLk7EXRx5S7nppNW4M7/l/AlwTm5yGZISK2w7y8SLJNtP+6xUv2AnDJqdPVz2MxCOityM08QF92bzWmH0QnDKBikC8OIornqDiTrls1ZJGB1d8EgNGoYoA+qiDCbhSh4ey7LOXWm4/mINL/vuShckTsMvpGvZGvxi8D+3Jrr+jnibolAfj4G6tkDfp+iQlVbtvToFGRsKaAxOxvm+vg3XKFuiNuPW/CDp0x7oTl03mhREEEyoZAjAoDKP6KF+0082mWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJN96SOtonnewU6PwW0Fzuo3fAgRQg7eaQpM6BqfQBymJYK7VWvf4c406JI6KPePxIuakFy00lDE9GanoaVHZtbb1tyKzfoDWBby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8fPd/Y2AL5TeQaX6XGIH1ORo+KlXbOJ+j2DOCw2PdT3NK0RjtJINLBLTVr8ikO3n6QNccOO/XLE6ACDwf94yKK6/IJ2L1uBdWA4S3ncqY12tJ6b+11OiNzFqPwv0nP0sP5W4fYsn4zK4EJ23uxQ2QhpUQvxTMwUD+sWG9buciYGFnWoUcqwNuVZ3JIi8mi8yGSLmdBWB580NeSJsKrpbXVKYb+v8Y2TKNcWfEoPBDPxdR+5UMYJvJVYNCbpYFM9ncR+pBQUd/IzhcfToHZ5ByWeUPQ5KkdgkjGiCdMx+Aj3kXFlznEg97cWMHvfg/hTcejM4iwf1oLOZLBGuKMrj84Dy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNsAfu4fjqbOnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRySpz0GsPGwEhziXlgLIuRL9V5vb0mIFuQc+fzBSU3OXD9Kh5oUnbOWD1VceMecD3u/XI6enqPtQzpSuOf+Qn9xcenq3SGECBO8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/Hz3f2NgC+U3oLFF05KgE4PTc+2J5/NvU8mS9kkii/K2J08ueDrquBNP8YS+Cff/RwS0xiBngYr5XcRiwtwdKjj+ro4JhRiFWAgotVE/6BHkPgpgeywSBMiRg0eF18pdwEue7H9bpqx5m0xLJZl22snz3q+rNCxNvrGBAf4OEaMnTfFb5Q2+efxgtEP0V+kpTVH19+VSNSzBP7rFS/YCcMms4LkgELa37/fqOkiVbwHr3jhhNk225C3LgszcVPCl4mpPcXOnTbefXC80ZqTn0uGG5ijMvAwQDKo1fNd3oasbYPhg6GMyuj81VkhtTh9oin65F/ApgNyE19EaZ2C7mTR/iMssJo4vn7X88nixuUVIE3lqWqamRuVv6Oj4VdSmk9BpfpcYgfU5GzCJron7p5vn6ADi5zKCB/NYthOnBhphQaahmzmemuDGFYdbq5YChhpE+OSviFM66g18ZZFxsrf/umSVrPD2sCNL2EtX5WUdRD0ExRs9ghbdwwqZv6zyy6XEYhV5OZR+XIX536bh/bUSJgdVLnNlZfPOVWO70dVHSgQi/8yIUikN3IFCzaTw3KSB0kgJQG/FKCDum0IEO27GGu+3/L5gB0S0xiBngYr5fdrABWlaMR8gypL2PvmW8G+iIYJGWW7VFRG6XgpwD6gZtf1gTYEA/Ox8PWGuMaT1pdHmN06ubPPQBa/VVA7W8OlRZQ9EDJG+ul02Us2asE3OiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZ/Kb8um8DAFoefA+bIGiTbmwExFCAxJYh6JI6KPePxIuakFy00lDE9GanoaVHZtbbSD3mvmJwIp2T+qGsY6m2I5T6VcfxlHAQFtXl/53HH8zi39mhiDpiBcI6xh3bsbOBDekw1gX0ZYvy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMu+RNAagucaKVFlD0QMkb6jkVVXz84g7lNz7Ynn829TyZL2SSKL8rYnTy54Ouq4E2g1uT5qIfGpcRP+C/1wxb106X0QbgInAHGPbG4bYuGlmwW9iiHlNjGUxsiS6w5TzrY07rcP8MzL7MABHaEHTv7iUoJf3Lz8Rmi86ql9T5WeGzrIzqfzMOSEPPl5PbH8grjzU9/c0Hc1Z8LjLxV4aFo8nr+ei788bEZAswKrW+p3NVZIbU4faIp6cQF8rEo9mRfRGmdgu5k0UTloJES88YVmuzqtwTl13MbqH3qqgQ2LcL9HJ40QoTvjAtCoWThn5wGrpekE/zBp7SXpSdj/z6B3HU4bFnMB+7HLeoO9GaC123gjXOEok0S2b38O87wDsDGPbG4bYuGlsXMfegnqYE+4JLCaXp9PTHj+8Z3qfmldDjCgNQSVdmT3X6Gpo1Ecw8UpcaByMV/KfpnYcUGthjUYimj81w6Dmzl4gXOzopOvp8LjLxV4aFo8nr+ei788bHboSUxH8NKAqvvciyv21W/vioiv24gbuGDiue/A6c+NupY+tBqgxbrCjwhkWzsEz4NBQUlLIPgxRj11ybcnTsfvzsxemkN7V79P3SaEG3GmpuGgiyYIJArmOPn+S+0DGi5YOX7gU6yaLHw9Ya4xpPWgsUXTkqATg/JQKNagKx+zjWRdmuPu52FH6kFBR38jOHT9cMkv92kqxtUITcVlKp3OBJt2vIZJkI/MGChbu+0GtYc6W2/xb8szzlVju9HVR2qu3dxEb2RCzdyBQs2k8NyLtByIixYAFmgg7ptCBDtuxhrvt/y+YAdEtMYgZ4GK+X3awAVpWjEfBac4htHVSbngihxWWe8JGUEIhjmoZMKesBYLB37rmkwhmF4u9UOwK+gczzEVznGKb2rBUoGQrMw43YVY774KSFYa18FP5By6aFOWhvQIMdb/umSVrPD2sCNL2EtX5WUdSx+9HIXJPPKLZr6hzUUudGeJ/98hFvjdXAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyMj1EomkBOXDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JqcaPVy+xEfDLDtqXO0KBr7e47YjfAI3Rz1VceMecD3u/XI6enqPtQwRXCjJMgCu0JQ9JVVkEDQ5+hzuLqeZjg+oEnKRDNvaBggzANOaTJRvY7JmxT5xAA5OLM28eBxmFaym0Pma3C4xPVVx4x5wPe79cjp6eo+1DFdh7Vv+tcqGqeJfESvt/thTICkvgs3qpx94lV4EiyWa8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAjUSjYfC4uFDlBO2gA/2F8Ezp6aycueeIKLVRP+gR5Dnh19obzwClQGjk/na9wIajtVylrfHRe3AWCwd+65pMMBYLB37rmkwOMKA1BJV2ZMMcppjA9Cl0v6vJjrxsKbfclm3bLTeGo8bmKMy8DBAMqjV813ehqxtGQLMCq1vqdzVWSG1OH2iKenEBfKxKPZkX0RpnYLuZNFE5aCREvPGFZrs6rcE5ddz7pTPnxlkJXnC/RyeNEKE74wLQqFk4Z+cBq6XpBP8wae0l6UnY/8+gdx1OGxZzAfuMHRKiVWorhuZW8Gn8vZC/dQajXlnLelg1ph9EJwygYowdEqJVaiuG5lbwafy9kL9S0Guq1FJHyvWmH0QnDKBijFNXd2820FOH1MVbgl0uWPUGo15Zy3pYMUgrKVu7yxRvkOHtvnsaz+zpuBjY2VybUtBrqtRSR8rxSCspW7vLFEr2R8N1Z4tWLOm4GNjZXJtPzoJLcMc7fFqh45JT0ecIpHPqrmw6kCTNJnuxRex9JY8oLDldgeuhlWmcDZt60tHLqIynEgHjSjMr0++HVT0C15V3ArZ8lWJzWLYTpwYaYVUoQOee4iJql82pIEH2bIPQmgvwJrWmnMQEqqYcFmbqLlg5fuBTrJo8G/YTAAVaBxy25srDJyDqIfuNho6mZBoS3bcyFj34MdboTyYFjhMlNvXpVJRtEcMCDAM8YgYDHjvaU6w36I5YFEAxF+JRlissfD1hrjGk9YETOWt0KBunDb9QuSHDNdeLcM29yBS0gtqgw9ADDPXNpqV2lm+2KZPRpo04L/I9Wcb3DzPhGSx6xALwey0QJPyhK8ME1s6ISebx5YDboEkQJhv6/xjZMo1o292Q3P32gUQC8HstECT8ly0YDxdzMK9W36t5Feex9KnPsJ7TwWzjMox5yiBbM5R8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+Td+E65KKgBL7mWvAnj1kYGjltCQFv7YKq/cDwz/C3OGLWtik83qahFyjS4Snukd6KkmqRRxoXb2Q6dU/zP5/JYA0TFyduL3b3qXPgh8X2M8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTzIvfbn7cn6wWVW0lhSZI/MMV0T8SMBWoZqzRz4JUZgmg1uT5qIfGpbKRdtogVez5GBZLF9KaZf6hkWxx090p8bCdTN1xFNl64t/ZoYg6YgU+4CClUL5U7hD8wPgQ7I4rsrI0o79d3HwlW7z7hm9iMv7rFS/YCcMm07OMBcXG9xSX3tdMOid564wLQqFk4Z+cjv3T3VnuhyxoGNLphMTV1UCGgMvrUkxxS2S5xRKA/eQnpv7XU6I3MWo/C/Sc/Sw/RjkU5vVrTtnvHm6kG96tzI93uu6lFqhB2/lkfrUwp6unNOR1VEMsPdS/uYXGyzsQvI+Z2ykUEdiCUGnKO+XO3RZVbSWFJkj8KgqfiL/8Z/dZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk5ObRzSM0cQs8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/FtMSyWZdtrJ0sDZ08pnFlqAi5nyDP1E0DJCY1ysKYHw/zyP/2JjkGQqHK6sWOC5+jy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPMi99uftyfrBZVbSWFJkj8TwAvW/GOR4EEyl7Jk0tKxqw9aDoVJ6fI6m3ZnKEGKjxtyYLJ2UTCoEIGkWjGk/dN2NO63D/DMy+TsRdHHlLuehdBvp8HaC+IDoB9whnnmD4nVgT0sSWwXGBMoG4F1/DFs6bgY2Nlcm0gotVE/6BHkDi/OO0O92Vu9215oa1VU9wnpv7XU6I3MWo/C/Sc/Sw/XpeXf1BiF80bVCE3FZSqd1uForwHiv5gTlJh3HQ/USYDDmo0qbnlti3DNvcgUtIL7wjmypMjbn3OVNoVzwn9NM7Y8Hd/UcbDV/Dycx34jdymNuCDaK9hoKbJDR6x5+oCExiPl2GBtgtleNlro7TPYMdVtoj3JR+qqISWRY85O5gS0xiBngYr5UAebsU8ZR7rQBa/VVA7W8OlRZQ9EDJG+j7rg1uuZU/dUG2DfJCuq4fy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNbwb5RoGmEZTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmHNadgaNZbXaByvXx8q+/QYphJmasRYuaowV/HkwsPCy6soU1Oc+1+NzNJkrs3yGNJYnxoB1kWmjygobzeeizJnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRy1qOiGQvRf+TrpDzHd8oOsh51Z9AaBJF3bN1CorWVibHBES0Mbd4vk8gIgRYEZiZBuo7IMYvjPym1nHdDsqfD1pM2TeZcsT0LJ3ow1ybKT4xgzCCGBflKmdEpX0cGoCbU+beGTHH2e+YRoHfVlH8TWCd6MNcmyk+M94yYSQwDyk0LQQf2XIS6XYwLQqFk4Z+cXBX9VO+RiPDci1cKIgfXaWRXZEp4UN23K2jqpFxOs9GiGZg07RJrMG7oZCQIRHOCh/Sf7KZ39OBmfs0s+9ZKEGpGPxRfAM1o5Gp+6lchOCaSSyzK8jRSyeL+qKSxS2MeCQmGKjdC1mVcKxAGdxrv7OBAg8JDou0Za/8wzBkrwCwo6crItFBuR4QuSKod9EjETUYCJpCW0hRQ6j2NnZrebIkJLTO3QsxL+t+OOFWOPa3ng0BEe+B2qnmptXwlS2yxEGavVPSi83WFy44jk47FMqZ4IPHG+DQH8+gwnPQ6KIJzeXSqrDQ5WLjzGEFdq/eyng/IP1kk20gX89NPrPpulNIC5/61ah9946W8a7hPk6lzXbt/ufjDdL4KOEGyxjmk028eMkOqhfcGYP6N/hbx1ag18ZZFxsrfVNpdHQ165KKG7NBAd3NJAkNhvIgnzBGTOnM/V5YMUuKoNfGWRcbK37PGvpLKJo2LW2fc4F7uH5r/Q7zpsr2o8RGgd9WUfxNYVEbpeCnAPqBm1/WBNgQD87Hw9Ya4xpPWMUHPCYaUlJiCUGnKO+XO3RZVbSWFJkj8oeVj/zANz1rVcj9aJHTBnvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk2wB+7h+Ops6cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHIubmRhqHvFkJNsYQxKFurCzc2icvd1bNFj26I8Y8vBzUxobaMEtKAI1tyKzfoDWBby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8fPd/Y2AL5Ter3DwGGOTePgfQFi+EaXvtJTOxVf6qMnZI4vTKyHBGc9sFvYoh5TYxuLXV/xCun2Y+ro4JhRiFWBNz7Ynn829Ty5LMadr0fltxj2xuG2LhpbjV75HjLUWU6oD9Hg89bFPdwJ2/0bXhnmaKFqcgCBWIkeUCxFioUi3fzR8aE3Jj7YgotVE/6BHkAqCpAcEzuEVLeunCj9lagooAoEm5Cge7xxHLifkb0sGJyOB5VW4JduTsRdHHlLueoWaelxFDnQYq+9yLK/bVb/BCooBKNUp7huYozLwMEAyqNXzXd6GrG0dK3Q9osuKHgLPP563bmahoq6LEWNoqwIwdEqJVaiuG5lbwafy9kL9rcxtJeIgD10wO89C+dp7igIuZ8gz9RNAHChBkRHlDB6CFfgvXHzSEdH7GmQwvAH5ZL+814w1rJY0gp4EJb87tWRXZEp4UN23hZ1rbaiayrtkGrgi5QFP91U4MDKnvD/ZL33eNzFCZOXqnqe7tkDQnGz8/3OvySf9oj0QCQIThh6MjytNhtsysivfikjTLMYb4J6kQ+Mcj5qm7gT3Uzcjb12Qg2Tnxxt3Z9/GABKylFYJWNMwJmm33EbQFv18ouev0+JeW8eajyGoNfGWRcbK3x5J+bZm07qZSwWzxdDa8rno268rga5UD48hz/Du+SoNpmFERzayw5MMvHoJrtpKj4i8oPtPoxRpLWM3ao0bLxS+uSw3LyOTo72T8Mvr/E4MwFgsHfuuaTDyOLQthF4BMHgnQBLyKdR5qDXxlkXGyt95iPr6syuvPfc0GxzRnJCmzTcJMLzhnQauuQ5+lUMUkhQy3bNosCBoenPTtAYOt1Zay9sXfxhZ5MUkSMtOha5KIhjfAIQdvZNi0B4Bp5BIlBEutQbNq7SE0bVche/0/U3AWCwd+65pML/hO2EdDA3tAAuJ8wpQLNMIV+I0T08S294EU5yb8ac20tzZVO2fSqDAWCwd+65pMEI9z8tyPfRN9bVb8PYeGSsKgqQHBM7hFfXj7OAFP4cDgV4MK3d8s+6oNfGWRcbK33mI+vqzK689QKYMtgWsYgHNNwkwvOGdBq65Dn6VQxSSaFwjASZ6Ard6c9O0Bg63VlrL2xd/GFnkgUgR6fLE+aciGN8AhB29k2LQHgGnkEiUES61Bs2rtISOQez8556vRMBYLB37rmkwdXpzL7f39xMAC4nzClAs0whX4jRPTxLb3gRTnJvxpzaNg8+YgYsDg8BYLB37rmkwQj3Py3I99E1xoz8oTOm6aAqCpAcEzuEV9ePs4AU/hwMaBrA70QjXNqg18ZZFxsrfeYj6+rMrrz1q3I/rgudS0s03CTC84Z0GrrkOfpVDFJIZ1KS9fO/ljnpz07QGDrdWWsvbF38YWeTnZ+AQgx2ovyIY3wCEHb2TYtAeAaeQSJQRLrUGzau0hJ2cB5gjwdDOwFgsHfuuaTCEYjk1HJ6S5AALifMKUCzTCFfiNE9PEtveBFOcm/GnNlgnuOfxkgDmwFgsHfuuaTBCPc/Lcj30TXg8vnUlwXTsCoKkBwTO4RX14+zgBT+HA4iV7dA29zlkqDXxlkXGyt95iPr6syuvPQGTPBpaWTEHzTcJMLzhnQauuQ5+lUMUku1a8gtert7DenPTtAYOt1Zay9sXfxhZ5BRCQRWg6Tl5IhjfAIQdvZNi0B4Bp5BIlBEutQbNq7SEhulFGsOWe5TAWCwd+65pMGVuIHKqil4UAAuJ8wpQLNMIV+I0T08S294EU5yb8ac2BwO6LPvtkYbAWCwd+65pMEI9z8tyPfRNXWxOMoBfj1AKgqQHBM7hFfXj7OAFP4cDLr26RiTh1IioNfGWRcbK33mI+vqzK689i3CJBDECr/nNNwkwvOGdBq65Dn6VQxSSyHBoYMjjH896c9O0Bg63Vr2rBUoGQrMwwWzRfs2dV621jYKECFFWP3FSA8dGCp5/3PrvpvZhM5d+K27BmNPaPAs5VGyYytarcyLHxo+Tln43hof78d/O3LWNgoQIUVY/5/30NCiF/HHR+xpkMLwB+WS/vNeMNayWL8TLnOCOek4Q9BMUbPYIW3cMKmb+s8su8xB7sp62pU2nNOR1VEMsPdS/uYXGyzsQvI+Z2ykUEdiCUGnKO+XO3RZVbSWFJkj8UAuCKeQIkbXkZJpKoL9z2PL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4Ull/LbH3nT9vq4kTJEDLitDbjdUkbb94bFiEQK5urj1ph9EJwygYpSBYRmj2zA6L90/v0Oz005grgujKbUrP8dYCA0bKI1vOF9KIYp+WdBG5ijMvAwQDKo1fNd3oasbeh1qQ2/ow+ualhR2xuroxkcRy4n5G9LBnPKxSUCjyIDk7EXRx5S7nqvVBp3gPhas6+HjxaB4B74rR508ZTGndEVEQXwYVOWpjDSY/eyTJK0BVA7arIErlklX26L3zEegzDCDFQmIOwZ1/PJ4sblFSBN5alqmpkblaFJimp63yp5yxcpQMJTtpE3b+h10OFk37Om4GNjZXJtSAVWkS8aK9kcEKnjbVUmOpL6FnCfwWq35iKqJZa0JmqC1yLxNPJliDjgq5bS0R06CqC/0emKpwkBYNAncoGkg5LFaicXcUrcRyTn9cOEr8iAbAWZCTK1uIMoNZA6HRxHFF7KRusJndFXrQ7OlVQkBwIuZ8gz9RNAridbypl26tkayBN1AGV5UfaT98RFxF5+BEzlrdCgbpw2/ULkhwzXXmCneg2fDdEd98yqiYko5XOp44d0tslT4H6593uYeK0iLH70chck88p41PNoccMihLNesFVE0RLxrHEBNYVWkOfy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JrcNMTuTwO/yimthJf9cGjaosMZZ5kmzW1nKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTTjVNpLzzzy5W+tVfWZG10F/wIG8QVFW+wElAv+IbV5SzZfqcOBG/ppDRDzKAm9d6wFgsHfuuaTDAWCwd+65pMMGeX39/rGN/M2vuo/UxB5xxX2xf0wa4oro4RcXixEUsA1xw479csToAIPB/3jIorpCBmYips0B8lBnDUMeY3ufm/fPgGiWhA5T45oE0FkHVHnOxXUsNyVZtaAmJPHytg882aMpvivJgky3wO2lkoMEwTXHnV1R1EmZlUP4sF28rW36t5Feex9JPTlGVkMDOhKiXIDk2erir/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHYO2fkMaHs6pDRDwuChd04SYu4KqWvjvGBna6Apbqv55x8tfLfHJerfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxH0ff2y5/aqubQodAFlJaNogjdfCYMdiQIe2amCghUb3U6tUPC7yY6WtFjD4NqZt0tVr5ID5f7EkbmKMy8DBAMqjV813ehqxtawR8GOrsKYmcia2nlyFYDvdteaGtVVPcG5ijMvAwQDKo1fNd3oasbUKum6teU2O0pAsce8A1ZdTkfcRwEJQISC7MoYZt3WznJ3ow1ybKT4znzu2uMSHUto/QVQVr/v286Zu5vfZMuusbmKMy8DBAMqjV813ehqxt3VEWkAG5j0ShZI3RmFz4q/FdVn/BDwXB8RBFcaRys7vnxVrQ0bPkLhuYozLwMEAyqNXzXd6GrG3D8MjB0QTMJL90/v0Oz005N4aH+/HfztwnejDXJspPjGDMIIYF+UqZW8DHVblvz5OMC0KhZOGfnM25Gciy7U+xA1xw479csToAIPB/3jIorjtROBJfLmguDPbkBzQdmF78n5Un7wD/4QNccOO/XLE6ACDwf94yKK5BOvtSdJmVOgGdEO7evJKa9215oa1VU9wnpv7XU6I3MVEQ1GYn2C6+XZCDZOfHG3dlcms3tP0my6A0QOlq7Ui3BXhXwPnjdQLr0Jr7PNO1GkL2TqHljvVfc1esvhvkCWazVzgLR/UXRjxpqnraFR1BwFgsHfuuaTCBg3892dJ3ZidQrN0m84Wjkh+vZ1RFSK0xfQfSHVsrqLEddF643SlE8Knkk2oup/20JprEbgTDXJDRDzKAm9d6YWaM3bdub3Dj5RcgwgjQhftC7lctD1rlISPML1E4zr/nQscv0J9FWd7WgwNsWJ3RXfJXyfehkB9L1ZlQy2vCPN1M02WG+cy09KUKeX69msxu8MzZDeX+JoutycULOw+ZGGu+3/L5gB1kjv3tpLEAMVrRl48WpUyYwFgsHfuuaTDP1xMkf6s/FlPs7tUKNMLbES61Bs2rtIQLihgwo+46jxhrvt/y+YAd6DoE+kLtHYUasmqulKUP5cwf0/YKm/V+ZXjZa6O0z2BK9eQ9psKy1t1RFpABuY9EoWSN0Zhc+KuANvWFrDmtlKBzPMRXOcYpb5lhdorn5WioNfGWRcbK3wTZmBjj0WyD3XYyQev/JUKoNfGWRcbK3wDy0piFYdZI7k/GB1YtTgC2QlcU0Sptg1j4WZkhe6YPGGu+3/L5gB3tJ1HzQxcqyRJ6e0BuxmJmSmjqyLPYB6d6oX+dtonMp9EWDFm3GSg5qDXxlkXGyt9bVYJxwK30C8IkvlgTzutEzJEucl7DC1hhVvIobLjnnOGNJuPv01Ucz9cTJH+rPxbYtUJqWqw4aTtROBJfLmguT7yWfHQMZqTAWCwd+65pMNZkHksjWl3Lwyhge52iavkvsTNisdrScqg18ZZFxsrfLcM29yBS0gscvViXJZL35M6Y0n7XqYAltY2ChAhRVj+dp+uGhmVtQTFnIRTgnaxPPtjExlWAHB33awAVpWjEfMBYLB37rmkwrTIP0x/AMDCmYURHNrLDk16JN6CzdglfB99rICNp8rSdC+dXQv00aeWushzlMVJxP8eTOG3K7Y2ICkiar7IDzHXUXy0wb/1S//ySbxuCBgL9su6TMtvxEzHiakW53PSIOCRa95Vj400x4mpFudz0iE/Jm1a0LM4cMeJqRbnc9Ii7GlmnqeOvn72rBUoGQrMw43YVY774KSFYa18FP5By6aFOWhvQIMdbnWj/g+hiLiQ1gkX/YMuNfXO+NS4W1p/zffqlppcnQWZDlBO2gA/2F7UCv9jAZMCN/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHYO2fkMaHs6rMLppaM2c+BLtUcmQpEQ929PAJsuVy0LBZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk041TaS8888uIZr3wF20l1qpX2t9XdoqhYqAxogQAo88mVvBp/L2Qv1hwPp/rG21j5h7XZedBf16GLPonSlUJLsh7ZqYKCFRvQ0bf3djsOF9k0D+UTm5vGuzpa8vIWCceKpgPjy26nTKIe2amCghUb0NG393Y7Dhffx80GuLNC1JAlZhMaIASUPrV76sflDlOePlFyDCCNCFIKLVRP+gR5C7R8nRAjOAozq2JQd4nTQPTHQDaku8kogh7ZqYKCFRvdl4QVY1mQmbsnMRARXKuj4KCNTTQuUYDBUjqW31aQvzIKLVRP+gR5C/txBcb/TY+PseEyrS1Tg8Sskg2k4ClR5TGyJLrDlPOuKMV9pwNoyeUQDEX4lGWKwgotVE/6BHkNZkHksjWl3LNrBKvbSWGzjHetHVooKpygNccOO/XLE6ACDwf94yKK7kY7HUX6r4RL+wWkWw+s+WjBtqTXhdQpknvS/Z5hBNupOxF0ceUu56aTVuDO/5fwJYBC3CNnLh5avvciyv21W/mlYqV8JzNNQgotVE/6BHkHMtXCRjlP6Sl0bajBE1p8zNzaJy93Vs0Ven4UCILaaxHEcuJ+RvSwZzysUlAo8iA5OxF0ceUu56Dk0UFQp8G8EJyS23yTu2xs3NonL3dWzRV6fhQIgtprE44KuW0tEdOkNxA9FrArjvQIaAy+tSTHE37Nk97b+6riem/tdTojcxURDUZifYLr5dkINk58cbd2Vyaze0/SbLoDRA6WrtSLcFeFfA+eN1AuvQmvs807UaQvZOoeWO9V9zV6y+G+QJZrNXOAtH9RdGPGmqetoVHUHAWCwd+65pMIGDfz3Z0ndmJ1Cs3SbzhaOSH69nVEVIrTF9B9IdWyuosR10XrjdKUTwqeSTai6n/bQmmsRuBMNckNEPMoCb13phZozdt25vcOPlFyDCCNCFUaHik/PTq/NKySDaTgKVHqAD0rdqQNfFws2OcOiCiVrBrSlM45ML6uQLATUJC6mfdMYIWZm1M+Eu6hrt9WoON7tHydECM4Cj+ro4JhRiFWB5iPr6syuvPVg5QRrrnN4GFjxv6zKMQVbY28sSJH97ZFegtTbhYyK7HmWvyhCceuj4mLcm8Rds6f2kAhdrEF6meoh/nD7AOs5JOdxG6uJZXag18ZZFxsrffpN2pfisbIcMhU7cKWORDGpQAz1rxM/KPdIWt/1GiPQuuKDMeEVk5qQHP4VQDraY9N3EtLgMdeVzLVwkY5T+klBGmxSbLRcDRwJRb7kHTYjAWCwd+65pMJdaByZavr6Yqee6wiB1Vn+WWgSCvNJaNonw1by4E5VnkNEPMoCb13p4Oyl8S5kmylo5e08NAzuUwa0pTOOTC+rCfeoAKtZ9K78MfJim5OdRWsvbF38YWeS10kqvJsPZ8l53Qlw6WgCmIAWD3mzrGzuMuDw1j6kUORhrvt/y+YAdUdtbDPzMjtK7n3/2AIYw6ONVAQ/EiHvdcFCXQb8MaNX4zSrs37+G7XmI+vqzK689GSg4TcxYEi0WPG/rMoxBVp5Ip/qkIkcoV6C1NuFjIrseZa/KEJx66B/LlZxyh4xv/aQCF2sQXqZ6iH+cPsA6zgubj6d7drewqDXxlkXGyt9+k3al+Kxsh/jGO5x9/oSwqee6wiB1Vn+WWgSCvNJaNhx1JU4jZ89qkNEPMoCb13p4Oyl8S5kmynXTsl4IcXqPu59/9gCGMOjjVQEPxIh73RZD3ziCX01Y+M0q7N+/hu15iPr6syuvPV2NzcLgpCnH0OGbUWpddRtqUAM9a8TPysmJ0alXzSQILrigzHhFZOakBz+FUA62mHlLb7oisLXwo/fytCe2lD/BrSlM45ML6iKbWGdK+z8Dvwx8mKbk51Fay9sXfxhZ5PQlnhUnstitLzcwK2ZYkc4WPG/rMoxBVp5Ip/qkIkcoRriuh3h0YN4eZa/KEJx66MVugnYKok7RlgkhBWyd7S1zLVwkY5T+klBGmxSbLRcD0DyJ7+iE257AWCwd+65pMOeH528NwAgyMmHf3extpKF8UkhzEaW2hV1wyyWXo5sBjS9hLV+VlHUASlQboJTlvl7TJuQ7Wnq8qDXxlkXGyt/7VEXBm1VyRLJzEQEVyro+4SSlnUTC2QhE3tygC005pNEFBPqBPlIHkdAtn2nlpC3fATBDECOXVrinvajFK68oSvXkPabCstZ6MITYtEeyOVS/OByfSKxS/GJjLnJs0Mm+OQY27/pgEFP4K/8MgfJgghX4L1x80hFb+kE84+RXOuQv3OCJL5J3MX0H0h1bK6ixHXReuN0pRPcqL0rSOl2NG2bhymYiei+JvNcwrG43Q4OiZaR9YS1r3VEWkAG5j0ShZI3RmFz4q1izx0rq4zjQqDXxlkXGyt9o+5jTK0ldzOdT8uEX7TAh5GOx1F+q+ER+iiHlSS6CcCYu4KqWvjvGsR10XrjdKUQXDzQ2rtmEAEKW800RllpNRtAW/Xyi56+YNTedzyCk1mQkS5VQoNqh5y0gNf52uF5rHng+ftP8ApDRDzKAm9d6UAbSjVcAROljxkwKDphL+zQ68/3TNPUeGmM340wuvpGzpuBjY2VybUr15D2mwrLWZBq4IuUBT/fWZB5LI1pdy0e2kAi0D/WF7Gfhw9lEZps2/ULkhwzXXoMqS9j75lvBvoiGCRllu1TFnxKDwQz8Xe5PxgdWLU4AtkJXFNEqbYNLcAnGSqED/MoFnr7X8il+6wKNvZXcJPSRjGUlDW9J9IKsSYdIp19SBMXQbpHQZoh+GbRxWNOKSWzdKQeHYiRcXm8WVmVKr1dabgZgHDnhf//8km8bggYC/bLukzLb8RMx4mpFudz0iDgkWveVY+NNMeJqRbnc9IhPyZtWtCzOHDHiakW53PSIuxpZp6njr5/HVbaI9yUfqqiElkWPOTuYVj74zqI4xqHasOuKOkW0gHBJnrnSFtVEm7Cl/JGm4dR5Jh7+id8RsVdyzdSCUW9Q1ugrRKjpvfLy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNsAfu4fjqbOnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRy2cglD0l5pz0d23OOOc6i5TUlCseUouyXOObwLqQ+MCTr0Jr7PNO1GpdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHy31CPaOtq8vX7rRLSaICkiqam7N0NVoQNrxW61GNIZezZfqcOBG/pjB0SolVqK4bmVvBp/L2Qv1hwPp/rG21j5h7XZedBf16GLPonSlUJLsh7ZqYKCFRvb4KOEGyxjmkQhQaHWyXaE/XTsWXSfnK7Nr9SXXkbQV6mVvBp/L2Qv2WWgSCvNJaNoZftVGNICmJMDq/2YwiEFyaVipXwnM01CCi1UT/oEeQ6DoE+kLtHYUY/ClpgC9udFliBO2/l/L+NmMm0JaOTmke0Oo9ZJ8VNSCi1UT/oEeQRbeIqZ6IjmuxbiwtjRn/vXcRiwtwdKjj+DyE0mbj/KcxTV3dvNtBTh9TFW4JdLljNzGIszx1/8cFumLOV0AfeH0La7jRIwW+Qg13joP1VKnXbeweNY7qyRXzD0fTmuMwtrDUxlZER58ydmgVrtpHYCgDAMvpvn5xzquoVBy1c33xwRugOJJ4Aag18ZZFxsrfOoILf9Ku8xeSqbONDs1eLYpuINZqYyRBQvZOoeWO9V97AaVpm3aMSfBOOZikY94suWDl+4FOsmhxaW+qjMrzqzyu7J799H0w4yI+9rdKR8O5YOX7gU6yaJHHobpjcJk1D23f5G3UlTIwTXHnV1R1ErOm4GNjZXJtSvXkPabCstYgBYPebOsbO7saWaep46+fFpziG0dVJueDKDWQOh0cR3ckiLyaLzIZm3t5LPWqDZO4+rfuZAHwHMYdkDsa4HYpGGu+3/L5gB1hZozdt25vcKg18ZZFxsrf0txNzmLMS2LCEyVo89VIMtHdHvTrpEi24SSlnUTC2QiRx6G6Y3CZNZajP9Stw42Z6alrjeeo4zF2cn2ZqVXC7gwrjVQlO79KzumJRJPoGAFz03ZuDCSed+EkpZ1EwtkIkcehumNwmTUPbd/kbdSVMjBNcedXVHUSs6bgY2Nlcm37cwsO5GXMRxpK5nLm8MCcmlYqV8JzNNTWLm3eKt4OT8BYLB37rmkw/svlj26sYrn5ZZc57rJAf+qBviJuKv7QkNEPMoCb13phZozdt25vcKg18ZZFxsrf3Dh93GlAL2IgBYPebOsbO/XpLehyluKynmWvwZgHfwqbSiTrhKqVr7C6M3JiYf1qs6bgY2Nlcm3zEHuynralTQKB52gK4D7dlTM00GfKTPHqlCiT8ZQpz+Lf2aGIOmIFcTk2kNf5UYKRR2sFbVXrHIWK9eVp0g8FdiN5TAWo6gFMEW3IaM8FXs/UMS6yM9kRakY/FF8AzWgwp+CRT6hA2s/g6GNg8GsSxyi9zcOSi4d509PVr4xpaUYiuUNV6itNL8VQN6IEW2hoyglypuIbeQ3+nyFHt7514Lwn2kgjW7eRjGUlDW9J9Jfvp1KNdrXQ6ZZrv6D4WWduz9MHEdbvNaXpiAQSMAKmSvXkPabCstZNQgUP9nS05j8Pk06CtQfz1XVfvxw0402Q0Q8ygJvXeug6BPpC7R2FGrJqrpSlD+XMH9P2Cpv1flCtASy1G9/aRN7coAtNOaT0AshkkhYDqKAEjYO/0klvPbbVbFC+fvSAzmx+qeIL9Rr77gjlOwWwWwLjA86VFcuzxO7EBtu+KMDkgWNUu3GLGcwHqst2z/p1jXfwXaQY4E9jmZX5rNVj2K6hMdSPTRz//JJvG4IGAj3MlDUftI0mKYXTmQMKxwu+YOX8ovzVo6FOWhvQIMdbajkcM0HTJMUCgedoCuA+3QWfWk3JRltaBLeuwy87CDPi39mhiDpiBag18ZZFxsrfJPB4LhfsEBWuFtdiuhrvFDl/R+s8OZ4S5iKqJZa0JmoI5HvehvWs2eksTDzC2lINxbanyvez7ZioNfGWRcbK36l8+09yWfa4dySIvJovMhmbe3ks9aoNk/qvwjECo0z5trDUxlZER5+ohJZFjzk7mBD0ExRs9ghbdwwqZv6zyy6HfTR5ca0q0sqTrrCT4sjJMsh7fPt7Lw9wRvkqg+qgS+pAOMlD32PVlXJ27XKaYaoZy0J0dq63E8dVtoj3JR+qqISWRY85O5g2UfFJj6Mr5CetGkdY4p7z1tyKzfoDWBae3p2HZyfx+zXZRCxKHjf47CaZA77djWHEQXXdm51jXVt+reRXnsfSMS4IH7UtZQXL4LoJ7AAs5pdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln5Ojh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFlxkhtePyRCkoYdb2T/ESwD+7VHJkKREPdvTwCbLlctCwWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNONU2kvPPPLiGa98BdtJdajYXtx1X2EmtA5bUdB+JOzs5tcEC/0813E/cHQBD+zjsh7ZqYKCFRvdTq1Q8LvJjpa0WMPg2pm3S1WvkgPl/sSRuYozLwMEAyqNXzXd6GrG0QgJrD97IYJF4Y5nUBAZoKO1ujAF54GXYnejDXJspPjGDMIIYF+UqZ0SlfRwagJtT5t4ZMcfZ75gt5NKr9oEMT5v3z4BoloQNL9I1RRP9vPELrkXX+HWfiSyNhgxLmo/P6H74q/g+ueJWzEJUWDeX1h1VhElid/3GCGwh01FTvH/IwXTI/4GlLME1x51dUdRIUUFRMWNwvMTB0SolVqK4brxcnvbzsaayEIXIVJEY3hMnCDe8WDYebmohV6hEoPPlBpfpcYgfU5KLS7aKQw5TPZmVQ/iwXbytbfq3kV57H0jEuCB+1LWUF0ePc+MKeFQGXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+Yrz7xR5vZrL0KyVEYCjTvuE5B2e4Roiw4bWnDTum0T3DsMHTjZeXWMRGgjptf/3NsvpGvZGvxi8D+3Jrr+jnia0gl4KH8XY0B+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7ceb9kf9ou0FunEd7oLfOMjkopFEfOCZur7e5YejT0xMiJfbXA7yKysEBTAa6bZhbdhaHEU7wa9vmJGyDGfAPnbv8t5sKA5ar57o3iO1GhsAMq5V9IKK+qZNnhGh578ay7T58qP7jfXrbMRSrTpupWcFmUMNY9FzR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/X0mFXQGDwUBfxxgLW/DpkietI52dApanS0ZwazF+DSia1Dv3sAhvWmfnNRqgv4UiYRGFaybmRCMZC/dfqF4dRbJ6YdRjDzAOeTI6HE24diUSVDOqZhdFAgiU2dFg3BcTQ+f9WA+wEPXz4emIpYW9nYIvd5WGTwc8oAxG2oU6OZ6I249b8IOnTHuhOXTeaFEQQTKhkCMCgMo/ooX7TTzaaMw98LvuzZj3CoqtxVnEmJPt8FKeAB5Wnrg88kZd64icY9sbhti4aWpfROrNVR+4+zNzN8dChk+45+LJbh+Zz9twDTVLbzJzRos15zAoco1aMBSJe7qIdqxj2xuG2LhpaUeLmv2Acxprg7fSQ3yHAQ1VkhtTh9oilg5rxIJ4tAlPhoiL8D6lHOdGBl+KB8WHOWOO3YyOCUu9ta4sVmII1I/JyRd77vY9sVw/kfraBEVHUEOxXUjh+ZAhNRP2BXtLthV3+GZxFyhYyKwQJITwh5yjyzpXwhGrlQqQm1J0ygC93weDPh/vl2as/WYVh76LxVxXZny2UoGXdmGxc1LSGuFlVtJYUmSPwVci0IpH5N/sY4Wrd8GuxqKklPVvhIMMBWkusaBbGR6Mct6g70ZoLXbeCNc4SiTRIjMiSwMMxFrKjPlC3rmZrfxUHi6YIVQgiMisECSE8IebIgOoSu2t46Trls1ZJGB1d8EgNGoYoA+qiDCbhSh4ey7LOXWm4/mINL/vuShckTsJcuiL3kkrXAiY0lEQFZDtr/9vLjhskEchEaCOm1//c2ly6IveSStcDsSW5Lvgxoxorz7xR5vZrL0KyVEYCjTvuE5B2e4Roiw09FOIbrUINm1EDF+eslQBKQHN4SSnUIgyorD3blmFjTALr+mDevBKTtMEoEICHI/3ng/rAIDuHgOMKA1BJV2ZPYyVp8Sr/Hd8Y9sbhti4aWbBb2KIeU2MZVxXZny2UoGaS9qYP+sefAimp2TZg4LRVt4I1zhKJNEtV47uTlp9NtJBDAd3faz0vD7PsrS7rJ6mgxwPOa+bCZn5irm3wPWUvZ1XWJAWInDx8X7HxOhyMdPr+LN6vnqEqPAS2iXIhuxSd6ekNIuEEQdyBsTm1jDkVOyaO+iDDjApY47djI4JS7hcS5/w+7rL4DXHDjv1yxOgAg8H/eMiiu6OpIWaTfNin30a9louFgO14Y7+Cn7apJBm7ERzGMJ3EKPCGRbOwTPg0FBSUsg+DF6SQqlZ/JIaokFZETg8+0GqIl1nMj+gMezzlVju9HVR1XcKCNrP6FqtGm0KX0TAtkHBCp421VJjrhJKWdRMLZCEr15D2mwrLWf8WT5B6IqhkxsyGJPT+0VN5gsAnZR8JdLqjoKmaa4CBgMmrP3mrF/Rac4htHVSbngyg1kDodHEe0EfTJMa6qIB/GOKNSVEIuFSVduAmgvOVn765kxnY8CJflSbQ/7r+gNv1C5IcM1169qwVKBkKzMKKQmR2vfjvxQBQaaXq1MbsBs51H26/Z+gahlXA/tK2OdHESNNBEBS0D25IqNMEG+nK6S8nT52GwpMgNlQbpC1BX2SE7VNdvUEV2JORbYTEFewOuTFQXEC836fokJVW7b/Wr9plpCs6BdB8KW+lHZr8AyrlX0gor6h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC5phREvPgpvHBpIYeA2rj5kBghSAkob+RtcYPplyneb5FgMEVi6IXblsFshSxqvZfeXR15LUBDW8Q9t/s4jiy19tVJMf5fqF0qOH/tgCkP0SSPXFdmWcYdtUPUy7bz2I9Sx4REdUg030yDo9yxQaQDLTGTCcLhx/z4ArzA5qdqOTH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LxrFahAkPT9XzCterMAWpOmg61dEmrqcrGh5U5irJnyoBYNAncoGkg3cEuzEuWPSs7wr+i+5ntM1vxmfrBcKifqbEW1/PGtVgPWu08ROnR1Qqn4zMQnkt1w8G5+oIPR9Y6qh1DAeJ70oBYNAncoGkg5+gA4ucyggfGnkhHOWLnddxX2xf0wa4olMzMTd2VbLANuF9Szb8bc+z9851P7X761CCcmaBVJKeAkgCwC5BKc0nUCoE+R7cwQFg0CdygaSDR2fVmEyqvVPW0WNAJ0Cwfk41CbBt0r7fJeg+iExCMrmHH8aTIeDvzX5MVJDRgr2AO2lIHFBSgNCklh+v8EDMafO5LdK+3b+OS3cdS8o8J0QWF+uipddfz+Ktywyzek7jUa0K3DhgdSUr5MLZhS3k9siq/Vdf0UZr4iaT6/CfvQaUzsVX+qjJ2Z0TyUy/Al6LMElkDr5B98jfErHC+0qu3MqvnBwhFB5sUzMxN3ZVssAr5MLZhS3k9rxVkKpH1/jYaxMfcx+78nY9zQjfrwajOKVqodDodiFlMsZX46ljmMxwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkziBgjj4KdLpWLrc8W8k5AfVm/e92CoVOcBI7DH3k5rqcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOHEvmurWIn62beZcvOjzS202GIUpT/ZJj8UnERL5ba7KZML55rMCzpg1JxA2QEztfm/fPgGiWhA7BvkETgs+XWmzXE6Su/2agpCbjHIfzrNblg5fuBTrJoSS9mBhKBT1R6rzqK5/ZPz9G1XIXv9P1N9xovJ2mxAzRLvnX2Duhfj3UWKJQ6R9GzprfkM6pnQKu/EUKWXiWm56g18ZZFxsrfsK5FJWwC8hD05wVcOT5CCHpz07QGDrdWrTIP0x/AMDCbsKX8kabh1EzM6jWgHkBNN/+tJh3oy3qaMASA/MemipdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Js7LxFjIAQ5ZENhO9insmxqqn36k551f/It7oX8asLxM8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEdxADbcr9THe05tXUsMiv/i5oyoIXeJbFuwNu9pJr5KepciTUmVl2NyLaph3YSB0q0NBQUlLIPgxU2EM6jlg+dX8wvcQ79a/M2OHAgZShzLsag18ZZFxsrfknrhHG5fERukhPdx7rRe8naoYn9Prc44o4RuG3gHBHIrjgGkXGDFCXqvOorn9k/PSc+YnhH5GrTK+nWq3cqxqoG3GviY1gpyjRBmQQXz8GWAbAWZCTK1uA/XOJfyF1XDY3sCEo28Fct8J/VrU9hea2suxKHYfDbF4SSlnUTC2QiQikNWOVABhrCuRSVsAvIQHLOro5RNCv2GtjkgpxUJ3JDRDzKAm9d6OdubC9H4RMubNcTpK7/ZqB/VS+a1SUsJaxMfcx+78nZRAMRfiUZYrMDLy3+Mdi3vpIT3ce60XvK0Gy/MgFhuQYa2OSCnFQncVn8hn0FpB/5KjA/NC8bR29A9MX1yFb7bH6kFBR38jOG+iIYJGWW7VJF+2OMZYkdNLM7YKWdMXREG8uzB6EnYmkSt62alONtI8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTiY1xyRj7Rgnq3YFFR2s4AFQEo83cZQQWB2LtnGwVQtu0gl4KH8XY0B+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7ceb9kf9ou0FunEd7oLfOMjkopFEfOCZur7e5YejT0xMiJfbXA7yKysEBTAa6bZhbdhaHEU7wa9vmJGyDGfAPnbv8t5sKA5ar57o3iO1GhsAMq5V9IKK+o6RNyaPbKgx5Dmkuk6FdqwYC9caZ5Y5+Um2utZi+wc2R+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7DDf+uMe8gUN484XrEbQGHynBJ8zx5c1D1FeqK9ACVP5ptEP7mnnShBhcHUGm+MHBqTTybj1KQHpgq0LWib305tJtLYbwcuF+UfO3WUUEQAIfbW5xlWyIij639AgtUFbpZgLI+Yp8uL5qr7N0RfswLXrN1j7uCq5790/v0Oz005mlwM6OUxR7etEZK7kisEEh2DWy5n0Tr/BMlZKI/I2EqsPWg6FSenyE7slFv/HsQ4HyC3GItNMeJxX2xf0wa4olMzMTd2VbLAOkoH8fk64raLK+21/PTqhE/840zD0CNxrD1oOhUnp8iQhOe3Rn12Au4OaKttStUS4q3LDLN6TuOl1wnSXp6wTUnIHb41QL9Mvt0W25erGIQD9tcnMj9RLqLq+pLFnqi87cyd9mf4kZkNs+RMmCND0sb2a3wBSeOcjC87P42sm04wO89C+dp7igIuZ8gz9RNAU9SKpkNZ/7fEGUh2bJugDNTSRCRalyta4cMmgMS30D0KDTzY6X5jNFnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZeTgn2ClOaSxLLTiw1XSH0u4JKxnBP4aZT9O/G2/kkc9PL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyBhIwYo4qRNHju25rmiL/V7s/8lKcx1TiZ/SDtPy6KROZ2MLP56m90YzpshkrQRXS8V8b58GG7aywKTkKJerd/ttQWgA0eu+ykJuMch/Os1uWDl+4FOsmhPHFCuYQBxjMi6d7xnQLFrJV9ui98xHoPTa9jgkAF3BIBsBZkJMrW4D9c4l/IXVcNjewISjbwVy3wn9WtT2F5ray7Eodh8NsXhJKWdRMLZCKb5N1G0dd0FhZxxkRSux4sNTCccUbasyqGxXAk6nycc8uuwB+yUmPFA9UcyaQ1b0+xjbVPe5ExNr4Ffkgc5vbuDPmhAtpi4ZmsezOrWWHiu9orqZYAgHpuDvEQyGgeJLO3MnfZn+JGZ/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMj18jBjNADgb94aJ5w0E8cEk7tUrZlVH1quVwFdRFvKNUrWVZsSF79FrvOgzPBTy6+g7q/hl4TBWpu4hMG3CBrDXz/9QgbnfGugCtMuwzpQuZsPEA18kKxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Lw77OF9d4rOWvl9lNkq+IdrX6T0NpFxbWIc83RD0iU+Wvu4K8NlLooedDa8/RTQEBD69i27DxUHP/OYV0R4td6r36mE7lWClZdLuAG7fM0+01lFoJxGMUvpIx0CS7zaDfWeKdmTkEiU3YLdOGkYIVwY24lfrlLE9SxJ3FHwuKI9vZtLL+yybWpx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7zhC1rRWGiQMZC/dfqF4dQAByi4Y+C90Y1qeF/3xLYVjbHasb8nNKb74TviO2/cKNep2m4JtoMo//by44bJBHKGMqnYXNKpFz5v2IOUDBbomml+w6KjXidU7TTGR6h4wnHj/Gt8G7RP99O/uKD1+pOLM2iYdad9RknyG/1KHTI10FBYAslSJ1lr9eDCYFmH8Zj+09kjcmNFdksP52LtI7Vpg9VCN9Fr9fifoxxjcwd648GcdeSei/lO5vKzHCw8N0e46mGOtMc0fBScgXRCZ2ZmFfPECuAdoJOZ9NVWVwgK4ZHVntcgEbOz4wAHRiqX5G2sx1pZ3PdoOtqfRq+Ast9OWkgbcNwpfjNteuhV8KLWNmRrKpqeIm9i4HI/NmS5i1CtKGqLmpTaWPCrRU0PtFpzfWju1MVcAVYbxWnrS7vaE+MzuKY9amSKSY22wp6dcp8DGFNgtD2BMj1EomkBOXDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8QGOw6IbIHiycUN+vGSD0iG+RoZsgfjhrp3E+b4VlDE1WcvLB4etVWny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8U3Ptiefzb1Pgt32UB3TPdJpJmSmcRhCxI3tJ0ixhWZt4mPiVsCvGBfvLBREZBsyKfMRCa9OZHwq3MsoLbO/P5NNz7Ynn829T27ujb3l5/Ve4MNMjb583UCN7SdIsYVmbeJj4lbArxgX7ywURGQbMinzEQmvTmR8KtQYcbQ7CXfDTc+2J5/NvU9u7o295ef1XrB0P6uKJghWje0nSLGFZm3iY+JWwK8YF+8sFERkGzIp8xEJr05kfCpqa3QvrayJxU3Ptiefzb1Pbu6NveXn9V7W/YlVNNnIF43tJ0ixhWZt4mPiVsCvGBfvLBREZBsyKfMRCa9OZHwqB3GqZHM1VDNNz7Ynn829T27ujb3l5/Ve/w4k5Ql72YSN7SdIsYVmbeJj4lbArxgX7ywURGQbMinzEQmvTmR8KkF2xZiXoP0pTc+2J5/NvU+DI9Rq4FPqikamOwvdTgylB6zgflin7Tx13xOEeKAfy+8sFERkGzIp8xEJr05kfCq/2FlDGmKnmU3Ptiefzb1PC0PGbnw3ifWxWyOSK05eZXnarYsvpvfZLlaEv1OfgYXvLBREZBsyKfMRCa9OZHwqe2pvD2SupphNz7Ynn829T4uKL9NtDuP/fRumwA92cdp52q2LL6b32S5WhL9Tn4GF7ywURGQbMinzEQmvTmR8Ku8a9jcOmwTKTc+2J5/NvU8wuy2fZjb7tWkmZKZxGELEje0nSLGFZm3iY+JWwK8YF+8sFERkGzIp8xEJr05kfCoz3E7PGE8ODE3Ptiefzb1P6ybPPnrvgaaOgvxMaPkQkges4H5Yp+08dd8ThHigH8vvLBREZBsyKfMRCa9OZHwqKUdgrVQckBRNz7Ynn829T6nv7HAFPaC+NIJjKfzTrTF52q2LL6b32S5WhL9Tn4GF7ywURGQbMinzEQmvTmR8Ki+nNZAcTx5ETc+2J5/NvU/OgiioHez9peYLunBaJS6Psffihgl2mtkHrOB+WKftPLz9Xyvy+2xa8xEJr05kfCr1vofQevc2tvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln5Ojh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2a0O4nWbZf6xYRUGhK9R58AOHcwwbGG4cvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHxE/4L/XDFvVpljzfsSBgtK4dTgHxwpzDefSuzBIKJD/AWCwd+65pML9X4crs+u5RewPNu32f/eEH8Gye4uYSMMRP+C/1wxb1aZY837EgYLTi+f54onteMZ1RYJjKrk4DwFgsHfuuaTC/V+HK7PruUXsDzbt9n/3hjj5EvJGDtdjET/gv9cMW9cpH5iHlem+Ex+wdG5+EvQ7AWCwd+65pMMBYLB37rmkwv1fhyuz67lF7A827fZ/94UQS1znI6MEqxE/4L/XDFvUIQRve/l1xDpEs3zX6/3IewFgsHfuuaTDAWCwd+65pML9X4crs+u5RewPNu32f/eGSSTIPlo0BkcRP+C/1wxb19URHQ+CkkDeRLN81+v9yHsBYLB37rmkwwFgsHfuuaTC/V+HK7PruUXsDzbt9n/3ha9sdJ8uLcFvET/gv9cMW9eOf7NZ9XQcckSzfNfr/ch7AWCwd+65pMMBYLB37rmkwv1fhyuz67lF7A827fZ/94Q9PL93HTWcmxE/4L/XDFvU2/fCtF9uEsZEs3zX6/3IewFgsHfuuaTDAWCwd+65pML9X4crs+u5RewPNu32f/eGbnes1mhZCncRP+C/1wxb1I0wk6TzGyL6RLN81+v9yHsBYLB37rmkwwFgsHfuuaTC/V+HK7PruUXsDzbt9n/3hX1odLVQAaK3ET/gv9cMW9YHXNoC/y8T6kSzfNfr/ch7AWCwd+65pMMBYLB37rmkwv1fhyuz67lF7A827fZ/94bFOR50Pd5NuxE/4L/XDFvV7qRXaI3enaJEs3zX6/3IewFgsHfuuaTDAWCwd+65pML9X4crs+u5RewPNu32f/eH3cT5Js0hnO8RP+C/1wxb1g596DlEbrNyRLN81+v9yHsBYLB37rmkwwFgsHfuuaTC/V+HK7PruUXsDzbt9n/3hbrQQ/nIRgtmXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZuyzl1puP5iDS/77koXJE7DN/jys/Hw1bJUzaieDhIg70ruTV91SZC4fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwuJKt7Kze/qfEg2GBGWdp6+ba4tYSGGu76g6WVlzc1l0pOTpOcBgaCoXHACojHgtWWxd7lNh/wwskDvGcVrJOJStW35N7S1tYN/XtlbBqfF9Pa2rh3gftwJY7VhrBYSvvzCIhsEgqDmKCXoCC1carmHs2AZsGdBy2wIMEmt5aG1PaxE9Q/Bl6fmP01rOY33+FoHX+qSeHt1XhQNnUhVa1lyg23vvwlFuhjoiiFVKiU9Uci8Z18ljzDoWw1kNChOLkjNKX6SOrau3rkWJgDew8VRaNIHC+mXi0OcFmUMNY9FzR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/X0mFXQGDwUBfxxgLW/DpkietI52dApanS0ZwazF+DSia1Dv3sAhvWmfnNRqgv4UiYRGFaybmRCQWc02j3u+2kOy44C5ZqFQCn5vz96kpWbDV8teH5GenKkEwb9B+/EJmjd0l7AcHpei++Ryg5I4/jZ1hd+V95nkAjqK/Yt6Um0La+WDqSMtRrpHCFgEF9jCJqOfUlpK0V+TlFZ1EWDqf8qn4zMQnkt1w8G5+oIPR9Y6qh1DAeJ70oBYNAncoGkg5+gA4ucyggfGnkhHOWLnddxX2xf0wa4olMzMTd2VbLANuF9Szb8bc805EtuKTzyxrCgt/GByzsK27wNWQR10PsMa7TfXeyjfwFg0CdygaSDn6ADi5zKCB8VSq4rEuTQlDAgLGi5HPbDIIvT+UNORMQoUXR6IDn/3ME2DcsMtfZlAWDQJ3KBpIOSxWonF3FK3DgddvbdX6MFbUXfYiX6zhRSORD7oAyhb755eJe5a/PXlM7FV/qoydkji9MrIcEZz51sEfC9MLmJ9bMpVXuOVT9YggAh2zYxKrOm4GNjZXJt3t81s5c/A11ipQ3jNDYXS8IKQH9xapKWakY/FF8AzWjNqyLGdo9RMoaELzFZeL6+QHV5xeL4xid7wn7sPvalYHHO1gemEq84IIvT+UNORMQYjDI2ctzIMI9onXBLEFsaUzMxN3ZVssA6Sgfx+TritiyBxu2/J+f+cc7WB6YSrzgCLmfIM/UTQBwoQZER5Qwea9CKQlY8TsI6Sgfx+TrituFUC5JyaHrvYqUN4zQ2F0udGlESu52O3o3MCALtK1/SLa+WDqSMtRq4TtEeILw6IqAzJs48yu0oxF5kW0MLn8lvxmfrBcKifjFYMcF+g/n5ipIACXOdjMm+3Rbbl6sYhAP21ycyP1EuORv5ew43Ht8RWyuwsUBZimEQAGals47Xmm20Jd5iXPesPWg6FSenyHeAIBdpfm+x/0ImPkJmWxowO89C+dp7iiCL0/lDTkTEQW6A1k/HcyPwi5b+modnlFMzMTd2VbLAK+TC2YUt5Paf1EW+8GYT06+HjxaB4B74AavDmDTROJGnJ6defzt03bvxG2g30EbbrD1oOhUnp8jm1YOQrl+E35wJ6kWNLc6Zl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZ5apJj9XwnyHT/O9OWBsaTWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMf7+dMeNuIteYnYRsMRz88KMnWfB579/6hYWAR161KjWdq6q+4iv7MalCoso7qGU4npv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWslaj5EDasCQBAV4uNyXBLaZDRDzKAm9d6zb0fxB8WhpiNEGZBBfPwZag18ZZFxsrfR56zibsJhlIvB2RBqE8Qg1dMh+6V41y3L2cA5cyiIMRHrJCQh8RyxWQ6arWa36ObYNTLRsAZTMhHLZ/lRM5hy7twcZyZxxott1OLXHeZwhiQ0Q8ygJvXemEf31XJNKne7TEbKty64h5s/P9zr8kn/aI9EAkCE4YeDCuNVCU7v0plzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZqryyz8VRV9SntLtFbFkjeK6WAhyHFIYu6/pegXl4NTmt6c9O0Bg63VroVbCVTu1DuSc+YnhH5GrR5oedj4PxwxnaoYn9Prc44ZjySmeLaPso3LeLlI0CMc+nLvhQObsjEYNTLRsAZTMilqmFVgZ1MPgPMMr/DPhRjAiwqbPT0HabMbIGcVH8k+TwYhfNYoFKi54MtvmMjULJCgdn9g6LifnVehHdXBAilfSu3iiju78GfAPOJZ5hkzG5gDe2xT3KzxNhphVs3/+yy/tlkJ/4rdmtuOIO51aZSlzUDFSbt8xjFosTdcpOMYxdrpjE2Io/UlBMp6HzCvmPsyqTD1boE/PfHK+wOUrreuBq8mjOt6AfMQT5ndyMiZ8dAsIJP9jW21JPESDv+/joy+8DjTEMyXGFwS03LFbZVq5C6U9EzXBYczSDxcOSOcrlg5fuBTrJo/0+nXrAtOe5D3jQjDnd4drhS4wj3wUsyvUMjnFDV4bTLpxbeKVdsmMBYLB37rmkwsQWmmlNblQ0P8yuqWk0co7y3ZrTToWSuTq5gFT31k3f93+VHVCc6R5mP5+TWtcwA27o9+AJt1b6Me39OvN8adcEHU2Tg6xBR6IohVSolPVFv50LWAgtlncBYLB37rmkwLW7uXzcC4bSkObYUAN2L7+EkpZ1EwtkIwFgsHfuuaTAcp4hvhbTsNnpz07QGDrdWpYCHIcUhi7qE8DVtppaTqHpz07QGDrdWb5lhdorn5WioNfGWRcbK33mh52Pg/HDGOJOPlfG5GDnAWCwd+65pMK0yD9MfwDAwl+VJtD/uv6C5Fr70UfGNISkJuMch/Os1uWDl+4FOsmiu/nS427wr6TWkPv8rdyGLqDXxlkXGyt+tMg/TH8AwMFVbcOIpGTPCIZVR/UTDmca3oHF4XEg2aYM+aEC2mLhmax7M6tZYeK72iuplgCAem8bc2MNXcGDL+IjdDJ9q+xjo4p51YmELEvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4Ull/LbH3nTy7MVmbSj0GZC4yqVudif6FWNVUbSJHrvBkmZ62k567U5f4b6u16m0yivXfiE+y4Y2r75Xq7KYVha4EjQb36tDvIlKFRFC1v8AMq5V9IKK+ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwuaYURLz4KbxwaSGHgNq4+ZAYIUgJKG/kbXGD6Zcp3m+RYDBFYuiF25bBbIUsar2X3l0deS1AQ1vEPbf7OI4stfbVSTH+X6hdKjh/7YApD9EgaSGHgNq4+ZnFb4VQbvyQ85CR3b7eb+cjCgwNA5DqFbjkGwgGfgT6lW9EiFfraz+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/SOUqXqc4IdsI6Op4SZut/nDzHsULEgQUFnNNo97vtp0uXiEffkxxqc/Jhw+MxWm4J4GU2KWCH2o7IgfUbYao66E0Ypsh6pbTKbtlqu6/gxhqfiesrmPWgl9BK0MsVDTVY1tXzOO1m7yvSCqDbzX+imbVrC4uDyJdep2m4JtoMoFA6vM2qPhqo180ffYo0kLjpYJZFHLSAli++Ryg5I4/jZ1hd+V95nkAjqK/Yt6Um0Z6aZwCSgsMYAQGjP89uJ4qvvciyv21W/mlYqV8JzNNR9giTzGNcK/gCGN6OvDnnfNrBKvbSWGzhGICsHLYYKtCqfjMxCeS3XDwbn6gg9H1ig0p2IaUHthcEfppvqcUz6AavDmDTROJGRubCehLyprSIpo+L/IexPrD1oOhUnp8hO7JRb/x7EOB8gtxiLTTHihgLnWkmJHXswICxouRz2wyCL0/lDTkTEO95IiZfXcDTT00i80nQXynFfbF/TBriiUzMxN3ZVssA24X1LNvxtz2SaY5iGH7r96QoGFUtdHnsdg1suZ9E6/wQE9l397Yn0DGu0313so38BYNAncoGkg5+gA4ucyggfXauXY8QQtzuSpqqKyDHMiKw9aDoVJ6fITuyUW/8exDiUyMpMFu/g+62LiTlmATyVMCAsaLkc9sMCLmfIM/UTQN8X6P4n8etka9CKQlY8TsIdg1suZ9E6/xVpVWDUN/+ETWxcDlor/l/BH6ab6nFM+q0edPGUxp3RqXINbESJTwlr0IpCVjxOwjpKB/H5OuK2NevrI21fTEz33vQVFlWnA3HO1gemEq84Ai5nyDP1E0C7mVmb2+QTluxjbVPe5ExNR2fVmEyqvVMgQLozWXkxVYGpLjXPf4P7Jeg+iExCMrkBq8OYNNE4kfwAdSaytepXH+VbvZ6pwOLR8jzVqDLOsXd/2KjKK2P69EB+b8grdruPaJ1wSxBbGs3NonL3dWzRKzXangPC1SJ4Z3eJFmVzXABAaM/z24nip85YDV7dex122ArGOOFvlQCGN6OvDnnfs6bgY2Nlcm3jYgY1I8DT8RVKrisS5NCUIGR/z632+sOlaqHQ6HYhZcmgRuZRQteWSiUiWog51c+ir2iOWZq+oJTOxVf6qMnZI4vTKyHBGc8+7fMKTrRNy1RWHJYQ/HeHd3/YqMorY/r5wehdIVIWOdbs/HwDp21crD1oOhUnp8jqbdmcoQYqPHPT6yNUvnsS4cMmgMS30D0fhcE4/+Cy3xLSFqhwq4BYTWxcDlor/l/BH6ab6nFM+q0edPGUxp3RqXINbESJTwlr0IpCVjxOwh2DWy5n0Tr/JWXjilvtWs7ipWeARDPSg6w9aDoVJ6fIkITnt0Z9dgLuDmirbUrVEhmIIIY4VdbrKt4Go7aas57WCqpp3lPw4r7dFtuXqxiEA/bXJzI/US7NhRrnTWoSgjyePkcjaHGB95KyKQDKl8tBboDWT8dzI0vLh2Lc3/FcppBg9+C3bxmqYD48tup0ytsDxyFjlO3cbSOCRWy11TQwO89C+dp7iiCL0/lDTkTEQW6A1k/HcyPXMbERwRon/MqbhWe0xtycAWDQJ3KBpIOcaiSB0pwUUyk//siOUjO5BAT2Xf3tifQ0YRGHlQeoH9WZoiiFN4qHQvjg2uKGm2zEMQgDNZms3Esm0JuZyGZSuuAHo1W8+UzqKt7dnBC6F85oHJfG1wo/K+TC2YUt5Pblsy++P37SHhVKrisS5NCUlM7FV/qoydmdE8lMvwJei2GiJIyLcU1+GyKKohN7Lcmvh48WgeAe+K0edPGUxp3RQZZGIhv0paHhwyaAxLfQPRSI6dQzrfsnEtJV8xwgsafhVAuScmh676w9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9FIjp1DOt+ycS0lXzHCCxpyJfiSqxiIXClM7FV/qoydmdE8lMvwJei7K6SAnMyYhqGFh4qNY7G7LT3UDwJBQZLAFg0CdygaSDnGokgdKcFFMdUnqwH69GR/PMtpsJZZrZrD1oOhUnp8h3gCAXaX5vsU9CnTVxY3vYIEC6M1l5MVUJ/HLEdzJ3hFMzMTd2VbLAK+TC2YUt5Pblsy++P37SHpnKcu8csCg/l7+OBOTMkQDNzaJy93Vs0Ven4UCILaaxHEcuJ+RvSwZFXGCifSifHEH10ILIM6PIGdUDaVDVGwTNTYZ8Q0socsIKQH9xapKWFIjp1DOt+yf+NMNrKex7vqODkWV7yhQilM7FV/qoydmdE8lMvwJei2GiJIyLcU1+aRW8cUxbqZU8Hfe4JT2CyZ0aURK7nY7epa/XkEGd4zccRy4n5G9LBoVVIPUUpxe0QfXQgsgzo8h50l/dgwUZBaODkWV7yhQilM7FV/qoydmdE8lMvwJei2GiJIyLcU1+4volq89Lfg2ym6TZ+4ZAL5TOxVf6qMnZI4vTKyHBGc8+7fMKTrRNy4J4fh36Dqz5QW6A1k/HcyPgTQAzGYCWz6w9aDoVJ6fId4AgF2l+b7FB9dCCyDOjyBHydQWgvelWMDvPQvnae4ogi9P5Q05ExEFugNZPx3MjOMHm+Q/+lsQwO89C+dp7igIexiXVXUV3EYGX9ylO4vlzY7WXoU7poGl/6bTjG8aSy/BJV9UtiIlbiYvUXNVjIpjNh4k5frRn1pEqQaFUe7oTyE4qkW6lWALBBjqHp9FK37cEVTJFRrSXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZt7lATO+fQUOyppQx01QgISJHggw+4pkqacnMu1L3SPEcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMk632GcagQytLnGvdljclOM6YTgOfBUyOhYWAR161KjZGADmCe/f7qlyJNSZWXY3L8QxfT+nk+N+b98+AaJaEDsG+QROCz5daOvroGNV3EmLT92eHYDCAlV5gHmKglRiBHQFnXjVGU4QAwcbwuXIsVZDpqtZrfo5tVW3DiKRkzwpliwFfSIl24R56zibsJhlIvB2RBqE8Qg+Vg2hDaiCKEbSOCRWy11TT2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTK3GgGumDdGP4SnxwPWBAJRdqhif0+tzjhHQFnXjVGU4SP1nBXwtP/N9qoHINnqNTQT1zWClEYtH4XLjiOTjsUytxoBrpg3Rj+yBqh5q+dahPaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMiJKspioodXhC+7dytmw+MV6c9O0Bg63VvOoYXf/L/aGXrdFSL68VgKnxG91hzMy4BvKpHIq8yAtpDm2FADdi+/hJKWdRMLZCMxsgZxUfyT5/E8WhcUBwubPPc5FBPOFcDk7mXP2p+dQ2ly6kYt+fJcveMOq1FeqVCP+77VB6HAZqTjwpWEMjv+g3Xa+6Y1DLQx9b3187N4RiWkCncOsPpTqKt7dnBC6Fw4lUt82goFOCcC/n8eXylhQD+a6MozVNGKc2i17wFLGBQUIeiP3IUDy4xKybdWbuACGN6OvDnnfYQQyiPLcTq58Scc1MPgfLZ8LkAubFoOawc7mYHRUR/f/CS3b9hr3I3hnd4kWZXNcAEBoz/PbieLhJKWdRMLZCEdAWdeNUZThADBxvC5cixUyNZtCbjGDoOsbBD4wDKXul+VJtD/uv6D+BYdEK+bzau7wl8QgYkVBQ6h98TuQu7V2qGJ/T63OOIMqS9j75lvBvoiGCRllu1RfgIcbEXWDEwQE9l397Yn0dq4mbHiBsNPrGwQ+MAyl7p8A84lnmGTMUQrZoM67hh2hH9pdAbvHUYKl9kZn9cgq99O/uKD1+pPND+QIaA2PQuuwrupyCFw2VzX04Xm89MpnppnAJKCwxgBAaM/z24niZGM9GzItU8NQD+a6MozVNL+1RAE+KJ5AqDXxlkXGyt+Pr2OBgqTqrld04W4wpo7k41O10RHHrr4Ya77f8vmAHeVg2hDaiCKEbSOCRWy11TQOUBICzFgQs3D3jZufTTGBMX0H0h1bK6ixHXReuN0pRFrWcRWBW8yoGFh4qNY7G7KaqJlJU1jdFS9nAOXMoiDE7Gfhw9lEZps2/ULkhwzXXoMqS9j75lvBcfToHZ5ByWcbfKdF9AnQ9p6iewCr2TfgmDbtbWCZRTKeonsAq9k34BUjqW31aQvzAxd5EwU8gX43LeLlI0CMc7o4TWGOq7a9qTZrPm9xGrOmxVNjopp9O6QG3kyTzDHT7vCXxCBiRUGq5oo6fqyaTAbrbHum4RqjVltyyQ2nJWAG1QDha/JMrUTe3KALTTmkirY9i21GUrClwAFiUQDmWiNDOWu8768V6gIFcFwuc36UyMpMFu/g+7TDWUEwuxNqodr0DK09K6ajsR/sBu021v6WIeNiQwBXzGuevNq2BAXf2ZfMmM0i36g18ZZFxsrfW5N2xteMiCTzldeans8+9l0S4wCHAjZhS1ZyzjNn3f2yDerzxkO6HR+pBQUd/IzhvoiGCRllu1SRftjjGWJHTS9udGlOlsAWlMzU7+QOu6CYmnGBzqxo2PL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln51cN3vRz6AXc1/85T6zUoShyXZQCIC2lpeb30mmomtpWc7jyWcOB6eb5i1OBd28aLUx1zwuoSsvJWPiNykRv14/ERKfyzaAKjbSOCRWy11TSscQE1hVaQ5/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxFUdp7p+cxlhSDh+JhZXj1cDyONhn10fiBLZc8CuCzO5wIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk94PmUCcez/2pxyd1LUdyLqklytWvAIW0IV/WU3qpuprBnFhjmmDxEr16dydkrPz1J3TUNlbZRD05CRqz7/gFKofUxVuCXS5Y9ScgHHXxjCJcoyu2wqIzs8RO5zafLLM3OYiqiWWtCZqtLBP58cOLnqd01DZW2UQ9DWkPv8rdyGLgGwFmQkytbgP1ziX8hdVw72Rzp/Eas+gdRYolDpH0bMD9bKlyQKyzfcGK6j7eV1Y4SSlnUTC2QiOTUFvulzbqYVGs94KMgGA4IEfocwT8sQvB2RBqE8Qg2FmjN23bm9wM1ILnQKCFfPmjKghd4lsW/gVzuJ+JsGkkD0Wvzzv53fkSCKtN6j5A/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8WlsSdjcKS3WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFlwEuO0+fAPHVDArIheVHLMLvZRSMZAkI2M/aU86MHqGMCFBs8ZB431pR9tmklx5bklnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTtPvTnl6ngWRfXDXEmsM9p/7nrjc+L9nP5oyoIXeJbFv4tRTJystVaMV3ivEv28U/Kj8tYIakxcxkV2RKeFDdtwfJ0qe1LpvI7H8KodNn21ZXmAeYqCVGIEdAWdeNUZThEfJ1BaC96VY1pD7/K3chi4BsBZkJMrW4D9c4l/IXVcO9kc6fxGrPoHUWKJQ6R9GzA/WypckCss33Biuo+3ldWOEkpZ1EwtkIjk1Bb7pc26lbk3bG14yIJHaoYn9Prc44vasFSgZCszC+cTnAo1owFGIKO/++klhwI1hFnYyfkJuowXOiQutLjzwwKx7gMCRC8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3Z/sInISWfk6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZamIuBW1zP7rS3p9431jslPTwar5gmcNMyj/OhZsCUtTNkV4iC7KdQDokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyESQOHfndbqhFUkw1ce6uQrBv4MqHVoNrJn9IO0/LopHzXL5Vsde/WzN8hwkaeXL9FU47DHWzeOzX88nixuUVIMk0flCMwg9o1dZ0prWwPdAl930UV3KhrmOfTLT3e9rBuWDl+4FOsmgDF3kTBTyBfgDkdK0NSoTvaDfN8yuJlY1RCWbeSOoaDeYkZzDDBaT79xikmyUKNrN/JBuYrBkiCao7hFXG+33obglCZfq9SqPKP86FmwJS1CkJuMch/Os1uWDl+4FOsmgDF3kTBTyBfgDkdK0NSoTvclW0zyz2/6v5LCgko+ER+khCbSbv2lPoY8tpHhCv+qGD7vKcI0rwkkD1RzJpDVvTtwa1lNNbSWZ2z+DYnDwqv4VGs94KMgGA7JlZuF+2zJROBgFo/zb+LiTxBGH9G9dZYWaM3bdub3AzUgudAoIV8+aMqCF3iWxb+oXdtYS0+fNV3jME9gKlQv+o6hWtmGM88v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTI9fIwYzQA4GlUgbrlPdH1t6kUq5gdfPbfUkE1t9T2KFuZ7wIVBB7TQA/bTlnLsNLZVE0IIzKXDI50s9YPmpnx8TSiwNEsSraj2GXuFFM61Sfk1AxrsWtWL5i1OBd28aLBMpRwFTt0j35LCgko+ER+gZlVMVVrrg481p4INTjNmb5LCgko+ER+tzo4+scB9LDQLw4iiueoOLy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR5mLge1gkCQqTydBziNYSbHpCgYVS10ee2gLnMoJSJnyWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJO0+9OeXqeBZB0GFY/oiK32ev3zcrwmkyPmjKghd4lsW/i1FMnKy1Vo4qGBiJ64m5/kPLlf4iuLNC2qYd2EgdKtDQUFJSyD4MVNhDOo5YPnV+Q8uV/iK4s0+VvqxG/F6K7hJKWdRMLZCMmgRuZRQteWSiUiWog51c8+PtLIAl07z2z8/3OvySf9oj0QCQIThh6B5vN6lMor7E04m/g0IngK3EiHSgIWVHN6c9O0Bg63VsSoai2FG662f45+DaOSPME0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm3EqGothRuutroPTioawmgi7TEbKty64h5s/P9zr8kn/aI9EAkCE4YeDCuNVCU7v0p8QyaTIpyFl7Y+n/vZaFAMuF0OMqX8TPvw+S3CeEs1VhE7nNp8sszc5iKqJZa0JmpiEw467AmM5sCLu3VTXAHWlpwAZIX2MBvYrqEx1I9NHIHm83qUyivsqKh5ysNCgDIVfhK1yE4xIBhYeKjWOxuyr2asQ/20rIuB5vN6lMor7AXkQQfNmGUxTVCXl9Ty83gj9ZwV8LT/zZDRDzKAm9d6d3/YqMorY/p+ihK4TVTFLmvsck9eipaU/g4C+R1K/bAYa77f8vmAHWETpzZc2/VMlvAmEYi0AhJr7HJPXoqWlLIGqHmr51qEkNEPMoCb13rxhA+nGH43aPTltnpmaj9/2i2F4MnGf/TLk+ksSBii9Bhrvt/y+YAdYROnNlzb9UzNfgAg5nDYHLtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXemFmjN23bm9wH6kFBR38jOG+iIYJGWW7VJF+2OMZYkdNXJPh18Qv+KcdBhWP6Iit9k+MCODvKVABOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHIyPUSiaQE5cPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxaaAnmoOVRXNmOR+P2/mhrYaELzFZeL6+p1sLjqTcO+Hy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTfTltnpmaj9/TVgcjkU7TuOFf1lN6qbqawZxYY5pg8RKumXPLHuMZeGhJ+dygceIfudtI/0UeRgdZFdkSnhQ3bdyErauFowuZqEn53KBx4h+xi1yExziaZRxCvea/bRFrO7wl8QgYkVB4volq89Lfg2NEGZBBfPwZag18ZZFxsrfzyX9SCyjrO8HbaHAM0lMvbtwcZyZxxott1OLXHeZwhgETOWt0KBunJJ3ezUKUQNvkSNzLiUetE2nxG91hzMy4HxDJpMinIWXke8MtH7iTbdxCvea/bRFrO7wl8QgYkVB4volq89Lfg1yutCtFkLjQ4gNIy7Xb5Q6UQDEX4lGWKx5DyozQXIMkyKGMZn2AOVqwNs7b3N6hD1xCvea/bRFrAo87QNhWHJ8EtIWqHCrgFiweSSCHUioFe2E3UGVHGNFGQbDERUKy5OoNfGWRcbK360yD9MfwDAwgz5oQLaYuGZrHszq1lh4rvaK6mWAIB6bVHw0ii+xUBwjT55PbmP2kjApRw+CA5eU8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3Z/sInISWfk6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZC3JEVpdpEDWm6OM5Gqn9Oo3ZwrW6BeD7OiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHI+b+PLlOZfNCDhR+puYCQteh7vTtA6Y2z8UnERL5ba7BqwbAwT32MxIoYxmfYA5Wq5QVYa+L9ezmRXZEp4UN231+hui0kVCNTi+iWrz0t+DZacAGSF9jAb2K6hMdSPTRwDiKW+ZEt1kCKGMZn2AOVqhPA1baaWk6h6c9O0Bg63VvOoYXf/L/aGXrdFSL68VgKnxG91hzMy4BvKpHIq8yAtpDm2FADdi+/hJKWdRMLZCI5NQW+6XNupJWXjilvtWs6hzzqlDrOrdC8HZEGoTxCDYWaM3bdub3AzUgudAoIV8+aMqCF3iWxb+BXO4n4mwaRYJlCGHNnosHAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsRyqznXagQA7cZZlMIOCnGIEihjGZ9gDlauNqxFSsuIt8rFGy3LU4fU3knY7kq9NuU/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx2Z1bAdeAjrKzZztQUvJ6wSZeaT/v8OS1YPDP1zxxfaincOAviM+2k9pLGDwrS7nlLaph3YSB0q0NBQUlLIPgxU2EM6jlg+dXwU4LgVK4+eeYUieJ1YegZdiuoTHUj00ciBz6eEcfK1ntaoYmNQeFPJXZg+ub6CpKQIaAy+tSTHE37Nk97b+6rmi6syZn5bD0l7deJwMlll+w9zAOf0R2zW4JQmX6vUqjhcv+0GNHQXIRO5zafLLM3OYiqiWWtCZqWUMS3Xqf10nKe9kjgiYRyySiXbk/kybd4volq89Lfg1MxA/8zyFC6YgNIy7Xb5Q6BFZjGzSvNg8H/Q3upe2BSyFQJqvh/liWLKvGxPV49nyIDSMu12+UOlEAxF+JRlisrTIP0x/AMDCbsKX8kabh1EzM6jWgHkBN8bcL1ESPzRi1uowg/jsLf3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcrpLydPnYbARTJ27vkeodiCBbbrUwso3fO6Te8WiyaHt6TR8HxZd624AKu3MThjjHJdlAIgLaWlkpDoL8UxvpMFs5QQx/G22WdTn5rN1vM85f4b6u16m04z+t1b5RIxZ4volq89Lfg3f29nOlhZNXYeoT8PZKa0w4volq89Lfg3JuHQ5widhwKxxATWFVpDn8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/G8tG2IGc9HiduyBK2DNHi0o23G+a5Thj477yCI4vDW4TokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRy5bTMREeIT6tJSpCCsaiAttqyNWqIi+hIJn9IO0/LopH66fLkuqiwqx8gtxiLTTHi3X5AT3IlYHEvFfG+fBhu2ssCk5CiXq3flyJNSZWXY3JGW8JzBFqqo41VxarjbYSyG3ynRfQJ0PZGb+OFFfiq+UBXi43JcEtpkNEPMoCb13oXAkyU+CdDppaC+Ni5NNHrdqhif0+tzjhmPJKZ4to+yjXr6yNtX0xMsHkkgh1IqBUlX26L3zEegzDCDFQmIOwZgGwFmQkytbgP1ziX8hdVw2QajirGavIYk8rBnyA2a2e6lpghXwiSzSkJuMch/Os1uWDl+4FOsmgDF3kTBTyBfl2gcFRnB/6dOMHm+Q/+lsSQ0Q8ygJvXehcCTJT4J0OmloL42Lk00etTHXPC6hKy8u9w00TM/K+UQvZOoeWO9V84web5D/6WxJacAGSF9jAb2K6hMdSPTRyB5vN6lMor7IjdCeCdiASumW6iHpTL3E8S0haocKuAWNWxV+32rY/VMX0H0h1bK6ixHXReuN0pRHd/2KjKK2P6wJJ2T/4TITntMRsq3LriHmz8/3OvySf9oj0QCQIThh4ASlQboJTlvmsezOrWWHiuajkcM0HTJMWiAiNHs4agN4V/WU3qpuprPRmDzGC0KjcXljJHaYnZh+jinnViYQsS8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCThSWX8tsfedPQBwpcmO8cUjl/hvq7XqbTz8Fb58oTtIrz2CFO7lpF2Wpu4hMG3CBrDXz/9QgbnfGugCtMuwzpQuZsPEA18kKxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Lw77OF9d4rOWvl9lNkq+IdrX6T0NpFxbWIc83RD0iU+Wvu4K8NlLooedDa8/RTQEBD69i27DxUHP/OYV0R4td6r36mE7lWClZdLuAG7fM0+3YEi4cAnb8S2bZXUjuWQOB4nYUgR8WpyA2FIgFREv8mr9O/e/erGsxSpHyxByx2B3e6iU6porcCj/vntd/amgABWM1emdk/d+81HlYleWfDocQ5WeS5NolAMq5V9IKK+rTc1BAUKC0PB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwty09P8htiA7a5WfCD8gy7r/pfcYVzcVjdk+/6CBSpoQ+9c4Zcw0m9czc2icvd1bNFLnqqfezW6ZZj0EJIIrJfLWBa/jGXMVR2l9JlDWvKVW+0bWTRss2SZ8HpQPe4SZ6bVjLqE7cxd49WDia41ibSM95KyKQDKl8tP32Qsz4x1ZmgxwPOa+bCZB6Ptd4HKe/xZoW/GvRb063sDzbt9n/3h93E+SbNIZzvSmqpTekqemjzhw+lgK6yXq+9yLK/bVb+e2eZLAFbFqEoGFXBlwsrjIDFLgXm8zaD7LP50KARLqiJz+49qRNFLrBxXQD2wvp5qRj8UXwDNaDgUxDvycU09BQuox4V67UBgPHSgvyImSmYCYVHcspp5wgpAf3FqkpabnAjLtURujfruUpkIJ2nllM7FV/qoydnBYUSx7a+c9sOnquJ1ZT5uMCAsaLkc9sMgi9P5Q05ExBLjxe+5KG4PcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/ZxbbU475oEKsPWg6FSenyE7slFv/HsQ4sfEoSEIM7uVeCQMHKUbNsNWZoiiFN4qHJQa2D2k/1ZDsY21T3uRMTZ+gA4ucyggf6lF4+lqJXDXBH6ab6nFM+q0edPGUxp3R6mdaDeTjPdNr0IpCVjxOwh2DWy5n0Tr/vRzFD1Ih1OisPWg6FSenyOpt2ZyhBio8nhp7AmtQlzrhwyaAxLfQPfj10qKusZM2eD0NOhcCV6ysPWg6FSenyOpt2ZyhBio8nhp7AmtQlzrhwyaAxLfQPSMMtLkbT32yfU1KG6V7Qq+sPWg6FSenyE7slFv/HsQ49kvbPLXWbC4qNxnjpd0MJDblq/hFE00omq4fKoPDMpRipQ3jNDYXS8IKQH9xapKWNuWr+EUTTSitCR/EK7KJ649onXBLEFsaUzMxN3ZVssA6Sgfx+TritgkiA0/iQMxTQhQaHWyXaE8BYNAncoGkg5LFaicXcUrcB6Ptd4HKe/wBP4Lg3ltyKuxjbVPe5ExNR2fVmEyqvVNFJZ6awgyw4EJB9PRMhOAPJeg+iExCMrmtHnTxlMad0WLNwFR20fl0ecZlzKNOXCo44KuW0tEdOm1F32Il+s4UESvn13ENqYDZdQdps8ZOyV4JAwcpRs2w1ZmiKIU3iodcBos8KZc6npU41/mYNZV8Np+ipJFgnO/C4OEyxUpTD+6iqgo/5TZNkbTZVWMn+txeCQMHKUbNsK8voH2jFdga+tyNk1P3TpukEwb9B+/EJl1YPKtcadHcCOX/tInXF1yROT71LE3gVQ18//UIG53xVbuKc9hHMQ6DZXXQAJLjiZt7Ud//wYYUbKHtxvXCpUAyxlfjqWOYzHzPFxTTWvuHZoOlDecgR6lOE8JKU7U8Ub/obgUrlrTAqkrfw71m0nJSRfq5O9pVHIJD8b73HO3EABiC3K9WHgQstsoQI1b/gubwU95hCTRJahhRZ4mHLfRQkVlLBF4H3hUtj/11qRVCtdZWz+hxs5o84cPpYCusl/Sy1YfM731qPfBeph9ewq0UEbVAuFkhHR2JoZE+6jouM+vr6PmT0MtDFvvpzeGkidWyKIbzMhJMUDR02VSSRBFq1Vsuhf2FdnedrM99k2UjbSKRD8qYg0/JHIMj965yulAPHiuHcPVLbbrrD+edxmRI1FeNwup/L8mgRuZRQteWrUkC7LYDZCNrH94qFsHdXN3VRd+PH7esZaXTxQ9QP0DkD0+5bMUZQSFAIJxhUD0L0KrIXGAtUK8Ya77f8vmAHcBYLB37rmkwT1nZXCU9vI2t/w2Aduk1E/kdYNCAtGp4AoHnaArgPt2z3MzWXtoojfSa5NP8WNXHexWzaab6KFAlGKNpa5yfwrfg+OFxvZPNn+YP4grcZBUlRxl7I63ZM53neQLiJuaPCOX/tInXF1x2IdBu8jtk4m+oxl8eQnuHnRFUoESi2wWU4FAd/tEDBQ1s8E7IYjG8E2Sd+2yQl1Y98F6mH17CrRQRtUC4WSEdHYmhkT7qOi4z6+vo+ZPQy0MW++nN4aSJ1bIohvMyEkxQNHTZVJJEEWrVWy6F/YV2d52sz32TZSP+n7KbXocN2rPYUPcrbRXbNuF9Szb8bc8t766baaDir9OGRz9CsCdVOkoH8fk64ra5aAljcDtU4tOKCkPqOrXqP/kD8Cxw7TdhfQeIFI3IYsI8R9UxTLrFcnLT90gppaod0XQ+KJVFODXR6dfO/9nfL51DMPqp5JUc7imwkX4OMaFcM9Yb44b2am7iEwbcIGsNfP/1CBud8a6AK0y7DOlC5mw8QDXyQrEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvDvs4X13is5a+X2U2Sr4h2tfpPQ2kXFtYhzzdEPSJT5a+7grw2Uuih50Nrz9FNAQEPr2LbsPFQc/85hXRHi13qvfqYTuVYKVl0u4Abt8zT7TWUWgnEYxS+6nDhe/thj1I8C5TsJcQtQXjtNlWkSC6Bh/phnzpTMTm6ky4dQaoOMjdmREWZQvqhtlxqQ+SrVvS5SjiodT2RZyba61mL7BzZH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LsMN/64x7yBQ3jzhesRtAYfKcEnzPHlzUPUV6or0AJU/mm0Q/uaedKEGFwdQab4wcGpNPJuPUpAd0tGcGsxfg0gGLdQeyYI73q47DanIsQyOuesPL3HrjaDjh33ZdFaPS7c0pt2RaKmEfKVl0mUo9TqPrf0CC1QVulmAsj5iny4uRIlIUxFkHzwz25Ac0HZhe49Rdw4YY69Xl/UKtaZ+/7eGNeHLuMDjlCi+E+3rirrLLcisHQG/3SYtxsIVISGqHnu2hyUEUHC7WmH0QnDKBivXhbJmtmkbM5JHQyonYvUq+Uv4lGNud8uZmUd9PwTNuad+WbYZY/O1oMcDzmvmwmbl9wsIcAO/aMCAsaLkc9sMgi9P5Q05ExDveSImX13A0+XS6JX6v8WPBH6ab6nFM+gGrw5g00TiREtRfj9IyqtU6GP0YiSUflzVmJzPpVUyErUHzjuIyseY44KuW0tEdOm1F32Il+s4U3PQklR7DhT4X34H2aAQeSDGFM4H4efwuGln+GR7Afdow0mP3skyStEx7gBn3LDygw1IMUJ5zDztzXUrUBDj67SqzwpefquLirZk23b3pB/JUBKPN3GUEFtb9ASa5UQIgWFjD23zL+cj7dkx5Hwxu+8RP+C/1wxb1hKtiNdPSCQxb9sCGAnn8yTawSr20lhs4lz50dlP/19nzbK6ANvtE18pJxVMp0yJQJdYoOZj2QO+JTxE5h6Vcj9Fn77dASp6JqEH4HU5T0HhNz7Ynn829T7VsGXSfEFv3n7K5SsmIA297A827fZ/94Vs1XCX0+GQ86icSt46qnX89CZQ7e0rb6OvJRE8fGHdIFgC67QWvNpeti4k5ZgE8lZ64K/wQvn7OGJQkVdzgUcRUVhyWEPx3h0FugNZPx3MjrhTDGlPrgTRByPWgy+P8ExI6YaHlgTxe4cMmgMS30D0cEwbZv3JZJHVQ6Yf4ZdgVxoFbhV09deC/dP79Ds9NOS0t5qCf9sEuDY/8nCQapr7MwP/CWhjSPzcjzxRVwwq1a9CKQlY8TsIr5MLZhS3k9ht3+qACy3G9P6FC7vZH6a4kcHKN9FQHLBREAt+7eGmp4Z5xKSDUJdQ44KuW0tEdOm1F32Il+s4Ub7CKGgQd+InN0MLwe8EQlaw9aDoVJ6fI6m3ZnKEGKjwKDpjRFY7VKjafoqSRYJzvwuDhMsVKUw/nSv/rNmDxCQWqkBy0jfPtpEC9P6LBYefNzaJy93Vs0Ss12p4DwtUi1MRa2IZWQ1EcRy4n5G9LBoVVIPUUpxe0BDlZGqZPqnYgeQFngs3DW/3+YEl8JkNJ1ZmiKIU3ioflGPuPLedAvAE/guDeW3Iq7GNtU97kTE2caiSB0pwUU7u0Mj6D3rb9/f5gSXwmQ0mlaqHQ6HYhZedK/+s2YPEJpewtr2lM+p3VCaIxs+10Sp0aURK7nY7esOL89vNiEXEcRy4n5G9LBoVVIPUUpxe0iEseqHI5ISdcJuTcNddNsaw9aDoVJ6fI6m3ZnKEGKjx6R47YbHjUfuHDJoDEt9A9Cg082Ol+YzSUO1G6ugToppU0PppPtSj3u3BxnJnHGi10eKHQ8KaQKJ56WEcoU4o4rDu2MDjYoqW7cHGcmccaLbdTi1x3mcIY9XH1gKupzdYSTu1StmVUfb8UASwL8w4Po9+A/OqXQtxZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWXUOKP3fiCNWnW+8u4REzHIDokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyzIv2fcuq7/Oti4k5ZgE8leaMqCF3iWxbLKorACqS2fQnpv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWshlj7bUb8Sjc3LeLlI0CMcyVfbovfMR6DMMIMVCYg7BmoNfGWRcbK364UwxpT64E0NJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpO8YQPpxh+N2g2uXO9FnjWKZPKwZ8gNmtnmNjZPrsSz73Lk+ksSBii9LPE7sQG274oTOxUb1lb40aqOXx3nNrXG7oVhN3kqhCwOVF5C+BkQx2oNfGWRcbK3zBrYnbzmcILPj7SyAJdO89s/P9zr8kn/aI9EAkCE4YeMX0H0h1bK6ixHXReuN0pREJuS805Uk+H/GW1voqCm7PyHguUDB3SUH4rbsGY09o8ajkcM0HTJMWQ0Q8ygJvXekgEw7YFL9ckXP9pLHdd8nopfZuT+neUKGo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa7sJpxVtDkruKX2bk/p3lCjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+To4dhv1qMaw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9lu1ZKE7sYMbfUU7oZD+AIKl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGYuatYSygaQE2ZSodoKWcmjBYQtlT4HBvMSBx+ApnC1dtyyQa5HMXQuJrZpNlGJw2hmUqHaClnJowWELZU+Bwbz9ASUYBCeDhst3RFoJP9wkAPjnNTabYevy8aXiejlooDq2XH2Gz7ZgM3NonL3dWzRNMdf0VOLQw7ymRM2m33Fbqg18ZZFxsrfnJ8Ci5MleCAIFILAg74Zsp0aURK7nY7eiKMAKkyVMvO7RrUDdWPIZd2kt3eo925JfSv41OLfC5kBYNAncoGkg5LFaicXcUrcFQRTQg1Qz1Ar6UhuhHB4PxT+D6NplXoUS3rGKaw8lmfJTwoPGW/kqUcuyxcVE9VcpWgH+DiJO1DS5B+HQuLItdxDu4MBCLEPLrzc7vG4bof0WRP9/7dMbG8VngA/qpziqDXxlkXGyt99QFCbsEdS9Dl4MXeNpD747z1eZWxDmhEtVDuLVhKgTT1N9d+fX7PwqDXxlkXGyt+WfTcDF5dBVCrYVflocTdqwYVIDFJRxvEr6UhuhHB4P2LX+CPbZuWdj0/592s/krZZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk0MSw/dqK9HHl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZMEaEGcGD5BKOCQ/Wta/Mur5ehiWYEzfDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8SB5AWeCzcNbVd4zBPYCpUI2jFsjiZ72mKZkUi6qw8jhtrLqfBnyQDMNBQUlLIPgxU2EM6jlg+dX8wvcQ79a/M2OHAgZShzLsag18ZZFxsrf/id2tyC4EWz1MOfjYH6b/Gz8/3OvySf9oj0QCQIThh4MK41UJTu/SmXMZs/QAAtMp8RvdYczMuBRY+fnLq7F/BE7nNp8sszc5iKqJZa0JmoFqpActI3z7Qb2EX1g657YxQAK/KaoBfdg1MtGwBlMyLZZzmiwPIDzxAHZv+4XFSw1Bv7tCWpq30LoEtw8CJtagz5oQLaYuGZrHszq1lh4rvaK6mWAIB6b9QpJmxp8dELUjJvBEBrO88TPB3CPV0+Ml2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGYZm3OeEG85u77dFtuXqxiEyYm7kPd+M9zmbDxANfJCsR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC8O+zhfXeKzlr5fZTZKviHa1+k9DaRcW1iHPN0Q9IlPlr7uCvDZS6KHnQ2vP0U0BAQ+vYtuw8VBz/zmFdEeLXeq9+phO5VgpWXS7gBu3zNPtNZRaCcRjFL5JfJT2nt/OywVqdALyGP3777UE666Fn1EAyrlX0gor6tNzUEBQoLQ8H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3LT0/yG2IDtrlZ8IPyDLuv+l9xhXNxWN2T7/oIFKmhD71zhlzDSb1zNzaJy93Vs0Uueqp97NbplarmDIzkr822b6s8qwQE970EPDmeXSehv1knBXlhDPOgjbPf3JibGSxuqimyh3chzP/GXOIAnlejc9ruZiEr/f+UN5Pq3V+oLjMPfC77s2Y8XL1EvNxXLYU6yiST+YAePvGEn8zV43XMjKCtCVdVaJ2gxwPOa+bCZ6gSoT9QrPPrApQSd0YuWARMEHsSu2CAyzY7WParh91YBPPa805uvte/JgsnaaCeDaZiZzWQhDGBAG/EfEl/qkONgsncp+v/amQTBejW2v3g9huH+44zQSbMU0mk17ArP0k3ChgsRduku30nI9zYFFybEtEOUOPLYW60BkabyZH4bEUa4ykaC+7p+vTuNojysk4CHfMgf4NRuXY+sCNd1Qag18ZZFxsrfaAtLJvDXGYMini80foEJI61LINW16fzDnZWfSQjdjbUgzjCOo/3lIbpMK+U2kO0glIIVXQGQjPUE70eaomHSXPkYAay/7HEWHn4UpoGMclkOgDx0d6L/Zd+UfsZauNDD7RD8QBrTnbvKdl3cDL3nACxTmf1fyIsp/xlrAcvVbtQTxOlE8M3lre0Q/EAa0527GK7NAXON3fTey8mWeXnmTkUXNXbtqj6hXU55l9oAocRCQFYwC9LxJoO+jQodlJ7WnWagUzz8bsO/BQuff5cp0kCTBzCUs/buhnVRff8x2u60H0Zg7zKUnGBoF5rPtH7/v9281ooBjDaJE/Zb6Hbk66c2f1VVmuUSE8TpRPDN5a3/w2FLUFcK76zrTZji625759zRccICf4R81RLeuFJR5BxzT7NM0Wt6qkQSA5V92Zg4JfynK9Mxxskko1qcSjzUYf4gLFcV7TE12hnVnvrqrvBbmLZtAZEgKew+SiQEfbSc4TT9YJje0xKTeJErnLzwoxvbTVzyFQ04ojn59kdZL0onMsT+Xt15VtZkmq9buPhHInH/G8pX0SScaidECqbfgodhhldZx2AUpzrbmgtzwdgtz4AvWr13+woIWP06rlTYz9m6BTUnFV1JyAFsvvm3Tze8USpQdXCEIcVjM2SmNLA3pP73E6/wsQrIW6nki4u5PBDGF0c6/pFfCeXQd2Gm2N0g3EFn3lNptIA2YuTc7ATjLEHKTMfmOCIZxRrkRFAyw2roHbwM0g75KFzTZ04K976Gy+uvbn0bEUa4ykaC+/BN/mM6hMbxaCAtfaSokd0trOJwnnVDn1sqvNyr/cEiWauofHjYq9vhv6cc7tP5gIgrSgztis4IrMmPsZj76dxkxelox8asYlTFTkfEvp74m02y+4RFbwmTbuSAGwXcUQ4FZzAioR19VHAI/mTjzB3774kvPYVlyNwPjuY1s2SpwFZQNVt1qIugetozNefMYMDTvKgAqp3v0BT6AZmfpUl3zjXtobNneFZcowUj58CMHkOgYfdUkGBuiioC+xWweNuINJn/xVh3hZsbyzM8XbOOEqnJ1VcChFlFOgcO0XJTAp58fxp2M25FFzV27ao+oV1OeZfaAKHE1lGX3YeJYp2JPdfW1JQ9npbmg1P6c9O1+RgBrL/scRYeH4rEGT/VuMVevZoBQ14kzXaf/opFwb0bIDAEaxf5+7/dvNaKAYw2MNV//4fepaoV3ikAsocgtw89BbCQ0q9iVlyjBSPnwIw9NAA//mYr6e7mP5C3hPnd0z7KyooCiOm5vGQlpP2aTRsRRrjKRoL7muK0febaj42NX8SSmljjU0Ab8R8SX+qQoj4CEiL+rFabm35VgN013alht1NYo93Co7KdVEu9A5ATBB7ErtggMqMb201c8hUNHbqqCDPGux71KM4KjsSLWRhrvt/y+YAdzhPy5WLVL5pfMxYTMgG9kek3SOpIjcczJJ7sSvFeigZY7GfGJXvVUbx1UxM/g1wzJhLEss7KIdKgJiXtAw758XamH/gDjO93hCHFYzNkpjRk8GJfbnl3SOfUPg+/LEG0G6h96qoENi2Ns4NBVtFnV645MGeQp/Jokd3rXe3ilhmEdRMGRdYD3AllpwxVy39gYUefu2/fBpuXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZtTiZMztTzKLJ+GRGEO4U9WUmLm1ZqCyDiEYU2GUilX0PWabvOQwxQh5nafVv2wVHKwVFlrSa4fnZ+NQ8IeUchEBbTe217ls/yDLnu4TwdG3l/4oVFc/5IoEyrp6E80Nb/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQky75E0BqC5xoA8M7MBdqNzOaD0aqz/P6VGCdAfSJQbfgYmABKohTdQLCLvgJmUs4yEHlVk4JZPDJR21zhtPqiFRwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+yzl1puP5iDP/GXOIAnlejc9ruZiEr/fw/tya6/o54mXz4emIpYW9lFN79dm5eVPJ+esGB8fwAJTGeu6K0lNTls2lJ26ewe1vL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZyoFMZWrhZk3HS0sFW/Gub0izfTW27Y1SAARy8hgXstCHOL+eo802L+LTQPUn6eOA/ZNH4bqOHFI8soFmqbETOmtD4F/KgD3CQnLeqDhtkvW6R4quGl2o/pdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm1EDF+eslQBLSXlGS7K5fkFFcZDqPf6s/HGc3e9sUZ2nkfcRwEJQISBLTGIGeBivlhP2l8bAAnxBPyV2GV/YmLSd6MNcmyk+MwUWZHyCBy9Jw1ldTe5/DDDc94ADxNcvl/usVL9gJwybTs4wFxcb3FJfe10w6J3nrhP2l8bAAnxAq5For5ln/meHDJoDEt9A9J6b+11OiNzFxIurGghkjiaW7AZH2cRVQhz1wVNvRMJoDDmo0qbnltlF3eSy6k0OCvM9IDKSSTtiQ0Q8ygJvXeukkKpWfySGqdi1rfWBr/+bgvCfaSCNbt85UIZCbh9wpkM+nJOcaRtjYI0g49L9yY5ROKHG0m4e4tY2ChAhRVj8IV+I0T08S27dHwsYS8hjgo1pWJmgkqwn6/c+xRed54FB5JnenTVIwghhVhdBMj3yQ0Q8ygJvXenlFTmHEr1hpeI9I+7yiZroAe/KElw75gWV42WujtM9ggypL2PvmW8Fx9OgdnkHJZ5flSbQ/7r+gliH6iLNHgScfqQUFHfyM4XH06B2eQclnlD0OSpHYJIz+tQwVim0IWlXFvxq60Zv4LH70chck88pyPXCr6PB0TOyHICzE5HxfCcSLje0H2Wzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNksW3Mb+3Jzg7DB042Xl1jX2GFVriH7Pzc9ruZiEr/fw/tya6/o54mtIJeCh/F2NAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu3Hm/ZH/aLtBbpxHe6C3zjI5KKRRHzgmbq+3uWHo09MTIiX21wO8isrBAUwGum2YW3YWhxFO8Gvb5iRsgxnwD527/LebCgOWq+e6N4jtRobADKuVfSCivqwGpkRC79t8iUuAH1jBo4g4VMZ8/4Eh00J67CWxSc/j2on6NxXP2f/lzyng9+sV+MVvRIhX62s/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv0jlKl6nOCHbCOjqeEmbrf5w8x7FCxIEFBZzTaPe77adLl4hH35McanPyYcPjMVpvtG1k0bLNkmZ5RRDns/Z1n8DwKRTyX3NLC/Akftdwe11rFNRFkT0e0y2MMpwoe9EBIlOUoh7DPDnU6W6ipCpMtn56wYHx/AAmXLoi95JK1wOxJbku+DGjG5elrM4Q2ayGFsfYaeB/EKeprxooDEabJyvR7VOaXDCTD9lqSuOVeLnrB9f+ubikYM0wKYLaIRvAiI30omj5uwjYw+DggAPAP7TBKBCAhyP/xaBuWUrhj6mO8wS+TYnIwb7CKGgQd+IkaXmHF1k8mnHPxd0F7ZZU0ZxHjVIk7Janc9ruZiEr/fylT50JpQ6IZBmmNrOWyAJ31YNB4puXDPq/jIpxUFunZIiN9KJo+bsI2MPg4IADwD+0wSgQgIcj/8WgbllK4Y+rBTB4wQehlNG+wihoEHfiJGl5hxdZPJpy97SL04EjNUAIyvvNAahmXn56wYHx/AAk65U3NQ3GzDDGfUzmQkKcXDJ9LeExL72SN+X5Qoeb1Fe7mlytUNHbR7V2TY2aqZZkAupHEAvr/j8oAxG2oU6OZZqjTTHV6cgoUlU5L/M5+MB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwty0FZSqHxxyyba61mL7BzZyM7HsuArKxnWKgQHJEW7mr+b1+0cFNq4p5R6wQtO5ErbvSeYB5Wlaoqq+DAj3H+611DFD/WjcsIsN0j05VF2845BsIBn4E+pXfnTACd7co8tUf2Bkgs2R3Kx9EvqNttpK0pub6IzwBdtGtQU15CxTGdqdYW/3K5vPGmM87YpdqeTgYgzk3cDU+p00MudCuQwYCjt+ZR5snEgjBkLRfibeoNfxJELxwGPFyASBxtXoUQiqHLlRyI367VPScSSDte2BHkSvE+pNC6MQRzpkwOn1cc2byXWxxM+WoQgOPAyYHcaedYlwjGXQpYRME7wDTEVMEYIEQh4M8ADSwUHORBcaj+94L6ft+sNhh8ZdEif0RhQg8CnWPp/Wk6NJIfkzf++2imZ1HdxrtavkgfnGzlcA4h2D1XiJ4sEN3Co9PiLr1p/yv/GIdp331Qh+nJ8YpcPyG9+8SzyeEuydG5UOuL9SBrLGU09kZcAvyMvOQGMG6G63hwq4PiB1eiRRDxm8LQMZI9Fpvu6q9AXyFJ9cP40xUyt1ibADTvstKWNH10tav41RtJNYUbU5mhXAYKQFft2f17ZWwanxfTRvQ+YFO5N12SIgV1sgWMeWsPLb3dhnlc+a37e9zPcsgfOnVu+8GOTaq5+B2jnlZINFniMvv3hgdvhS00oL+KEFeNkqdFZTJYjNePsL6IxC1lfWzpFP1CIb5a7LkaX2IID1wj5rVvW1PEoGwaJlpMcU3rtVsp6HQnHzgB2pXDwa/PDL3JFHEMVz6MUESbHZ7T0wAIi33AP95IIFX2mInntvjEGIa4q51PNqyLGdo9RMi2oo+yP+BYmOFgEJPnQZAWuoAXdJrbeaaGMJr/RgsKq9FlqC5SJHKDjAulTmNO9e5hvgntd6t+gWqG8lmRu0dNd+jCm87kHB5wWZQw1j0XNH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8L9fSYVdAYPBQF/HGAtb8OmSJ60jnZ0ClqdLRnBrMX4NKJrUO/ewCG9aZ+c1GqC/hSJhEYVrJuZEJBZzTaPe77aQ7LjgLlmoVAKfm/P3qSlZtquYMjOSvzbZvqzyrBAT3vQQ8OZ5dJ6G/WScFeWEM86CNs9/cmJsZL0oCK5Nw7o/HWScFeWEM86J0oIAp7uKg8sFAU5C9nfKJWNbV8zjtZu0mLyaje7hfOo1Rt6Fw6V9fqk62RHlAjuueTI6HE24di+4qJrPJDTsLKAMRtqFOjmbXyY4p3wSQhwvwJH7XcHtf1YNB4puXDPvd42g6CTnXogngZTYpYIfZh/AK6jyUPsZ+esGB8fwAJly6IveSStcB532mKjRs8Ag1fLXh+RnpyvobJNK15PSU8tc3YQOrzztJCZTW10xy+0kpBS5r4LY4+/8gGLek9mp3E3uavtjBHa6sMkM+revdIECM44M6zSyTns76LF6di+5w6DyHzunJHqlF7ubtva1h5E0gkpomTYDx0oL8iJkpmAmFR3LKaecIKQH9xapKWm5wIy7VEbo3tIPi8/JGwoF4JAwcpRs2wpWqh0Oh2IWULQ66nxKXucTrs7IZ1ypQh3Jw9PGjYEhWUzsVX+qjJ2cFhRLHtr5z2lMrT3GRkm/U3VEkFOPxs0V4JAwcpRs2wpWqh0Oh2IWUcyI5pET4IalzGchwav//MwV5kUMSlBLg/AaikY3kVDlKUnG7T12N5i0kWLnusckK6maR0RWksW21F32Il+s4UEtRfj9IyqtXPgXetxsYfRR3bcYOqDhgjKJnyGPmNyWbhwyaAxLfQPWpGPxRfAM1oUcfJNDRFkYxQgnJmgVSSno37qMTokd4LNDt7WTzRCmcfSSbQfgTQYg+w5CPuIzPya9CKQlY8TsI6Sgfx+Tritgwdk2R1rKY9KyiyGAu62Zo1Zicz6VVMhCi+G04JfRlATHuAGfcsPKDDUgxQnnMPO9kTlmHI0o6TIdgmsrSlvKHkjghcGjiDYSjfqPGNwc8LzeBWtZqC043c9ruZiEr/f+iNuPW/CDp0s2viNXujF4FBSmLbge19npwRI0iJkowNK1itPE1WJx+541HACg0JsjpHZex+pcjKVHradYcWh6s/auhmEWhjBcVuQ3556WeSvJ5wdRfQYQaMw98LvuzZjxcvUS83FcthRoT1ujn527CRrsOe4wGmcXRC9BQrQSJ4g5gqzDThQDlrMd5VsR3PnSDFEXspuZugTrKJJP5gB48KNuDTzDWbKm3gjXOEok0S6vEkxNeBBm5pjtT3R1NdwsY9sbhti4aWnGRy423rjn4yJabVrCkUkXcKW6+dKgEYDp29fNwR3gn5mIpPSMlFCwSoFZbQkvHu3hI1zvf4/zeLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhRvsIoaBB34iUJD9RYEgn3vkoejOOHQ5KMomfIY+Y3JZuHDJoDEt9A9FIjp1DOt+yeysXhkHKmrsPqesaXJsluNi0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+In52yY94aShOzGTzC+tFdi17GNtU97kTE2caiSB0pwUU/VvfHslr74/+dsmPeGkoTsxk8wvrRXYtexjbVPe5ExNnGokgdKcFFMPersQfH6Va1bLmetxGx9zq+9yLK/bVb9SUGx8Ab27w+w8b997gxGgFIjp1DOt+yd9am3/OvHnzqvvciyv21W/UlBsfAG9u8N68qlQJLzMWPZSw9kAR1FocwdJmPvf4L4U4gAMoeB/kOLB1ganHNIpghX4L1x80hEYc/mEl1wDHrTP7k/Crfx1WIIAIds2MSryTKIkUcCMHWKdV79OQM270hWS+9p0SADV3amXOXEZSonXxmFhT0zanGokgdKcFFMg4wXD5mlLkNIVkvvadEgA1d2plzlxGUqJ18ZhYU9M2pxqJIHSnBRT64pLFBtl8CUNGJBfAmFVQ/2YYgi6qQBhzm2wZnIT5MfhwyaAxLfQPRSI6dQzrfsnQlrkXNs7jE9udQuF8S7kS5KHozjh0OSjgQnjE8gCmM3hwyaAxLfQPRSI6dQzrfsneiHyb/5OcdVWfUwRq12c9GMF9WizK2bjHCmANQf1H19r0IpCVjxOwivkwtmFLeT2axhN9NnEA2u1wapN/sxdpzBuOxooRq5OWIIAIds2MSryTKIkUcCMHco4acBHHgDeCB/Xbx77ZFmLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhTbA8chY5Tt3EaE9bo5+duwjEw96mKSyO+IhdTrbbAMB1RWHJYQ/HeHQW6A1k/HcyOMHf8CIdADG+hIWnndeRrgiIXU622wDAdUVhyWEPx3h0FugNZPx3MjBTQ/eOUN9k3zmlPnVztZ/76vp/Wlrty7a9CKQlY8TsIr5MLZhS3k9lp9zaVRPi/Y4whKhojeXZ2Sh6M44dDkoyiZ8hj5jclm4cMmgMS30D0UiOnUM637J0rtiOc50uUSNuA1T29vGtnCCD8Qa/jQUE5Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCT6ovuNWQ2fynSIhbYck6hU1Zicz6VVMhCi+G04JfRlAVFYclhD8d4dBboDWT8dzIz1fALIrSJM0waC0+B0LF+mLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhRe/3IFH7+KMEA5qv8I5YVt/pLtyZcLyDV1YKbw3tpRShxHLifkb0sGhVUg9RSnF7QEOVkapk+qdsyGWQquamDBPS2honXOFi8RaygtE5naOViCACHbNjEq8kyiJFHAjB0Lj0mYYo9g6KuJrP4Ul/Z5ciwtx2yRK2IQ59kSE4goE+dK/+s2YPEJJgGuAYBghdiz21yojlDyZhJff4DZ0CW6nZkh6++iwO4r5MLZhS3k9kM4o5uTlB89Vn1MEatdnPRpKqP/7DJnXQoI1NNC5RgMoTg24V9jXfozz39o5xxx3EsB2DYr6xqhfM4amjHtWCAmrE1CkbN/Yd+Vi/JNyV4hBLRI3+DyLvnUjJvBEBrO85KHozjh0OSjKJnyGPmNyWbhwyaAxLfQPRSI6dQzrfsn3b+3M0b5yi925uOVPuyY8XVgpvDe2lFKHEcuJ+RvSwYPC3wxD/VREBGBl/cpTuL5OiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHIRFJnE6Dc1pfpb6n37APDoamIuBW1zP7ooSCx692z/0+ENbGpoR1eDl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGau8gT8cx5ihtlv37lTTc/yJhKqbAPrHo/8UnERL5ba7Bw2TEYBX3tTqxiEouaRpssvFfG+fBhu2ssCk5CiXq3flyJNSZWXY3L5W+rEb8XoruEkpZ1EwtkIh5qeR1uvF29IrieUBknEVxt8p0X0CdD2I/6fI0QRgF12zDobzDo7Yag18ZZFxsrfExjs5JK/Inbx6uW325OK0mz8/3OvySf9oj0QCQIThh6SoGtWHrMQoF8Zp0AYsJN5NDrz/dM09R4aYzfjTC6+kbOm4GNjZXJt86hhd/8v9oanGTQoBpT15m4JQmX6vUqjr52FJW9ZFldXmAeYqCVGIMxBPmd3IyJnOyxQZ13Y28ciwNAP34iStikJuMch/Os1uWDl+4FOsmiHmp5HW68Xb0iuJ5QGScRXGGu+3/L5gB06k+0KUa+B4uRpYN5qRry4fituwZjT2jwxnN5zg1hvpmKARRcdxh2ubEegyaglFcoLXkwTLBM2QP9VOEEPlSHPQkP1FgSCfe9rH94qFsHdXGWxPwOOlMm6qDXxlkXGyt+pfPtPcln2uJl+ArswASgGTVP9cq4atqRKrj66insYQ145BQ+wFcZ4JemFYOlJLhlXlwbgmXVaZVbLmetxGx9z2EUZMhFlD11Wy5nrcRsfcy+qjnbpvRI7C7fC/pB1QEsQ9BMUbPYIW3cMKmb+s8surTIP0x/AMDCbsKX8kabh1EzM6jWgHkBNdvgvANcb9+1KLpKtGGwQ3nAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR+Qi2V3pcu8vi0ObZKSgLuYiqp5DnfY4FjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyqf28mTmm3ajORD6cTjZ/wSZ/SDtPy6KROZ2MLP56m91/Q3YtcqFzn9fzyeLG5RUgyTR+UIzCD2jV1nSmtbA90OzKeOakhOUTV5gHmKglRiChKlCAG3SxEo4v0hUlM0ywfvOR2XnFrlVs/P9zr8kn/aI9EAkCE4Yeslcs7/TDgkL2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTLWW1EiILdaodZYyOrKEyrgUQlm3kjqGg3mJGcwwwWk+/cYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaKPt1+NzKEkemQuDrbCd8gTbcimc65tP3FeYB5ioJUYgwFgsHfuuaTCRkfb+deNGY9GFYs/U5H4LiE51hQfB+RfhJKWdRMLZCMBYLB37rmkwExjs5JK/InYOekTqZfSz50JD9RYEgn3vkNEPMoCb13qb4UE/n9X7qxhrvt/y+YAdN+plWTQJSyzcLmzY0YOPT2BscT8ZbRQBF4AjPNeCbtmDKkvY++Zbwb6IhgkZZbtU/1U4QQ+VIc9nrCxK0k63U44v0hUlM0ywTKVS+fDCQUJqORwzQdMkxZDRDzKAm9d6QHz0jGxd051EOl68b8i4nYM+aEC2mLhmax7M6tZYeK72iuplgCAem/guu0FDrIs+f74jSUDzvLGXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiY7+SuqaCode+zu3no+i50PfZB5ZkedC8ny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8S9BuRSyO60yrZolxh7PHEPmjKghd4lsWyyqKwAqktn0G5ijMvAwQDKo1fNd3oasbYAonLDhVfq5i0kWLnusckICca2Mr6/QFW1F32Il+s4U0kfhGIVJ+sp4LB8SnYnkWKcZNCgGlPXmbglCZfq9SqOvnYUlb1kWV1eYB5ioJUYg+QXlou2+5t6luwGR9nEVUIc9cFTb0TCaAw5qNKm55bbJZIJ3xSMlNzI2uIlbK1BwbTBt9inE+0WawCCQAbl/Z8Qwhr2xk7+pPoez99LOs5SqFPCWg5/NPjiKfefDbPYZtJelJ2P/PoGQ0Q8ygJvXevaLSfHmqIyxEdZ4f8IGfUHEMIa9sZO/qbJhmqdyUVDjkNEPMoCb13pYa18FP5By6aFOWhvQIMdb4axIQeSuScHVwtYmcO0O7PCDAdI6K1zorTIP0x/AMDCbsKX8kabh1EzM6jWgHkBNgZB7BiR2GnQVDR0wpi/825dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Jn0P/l3tv2QupHX/7psnIxumrIyMmM53oPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyBhIwYo4qRNhyqqIMZwKRImXmk/7/DktWDwz9c8cX2oM3yHCRp5cv16eTMFa3S0myHtmpgoIVG9A8prdwdBC/jSFZL72nRIAMFD/wr6SBxXKX6FkM9GFm4BgJmCwtDu5m1F32Il+s4UIe2amCghUb0uwY2ce6+DxxBP58I61nv5UwM17ovWmnI1Zicz6VVMhJEjGY8/zfpUVFYclhD8d4fm/fPgGiWhA7BvkETgs+XWGnkhHOWLndeYUieJ1YegZdiuoTHUj00c+tO9WaI/1O2CoUVSF6OrzeOnUlXGd5qDUQlm3kjqGg27cHGcmccaLau89FjbHlF3E9c1gpRGLR9qkXUdqyH+T8ABapzRGOwDl0ZJAso0G7j7rF/xkd94BDQ68/3TNPUeLF8Yj3+jKids/P9zr8kn/SVfbovfMR6DCZrVxtmjyhmzpuBjY2VybWCtwhOHF18XCJvvwm5Ml1YlX26L3zEegzDCDFQmIOwZqDXxlkXGyt8MHZNkdaymPb5zxI7TXmNiUQlm3kjqGg3mJGcwwwWk+7vI+FEkJseP/gxqQLfDQTr2qgcg2eo1NMOTyNLgcNdkQIaAy+tSTHGq/E96ZInMfqg18ZZFxsrfW4lF02g4zIcN4iZMez+iFzQ68/3TNPUeGmM340wuvpGzpuBjY2VybUzVQvBu8/R3Vn1MEatdnPTx6uW325OK0mz8/3OvySf9oj0QCQIThh5tvMG837M6c7mUbQZnv0hfu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6Pqi+41ZDZ/J1AyOSpe+YWDQ68/3TNPUeGmM340wuvpGzpuBjY2Vybfw6f250hdVyNuA1T29vGtk0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek6En4vhJZYh5qYtNbAysCwf9qoHINnqNTQT1zWClEYtH4XLjiOTjsUyO410o0DKE5eAXTsdYWVnwH7zkdl5xa5VbPz/c6/JJ/2iPRAJAhOGHsJ+MHSONXBWN5kVkgqLvuRfzlp9Qg9NWVEJZt5I6hoN5iRnMMMFpPsDUuqo6zWRC8yGWQquamDBH64dY+z+8hJAhoDL61JMcTfs2T3tv7quG3ynRfQJ0PbSUoEq+NKnzq9oqnTXLVq558Va0NGz5C7jqS2b4yIpdmoHFWraxW1GwpO3pOPxV1mHHwGW7ErLXo0vYS1flZR167Cu6nIIXDbISx9BdF4ZgkyfiZMSzGFCsDBYXILUH7UtmJaBJcfH6g5QVL/BuwBLISegBf2ypJK2vJPqiQo57Iu0xcAZ+nMEgGwFmQkytbgP1ziX8hdVw2N7AhKNvBXLfCf1a1PYXmtrLsSh2Hw2xWbvhUt/OZE9RN7coAtNOaQ+JSMIiVeI2UVPA3bfKsDPGx82ThwHw/VwQ9XNkx+wnzQOaQkC+0Z0Q098R6xZWnvzO5I80BpoNW60EP5yEYLZQvZOoeWO9V/RuN+zBfi0eM17+agt1qmn2K6hMdSPTRypKYWU3R6ZbCcgJfMYV6lho810znO5IsoAWnyLD80cW85x44xaDmPTTrCUc3nn2fBU7zspTuJgGlyrEwA3hrVVidfGYWFPTNo8Rp9SfcLUH6g18ZZFxsrfze5FykcdWSY1FvD0r62eQCWzqJSeg37mLOVyEv2xjpqQ0Q8ygJvXemFmjN23bm9w4+UXIMII0IX/VaSxankcdm51C4XxLuRLje42oZa0ePviKwa24/UsHaj6DzhqWt0p0C6As173b7Dpd8Sh3Famxv9VpLFqeRx2bnULhfEu5EsWQjte9/SsM+IrBrbj9SwdlEzuUcQChQHQLoCzXvdvsH4rbsGY09o8GqL7zgrhAFrISx9BdF4ZgkyfiZMSzGFC/5MkbzKdlzrAWCwd+65pMFuJRdNoOMyHDeImTHs/ohdhnzKtQVN2IoKhRVIXo6vNF9VwsBAq6Q2zpuBjY2VybfcaLydpsQM0W4lF02g4zIeIzbG+JEb+nlnIPOi/OFb05iKqJZa0Jmr6071Zoj/U7VZ9TBGrXZz0h/9/eVSu7RcnICXzGFepYScjgeVVuCXbm+FBP5/V+6sYa77f8vmAHSYBrgGAYIXYqRVQDWRKrRyo6cpw9AXIXIKhRVIXo6vNhgKfsczLG+KzpuBjY2VybWo5HDNB0yTFAoHnaArgPt0OUFS/wbsASyEnoAX9sqSStryT6okKOeziKwa24/UsHVz1xIy74n4cG6EP0zkPl7eblGqqo1E5zIL+6S3WR4x8SRfmKYAp9StPUa9cVNYyUvLjErJt1Zu4Aad5VnW3MWqIzbG+JEb+nhqWmfBNaDlHGGu+3/L5gB1ZGCWJsTZkMG51C4XxLuRL9qoHINnqNTQT1zWClEYtH4XLjiOTjsUyb5lhdorn5WioNfGWRcbK30zVQvBu8/R3Vn1MEatdnPQLKxBAUy6zhJdGSQLKNBu4DoqPZV6l5u/ZNOzgsBdJGIMqS9j75lvB0/XDJL/dpKumYURHNrLDk464eaCCUZTwRsSBNiRSt2XvXPm97zBlmxhrvt/y+YAdNmKt02Bl7v3RdlEeUweax8BYLB37rmkwPVkGDmtZH5ZIwaRpgISuRLWNgoQIUVY/pzJyI4BKxS4Sc4euQO4jt4sgXo/zLRX3mSwmtAOohQT2IOLpAEyxNchLH0F0XhmCikrBdE183dfAWCwd+65pMPN0eLAOXXJz0hWS+9p0SACY0t/+1Ijsb1PE/sgT7J/pmceagzYIXt1cqxMAN4a1VYnXxmFhT0zaYvsolD27kpSoNfGWRcbK33mI+vqzK689HK4J4v+hznjAWCwd+65pMG0tBOzulMIx0hWS+9p0SAAf6NiVFXsIpf5Y1Tpf4O5UqOmaUV49yKkmAa4BgGCF2InXxmFhT0zaA6h4hIo1ccOoNfGWRcbK30r15D2mwrLWXKsTADeGtVUSc4euQO4jt86bzEKTHmug2TQ2S3XJ9s/53/e3dBzVMshLH0F0XhmCikrBdE183dfAWCwd+65pMOeH528NwAgyDx6hfzAOp2jAWCwd+65pMN6dmOV1R27i/bcV14ilCVqNe2agDQPBRC2yWJJ6HpAO+UtuVdqoNh50piTdNFHVcRnTKHp+eudmZ5wVn0GGC8Adv+CffYE3kcBYLB37rmkwyM/eT/vvYQEQT+fCOtZ7+VMDNe6L1ppy/ljVOl/g7lSo6ZpRXj3IqVkYJYmxNmQwGdMoen5652ZDI3OjB5QrsB2/4J99gTeR7Gfhw9lEZpvG4+SZ6/62xqg18ZZFxsrf/1WksWp5HHYZ0yh6fnrnZq42YXW6iBFoQLNW2v0RlFgZ0yh6fnrnZlrzBFLlvN8qAYCZgsLQ7uZgKQCidZsjAFuJRdNoOMyHJMLejpnt+qiQ0Q8ygJvXeg5QVL/BuwBLCZ2gL/8pNVN3DbuM1kCXJyDtoVjunTXW0hWS+9p0SABOfUTJvCYpZxHSZZkqSsKs7chJaFAGYb7XC2r55NXyEAmdoC//KTVT8SA55FGDbLAASlQboJTlvhLubMjDCne3qDXxlkXGyt8F47xEMxrtngs34PdN1BBatP/8iyWTRROhG37csGjubrmUbQZnv0hf+VeIlTrTM+5qBxVq2sVtRsp0L1GaQUsTbWqPf/e7KegnvS/Z5hBNukK5oDZ7hM+0+B3ElgcNhzMDCX4eEODRaJZPS1/oJxSYqzUqO96X8MWoNfGWRcbK3xS9+cdPvQDIZCEv/049WIweZa/KEJx66KYCR9FIteE2qDXxlkXGyt87jXSjQMoTlwaILs5SWlCyrKG5K/BdbcHuX4Qmk8dgjsBYLB37rmkwQoDhL/tAYsRIwaRpgISuRMJ+MHSONXBWOWzy0Nx5asGWJJBxr2B8ui0AW62GiphKGGu+3/L5gB1OiHWQHxWMsEv8MthD2qTcA1LqqOs1kQvEwjKBp1lR/qJKVWyyihRgIZWeROrGVeKoNfGWRcbK39GgdXy+4gfpkDDWQuD1gJbAWCwd+65pMD1fALIrSJM0mnLUpQStEK4fV6Fy8mFeJkhlkQm3ExrseYj6+rMrrz2LcIkEMQKv+Uv8MthD2qTcL34jfyAKTSye3/v8nWoHdO/HV9gw8h0RCTRxMgdUGTvMQT5ndyMiZzssUGdd2NvHczq9vXegaJ4pCbjHIfzrNblg5fuBTrJosG+QROCz5dbDHzwZbJ7YC6ZSXhw4JRYfvxFCll4lpueoNfGWRcbK3zGc3nODWG+mF5TvcqXOBv1Mpsmp4wz2866MGUd0v7RjqDXxlkXGyt8xnN5zg1hvpiggprp1pzOUTKbJqeMM9vM4mYBN5SukVKg18ZZFxsrfO410o0DKE5czz8ckyViae6ISItNWpOCYOWzy0Nx5asGfmmS/7b21ALxDUrSDsZSCQDmq/wjlhW1Atle3BsPd5j1fALIrSJM0wlrYvtwE9H7AWCwd+65pMKl8+09yWfa4wFgsHfuuaTAMHZNkdaymPeCEsyAb0kcwzIZZCq5qYMEXgCM814Ju2cBYLB37rmkwDB2TZHWspj3lTdi5zjJiVMyGWQquamDBuKPqxC7RtK+DKkvY++Zbwb6IhgkZZbtUAEpUG6CU5b5rHszq1lh4rmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa8KqUVY8Z8/lUG2DfJCuq4fy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOFJZfy2x950437qMTokd4LkIbDI91ni1wuxPUN2+8SQheAIzzXgm7Z/id2tyC4EWyd4/Q3+4GQ8wwdk2R1rKY92WaafzXNgCKXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZqj/hYUlbLd7JWttJIIaWmW1SDjomtrsiLcJYGK8HkqvC6aKeiD68NA3lTjMbfbReIQ2YROC9cK5srylMMcxKxwkG2HUVfrdqq6H1onROXnd1B7ulwg9TIMinJhsEsMEyFDsTaK2LyoCf8sEkm33TSjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2Q26j4q+VAd8HG4tIo5YEpurKbRDLBZ59moUX5Omw+pt6vEkxNeBBm4kcueB1sYHofqXQWapejhd7/wdIripxs6P2Y53F7m+a0CAuwH0oe4Q2zOL0ipploSe9cCWsav7W5ELeDiO4EYRG+4V5eP/GKitvZvcz7NvWBIRvupT+fBRegvh1ja3Ig0+EJ7MuzrICsLaZdYiWxj6CDAM8YgYDHjvaU6w36I5YK53VJAQUklVDbqPir5UB3wcbi0ijlgSm/03qOIzJ5d08v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3Z/sInISWfk6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZJxySuyuWh3uG2wQmryA5pfaoV1U/wv+YeQNK+vHa1FwL39q2OrdvMfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxX7OEBZWYvk346SZL/SDXx6z2YvovkAtYYAcQM8A6deifnrBgfH8ACaMde5OBYCMAaAorIsEFx+Ckf6Jhc3anln+gJk042NZfA2JbNZXiTdJq62he6O2yeTi8sDixjycgKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTyNOGBYR8d3lONOQJDgAgCarT9KQ3pbn9GesH1/65uKRg0DDZRAYBhdE8aGoZki/xCLEXGmfgOzLOEuUcVIElGxfZf1NxPMwd60BiPpbsi2boF1EJV5+ymbqPA8XIE0tuMKaIn7NYNLGIL5ZgXVjx77J6uDga56J/0QkP1FgSCfe8L1TEereSyJhpeYcXWTyacsVty0jvqyd7UJQM043pMr14eOBK7vhtvwxXRPxIwFah9jI452is3oTo76zuFDULSeF4C0mUbSnUPyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoPBJmRrhKB5X9sqKEd60d2x2N71FU5195hOXwpBrxr12isR4oKvE8eWOhqVPaMD2KgJDYB2RmqX0HB8UTeMQO7rnswU3AY2t2pCkjmt314ynwirMmvQ7qtlJ3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb4MHZNkdaymPYNZnRYrjGgmv6uQ1bQ+V1P5g+3VUkwsBNEUaFVzusiycCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMMihLJdAxE+aIc/j4NtRsPsNMwfWlh5XJmqNNMdXpyChSVTkv8zn4wH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3LQVlKofHHLJtrrWYvsHNnIzsey4CsrGdYqBAckRbuav5vX7RwU2rinlHrBC07kStu9J5gHlaVqiqr4MCPcf7rXUMUP9aNywiw3SPTlUXbzjkGwgGfgT6ld+dMAJ3tyjy1R/YGSCzZHcrH0S+o222krSm5vojPAF20a1BTXkLFMZ2p1hb/crm88aYzztil2p5OBiDOTdwNT6nTQy50K5DBgKO35lHmycSCMGQtF+Jt6g1/EkQvHAY8XIBIHG1ehRCKocuVHIjfrtU9JxJIO17YEeRK8T6k0LoxBHOmTA6fVxzZvJdbHEz5ahCA48DJgdxp51iXCMZdClhEwTvANMRUwRggRCHgzwANLBQc5EFxqP73gvp+36w2GHxl0SJ/RGFCDwKdY+n9aTo0kh+TN/77aKZnUd3Gu1q+SB+cbOVwDiHYPVeIniwQ3cKj0+IuvWn/K/8Yh2nffVCH6cnxilw/Ib37xLPJ4S7J0blQ64v1IGssZTT2RlwC/Iy85AYwbobreHCrg+IHV6JFEPGbwtAxkj0Wm+7qr0BfIUn1w/jTFTK3WJsANO+y0pY0fXS1q/jVG0k1hRtTmaFcBgpAV+3Z/XtlbBqfF9NG9D5gU7k3XZIiBXWyBYx5aw8tvd2GeVz5rft73M9yyB86dW77wY5Nqrn4HaOeVkg0WeIy+/eGB2+FLTSgv4oQV42Sp0VlMliM14+wvojELWV9bOkU/UIhvlrsuRpfYggPXCPmtW9bU8SgbBomWkxxTeu1WynodCcfOAHalcPBr88MvckUcQxXPoxQRJsdntPTAAiLfcA/3kggVfaYiee2+MQYhrirnU82rIsZ2j1EyLaij7I/4FiY4WAQk+dBkBa6gBd0mtt5poYwmv9GCwqr0WWoLlIkcoOMC6VOY0717mG+Ce13q36BaobyWZG7R0136MKbzuQcHnBZlDDWPRc0fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv19JhV0Bg8FAX8cYC1vw6ZInrSOdnQKWp0tGcGsxfg0omtQ797AIb1pn5zUaoL+FImERhWsm5kQkFnNNo97vtpDsuOAuWahUAp+b8/epKVm2q5gyM5K/Ntm+rPKsEBPe9BDw5nl0nob9ZJwV5YQzzoI2z39yYmxkvSgIrk3Duj8dZJwV5YQzzonSggCnu4qDywUBTkL2d8olY1tXzOO1m7SYvJqN7uF86jVG3oXDpX1+qTrZEeUCO655MjocTbh2L7ioms8kNOwsoAxG2oU6OZtfJjinfBJCHC/Akftdwe1/Vg0Him5cM+93jaDoJOdeiCeBlNilgh9mH8ArqPJQ+xn56wYHx/AAmXLoi95JK1wHnfaYqNGzwCDV8teH5GenK+hsk0rXk9JUlaeKssDXG9Z+CulQJw8O09JiKzD8Imx+Hqxs2JxBciGPwpaYAvbnRZYgTtv5fy/gbJiAeHyu+YlLgB9YwaOIMXjIUSRp5iLOqYLJ9NHkvPVCln62da3lgmpZsQwb0+snFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/5uhHwoq8y0TZgJhUdyymnnCCkB/cWqSlgg+s3mBdZzXmQuDrbCd8gRxX2xf0wa4olMzMTd2VbLANuF9Szb8bc+z9851P7X761CCcmaBVJKebEegyaglFcrBIhwyo2i2bjVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3h5V3hyOyNkFbVNq16QQ5YAQd23GDqg4YIyiZ8hj5jclm4cMmgMS30D2ncXb8pkNlLY1eLN8gFb0Bi32YOSX61agxk8wvrRXYtexjbVPe5ExNn6ADi5zKCB8/AaikY3kVDkDhLSa4JNSDdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDSQAYMCrv5UBy5MK0fr/Ekvj10qKusZM2UtVYLGusEUFCFBodbJdoT6qQD3q+pGjRHEcuJ+RvSwZzysUlAo8iA437qMTokd4L/R/M3OKuO2K5DrFj2qvbOe95b3xuiqJ14cMmgMS30D349dKirrGTNg7mSHva6dxXQhQaHWyXaE+qkA96vqRo0RxHLifkb0sGc8rFJQKPIgON+6jE6JHeC9z/BkSUmEwOuQ6xY9qr2znveW98boqidaAzJs48yu0oxF5kW0MLn8nqjfeSSZh8UTnPjBIJZ00gnTLGBsENvg1Ldx1LyjwnRBYX66Kl11/PeA9CCZgqZJGJPW1XcIzx6POdE8vmZvuYFhb8ufRX5WPhb7aPzDOIdGc9zFDouWxgDt7YlkeJWPelXB2CrM4844Vln4aeijNFOnkRQ0EFx9waNwtccnXh+bSgrDKZFC2O0e6g3s0CwG1JoF+NBx45uLDl1Bw7HnEHrbAILbb24aGCYxw5yUtCpARtQRQh4tEFn+EnEsMe/bGKAEJjHMmaFp15py/8Y1MDPh09EGhq73BfnkI5Bo5EwAy4dHIC0TIQBAMmJlrRzaZNz7Ynn829TwlSnl3Qx+dwlo3fyzz2+XS8ig6NpXLZ/eRaK+jVTVinX9+z5o2VVRKd+PUEHlV+nsdVqYXWvVIvg25hq63YzbgVgrkjnb/QmbU3CQ59Q7oH8KCAxM1CeXCRohuL8WB/hHchof7A9tqsHO9FcwUlYu0O+z3TIorV+eHbonLmuc8Ea3t2nq3CirttY9L7Go8VjP/cjR+QxC6yJlQmvozb6vAA1+8fjJGguZ4Cfah0eHXQWJ58OqDN5d+EWtV+XTBRAViC45K5VR0bcaLx54mnbZ8m4Olu28ijPBsRRrjKRoL7oLnN2gCsPuZem4qWpsGiCUe4iM0H21Y6Ek19laVEoLwYQw1GPBH1QSTIi3d1F+AHf5ZqjnBY+iuyiJ+CI9ePduPUTc10Cws+TOHS8MWPAZUCFReMAR0LSPnpIl3Q/lMedlJAD4jO2IoRMXXX7W1IccHI7LaUnBArpnqIHQI6XjxdBi8ahMoUJRDnDED+DY8pGkgvKqYG5M1eCTa5Sotc2n+lHELMaANRhJw2i2oF+xGiolr/ta4VTtitSxOx6LSm1ngfALF2sPycVcLAF1MMVyI8XQoy2BqI0/V1T+XTxq6wdKFZiBiDlPaipube+GnnrcwHu5gS1vK140mCRc7vSWGdQGR7Fmlr84XGe6EEjYiq1H4gHDRrKP76MBoD4WK6DUNvifqyWwlcLmBHYSao93EcQuaPE6ShtKXxAi0+WtdS0XzUIa6BvTndIcmrrctBTRU6KgQr0ZUQZYrxVtXQgCerPndV1LXxYkA1AoGOy5h6jMQSACjA7IY/Ru7H9kWbsoifgiPXj3ZXrlhhA95gwwEmRmcFdDBZEGWK8VbV0IBD/zn4C/Ux8WJANQKBjsuY4/ObbSy9m9mcsumyMmIxkg4FZzAioR19RoSZ3hFIy88E2ZgY49Fsg+v7ZDPIZj5C+VpCcMwhcDYugPLosyYZTT6RmXHggkwMqd42Pjm38TYHaNQ2y7XxdbVAv9+1wyjcgzjQFFAq6vDhGVl4ORyBSB2fsw7CTQN2VsVsYuuTCO/sGGVMDYqF0tTYErX67tvDcICN93vFAvYwJ4EETcBLLI/Aod7Q1SgfzdcZ7Db3q+GmP7bmU3mXKQAB4LgJfBifX55COQaORMCBrN6pe3wvMQSEjmjIXHlaBISOaMhceVoEhI5oyFx5WhTrxifDjJVwxE/4L/XDFvU5wZX1g1wD5weT3VBaTlQUZ+n066+JUgaQwAFBTTMvyyrvwvNVuPSWrMZL4PvkWqqzbOA+KFFxN7Ns4D4oUXE3s2zgPihRcTfI81TG9lnq4MRP+C/1wxb1HiI6cfs8sU4uK+PwVNIwjDawSr20lhs48PALAn8jHo4expClmtLdd+dK/+s2YPEJwJQiQW/mp7cjTD0h9C086g+w5CPuIzPya9CKQlY8TsIr5MLZhS3k9of/tQ1TnyNOBKdnBX/pvPkRaygtE5naOViCACHbNjEq8kyiJFHAjB1pQKpSyhKwaaWFVpJ0g2P5i0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+InLfoZr3JwgyMIIPxBr+NBQTkGSJu/s69jC4OEyxUpTD+dK/+s2YPEJwJQiQW/mp7cFUPI9CR2jkhJ4GtAsMnHhOAsiQSggdl2CeH4d+g6s+UFugNZPx3MjYSBlwfxDgEFgbaw7GcYS51TM/LO5RPzdAYCZgsLQ7uZtRd9iJfrOFG+wihoEHfiJJ+K7bVNLNKg4v2za4HkzQPIgzia1FgSK/wHRTIPKtp3xGnuR0P1b1yvkwtmFLeT2RWLIkthUexk1Zicz6VVMhCi+G04JfRlAVFYclhD8d4dBboDWT8dzI6wA54XoKjzlIXPT22KgGxZa9Sh843vJFuxjbVPe5ExNnGokgdKcFFO+TTt0tEZq+7/ux4kGVmNUUzZu75YUdPWuQ+RKuafW5MLg4TLFSlMP50r/6zZg8QkHAZRyjFo+ubnVjHj7Rdt/AhvdyTLloBFYggAh2zYxKvJMoiRRwIwdSXFnkheyCSVTEW0+kmGFFjawSr20lhs4/OYyC6BzaD5g7ihwIejMkJuWjUz+uQit51tNIpUD1d8ib7252sczrfjPK/2Pd9KiWIIAIds2MSpcXFaU77b1OzO49cI1zPwMOOCrltLRHToxrpe6CThe1+dK/+s2YPEJJgGuAYBghdiJ18ZhYU9M2t2S1Yr5CIUpHSMNywugcshaUSRYR6f4J3oh8m/+TnHVgqFFUhejq82WjuF0pMCBqyqzwpefquLiFIjp1DOt+ydCWuRc2zuMTy5CroRa+KGQdVbekXCanteeFO+rSdcfihxHLifkb0sGhVUg9RSnF7S1Ut3ldwINVZdGSQLKNBu421MolEyZoJ/zmlPnVztZ/76vp/Wlrty7a9CKQlY8TsJuVjd/BSO6YcVNzNk/5DKQW4lF02g4zIckwt6Ome36qLMKZjxaW7VpbcuKYkbpcAjsY21T3uRMTR6upvwO+xTcT0KdNXFje9ijprU6DGn78i5CroRa+KGQdVbekXCanteeFO+rSdcfihxHLifkb0sGgK2O/wyEwTNBboDWT8dzIxl1r2Rqu6xmCZ2gL/8pNVNiamlU6AXXnehIWnndeRrgiIXU622wDAfgi4lQdJwJD1pRJFhHp/gnPzqlayH/zDKXRkkCyjQbuNtTKJRMmaCf85pT51c7Wf++r6f1pa7cu2vQikJWPE7CK+TC2YUt5PZDOKObk5QfPYKhRVIXo6vNWvJKkqbtOlkh/4xmHNo4QZ4U76tJ1x+KHEcuJ+RvSwaFVSD1FKcXtOW+iBe0HI8E/bcV14ilCVqyCArkcE/Xj/OaU+dXO1n/vq+n9aWu3Ltr0IpCVjxOwivkwtmFLeT2mHf3VIygpZMJnaAv/yk1U+NUPNETNEP5xh1RiIaPm0zcFWd01q9Ao4HGXTL4rBS7bUXfYiX6zhRPmMvpT+7RNwGneVZ1tzFqV79JGu1p7k1xCEQ9J2jli4610hrQflL6WIIAIds2MSryTKIkUcCMHWKdV79OQM270hWS+9p0SAAGqhihxL4Kv8IIPxBr+NBQ1hAIlb2xXDLC4OEyxUpTD+dK/+s2YPEJJgGuAYBghdiZTpXb/7goNd9jcx7OO4uWOIzwpEsi3BFYggAh2zYxKvJMoiRRwIwdM89/aOcccdwQT+fCOtZ7+bYY6oUv3wG/koejOOHQ5KOBCeMTyAKYzeHDJoDEt9A9FIjp1DOt+yd6IfJv/k5x1YKhRVIXo6vNtSa/p0vVFfYpfoWQz0YWbgGAmYLC0O7mbUXfYiX6zhRPmMvpT+7RNwGneVZ1tzFqjmGT+9BfA0VSZJyeIAjc/yLhDy3lF9cj7GNtU97kTE2caiSB0pwUUyDjBcPmaUuQ0hWS+9p0SACSJnKM0p88PMIIPxBr+NBQ1hAIlb2xXDLC4OEyxUpTD+dK/+s2YPEJWRglibE2ZDAuQq6EWvihkLrOnDbrhW7+CzKMGFbWp9ccRy4n5G9LBoVVIPUUpxe0tVLd5XcCDVWXRkkCyjQbuK+f1bMKiqFfxuW/DlbnzdscKYA1B/UfX2vQikJWPE7CK+TC2YUt5PaYd/dUjKClkwmdoC//KTVTTzB/0Ooyj041Zicz6VVMhJEjGY8/zfpUVFYclhD8d4dBboDWT8dzI9G437MF+LR4HTPQq2JsZnIzuPXCNcz8DBxHLifkb0sGhVUg9RSnF7TlvogXtByPBCQ8jaUoRpmEc3Tiz3WyO2ILMowYVtan1xxHLifkb0sGhVUg9RSnF7S1Ut3ldwINVZdGSQLKNBu4HWGa0srxhnopfoWQz0YWbgGAmYLC0O7mbUXfYiX6zhTzqsUZ4hmxNk3DgPAP7CPmqC9rh3i48KzcFWd01q9Ao/WCKtFaAB0pbUXfYiX6zhTbA8chY5Tt3EaE9bo5+duwjEw96mKSyO+IhdTrbbAMB1RWHJYQ/HeHQW6A1k/HcyOqtTZBK/sz1g1kl9fhw5akbcuKYkbpcAjsY21T3uRMTZxqJIHSnBRTc23KWnbOQ/RI5fkpKwBOviBV85vnPyBcdEL0FCtBInjC4OEyxUpTD+dK/+s2YPEJaU5KmyApi7cgVfOb5z8gXHRC9BQrQSJ4wuDhMsVKUw/nSv/rNmDxCVi8lA5QkSZMJ3lAqaRgjfgKCNTTQuUYDKE4NuFfY136Yp1Xv05AzbvISx9BdF4ZgkyfiZMSzGFCtsFlF0j88uWRlfxxXErOXsjbiI4yTVEYagcVatrFbUbCk7ek4/FXWeuUfkMltpiAEOfZEhOIKBPnSv/rNmDxCVkYJYmxNmQwbnULhfEu5Ev8rfc8UUu5qHDV9V6q7XQ5FIjp1DOt+yc5Cyde4BY3XAEbMptBX037NgmrLZ+Lschw1fVequ10ORSI6dQzrfsnOQsnXuAWN1wBGzKbQV9N+ybMsk72AexicNX1XqrtdDkUiOnUM637J5znrovwNLCaSrNyZ2O9qeDlGiMDSAu4AuxjbVPe5ExNnGokgdKcFFMXyaEm53u+WP1220h+rjcJqpAPer6kaNEcRy4n5G9LBoVVIPUUpxe0xvZrfAFJ45wUkLvcsBBlJ7BiobIKCIscGa825ZkoTmccRy4n5G9LBoVVIPUUpxe0BDlZGqZPqnYgeQFngs3DW7QcfHZn8xcY9Dyfl9n8vc84HXb23V+jBW1F32Il+s4UXv9yBR+/ijAQHdSJbvZcddQ6blVvwKnwuDMwYXLoEPg+7fMKTrRNy1RWHJYQ/HeHQW6A1k/HcyM9XwCyK0iTNLK3DzyiG45zxMUzSIq7Wq4oco184hoJLMLg4TLFSlMP50r/6zZg8Qk+qL7jVkNn8sdgzGu7iuuee7Xdkc5z3yRZvmYggtqVAuHDJoDEt9A9FIjp1DOt+yfdv7czRvnKL6+7HokwiEStFLE6gy+KXP1YggAh2zYxKvJMoiRRwIwdaUCqUsoSsGkaXpoZ3OyQfjVmJzPpVUyEKCcjwbuij8hUVhyWEPx3h0FugNZPx3MjDB2TZHWspj2joXGnl07ulSmKbl2BmuF0a9CKQlY8TsIr5MLZhS3k9v2s1D2kyMWn0iOPfk+CJxqqkA96vqRo0RxHLifkb0sGyPNUxvZZ6uD5WqwcrJXfVKG3vUvHTcFVMMM87GZruLMOgH3CGeeYPtkM1JKfl+0h+FotoRIKEsjtsEHD+pcpuq+jZ7tkca7jagcVatrFbUYxw/B9q50PNFl5PkURucEw3wAJDf3xiMz4j5eTImYULtkM1JKfl+0h+FotoRIKEsjtsEHD+pcpuuC2sOEpIU8dAad5VnW3MWpXv0ka7WnuTeNGSamGp+r6JnWyFGYcxASC0NOGP9KsiLOLgppTO0SoAsL4eW2jSDZKnpQbBzpqXPmLz9on08CpW4lF02g4zIev1LqOVaAsXLsJMx24riqme3e9qzTxDx7NqyLGdo9RMhhDbO2fqMew0GaT9Geh3N1y6SUn/IOb9WPC5sDZ9s7TJgGuAYBghdiZTpXb/7goNd9jcx7OO4uWxV/6M5p/R7ATFaj6L4K6cPicEoCsjB16ZdsjXDviZ5zzIKTcp0JivuO5E563YAuSux1xW2FKV9CCoUVSF6OrzZMVKl0z/1hUWxlmFzUcFasOPiXyJSi3c6zM7/X368bkCrwi/h0gOmiBPozgbBitCvGpW9+dwQiu+BX1TLYqBQbSFZL72nRIABYPBSNu8LHp5DHa5eRNiiRlur3T//WRN977PGJXF7krafAXapYNs5udCClQjtkLmgOmQJqWoxifr0B8l9ohbmSXRkkCyjQbuK+f1bMKiqFfeE/r2e+TbD0mdbIUZhzEBILQ04Y/0qyIs4uCmlM7RKgCwvh5baNINkqelBsHOmpc+YvP2ifTwKlcqxMAN4a1VWpk6jHdQaYkMHL8fOHTBcPFX/ozmn9HsBMVqPovgrpw+JwSgKyMHXpl2yNcO+JnnPMgpNynQmK+47kTnrdgC5K7HXFbYUpX0IKhRVIXo6vNuVB4J76HlwRbGWYXNRwVqw4+JfIlKLdzrMzv9ffrxuQKvCL+HSA6aIE+jOBsGK0K8alb353BCK74FfVMtioFBtIVkvvadEgA1AcTYxitBR7kMdrl5E2KJGW6vdP/9ZE33vs8YlcXuStp8Bdqlg2zm50IKVCO2QuaA6ZAmpajGJ+vQHyX2iFuZJdGSQLKNBu4HX4WogV+u1wjTD0h9C086iZ1shRmHMQEgtDThj/SrIi6cWmkkLq3LJwJ6kWNLc6Zl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGaM5YIlEkpSTxuCk22UP74wAjpnoJBn29A0AJGzHDO6CCPL/CaaqnEGOrTlqFJ0CO0A50aFcFGB3i/RAXejHHxz1ZfFjEE8emLKP0xWJFtBKIBKVz0d0HCjIqcpI2SOkFIXGE9AgV6ngq3vAPCmghKL8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEf/oLRBc1dmeZHrf8s6sqBUNoxbI4me9pimZFIuqsPI4YDrXOrkvJEoAM0VMcNdjM/m/fPgGiWhA7BvkETgs+XWGnkhHOWLndeYUieJ1YegZdiuoTHUj00cN+plWTQJSyyhjQtlQP58ojSc3R/HQ5ndZL+814w1rJYvxMuc4I56TjfqZVk0CUssBA7GkL0TsmRAhoDL61JMcTfs2T3tv7quYVxXqkpAiBjJOUy7k7ErcTSc3R/HQ5ndZL+814w1rJYvxMuc4I56TjfqZVk0CUss2HZV5cBN5+5AhoDL61JMcTfs2T3tv7quYVxXqkpAiBjLfoZr3JwgyDSc3R/HQ5ndZL+814w1rJYvxMuc4I56TjfqZVk0CUssxCiRyLxH8wU0OvP90zT1HixfGI9/oyonbPz/c6/JJ/0zJ/bYDVRTMKEqUIAbdLESC/aD28SwXa+T8VrTMwIBqDSc3R/HQ5ndOSHV1ZqHYJlRCWbeSOoaDbQLbwE2vp5paLqzJmflsPSXt14nAyWWX0NaRZr5dtq7lcwbKRQEQlmWnABkhfYwG9iuoTHUj00cWmZy3pVbVk5Xm1D9kTN8cOI3sv05ME8NsG+QROCz5dbDHzwZbJ7YC0JgWLIeqDPpcQr3mv20Raz/VThBD5Uhzyfiu21TSzSoTVP9cq4atqRAhoDL61JMcTfs2T3tv7qul+VJtD/uv6D+BYdEK+bzapKga1YesxCgKIDDWJwVSi2j1LPZE6uc4iiAw1icFUotRh1/dUe3fOODKkvY++ZbwdP1wyS/3aSrnwDziWeYZMzX8AjISKtMcDhszRjqw8t8fSMyXoLumZf8DWxmzGd+ycxBPmd3IyJnOyxQZ13Y28eB8SJ0Eoctp8uT6SxIGKL0GGu+3/L5gB3AlCJBb+ant+KQsqKX7jOl3Hby68hWu5GoNfGWRcbK39boZH+dJQSklVceTXqIAKhKohXig4QGZJDRDzKAm9d6N+plWTQJSyyS/XOe+7bfPD8BqKRjeRUOb+qlMDhdrCQxnN5zg1hvplFnSrFpTE5RFQRTQg1Qz1Dh/ynDAobVPQwrjVQlO79KwJQiQW/mp7e5roVMTJe1k/w8/5AeSbpDKIDDWJwVSi2e3uIFbhG4EiZeXR2jc9w3TbB3mVsru2mSZCCuzeFXVKg18ZZFxsrf1uhkf50lBKRJ6shrRPWUp8smgqJhmepjGGu+3/L5gB3AlCJBb+antx0/XhGDCcxKiQ4zdnNltTPAWCwd+65pMKvV8ZIoYFr4s/IT2ZPQHhlTu72xtSK0P/9VOEEPlSHPy36Ga9ycIMg0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4Q9BMUbPYIW3cMKmb+s8su1uhkf50lBKRSQiTI9fxSysCUIkFv5qe3jMLLxsQny9yIrH0FI6EKS1oXwe405BMXo/WuDZEL1ulv8q8EUehCOo8x4eQWWX4LkqBrVh6zEKAogMNYnBVKLb1tbidPYvITYGxxPxltFAH5Rba6jvPVT3Fw+X4Dn1Z+PuO2z0P1V/oWu86DM8FPLkGK0kCQb+z+JuArOjbYDxHAlCJBb+ant6icXrE9H7kEvasFSgZCszC+cTnAo1owFGIKO/++klhwU6SbMn64d6oSPrFIJZWI1eRIIq03qPkD8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLc+FSKon89memdnV7G92gbdhN1BvCANmMngDx2Hx3qICy5VaKJckYTL0fVH7sA4C9ZgbHE/GW0UAd/b2c6WFk1dh20VhKqnFtwEA5MlnbvkHmBscT8ZbRQB+UW2uo7z1U9+3/Xmuars+cMb/Nwqih1HV8dTK5J0h5Ca/sbTdmm9xeyLyQODB5SpKIDDWJwVSi3wqOHo8r3gqqP8Svci7BVicdmIiNk4jAg6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZ1G10OVJSLFZP1wwePcB3niMYZaUaRmBG6lgWozxo8h6DVq0jCvH3W/zRiUhLgJ8PcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJO68WUMt5UCDDRKfJhTPauSx5P0MnjyBFn8UnERL5ba7I/2fb0QO6SXk7EXRx5S7np1p3ZkMs6b8QGB0jqzgJ02CeYwq0F7hzdr0IpCVjxOwtfzyeLG5RUgyTR+UIzCD2j3gRvClmu+NJCsWg2rHz6bYv0GcUwNsoIpCbjHIfzrNblg5fuBTrJoHTyFicbK0d5njDF5GcwuOMHKH+bXLzARqDXxlkXGyt/9A8k5xBohHRHWeH/CBn1BQcN+BBMMcz5oSaLpq3FPRw6dggFDDYz4I/6fI0QRgF0cw7FaFR6fNepCD8amLUG6skijOumT+0e+rgCQwqT6QcRKML+TgQz/EdZ4f8IGfUFuLI0QnMD9a9+4z/c88WUgdlB2sBpybScR1nh/wgZ9QcQwhr2xk7+pp34gAL0xItQdD/YDI7meaLT9o6IPjbYyVEbpeCnAPqBm1/WBNgQD829veL2IvA+sNPXKOfESRK9AZHhW/oOWGL2rBUoGQrMwvnE5wKNaMBRiCjv/vpJYcMx5gbgG8/5v85bItEi16fH/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk1vBvlGgaYRlsoRPQUor1JZBJweTZ0cU5WsWIuqa+R+hF1+w0J386bKG55N6vU5ojiuLI+nVqGOGCXjktoi0g9UvvTazxYAV5sEtpKdRPXl+OdpHvlipyiBbYQAZh5KRfAZae2YfjgYJHpar/ooZ0cFaCEihUNo2NYu9JBHxykHNBvtdZhlL105vPvscxb89PM0PCSRKK0oE/vEgZ9zWfrAL9oPbxLBdr+9z9Qe5ieDYyKgx14rCZ5SICFg/Ipz16Yj9DcF+tcmG0bjfswX4tHh9v6KkB5/9VSEnoAX9sqSSKiNB//SHf3DISx9BdF4ZgvOULQg9Hit+JHxc1axEYHhG29kNKBrGeCtgapqcTDSgiC8dQRZ042ENP6X/OH3jggwNv8MNhF9K9X0PJ0frpVuirr9WB3KhzBWw217nLmPwC/1YwoX2QN+5gBP98rq7vlDodqjtdsyQkkgl9/s3LB3Y0xOswq87CmhznxziNiCCcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JuYCF8aFffEfRPASFTGAlbH4Dhr1DSA590ChIjub3THD6637rD1jOjny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTYcqqiDGcCkSJl5pP+/w5LVg8M/XPHF9qDN8hwkaeXL9enkzBWt0tJsh7ZqYKCFRvWatJv63NJHSu/f2jwP5f1/CCD8Qa/jQUNYQCJW9sVwywuDhMsVKUw/Bnl9/f6xjf8mAMeTsncOjENjLjRk4j58UsTqDL4pc/ViCACHbNjEq1qk6FYBnBqZs/P9zr8kn/aI9EAkCE4Ye5v3z4BoloQOwb5BE4LPl1hp5IRzli53XmFInidWHoGXYrqEx1I9NHBsfNk4cB8P1cEPVzZMfsJ/5RqxiEiLZGS2YloElx8fqGx82ThwHw/Wi0aAHXIcx7rtwcZyZxxotq7z0WNseUXcT1zWClEYtH44v3PQhoFfM67Cu6nIIXDbISx9BdF4ZgkyfiZMSzGFC2izoChY4j6wtmJaBJcfH6vrTvVmiP9TtVn1MEatdnPRpKqP/7DJnXRrA/senfGGrkNEPMoCb13omAa4BgGCF2KkVUA1kSq0cNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpODlBUv8G7AEshJ6AF/bKkkra8k+qJCjnsi7TFwBn6cwSoNfGWRcbK31yrEwA3hrVVqRVQDWRKrRw0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek61/rmJlpZgcFEKeiZfADjpkaUa6iPBqaR7IbirU4mKIqg18ZZFxsrfR9qdNNHkoE8m2Fqa/z6XjPnnmviumZaqjS9hLV+VlHU+DGFHP0RzNfpsDMN77LRP4RrstP++zBxs/P9zr8kn/SVfbovfMR6DCZrVxtmjyhknaHfzp3fCq/rTvVmiP9TtgqFFUhejq83jp1JVxneag1EJZt5I6hoNu3BxnJnHGi2rvPRY2x5RdxPXNYKURi0fapF1Hash/k/rr3MUWOscilyrEwA3hrVVidfGYWFPTNr2qgcg2eo1NMOTyNLgcNdkQIaAy+tSTHHkQK/WNyYU+xpjN+NMLr6RHJ7TLaX4iiJWOlUA/aj4U7B5JIIdSKgVJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfRBBK7TczA+v2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTIA9ep8vX5pO4VEcGIIZz8GNJzdH8dDmd05IdXVmodgmVEJZt5I6hoNtAtvATa+nmkQQ5ha4ATz+BAd1Ilu9lx1R6FaXHcMmawlX26L3zEeg4h4BdF8CI0lZL+814w1rJaskPxLL+8gfTuNdKNAyhOXDB2TZHWspj1Zu0xVYcwPZ2z8/3OvySf9JV9ui98xHoMJmtXG2aPKGZDRDzKAm9d6Pqi+41ZDZ/KmxXgTmYlxnDQ68/3TNPUeLF8Yj3+jKids/P9zr8kn/TMn9tgNVFMwA1LqqOs1kQsgeQFngs3DWycN6Hd9SZc6QIaAy+tSTHHkQK/WNyYU+xpjN+NMLr6R6NLvPlfAjkYiEFgcKS80jEehWlx3DJmsJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfDB2TZHWspj1Zu0xVYcwPZ2z8/3OvySf9oj0QCQIThh6SoGtWHrMQoKbFeBOZiXGcNDrz/dM09R4aYzfjTC6+kbOm4GNjZXJtYK3CE4cXXxcnDeh3fUmXOkCGgMvrUkxxN+zZPe2/uq5ourMmZ+Ww9Je3XicDJZZfQ1pFmvl22ruVzBspFARCWZacAGSF9jAby4bWViPLkGuRjGUlDW9J9Pux3ePJYNj+ahWL3eRIq6HN7kXKRx1ZJvIBDOmKt3Sa2SwJDK/Ezt25roVMTJe1k6HtPoHk3bTbTbB3mVsru2n0M4AtCcGdF1DodqjtdsyQVpIewvJE6DHYGRDsmjbJQrJ0xnZnSIbqs8TuxAbbvihbdWFcQQ+Y4vIBDOmKt3SacQr3mv20Ray1jYKECFFWPxE29TrP5Ai/hVppLxC4y0Pg5w7xuhod93V0+5KmdlH7IDciwWCFEt2z2Pcjytgf41ipdOwNObxmWRglibE2ZDAuQq6EWvihkCNLZvLRkPSKCjztA2FYcnzSUoEq+NKnzvXuu1KtRcY0JyAl8xhXqWH1girRWgAdKWApAKJ1myMA0bjfswX4tHi3pdqkk+LLARD0ExRs9ghbau/FRvAupn9E3tygC005pGQSZgj4ECnQ4gqPO/TyKVTjqS2b4yIpdmoHFWraxW1GwpO3pOPxV1n3+H7Lk5EA4IjkPMAqjtJnVHbwYEeTdWIHAZRyjFo+uZXOMNATyXaIthjdCeLkmn7Gw1V3wxTLxnydKb4opoMSwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwQ3D2Q5Kbjw65roVMTJe1kzBgmJULdk6vUOh2qO12zJBVAGpeCbzmnNgZEOyaNslCnt7iBW4RuBIctas+oPi1vMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMAcBlHKMWj65+a8qWT/jqVi2GN0J4uSafuvGVOcTC19Qoe0+geTdtNtNsHeZWyu7aTMfZpkiXy45wFgsHfuuaTDAWCwd+65pMMBYLB37rmkwo94iATDrtkNQ6Hao7XbMkPXDSXil0gFk2BkQ7Jo2yUJPkdZLtgU8sMYDsdHTlX9WWUsZoZ0EBfiQ0Q8ygJvXeiYBrgGAYIXYs9tcqI5Q8mbnzOUaGTzpYwcBlHKMWj65FSIo19rZmLm2GN0J4uSafsbDVXfDFMvGm9oCwLODrdFNsHeZWyu7aWq4zPXPdCQ+iOQ8wCqO0mc/2UGn8SCKHsxBPmd3IyJnJgGuAYBghdiz21yojlDyZvkSZlKfupvguWDl+4FOsmhQJ31G5nUyPSEnoAX9sqSSiBmxUPf3zDokfFzVrERgeMZyfDAmTwNRFpziG0dVJuelDy8rLqxLOSEnoAX9sqSSYil8lt31eSxxCvea/bRFrM5UIZCbh9wpagcVatrFbUZhfFi2FgFwyli8lA5QkSZMNNL4R/na59+X5Um0P+6/oP4Fh0Qr5vNq67Cu6nIIXDbISx9BdF4ZglpQUak6jQ9fagcVatrFbUZV5hgbj+TkEXE245fgOSRjajkcM0HTJMVxB4J8Y8cmvJGMZSUNb0n0Ncvy1Fl7TZbiCo879PIpVDye2Fuyx1SgAad5VnW3MWqIzbG+JEb+ngX0lQJfZh8bUi+UbV4XaYtfGtVDrj+9MJDRDzKAm9d6CgXjU6hDwfzISx9BdF4ZgshF4aS5pXsa4SSlnUTC2QjAAWqc0RjsA5dGSQLKNBu4YXxYthYBcMq7cHGcmccaLbdTi1x3mcIYkNEPMoCb13q9t3/R4rnksue7kTKg4X1cAad5VnW3MWoN4iZMez+iF1u/wjhN+ETgCZ2gL/8pNVMF2JeqqJQbC5DRDzKAm9d6YWaM3bdub3CTm0c0jNHELDjYx7mq6+rS8WxXpySov1u8IIV9Dbqn0rX+uYmWlmBwUQp6Jl8AOOmRpRrqI8GppAcBlHKMWj65FzZU3zYUKXTGA7HR05V/VtznV8bba/bZthjdCeLkmn7QLoCzXvdvsCJ3mG8Pb9NnTbB3mVsru2lhhxFAxerl21FtoQJBI4QNE6VZWAUpdcEWQjte9/SsM5HC6CQ1hda/8E5ZjCzjPn22GN0J4uSafte0EO3Z8OWas2VRFtFcBYm5roVMTJe1k3ydKb4opoMSwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwZM+IqpfDYgaYtRaReIvRPrNlURbRXAWJua6FTEyXtZOHHhUgnWFaY1DodqjtdsyQXFsyrNUaL64Ya77f8vmAHcBYLB37rmkwwFgsHfuuaTB9C2hGWrbjH02wd5lbK7tpH1+7mNunDj2I5DzAKo7SZ4tvNQPRihP9BwGUcoxaPrn4uNI7dF/dfnAFyDnvuOjewFgsHfuuaTDAWCwd+65pMMBYLB37rmkw2BkQ7Jo2yUKk6WJ4Srd4PsYDsdHTlX9Wz20RHOVQvoSzZVEW0VwFibmuhUxMl7WThqeiEGoiTAo525a2KTMEeCR8XNWsRGB4NXjoaTKOL7FxCvea/bRFrJG7d8H0C1ozTcOA8A/sI+aOC6phmVYupWGfMq1BU3YigqFFUhejq81JjZl9O8q//MBYLB37rmkwR9qdNNHkoE8nkMrSZARhKg/vQP6chh4CCZ2gL/8pNVOjYRNNtsT2oRhrvt/y+YAdWV9bOkU/UIjE6Qvm6OsJaiDtoVjunTXW0hWS+9p0SAAbcsQkHtqFjqg18ZZFxsrfv5E/GH60cQkkfFzVrERgeN21ww6EJiGccQr3mv20RayRu3fB9AtaM03DgPAP7CPmjguqYZlWLqWk8IB+IcARtwfyNHlccJhXs6bgY2Nlcm1RbaECQSOEDROlWVgFKXXBMFB2sJ3m6F1Nw4DwD+wj5jE120KBt0SxGGu+3/L5gB1ZX1s6RT9QiMTpC+bo6wlqGckRWJXZYkETpVlYBSl1wSDN5ixMJnQvvasFSgZCszAqD/TbGbMx358A84lnmGTM5gIXxoV98R9E8BIVMYCVsfgOGvUNIDn3QKEiO5vdMcOcttEH0AG40x08hYnGytHeZ4wxeRnMLjjByh/m1y8wEag18ZZFxsrf5u5P14gcytUoxhHq1tfLkMBYLB37rmkw5fYb0A4LGJtL/DLYQ9qk3MBYLB37rmkwW4lF02g4zIckwt6Ome36qEe8k73t3zA7ZVn8Et1InyuTZN9cXlWRmyQ8jaUoRpmEQM8Ef6sjjjTAWCwd+65pMA5QVL/BuwBLCZ2gL/8pNVNVQVOzjNIQMIXS8Z9Ju6GQqOmaUV49yKlZGCWJsTZkMC5CroRa+KGQYgii5knpzSwYa77f8vmAHXg7KXxLmSbKBz08USkNXKjAWCwd+65pMP9VpLFqeRx2LkKuhFr4oZDzEyOvnDD8kzT1yjnxEkSvmceagzYIXt1biUXTaDjMh1e/SRrtae5NFCz+c/tzQDjAWCwd+65pMA5QVL/BuwBLCZ2gL/8pNVNVQVOzjNIQMIXS8Z9Ju6GQqOmaUV49yKlZGCWJsTZkMG51C4XxLuRLkNEPMoCb13qkBz+FUA62mJcRaHwDcIfmaFTnpZKiSGfAWCwd+65pMCYBrgGAYIXYEnOHrkDuI7cEMg3yvjt2+YehLgG8dZzZNBR9H7I9lXdqBxVq2sVtRjHD8H2rnQ80sFAZo7HDX7GoNfGWRcbK38ABapzRGOwDl0ZJAso0G7jg2j4oeMuRzBHWeH/CBn1B2TQ2S3XJ9s/53/e3dBzVMtIVkvvadEgAVrk0Qt7WJ7lQ2w/oA1nAlMBYLB37rmkwlhOdkPAYuVcnaHfzp3fCq+uwrupyCFw20hWS+9p0SABOfUTJvCYpZ8nMmVMIGdEl0hWS+9p0SABOfUTJvCYpZ825+94HaEtyQ3rlTdTGOiEAVplKQwPKfdIVkvvadEgAvQh6UiXQPX+bnVrEUTBOFee7kTKg4X1cAad5VnW3MWpd7KO/+4hdexHWeH/CBn1BXKsTADeGtVWJ18ZhYU9M2iCWkfLZMXLvHEcuJ+RvSwZoFT/zJseJVKOmtToMafvyLkKuhFr4oZCFZ6ABgRBrdqg18ZZFxsrf8xB7sp62pU0VfCSULxcpWZGMZSUNb0n02YoZ4D17th7pVZV7cMebZ0lG5W2yqFa+Pq2HT+b5sQjg10zOP2Nj7NIVkvvadEgAvxTasE+toySV3x7u7HaI2QbdIk8JrCDe+oFv95X11+eRjGUlDW9J9CDRaLYPhCEr8YvKH0AvA/DubG8dxB6p2Vf+b5SEvOjF6hWD4T5dDCq6of3JjiVuSTran0avgLLfCNLWMLgXR5tQpqjtfsGDVoSUE8Ofu8VlsXKfUFlRz6eIlIbyK5hxp7dioAahW9MfagcVatrFbUbbUyiUTJmgn6jpynD0BchcgqFFUhejq81HEWLf/jjL+KOEbht4BwRypRdgl2+7HtwuQq6EWvihkIsJMzummSZgpzJyI4BKxS4Sc4euQO4jt6iYQd/hHEwRJbejIBEUWm4Bp3lWdbcxaiTC3o6Z7fqoIO2hWO6dNdbSFZL72nRIALNHLBVwULm1669zFFjrHIrCQY6EvQFssNIVkvvadEgAqLLN5A3M+uuVRGnMsTVoKtIVkvvadEgAs0csFXBQubWoNfGWRcbK3wXjvEQzGu2eCzfg903UEFq0//yLJZNFE6EbftywaO5uuZRtBme/SF/5V4iVOtMz7moHFWraxW1GVeYYG4/k5BFOSnlK3EwW++OpLZvjIil2q43t51BTNhhscGRP3anPN6a07NRbnjx0T9gx727NHxdAvDiKK56g4u0hvUBC+7PROW2o4CjsVujfBTCEmXgOSlGpvdtHMHKY7BC1zngkMKvLbMWGDxvDKNlQ6Iq7SaR2YIQmwql9MYmSHPgP+RzESyiAw1icFUotcYe+2HVB3n5J75lJu2/Cd41VxarjbYSyGGu+3/L5gB3e2+IB6jW2q8i6d7xnQLFrRBBK7TczA+tHrKWdpHDYSs4Rk+39YEMdzkyQmBmQ0joOgngeRpQU+6P1rg2RC9bps6bgY2Nlcm1qORwzQdMkxQKB52gK4D7dPoTs5dyOyxkxHcxmNOM+mO+wSIJbTAkQNJ2PaF6xlXHMQT5ndyMiZ8CUIkFv5qe3oO8p6vsn42Ep+4baVXgBLLGcsr0LskPbGGu+3/L5gB0+qL7jVkNn8r7tMMLS4kWrdfYEVXFgVcEKpPFl5icPe1iCACHbNjEqs6bgY2Nlcm07jXSjQMoTlwwdk2R1rKY9aKBTwUEcC/EkXFK/f52xBoiF1OttsAwHNHpy8+pZSlu8Q1K0g7GUghAd1Ilu9lx1QyyEUB36RzTZW9Tc6xei2092CaJGiDpYLjX2HVkz/xWQ0Q8ygJvXeoSfi+ElliHmZ6laVXeHlsszqzFeKqpMDz6L6dlTtuNwKL4bTgl9GUBNkdqcAwI8uhac4htHVSbnJleF7SWM2DU+47bPQ/VX+mI89vHdwFrMD3Vtl8iFR/y/J8/NB0ZItnEK95r9tEWsvENStIOxlIIQHdSJbvZcdUehWlx3DJmsn9dIJIMsjuw+qL7jVkNn8qx7b49u2rsEEB3UiW72XHV/KZ321NwC0G0ikQ/KmINPe3hqEB2OSd8DUuqo6zWRCyB5AWeCzcNbZjDOqQme523/G/tIH8aRKD1fALIrSJM0NdTIXDtlGaQgeQFngs3DW434BwZtN4oZHEcuJ+RvSwYnI4HlVbgl28J+MHSONXBWtlnOaLA8gPOUbgpAAq5yjF17GQn6snScEB3UiW72XHV19KWHLXaiV7ZZzmiwPIDzdG2W8z39Rvuj9a4NkQvW6bOm4GNjZXJtO410o0DKE5cMHZNkdaymPY0em2vJ8o/+4B/DQZhqEIEgeQFngs3DW67QmtLrVR5JDB2TZHWspj0rlyMl5V3mKbcGtZTTW0lmkNEPMoCb13phZozdt25vcOPlFyDCCNCFPhUiqJ/PZnp8kLRuoH4gSQAJmulweyOMayibrln9UraLe6F/GrC8TMRsDYxocx/qJ+K7bVNLNKiLNBPoJTQF2YIV+C9cfNIRt6zmj22E+gCoNfGWRcbK32CtwhOHF18XRAhxwjblPwUQHdSJbvZcdXaCaeVk2AM+qDXxlkXGyt9grcIThxdfFyLRsOqBA9RREB3UiW72XHVYNEObgle7Zqg18ZZFxsrfYK3CE4cXXxdy/hXdBH8CexAd1Ilu9lx1coeG05lg7M2oNfGWRcbK32CtwhOHF18Xcaz1hl0RxK8QHdSJbvZcdfMpj/Dwd3MNqDXxlkXGyt+tMg/TH8AwMIM+aEC2mLhmax7M6tZYeK72iuplgCAem2HAMBrFOGQZYVTZrspcECWXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiaX8QM59V+jqhZrN/Jo2nVInAp77gCTU27NqyLGdo9RMmyVA5YWJtbGngPNrBqQHVbMlzDoYcoiT05PUQF8eqGh4Y14cu4wOOVWRbMn7tAZ/L8fHec4SQHeeWcZErNX4Fh97Q4YLVT3ubnhN/xhR9S4zasixnaPUTL79lR5CFqdQlQBmbODaIcJsoBAc8MkwMuR80rvFnXDir6a0G37caWPl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGagP8Mxne+ejF9h9IOivGxLzasixnaPUTI0ijJYlkY2uZObnKdFJVypBRcpoz+aVLk98F6mH17CrVAnfUbmdTI9CZ2gL/8pNVO23mvmx4x7LdyyQa5HMXQuJrZpNlGJw2gavUEGp5IL3M9nhlXRUrw720UfxrAW9Z5oMcDzmvmwmbMJCajeGgtgqY3O8XQNLMWLGTIcb5Bh2/uzNxSojBuR/4NLKfJ++hCnMnIjgErFLrURSqqm1aeVSnsbRkVzEj3a1Zni5uVvKw6OyG6bnoLJwFgsHfuuaTBYt+40/kUJWGf52OwzgI9tGGu+3/L5gB0fILcYi00x4h991K5Rjd5QAgRr7UzjYUyoNfGWRcbK3xLUX4/SMqrVVFrs+/25jsn9txXXiKUJWnAlDQ+W9YT+j6LoT4+u5D9mPJKZ4to+yu4ZC1Q/KF70Iy2e3vjX/4qCoUVSF6OrzVrySpKm7TpZYZG2YvHFvHUCgedoCuA+3VkYJYmxNmQwGdMoen5652Yj9fl/m5CT7I5wsN366cbVyo9VqbL6rO7rEML7AL6j2XPpFBtQkSMfqcJVNzczxRKoNfGWRcbK35R0IgKgw3cUOE4R8f5vSSCoNfGWRcbK31M88Tq3odGE+fl4Jzeg7noBp3lWdbcxata2GmZNWhGjgQMstZ/zZTAOoV5ciNV9Q4/ive0PzKRfYu5mMV9FnqTjo7C3kNP3INLkH4dC4si1wFgsHfuuaTCXIk1JlZdjcpMRkOQ5VOTcOtykQczYjX8Ya77f8vmAHWxHoMmoJRXK7czDPliizRMQT+fCOtZ7+XAlDQ+W9YT+j6LoT4+u5D9mPJKZ4to+yu4ZC1Q/KF70GDeCzxBtH1MJnaAv/yk1U+NUPNETNEP5yk7d03eqHkVmZVD+LBdvKzXR6dfO/9nfk5vDWDoY7XBYWMPbfMv5yJu/jTnzePw8LEs7wHa9mjny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPFpbEnY3Ckt32nQKBOgs+dwIu5oG++L0eGqUxWEUwxjMeT9DJ48gRZ/FJxES+W2uyJSqCvee3WvmRXZEp4UN23eQ8qM0FyDJNmzfnCvpTk9bhdDjKl/Ez7cEVQvmZs4ZhxCvea/bRFrOuwrupyCFw20hWS+9p0SADBcR9+1LSQ7MnMmVMIGdEl0hWS+9p0SAD8IR2ex6yAU1gWIvmbRDqwqDXxlkXGyt9biUXTaDjMh1e/SRrtae5Nt/JhIlQPb+BbiUXTaDjMh7wgl5kPCv8Skh4zjHe3HYcnI4HlVbgl2/rTvVmiP9TtgqFFUhejq81CGB8z29RQVqjpynD0BchcgqFFUhejq81a8kqSpu06WeNnDqELVCwE+QXlou2+5t79txXXiKUJWhMkTNpZjbuTOX7gg9Mlkun9txXXiKUJWl+SeOtU1HJ0tHNobvDzG2WQ0Q8ygJvXeiYBrgGAYIXYBaUg66Mg/LGC2Gsng0c8ZSYBrgGAYIXYzX6feb30SdAITcG8nDE5TKWoNek0fwRjUCd9RuZ1Mj0JnaAv/yk1U6NHqLfhDGbjOORmivZIvPYJnaAv/yk1U+NUPNETNEP5Z4VAcGrTdH/jqS2b4yIpdmoHFWraxW1GMcPwfaudDzRExd3+dX/+32oHFWraxW1GA8bLz49YRl2LBSy5zaaQcrOm4GNjZXJt/1WksWp5HHYuQq6EWvihkMxvZgSwlS+tW4lF02g4zIe8IJeZDwr/EpIeM4x3tx2HMosEwBjbwnL6071Zoj/U7YKhRVIXo6vNi9sCWg8jpBgmAa4BgGCF2JlOldv/uCg10BSf6LEKTR1QJ31G5nUyPQmdoC//KTVTSvrZVi0OvD045GaK9ki89gmdoC//KTVTF1kX6jGtvMmmYURHNrLDk1kYJYmxNmQwLkKuhFr4oZD18i9cPMJ5FlyrEwA3hrVVzX6feb30SdAITcG8nDE5TL/gSNtnTmQLnYUCvTflwMzSFZL72nRIABYPBSNu8LHpD+9A/pyGHgIJnaAv/yk1UxT7W5VwEmYKPJ7YW7LHVKABp3lWdbcxao5hk/vQXwNF17QBeNIO09KXRkkCyjQbuK+f1bMKiqFf6XfEodxWpsZM1ULwbvP0d4KhRVIXo6vNgfD9L+YU4qBZGCWJsTZkMC5CroRa+KGQB4UD3bL7YX1jVzfHpaQnsxBP58I61nv5bbelGUC2qG8g7aFY7p011tIVkvvadEgAStsjSkndLbeoNfGWRcbK31yrEwA3hrVVamTqMd1BpiQtMrwywRkQfwGneVZ1tzFqjmGT+9BfA0Xs5Of95XYZ6g5QVL/BuwBLCZ2gL/8pNVNybppH6fKCimGfMq1BU3YigqFFUhejq81GUA84gdgyi8ABapzRGOwDl0ZJAso0G7gxw/B9q50PNPycPm+8FtLEAad5VnW3MWqOYZP70F8DRXmPQy2X4xSaDlBUv8G7AEsJnaAv/yk1U03q4kFKw/ZGIO2hWO6dNdbSFZL72nRIAPwhHZ7HrIBTZ7/voeDHk6aoNfGWRcbK31yrEwA3hrVVBaUg66Mg/LEvlOXLT3XBjlkYJYmxNmQwLkKuhFr4oZAsfVugM3nBzjL6aoGu7kGFY1c3x6WkJ7MQT+fCOtZ7+RMkTNpZjbuTptJgn108PNCXRkkCyjQbuAPGy8+PWEZd8GuSrbY01duzpuBjY2VybUzVQvBu8/R3gqFFUhejq80YshrI/jVrEw/vQP6chh4CCZ2gL/8pNVPjVDzREzRD+UE4EKHoguOUPJ7YW7LHVKABp3lWdbcxale/SRrtae5N6dXmG8ydO0VcqxMAN4a1Vc1+n3m99EnQCE3BvJwxOUwYRttBf5DujJ2FAr035cDM0hWS+9p0SADxL+uhYI7D2qYwfd9h+fUkEE/nwjrWe/lfknjrVNRydAn9h1u6+vPekNEPMoCb13pZGCWJsTZkMC5CroRa+KGQypoJBfQzqklhnzKtQVN2IoKhRVIXo6vNWvJKkqbtOllvyxVBL++h+b2rBUoGQrMwvnE5wKNaMBRiCjv/vpJYcGbjNZJwnSwMZtgSPO+3yWOh9frKj2o4oxhpNQC36zt1jfuoxOiR3gtHoVpcdwyZrAwdk2R1rKY9Bslab2P8omcMHZNkdaymPR0/XhGDCcxKeppZo8RsuOzTmYJPsMg+Q6bFeBOZiXGcJsavxjE8f2u0vHvd+5v00/4ndrcguBFspnhPA16MAjVnqVpVd4eWy6xxATWFVpDn8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/FISXPcEbu9lxnTMmIRq4lhdQ4ka7YhB8iH+mGfOlMxOWc0r+BO1+aIrQI1vzPx3B/HDAE/DccCDbOaS9bg3aDIhuS0i7MtH1UYzxOZ2iMHaQTYtOoT7nIVf2CcPL9BVMWsdvkInikv0HAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAW4EXs3c+9NcIJECOL9wK2g3G/JDxBbWRbG2/Dx6otjNsLDGQTJXEeQ1Hx8fLTKS72wkBs9x5ieHk/3YY5Db0vBv2EwAFWgcOzbOt5VoinonpitYp+OhFaSwCs1OSwqFagvm4o0bp93Ks7f1SokZXxHIdG8dE+ZW762MrPyEN6kIq/p+2dn/GtvmIBc9yfI+xWNEy67WY0YnsD6jHXeugBgx8BVnJjwbcBnBVugccWsBbgRezdz701wgkQI4v3AraDcb8kPEFtYmyODlNNZJBvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk2wB+7h+Ops6cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM1ydMezGn0ONdcHL6gJIlARJpt8QnfDZMEmHeRpJAJgRn+GJxGkvbcbNpSdunsHtby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2Q26j4q+VAd8HG4tIo5YEpurKbRDLBZ59hpcOkpH2V6WOc+MEglnTSDqKE4RheWwcTO5ChtnyodHKCplXICzSMV46VmLu8LHZaz/XSn476O8cHef11XI2sLVbv6OWqQ4Yzry0mXrQk9vQEYjgY4ueShBmX7RArBPiKuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSE7UK/CN/hKc+X6yPE1Wuj6uq6+quZIILtz2u5mISv9/ekAOCaaxKJd4A9eqSnfw53ARTTIGopTtTQ+EHwFInoSUjIZoS0M39+he2MtA9cqAf+W2aDVBLZXwOE4Bv05OIEOxn63eLV1IWDiA6bJiA7/4aIi/A+pRzjGWibpKknJBy/BJV9UtiIl8aWSUg45QJ+EUY5Sut27RYAcQM8A6deifnrBgfH8ACdRM/X1FJBp8PRmJidn1y5Ckf6Jhc3anln+gJk042NZfTYP2BaKjE7bRp6MwmT5LXEoYp4EPFfJu7Xg9FghskJKo0RNRq+2Ge74C+AGhK0QLKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTyNOGBYR8d3lNDEhTGGbKDibi6ANeDp84/9WDQeKblwz6vMQ9YIshs6YlCbGJ6SQuuZeYrvFxsVeMzeSEjdtf7rmSiJFjvg31QyrO39UqJGV+AWCR+RqhhKxeKgUkY0hME131YbqelIVgky15w/MTbiz7fBSngAeVpmkFWFrOe10MVdf0sP8GLr5jSWuuVaacATJaMT3Qze5C0/SkN6W5/RnrB9f+ubikYDe88hbOmTag2vo81yisCMyxFxpn4DsyzhLlHFSBJRsXLjBku5s3rEOeDQER74HaqwuQe4YwbwdaT1PPmfZb2wyfiu21TSzSoNASber4fRi+jwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+zsi8kDgweUqSiAw1icFUot2N71FU5195hOXwpBrxr12rQY5Xnh4FP5Wbpr3Uyr8BAACBDauxhAM3B8UTeMQO7rnswU3AY2t2rWmH0QnDKBij6sAtl2NY2EWfICnSDcVrcx5Q7BVE+WFpHyq54BIBi8J3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb5EEErtNzMD6wvVMR6t5LImGl5hxdZPJpxwB4IzSaZLu93TTEmMqmKLXh44Eru+G2/DFdE/EjAVqH2MjjnaKzehhCFyFSRGN4TfP7KQ4FWvuQrzq6BX7MnoLsT1DdvvEkLHrOV6uonxVQ/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8EmZGuEoHlfUtVYLGusEUEL1TEereSyJhpeYcXWTyaccAeCM0mmS7u0AF6cV6CwbV4eOBK7vhtvwxXRPxIwFah9jI452is3oYQhchUkRjeE3z+ykOBVr7kK86ugV+zJ6C7E9Q3b7xJC/a/B8zGDQT0PyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoPBJmRrhKB5X5wOnAF3tgJiC9UxHq3ksiYaXmHF1k8mnHAHgjNJpku79bNJH2HNbSJeHjgSu74bb8MV0T8SMBWofYyOOdorN6GEIXIVJEY3hN8/spDgVa+5CvOroFfsyeguxPUN2+8SQjoWQg/FEvRyD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDwSZka4SgeV8O5kh72uncVwvVMR6t5LImGl5hxdZPJpxwB4IzSaZLuzTZieecEgPFXh44Eru+G2/DFdE/EjAVqH2MjjnaKzehhCFyFSRGN4TfP7KQ4FWvuQrzq6BX7MnoLsT1DdvvEkJ9e7PSi83Rgw/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8EmZGuEoHlfZ6laVXeHlstCeT0qBtJk/TGfUzmQkKcXDJ9LeExL72R/x+iCgxSc9pdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmGZtznhBvObu+3Rbbl6sYhMmJu5D3fjPc5mw8QDXyQrEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvDvs4X13is5a+X2U2Sr4h2tfpPQ2kXFtYhzzdEPSJT5a+7grw2Uuih50Nrz9FNAQEPr2LbsPFQc/85hXRHi13qvfqYTuVYKVl0u4Abt8zT7TWUWgnEYxS+luIkqfpKTTgsNtEsSEq+RWAL+BJNbGGCro7OtOahbcou0+fKj+43162zEUq06bqVnBZlDDWPRc0fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv19JhV0Bg8FAX8cYC1vw6ZInrSOdnQKWp0tGcGsxfg0omtQ797AIb1pn5zUaoL+FImERhWsm5kQjGQv3X6heHUWyemHUYw8wDnkyOhxNuHYrGs3fCXspGa6pOtkR5QI7rnkyOhxNuHYvuKiazyQ07CygDEbahTo5nXqdpuCbaDKP/28uOGyQRy9yn94RlE9ZSgDV9FwUx4wJcuiL3kkrXA7EluS74MaMaK8+8Ueb2ay9CslRGAo077hOQdnuEaIsM2ev42Ezam8IpAdCTzoILu4nAtkrelFxuxk5s5HEOA0DNMCmC2iEbwIiN9KJo+bsI2MPg4IADwD+0wSgQgIcj/8WgbllK4Y+phEA01UtgKDedK/+s2YPEJ5GrzCGYjXc+9/93mZ2TR9HPxd0F7ZZU0C8IzVw9AQMKMD46cGrXy4hPLwbb4PU/WFIjp1DOt+ycoHMCwDGMAsowPjpwatfLiq/3yDA5sixkkQU3a48Xf2gfiENe0Oug9OImUKXJV+UAr5MLZhS3k9kKmiUYuNLmVgr0VuPCER2USNujLFNzqCzzF7u5zf3I+EUTVH31rEZ73hiwWsip3UylT50JpQ6IZBmmNrOWyAJ2SZuYxABixyiMDhSXtJ91aKs50dX2dBVAiI30omj5uwviiFGcBNEXi7TBKBCAhyP/xaBuWUrhj6mO8wS+TYnIwb7CKGgQd+InicC2St6UXG7GTmzkcQ4DQHJfMicyeYvaWOw6d3mfY4oK9FbjwhEdlEjboyxTc6gvgGj5hwdWGvteCiZpZemRCQEl4tQOBzxL1h2+Z+wg/MY+XytddD6F4yd0IPT9GBmxdT1HB4EEopbKWybNcdnPHXhjv4Kftqkn8yqqCuYL0U+dK/+s2YPEJ5GrzCGYjXc+9/93mZ2TR9NlQBwD3jyrD1ntb3VK7iqiHMMQM43aeF6ANX0XBTHjAIOoc04mT1XtU8aqrXQC9Q2+x7ws0qUSn6mvGigMRpsmTRl/lPGcXmkCp4bzFMiodgr0VuPCER2USNujLFNzqC1NXU7Djqa5yMMoZvruZn7HXAfbv6lmCUB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7gcnfz73q0BWqkud8wbS/IZy13SH1ztbzaUEFn+R72FPnqGuqxTSbv0Eh9mGRVt8RXhOmcqaGhX21pscx5UvVz4WPsQDweHd5IIFX2mInnt8u9xW37AAlntVCrxgQXaiOs4tt7QBeozyqKLF5ZhqmfZtLL+yybWpx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7zhC1rRWGiQMZC/dfqF4dQAByi4Y+C90Y1qeF/3xLYVjbHasb8nNKb74TviO2/cKLXyY4p3wSQhQun+fadIqyRtOCB1pVP/YIVe74nJ6edzid0R9SwaTlvBBQDkg8Q3rOQ9zsKk8AIidXQoFv1vZWB532mKjRs8AuQ9zsKk8AIidXQoFv1vZWADlhEDka/jouqTrZEeUCO655MjocTbh2K5BAP/YCJG9jNis1qs5hxNgngZTYpYIfYyWpHpKzStajg61AfCh1iQ3vOjK80/wlw0bOxDv8HmnztPolD6Gk0Rly6IveSStcB532mKjRs8AuQ9zsKk8AIiLUyStkLsQpg5PbiRLXQkHAm5qCV94BibIqrp3xKIxtDtG1k0bLNkmasdcs7DNaVYgr0VuPCER2WHKqogxnApEmfgrpUCcPDtPSYisw/CJsfh6sbNicQXIi5WhL9Tn4GFRg0eF18pdwFF/LKGsCNOeALfEAoiKF8CuCNt682259vQPjRxVXbyJjpAfkv3Xezi1lfvX7UiJ2VGDR4XXyl3AagpBp+LCkduEREJN+TVUs8dmQhiTjlddSPlEkw7f55TrRGSu5IrBBIdg1suZ9E6/wTJWSiPyNhKrD1oOhUnp8hO7JRb/x7EOB8gtxiLTTHiGvuCZChpPFyUzsVX+qjJ2cFhRLHtr5z2lMrT3GRkm/VdqbH09M40Sqw9aDoVJ6fITuyUW/8exDi2iW8nonK7E+dMGZISrr1mE4CB0rbYpEssW7QMt5W+N9N1GoDN5COpEtRfj9IyqtXDHdoXX4sTnXFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/xMY7OSSvyJ2J1AqBPke3MF1YKbw3tpRShxHLifkb0sGc8rFJQKPIgNsR6DJqCUVytkjreHqRxKOnvPZszYH98tOQZIm7+zr2MLg4TLFSlMPXOLFD8ojL7/gLG/13Fj1hfn7t0tzKCww/id2tyC4EWz5kLyfxrYOao9onXBLEFsaUzMxN3ZVssA6Sgfx+Tritgwdk2R1rKY9gJnn4ZpykqA1Zicz6VVMhCi+G04JfRlAVFYclhD8d4enC3EK7+Fb/ExXPmRW2GhfTCIv7ttHc24RaygtE5naOViCACHbNjEqs6bgY2Nlcm3sraSRM2ri+BJb1UXRUP7vcNfEQ6t0qItIOVQD30rVj3HO1gemEq84Ai5nyDP1E0C7mVmb2+QTluxjbVPe5ExNR2fVmEyqvVNBmcX0e30+UpJjA/vwq7npSeCdmyU1jT+DcSDGIc5qe6AzJs48yu0oxF5kW0MLn8mjqGZ+HZ+yEb3/3eZnZNH0IdgmsrSlvKHkjghcGjiDYSjfqPGNwc8Lw0TuGQVpDZKMD46cGrXy4jy1zdhA6vPOfo7z4kSyXGjyev56LvzxsVRUH+dXRbsnq+9yLK/bVb/BCooBKNUp7sGOdbJ9JQtTsQYLI+YZ9y9Is301tu2NUgAEcvIYF7LQZmlHHhYQb2zI6AyniWV02S5bYlRd8WtlUIhTjrAFHFqMw98LvuzZj3C4ZTnP7g5hHeJhhcI+4kaAKJyw4VX6uaZh+0snz1uVC3zzBCPUeV2Ns4NBVtFnV0ZubqnDdgkq2pCa7pt7BW/4SlMrg4AeN2TE1xI0cZ48v9281ooBjDYJhM6ATqvclfpRTgXgaovpyKfPWlI16cfNq16wGOeBAH0lXCWEsSnICyPety8zSXbAWCwd+65pMMBYLB37rmkwFWggZOTzsP18gPwsN5c8KiRYY2lKl+qZ3ChCKiQn77YtWfJst5SQe0bYXmHqYV8eGc2ZixzV8RUB8MhZKyq/94T3EQeeMd+6xKglXC65iKEuZLJ9gvip0pppfsOio14nYisbvJM8edTfPqAgtpxAQZEcis9l2mFGCIUVT4aZAAkPW02ZtLS4NEi2ctFjXprcY8okM2833tnrMqttSfnW3isS3fmNorx5BNi06hPuchVDPNnUCa7zAmAcxw8jtEguwnGUHq79TgsND1VXHf5yJeGncZV2xvcgLD3MVmnwftB58fzTz3GjMqSw9saJrXoqFOp7cEeiX73KScVTKdMiUJyL/HmTQUwmgKSTbJUGb2I4woDUElXZk7Qjjfohfga0PwGopGN5FQ4XX7DQnfzpsqvvciyv21W/usOSoQzrQ4dQiFOOsAUcWrk7lnXM++/tjMPfC77s2Y9wqKrcVZxJif0Ck0YO2UEFBEeVTjD9L6sEtRlE/0rodpHd613t4pYZfAEKT8GZ52B0SUzYuEhRYfRxZobh+MtZXiu5UQV8FEMIeHeJyIgr0xNdnFsInRFoVMz8s7lE/N2Bxl0y+KwUu21F32Il+s4U2vT/xxzABuHuxsvB00awOFM2bu+WFHT1/jJ9evvwc5rC4OEyxUpTD+dK/+s2YPEJwJQiQW/mp7cFUPI9CR2jkhJ4GtAsMnHhTd/Um3SPHHDNKCniTOYKh0nMIVVZcTIUWIIAIds2MSryTKIkUcCMHWlAqlLKErBp2pfawjjb5jmym6TZ+4ZAL/SjPdZPbMmLnDpjVDYkKfkFmBxB7jjoLuxjbVPe5ExN5LHyHWE5nWTyev56LvzxsSlr35TeoRtZWAQtwjZy4eWr73Isr9tVv1+aenYPyLLrWF3ZgADZMqINRUOOt4BkFObMkZ2fEVkDspuk2fuGQC/QSVDkiTbSp2imZxE5WiPL0ph/U5mIC2ud8tdJ2Vfe3GvQikJWPE7CK+TC2YUt5PYNufPu+h+TiI6nlJeJqL0d1ZmiKIU3ioegvG6Gn9kH3JUYE55YHeIoOOCrltLRHTp7eGoQHY5J32+wihoEHfiJBUpe48G8Uie9P28sza+jCjA7z0L52nuKAi5nyDP1E0Cnl1V+fItZiSA3IsFghRLdLad8u35k2XUw0mP3skyStFRWHJYQ/HeHQW6A1k/HcyOPkgBJUwhBsoza0vpMbdC0AWDQJ3KBpIOcaiSB0pwUUwSoFZbQkvHudU0R33f79RnqbJw4U1eyg5TOxVf6qMnZnRPJTL8CXouYSkX4kZYszbh7N1Vpa3I1e7Xdkc5z3ySeK/7WI1Ktf4TbSNdaFblRWIIAIds2MSryTKIkUcCMHSyEiXTMY+JIioFx3H9zRjg6MAILecnH7NuvDz/TZisvlRgTnlgd4ig44KuW0tEdOm1F32Il+s4Ub7CKGgQd+In9FHc1iKADHJKHozjh0OSjKJnyGPmNyWbhwyaAxLfQPRSI6dQzrfsnsrF4ZBypq7A9LaGidc4WLxFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHWlAqlLKErBpYxK9uLmj5jeSh6M44dDkoyiZ8hj5jclm4cMmgMS30D0UiOnUM637J7KxeGQcqauwTahUVhmB9Wuvh48WgeAe+AGrw5g00TiRb7CKGgQd+InaFiEijCCt1AIdm/n83bxcAWDQJ3KBpIOcaiSB0pwUUwMktyv9CSekV10i/YyK4kqM2tL6TG3QtAFg0CdygaSDnGokgdKcFFMDJLcr/QknpBKH3bFKkOIhwgg/EGv40FAklzBjuRjYD8Lg4TLFSlMP50r/6zZg8QlT84Msn/lKHCR37x+u6GKDdWCm8N7aUUocRy4n5G9LBoVVIPUUpxe0BLRI3+DyLvl4OKyPlCtndtEMoXwrc0LWwgpAf3FqkpYUiOnUM637J3R/b5Q1kQVBI0w9IfQtPOoPsOQj7iMz8mvQikJWPE7CK+TC2YUt5PaVozXmjYIfHud0RWGVAUyxMZPML60V2LXsY21T3uRMTZxqJIHSnBRTBKgVltCS8e4pnbDF2asKJDVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3h0FugNZPx3MjxQAUrtvuvYN/rmlOCs+pkTGTzC+tFdi17GNtU97kTE2caiSB0pwUUwSoFZbQkvHuz8orPTCpWIeLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhRvsIoaBB34iauU1oTSX2YdkoejOOHQ5KMomfIY+Y3JZuHDJoDEt9A9FIjp1DOt+yfdv7czRvnKL5UgdgGX9/YbOU8GPMsjGFEBYNAncoGkg5LFaicXcUrc9YIq0VoAHSltRd9iJfrOFG+wihoEHfiJ2yooR3rR3bFjBfVosytm4w+w5CPuIzPya9CKQlY8TsIr5MLZhS3k9v2s1D2kyMWnMdwO7xcwqNuLSRYue6xyQrqZpHRFaSxb0Yob/G0Ph73qQ6X+shkHMWEgZcH8Q4BBdqyImDHWmkxRiHun/cm49/l6fg1baCEJvfmh4dukp6zB8apRO0SU/GUbqP+qO9rZIzNO2IT5rv+m0ALJ9DE7QoxngX790NXvyOwislSfVc0f9/gCQHLRvIzD3wu+7NmPM9AlMnkIs4pU3vS85A9zaVkP0muh7dxwv3T+/Q7PTTnIaEL4M/DUtk3f1Jt0jxxwzSgp4kzmCod4Cf9C/mocu13OZzYTAfDJK+TC2YUt5Pa/8/T/TJskFHwVJOu/RyyRrD1oOhUnp8jqbdmcoQYqPFC7qAkcRcwYwdImJ6g0sGVxxa/ul5oI6GvQikJWPE7CcrpLydPnYbCkyA2VBukLUFfZITtU129QrPZi+i+QC1gwJ4EETcBLLL5FmcwFiLIa/6ctvWd+zIsB+D15OUZZzmFW8ihsuOeccHef11XI2sIjOFuc2r7u2U5/qQ1p3rDjMU8QSEFTD3lU8aqrXQC9Q2+x7ws0qUSn6mvGigMRpsnIeB4p6fOSuAUUd1BPN1gS8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEeg06jUQ+Vkdiur4JmK/s+2xSqlDvFoY2zy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR9t8viD2PcboLE2o2qgPPbdUzPyzuUT83SpYJhAYmxpy/ZyYvbWLmU53sJTSVDJyXkvRQW+44mEHhPfamvGZc9cKQ3fbP9hK1mODn8XpikSYWpoJfdxr4eb6YPY4MasHhYd4E1Rl7VhXAWDQJ3KBpIOSxWonF3FK3MOhoPLkzczEjqXIExYfdqsCLmfIM/UTQAzOPu2gz+moZ5Yau/i7n7OXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZu/CBLhW1GONHBWGl6/WaiUsTajaqA89t1TM/LO5RPzdG2hWxGS1no2aS1XOsRwGlTo4dhv1qMaw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9nM4w2JNJ+zgeLiSu6qx3woNx0vrInbhVLyBN1K7j5oqNVzCs1YNZ8N3fbCoZ6u0pU+Zhk4Hg7bt6lBskglapV+OIHaUl9UXi/S/CwkHqg2zAMpET5IJFibOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHKx1f1+XtgrTuFICD2nOHqdM+Ge4IUSMDog8QQ46zmxgkWGz5Pqa8LcGnkhHOWLndfkJGrPv+AUqh9TFW4JdLljfY+SK17iu0YpD1cpko4vTY1VxarjbYSyYVxXqkpAiBj9FHc1iKADHPaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMjGc3nODWG+mfR3I6JJgq1e7cHGcmccaLbdTi1x3mcIYkNEPMoCb13rAlCJBb+ant12IRp2JELQfJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfGiMFB2SyS1+j9OEZwp0HMS9nAOXMoiDEkqBrVh6zEKA1epxaUq4HuAp9nz11sp+MkNEPMoCb13rAlCJBb+antziWjcATlXd93O7dk5YeTiJ6c9O0Bg63VvOoYXf/L/aGpxk0KAaU9eZuCUJl+r1Ko6+dhSVvWRZXV5gHmKglRiDMQT5ndyMiZzssUGdd2NvHgfEidBKHLafLk+ksSBii9Bhrvt/y+YAdwJQiQW/mp7fukZUgm5l+TxMY7OSSvyJ2UQDEX4lGWKwxnN5zg1hvpn0dyOiSYKtXbEegyaglFcpilMPUegvhbv9VOEEPlSHPBUpe48G8UifjU/I4ewwbiD8BqKRjeRUOS8m86eC3M/ODKkvY++Zbwb6IhgkZZbtUQvZOoeWO9V+UytPcZGSb9SpJ294uylbYV5gHmKglRiDAWCwd+65pMBMY7OSSvyJ2DnpE6mX0s+f9FHc1iKADHJDRDzKAm9d6N+plWTQJSyw73cMtbcySBzWkPv8rdyGLqDXxlkXGyt+pfPtPcln2uKEqUIAbdLESji/SFSUzTLA0UACRRuiCGcUXTGWfYsZIGGu+3/L5gB3AlCJBb+antwScYc3doVCqdqhif0+tzjiDKkvY++Zbwb6IhgkZZbtUkqBrVh6zEKBjEr24uaPmN8MqztNYZUr1YGxxPxltFAH4Fbsq/pafJ4M+aEC2mLhmax7M6tZYeK72iuplgCAem+tgIIc8dSJLhbRlqAPHg567O2x2dtxztTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyMj1EomkBOXDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8ej7kOjVyC6Z+lJc3Iqn+DLfPV3eKfHu/PL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxPs1XzEObJXP1h2+Z+wg/MUmHqaCdUVS0oWFgEdetSo1OgFKyacnuLyHtmpgoIVG9Gqu0gl7pG4qym6TZ+4ZAL9BJUOSJNtKnaKZnETlaI8vSmH9TmYgLa53y10nZV97ca9CKQlY8TsIDXHDjv1yxOgAg8H/eMiiufhmCh0/sNB3CCD8Qa/jQUH4F5d6D2LdwwuDhMsVKUw/+6xUv2AnDJrOC5IBC2t+/HBWDTpuhP4qLSRYue6xyQoHGXTL4rBS7bUXfYiX6zhTSR+EYhUn6yngsHxKdieRYpxk0KAaU9eZuCUJl+r1Ko6+dhSVvWRZXV5gHmKglRiBE3tygC005pNRtdDlSUixW+gZZ7FiqYx98gPwsN5c8KtvLh+8KncpTGWOEPCi6UoKjIryX2ZXEFiQa4O+SuQnc+X8LkzPjmcf7dx1PZm9Lt4nNKM5HedM50iE/rsSViFSfAPOJZ5hkzOFVnJvCZ8BU+uM4WFVcntDKh1luOR66oDInjIw3gT6rYMfJliQueLHML8H3LkfDQdN0sZE7NCmBTQTA4TPTF4krJgj0vjeWlGDtn5DGh7OqOQqcgg5eUSYaDdzczqiopS45CVLQyni9RM048tBsu7cLjrgV9vZUpeuwrupyCFw2Q/i9SenvYJ+4QHkjGNhy5oTbSNdaFblRAw5qNKm55bahKlCAG3SxEn3O9jvVOYeE4s72vXM/l8Fm0HUNMK1PfYisfQUjoQpLUKWXU6NLN5CvZNE73Oyv7DSoABMgJpjmkNEPMoCb13pfNHiadfmgKLbp+WvagYMoKbmMuXjGRlD9ApNGDtlBBQ6VNFAG5w/Ves++RXBqbpbvfrVTW4P1EO8Nu5cNDjN+9pffkpP0ECAOCIMlvPkFju/N8uCHBPv/1lDgjrYx3nJL28NUmmzwwgMjik5mkGFB7Iyr2PhVCCzMjIDwpMqAJyDJaCGx+54iO5dZt1IpGFuqe1mKbAb1xbOm4GNjZXJtx1W2iPclH6oboIi0Ic7RFJGMZSUNb0n0PPhZFc+mQ6IugPLosyYZTWCEJsKpfTGJ9+WyD/RZULkqOFPmIUduelNiZnUU5GjW8r5tgv0vPLlEVjr8yfq4Iye9L9nmEE26loS5jcYy6paGha5pqfgj8Da+RfpS+7GBK0i6ZHemGqOoNfGWRcbK35cRiFXk5lH5oWsyIbephpNQiFOOsAUcWrhLmDiLqTUvGGu+3/L5gB3UuB0qNOIl0Jwf+MK7hPDW+GRfVPy9wQTwME/lkxplp6g18ZZFxsrfag6rbpJO0yA7xGUYKaSuKP93ii+Ghct3MnHjuenUQZMAbDeNMssDyJ+DaKO+HfWWPJ93tX7LVdh8stuuPVvalU/VtY3yqMaYU2CrIiYLyP+k+WE1uD4+xUTe3KALTTmkW3ZQw/bXVrDjZkJE6PFdRWeTUUdq8qe7tK24SEreA0hDBSvaUNFafoprmaMiGWgzIU+2ZYn19aSVabdsv7VDk7pDSUijWN5iJkTxgcL2OpUYa77f8vmAHVw6EWxEjWq6EDkjTEklU4+fIBGkq7jSxoboK+FZF6apZq5iYBpEaOktPO4b+X1DXq6E6k0oCYu0ULhE3PN1h099UH2kDQdBe4yrRPgF8bRio8ZTxt8u9yvu+49+N5j8NUx7gBn3LDygwFgsHfuuaTDhTPMhItoc6Ta+RfpS+7GBv+CzUFE4PRGyBG6pf57Gq7eHBAkxxdcXIow49YGT/zfTrNlbZwrN4U4vKQvMYe4Rj/CrqYSvtqGQ0Q8ygJvXepaEuY3GMuqWBslTRynrC52Jmstn2WPnFB1l4Ax8JN77XDoRbESNaroVOon67fE2o+HDJoDEt9A9GGu+3/L5gB0rbCHrVgTCL4aW6qSRxOhIhen9flTl3BmWJu5uUQDyE7WNgoQIUVY/fhmCh0/sNB1lIC9xNtA9HxP/npIZ8Jj2MFpJqr5X59iBxl0y+KwUu21F32Il+s4USvXkPabCstZPAB/XLCNENdIb3b44E1ApVwYk6rTBZturjI4RGnWdkoGQE2LVUa5BUH1QSdhfNqSXx4uKyktAfXU5mIdmUsuYkNEPMoCb13qWhLmNxjLqlgbJU0cp6wud4qH3E3/glyjhTPMhItoc6btdDpSOynH3Wt1/BG5Whz7sY21T3uRMTRV8JJQvFylZtY2ChAhRVj/721PjSI4KWxv9wSpfkzOk0hvdvjgTUClZjdhDkLHxMCKMOPWBk/8306zZW2cKzeHO7JBa88Q6xLWNgoQIUVY/+9tT40iOCluIZcgqOrwdjDa+RfpS+7GBv+CzUFE4PRGzpuBjY2VybcdVtoj3JR+qG6CItCHO0RSRjGUlDW9J9M2rIsZ2j1EyO8RlGCmkrigWX4Ha/KFuzNboZH+dJQSkUkIkyPX8UsrAlCJBb+ant4zCy8bEJ8vciKx9BSOhCktaF8HuNOQTF1iCACHbNjEqb/KvBFHoQjo0jQIffM/rU6g18ZZFxsrfKWvflN6hG1m1Xcxljq385A60nEj7rYiBgz5oQLaYuGZrHszq1lh4rvaK6mWAIB6bBxbMmPtT9FeMD46cGrXy4hPLwbb4PU/WcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHXVg5C/HSbgq1fAMI3AK3KTzjNU2ErTzvKkpekv6EBYqXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZg1/2lG9l/YWMHiwATbD+KiEfmlFUJmC7iZ/SDtPy6KROZ2MLP56m91/Q3YtcqFzn9fzyeLG5RUgyTR+UIzCD2jV1nSmtbA90OzKeOakhOUTV5gHmKglRiChKlCAG3SxEvrulmFJfXtIIC1mSktdDCA0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek7xhA+nGH43aDa5c70WeNYpk8rBnyA2a2eY2Nk+uxLPvcuT6SxIGKL0YVxXqkpAiBgFSl7jwbxSJ70/byzNr6MKs/IT2ZPQHhnDHdoXX4sTnbSsIYx4qDmZ+u6WYUl9e0h6mMbAKVhUekD1RzJpDVvT7GNtU97kTE0O7YqpQ3d2HeWSghY9KOODFT0rj25CVXAQ9BMUbPYIWyzSrZCTRoPluBJBuMQkbczDW1P3Omk7cjB4sAE2w/iowzyOGNtmZ8ny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+To4dhv1qMaw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9k0wVYUxRmEITbLz5OIBJLeA6TshBXMkeKg7TSb/dl8EMyetzvpYcpWXRcttFc2rqOZoZjy4QDDmf2gvcC/wtnUxJtA9ZWE5I1gIInv/0WxLIA7j8PfMnuZ+5cA7nYviOOekoY3Dr/aBdeeSdWsmat56gkUc2oa1BG7hq6WZGYOeGxkET/s4ySsH+HtOqV22zkSNVOwHTS/X4SqR32UWvDOWSDF6Maph9NZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkxLIL9TF1yaItfNaX9JCLjgltvwaKfnW3SDxBDjrObGCRYbPk+prwtwaeSEc5Yud1+Qkas+/4BSqH1MVbgl0uWN9j5IrXuK7RikPVymSji9NjVXFquNthLJVW3DiKRkzwsDcSZ7I1QsZ9CTgLGddiM9RCWbeSOoaDeYkZzDDBaT756ZveXfqotOBBgvxoLr2hVm7TFVhzA9nbPz/c6/JJ/2iPRAJAhOGHqEbftywaO5uYx9hM3pV91lHTf8B3+//fS9nAOXMoiDEkqBrVh6zEKDFDV+9J/wBRiVfbovfMR6DMMIMVCYg7BmoNfGWRcbK39cQmC1z9CjGNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOVEOai1ni3uOP9XyPPsAvwWQ6arWa36ObaLqzJmflsPSXt14nAyWWX0NaRZr5dtq7lcwbKRQEQlmWnABkhfYwG9iuoTHUj00cqJRIh0tydLOBzQEh681GqtIVGUW7XnEliuB6xyQBZz1g3folm8Hs8CXH0HK3z8hbbTT3o0xwnyORjGUlDW9J9N1Ec48yadOuk/v3XpfyTq5r2ZfyF9qvXJ1PbkeQjXTqBw/1fI2CvuKoNfGWRcbK35ZPS1/oJxSYtXSMEJaizuWs9D40Ir1ocow6dlAUb6swzs/RQynj5v6VGBOeWB3iKHU98MqCvYcVBviG/kNVfGioNfGWRcbK35ZPS1/oJxSY+eoeEhtfCBj9ApNGDtlBBYbd/hhOo6IV65/iDMVbGEDLyMZ3ZcNv56EbftywaO5uYx9hM3pV91lHTf8B3+//fcCUIkFv5qe3q0oMMMiW2kmG3f4YTqOiFbxiooMp8Wxa3KjZPqsRiGCJEjvoFiBQ9JGMZSUNb0n06sQ7XfRpjeXdRHOPMmnTrgOoame3YhJKx+K1a7voG88OiOyiZeIxq53GrM7Tio95e2Jhhfq0OBvVxH5RzVBk/YmbEZZxuEH2nwDziWeYZMxFT60IR7KgAXGKw5qhIIY+TGx1xlIdeGK6rVpsXNMJFo6FjIdBo9fmrs+PSq35QfthXFeqSkCIGEDN3yDNZaLqijqFd9gfTUR1qzNemUw2QayvLeiQ+SC4TlFZ1EWDqf8xnN5zg1hvpqn/IWTaO7XHAwl+HhDg0Wix++YfTkoVPYGTgZeRb0rMccDLF+oDK4SzpuBjY2VybSmZmffsd5rEwyrO01hlSvVBM/P8u20+93g4rI+UK2d20xf1dm3aO3xhZozdt25vcDNSC50CghXz5oyoIXeJbFsoUHXs3/w08ElL4YuPHyJbWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm/AB1JrK16lcpqhuNAjDDDjOCZtXQttM8yQjG2JLz8lRfGDwa/YgAz0Lr46t7hLCmt7KHJ4f4HgN2woXz0TKgO/0wuRZnVU8ArDcDh/vwCmZvv9rvsLTtvARhHBtsdjRsc4EDOqBnQon9ApNGDtlBBU1iFwsBvacqh4Eqf6OFsR9X5L6vqDdD4juRqmrknC6B8Sod9zHevvFNqFRWGYH1a8pd7uUFOsJ+GrGD2Hb4WNN7VvTah2RHIJxQRjqv6t2XnUUwFY0vVbtwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk1yBfqvVQn9jMMiNBIizGt96Hu9O0DpjbPxScREvltrsHDZMRgFfe1OrGISi5pGmy/7rFS/YCcMms4LkgELa3780Mg70QREKmPkE77jC6kROnRpRErudjt7iWWJBHoCpYmkcovS8Ughq/Vu4MN/18OfsY21T3uRMTTFNXd2820FOH1MVbgl0uWN9j5IrXuK7RikPVymSji9NjVXFquNthLIR6UkUZS6J2TQyDvRBEQqYaDfN8yuJlY1RCWbeSOoaDeYkZzDDBaT79xikmyUKNrP3gRvClmu+NJCsWg2rHz6bYv0GcUwNsoIpCbjHIfzrNblg5fuBTrJoev8Vy9JoCvWbmzzPUPBXvaB+zkuwLOV1Q/jWzBuvjX/AlCJBb+antxLmTerGNq7KEelJFGUuidk0Mg70QREKmMsCz2sxeKgezE2CWteJ6YcNUu5S0LRZXzDIjQSIsxrfrDVmeF0AhpWf2tnZsJ2p021F32Il+s4UajkcM0HTJMWiAiNHs4agN4V/WU3qpuprhMEgyt44zCr89nZhYcsvK3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTe3iOGeUsC/kc/Fu6y1gms7MacMvqox5wNDIO9EERCpgoTXZ+7b5T2wRWYxs0rzYPAiPNmJRuMedwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyOYkaacOUflhYMY+n1HoeHXXBy+oCSJQLCQfKeMfpcFuYvb7Ueb1+LsDR5sG2RgC/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxDrgzq2MKWHGo5FiHNy2C/uswNMGaW4iR/FJxES+W2uwcNkxGAV97U6sYhKLmkabLLxXxvnwYbtrLApOQol6t35ciTUmVl2Ny+VvqxG/F6K7hJKWdRMLZCDGc3nODWG+m0S06RiuTZys0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm0pmZn37HeaxBbxb5+Nq/QPJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfsqhNWCzrW4Px6uW325OK0mz8/3OvySf9oj0QCQIThh6SoGtWHrMQoKOFM3vPrWmZNDrz/dM09R4aYzfjTC6+kbOm4GNjZXJtYK3CE4cXXxcIm+/CbkyXViVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3wwdk2R1rKY9vnPEjtNeY2JRCWbeSOoaDeYkZzDDBaT7oSpQgBt0sRI8UrTlyyOsfL0/byzNr6MK9qoHINnqNTQT1zWClEYtH4XLjiOTjsUy9xovJ2mxAzRLvnX2Duhfj3UWKJQ6R9GzprfkM6pnQKu/EUKWXiWm56g18ZZFxsrfnDmt+KZ4Mh1VWzUdziaqoxr0jRh3Dlj2e26IMgzJNWmQU8dw7feh4jgJ6ZmFH1r9twboZi55jEGoNfGWRcbK32jqtGKczLXhYhg/UIOd6cyWnABkhfYwG9iuoTHUj00ckqBrVh6zEKCL0RV+wrKe+KfiqBihguvh/S7x1rlSv82SoGtWHrMQoBcTnoqAAyXdp+KoGKGC6+GlZdKbZiRX8hD0ExRs9ghb0uwTtBtpz0T/T6desC057u3m7P86uO5uLB2u5nwIp96H6AzzQsMsD0s430bqnyAEyl5/tIagyVitr1oAQUPw4BqGgTFCbJiQUQDEX4lGWKzKXn+0hqDJWJqxY4lWWZMXoQ4aBSpzwGumYURHNrLDk8ffPy3ykWGRkU/Wu/pO/t7lzhRMhUwT2eEkpZ1EwtkIRN7coAtNOaRQ9ISXbmEENqc5pNmDRQaQ11dmm5vyS3m1oGx8AgVTGd3JflbH5MMKRN7coAtNOaTYKu5maVzQwq10g7jIlhmIsohlQOPzlxx4ud2ifpytOyG/zMuttlk6ZFxltn31g5bWfIs/JKfT5+xwq84wErVKuCfi9rWJR5aSoGtWHrMQoMbXe09SFZZkp+KoGKGC6+Hsaf2MkendEcBYLB37rmkwDB2TZHWspj1JqWNRDiSJdEQNQLTZeyIoFpziG0dVJueDKDWQOh0cR1zixQ/KIy+/OEONYiYwWXWTQseOx3I/54QOgo3F/ehSwFgsHfuuaTAMHZNkdaymPVcIaOmQsF950bvMLKa0xpaoNfGWRcbK32CtwhOHF18XneP0N/uBkPOAXTsdYWVnwEylUvnwwkFCajkcM0HTJMUCgedoCuA+3Sxqu9nXfz0fVCAOBDojWhA7LYcQYl0OOL65j3Lu4pRvHaY8JecNSSkz0Z/v5WXOY91dVSReGT08l8NuPit7afpTvXeA+EzUi9biHbGth/vbkYxlJQ1vSfQUT2J90ec00YM40BRQKurw+YbHwIT40zfWd4V+hJ7yXh0pubUaT2VbYVxXqkpAiBiIxKUD+YXwlQp37lscs67vo9Sz2ROrnOJ7roE+YpEbxRjw3rHtyzD6DB2TZHWspj2rSgwwyJbaSWxIXvOJu4IsOOCrltLRHTrxQq7F7a7w3ng4rI+UK2d20xf1dm3aO3xhZozdt25vcDNSC50CghXz5oyoIXeJbFsOuDOrYwpYcajkWIc3LYL+RK3rZqU420jy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOFJZfy2x950437qMTokd4LD//YU7iEetmz8hPZk9AeGSKcIW0S4ke4FXzu693lZFSIxKUD+YXwlQp37lscs67vQwh9hDMyBQfQ57pjagUkkdSMm8EQGs7zs/IT2ZPQHhnxiaFR/tfzL9OZgk+wyD5DTFc+ZFbYaF9G/RZgc5jNm2Z2JKG1Ab8BWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFl08nQc4jWEmxEWirsvf/0zOLt7Yp1VWFUIJjubSHeqZ2fPFJUI4vifHy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Jse6E5dN5oURBBMqGQIwKAyj+ihftNPNpri6ANeDp84/kmbmMQAYscojA4Ul7SfdWuooThGF5bBxwtZ0QBNEyPNwEU0yBqKU7RmOYgTRnNP30iQ/6mZ9pEFTfNmEUmqMgcFqtQFTH7C9Iyshl+2ZnBkPyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoMCqmU3dxUTNT8BqKRjeRUO3gy+nTaA/6/kavMIZiNdz73/3eZnZNH0sVty0jvqyd7jn30dsLXUp14eOBK7vhtvwxXRPxIwFahrxORbj2DDnLVRbMaU9R3EaHoIXpunfjtCQ/UWBIJ978fLpL/P9hSAPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuvmNJa65VppwDrVedGrotX22kYId6HEltNdZ0wkesP4yFWjquXsqsGtkP4vUnp72CfuEB5IxjYcuaE20jXWhW5UWUNpLBUAVv7u0ekMY82N2FASXi1A4HPEvWHb5n7CD8xw3jAwnCbrr9rnU4xMwhhXQkNgHZGapfQcHxRN4xA7usfl77NJjyw0enRjNxs6iZ4MB3hZUJQ5OkDI4pOZpBhQW/jxpmwgjWW54NARHvgdqpb8lZHdGhSIqcnLVu656ddo8DxcgTS24wpoifs1g0sYgvlmBdWPHvseWX0sWWA7rvHSk34WIXHAhye0y2l+Ioi9wPYj0gtnsaMD46cGrXy4isR4oKvE8eWyo24N/V7MkQi5Hd0uVs/QmXmK7xcbFXj52NFPl31wE3Vky97a5W3s6EM6PsRQw3riFct+CLnHGHTrNlbZwrN4U2D9gWioxO20aejMJk+S1wjOHP0uzGnHo2iEt8BRUs6KVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTy7kZ9lmlW+P6gJaNwQWSsShye0y2l+IoiQmYYXfngN8q7oVVs+9lAazPGIAtzsAXzTj72s1kXJKF1nTCR6w/jIXNu8mA6BEu7Q/i9SenvYJ+4QHkjGNhy5oTbSNdaFblRZQ2ksFQBW/u7R6QxjzY3YUBJeLUDgc8S9YdvmfsIPzHDeMDCcJuuvzOeFTUZsDMEV+1MHGRm5vQiMeUPsFfKzzUTC4AFRZ/n52NFPl31wE3Vky97a5W3s6EM6PsRQw3rDBTzW3u6YLjeOLHjm8vNd9aYfRCcMoGKPJwZXjsJVV1yuxb7cV8hF7wPLueC2ZXK+GiIvwPqUc7IeXjNT8tSYsBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwu2TXWro5hPL9cehfR54gyffgbefuh/1M6NLvPlfAjkbkavMIZiNdz73/3eZnZNH0sVty0jvqyd5GI4qA6CI5342zg0FW0WdX3cB+INvxpLpeHjgSu74bb8MV0T8SMBWoa8TkW49gw5y1UWzGlPUdxG/x0uNED2jcnwjlW3HkivtNg/YFoqMTttGnozCZPktciGXIKjq8HYxhprdQ1vh8+g/IYWiIqjyhXlB9PcWZIkk3FsTkwJY81cBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMB96kY8IIjl1L0NCG4eImb4pa9+U3qEbWfFsKlx1mfqPZmVQ/iwXbys10enXzv/Z3yf/lIi5tAjPt5/UnNypsJ24ugDXg6fOP5Jm5jEAGLHKIwOFJe0n3VrqKE4RheWwcRcP+fZBeE1wHRhm2epZiYheHjgSu74bb8MV0T8SMBWoa8TkW49gw5y1UWzGlPUdxGh6CF6bp3472yooR3rR3bEoUehIK1LLSaPA8XIE0tuMKaIn7NYNLGIL5ZgXVjx77OyLyQODB5SpI4ZWjlaWKT3DFR0jIQgdxEBJeLUDgc8S9YdvmfsIPzHDeMDCcJuuv59Q22YdNV+XqWSbC1Xw9h5b48tYcnBx2ygqZVyAs0jFLKSKzKkaabfOuiB6J/O9FHyNEucKocBuLsT1DdvvEkLgS7psfl3kYg/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8EmZGuEoHlflYarIpZQJ1Jg5Lf+K6r8Q065bNWSRgdXfBIDRqGKAPqogwm4UoeHslnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTKoMmaxH/2RaiHP4+DbUbD7DTMH1pYeVyZqjTTHV6cgoUlU5L/M5+MB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwty0FZSqHxxyyba61mL7BzZyM7HsuArKxnWKgQHJEW7mr+b1+0cFNq4p5R6wQtO5ErbvSeYB5Wlaoqq+DAj3H+611DFD/WjcsIsN0j05VF2845BsIBn4E+p2tvXwJlKpRDFAFR21dSD3prZsMI5If2PUZWRvRhR8T+dnWUc0rmwGbEh4ZYMZnP+J8INnicMgBu/nfIMm83p+HzHdP6daf35EzYWBrk4CmlNmcjidK2GUszmkN4NvJP45rBaSix9SEwMZWQ/t+vjg24S7MtAeUHgua9hF2AWlHqMjXUlPGluXsHdA6JnAJKc4JppTCIZXB2xAc0k8FOSJeOJzN1aWbkWul13NcfrtCt6CFTH9NElHHLKVEcAzrpp14gOZlIYAvylVI5U9r6HGuzaskJ0t8DF4Y14cu4wOOWOFXZPAKpZADnkspgM9yDOLWdTihq5fNsUfyNj3fdwuL0LKP82o7u7JyuEjckbVktW5TwB2gV6RRNJu74PkAwaW3cu57R+r0QAyrlX0gor6kt07wCLvaFL0sjHjPOUb0zcUECgwZXCjE1yGHQHFsp1jMdMjFP6oCH0KWvjiqZu2f4QQY2ggkjI+4Thz2RZWraXcjdROOYkivQpa+OKpm7Zu3wi7RwaKz2XPav8BEGLU3YAdZrAqa9Mwg+SFO4YWYS4sHs5YKNom+QJ2hHn9a8aVS7MXWCJPL8lG/wQo8u2TW+pbmcnCDUJaRJEXOL5s/3my8G10yS4nHEx4kZVvK4LPmzJjv0jbyHoEixDSOaunbw8yrBlALsZk/l92SRuPTl836aGJ6c8Fb/5eWNM29TOkggVfaYiee2LGLbTW5DQLQ9f5MSqbLD8CMnlLxQHHMfA9nJ+iH6Y1aG92mvSKuyJRPASFTGAlbGHJE0BCHjrbBmxANNNUZAyw+X/Plo19sJ5Tb+spHGP86Optg1IoOK/UAnTvq7uXQhPh+vqqcWlNP2r8TIH2uO0kn3sgcdrMwsNz4rRwjBiQZE14vDqwgyyR6R2Io1Apt6iQ6J/V1vTdYgGMQTaPjz4XKMWHy5Xllwm2utZi+wc2RRPYn3R5zTRnGuANZTsWW6wKiLOWMEK+Rph5S9PiMfC+R9U44PrDq7mlwjuN09KXnMTnspNe37kjDz18Ia764Xp3v9OgOxUf8gX+lOdzu8wQW6A1k/HcyM0PjlidWHKnzdCSRiEUsATFKZjcaqZgVuRWJoAkfDaqblrCFXfVz7+ZNChmFOPz7M81+yMnQp2Nyo5ozFHJQV3+4yNGfFXJqycFmUMNY9FzR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/X0mFXQGDwUBfxxgLW/DpkietI52dApanS0ZwazF+DSia1Dv3sAhvWmfnNRqgv4UiYRGFaybmRCQWc02j3u+2kOy44C5ZqFQCn5vz96kpWbarmDIzkr822b6s8qwQE970EPDmeXSehv1knBXlhDPOgjbPf3JibGS9KAiuTcO6Px1knBXlhDPOidKCAKe7ioPLBQFOQvZ3yiVjW1fM47WbtJi8mo3u4XzqNUbehcOlfX6pOtkR5QI7rnkyOhxNuHYvuKiazyQ07CygDEbahTo5m18mOKd8EkIcL8CR+13B7XkmbmMQAYscojA4Ul7SfdWts7gbstDN5asFAU5C9nfKKmCrQtaJvfTpSneC5GunO6sZObORxDgNDJWLkF3ibwC9JCZTW10xy+0kpBS5r4LY4+/8gGLek9mi+nta1340811ph9EJwygYrzD7h2IUGu7wLfEAoiKF8CuCNt682259vQPjRxVXbyJp8DpgLoxhi6Ik2IJ2hGPYqcLahDynC0qMEfppvqcUz6AavDmDTROJHSgxLdGV0Lwmm2mMkhPMtOrD1oOhUnp8hO7JRb/x7EODssUGdd2NvHIsDQD9+IkrZmAmFR3LKaecIKQH9xapKWCD6zeYF1nNeZC4OtsJ3yBH/IpES0LQakrD1oOhUnp8hO7JRb/x7EOLaJbyeicrsT50wZkhKuvWYTgIHSttikSyxbtAy3lb4303UagM3kI6kS1F+P0jKq1d4SNc73+P83Hdtxg6oOGCMomfIY+Y3JZuHDJoDEt9A9p3F2/KZDZS1CQ/UWBIJ97/83YxNodUb3EWsoLROZ2jlYggAh2zYxKrOm4GNjZXJtVBRdCi75HEfNReFosymZhGF9B4gUjchi1IybwRAazvNCFBodbJdoT3VgpvDe2lFKHEcuJ+RvSwZzysUlAo8iA437qMTokd4LMdwO7xcwqNsfSSbQfgTQYg+w5CPuIzPyroTqTSgJi7T4SW4WqIeN72vBAGOel1nyjA+OnBq18uJvaTYvfvLB7J7Jpks72RHCvt0W25erGIQD9tcnMj9RLkRYqq/gjr8D9YdvmfsIPzEXbRnl4L0Q12nwF2qWDbObnQgpUI7ZC5rnMUy2k7tYkVMbIkusOU862QzUkp+X7SH4Wi2hEgoSyP0QyDeUmpFxLCeQNVV2pHjRhWLP1OR+C51/qcGxeC8O1635+2GvFBT6g8kyTnTtOdBmk/RnodzdrZ+y1R+IOdIY6Vc+Q2OYPpkLg62wnfIE03jce2p7lxHFX/ozmn9HsO/MErbF21mpFIjp1DOt+yeysXhkHKmrsA5XrNsX18DpEWsoLROZ2jlYggAh2zYxKvJMoiRRwIwdaUCqUsoSsGnvfAdTI+c+lDVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3h0FugNZPx3MjExjs5JK/InYm/iT4JatGqhFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHWlAqlLKErBpscySv1+2J/itqwjWtdgaSxbvLaxlKjRTHEcuJ+RvSwZFXGCifSifHMb2a3wBSeOcPMCck2tjnuviwhw0QQOyYaOhcaeXTu6VKYpuXYGa4XRr0IpCVjxOwivkwtmFLeT2GgallM90IE+MqGLRaexoCn+5OB75NeKcNWYnM+lVTISKQvleug2OFFRWHJYQ/HeHQW6A1k/HcyMzoX/kY9emE0fanTTR5KBPY+hjyRwMfUD0PJ+X2fy9z/WCKtFaAB0pbUXfYiX6zhSnJ6defzt03ULKtEsT5F1cCxxfhOuc5BRmmEIaj2s5WOUaIwNIC7gC7GNtU97kTE2caiSB0pwUU8nghxtgSf/dxglGv1riOPHZPbL0NbZsycIIPxBr+NBQgrlhLggsqd7C4OEyxUpTD+dK/+s2YPEJodQ61vbxLBOJ18ZhYU9M2sTx35SW6QjngefAXytcIYkcRy4n5G9LBoVVIPUUpxe0xvZrfAFJ45w8wJyTa2Oe6+LCHDRBA7Jh7Yvb+s7pzrexPs6payz5TFiCACHbNjEq8kyiJFHAjB3u0V+ntFmUQReUb/rApcMwb7EyD7ylLauSh6M44dDko5SeTYBFa4Rc4cMmgMS30D0UiOnUM637Jz3hEYkg78NmOSD5Z/3G+J4nQyL0GMAaKaP33I5QEiCsupmkdEVpLFttRd9iJfrOFKcnp15/O3TdQsq0SxPkXVxGB9EArYhg6eO9Lgf1mcX0ggkQSYew5vUcRy4n5G9LBoVVIPUUpxe0xvZrfAFJ45w8wJyTa2Oe6zP9pETYL18Pz6X3yCyT/csYGXhDpCZo02vQikJWPE7CK+TC2YUt5PYaBqWUz3QgT4yoYtFp7GgKGyObHvsQT+s1Zicz6VVMhPOT0CnDw3pwVFYclhD8d4dBboDWT8dzIzOhf+Rj16YTR9qdNNHkoE+viFskT/G0eg3NAS0x7zxnWIIAIds2MSryTKIkUcCMHe7RX6e0WZRBF5Rv+sClwzASAdKD3JZybwIS6f6GLoP5g0cDMgQwDJ3sY21T3uRMTZxqJIHSnBRTyeCHG2BJ/93GCUa/WuI48XkGSt8JC63kwgg/EGv40FA9fZwWGKnHe8Lg4TLFSlMP50r/6zZg8Qmh1DrW9vEsE4nXxmFhT0za9dLVYRpNglekWh/Hpoj0SBxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnDzAnJNrY57r8W32jf1Y5gN4T+vZ75NsPaoKuQ38HJrla9CKQlY8TsIr5MLZhS3k9hoGpZTPdCBPjKhi0WnsaApO5U1W9cQH+jVmJzPpVUyEKCcjwbuij8hUVhyWEPx3h0FugNZPx3MjM6F/5GPXphNH2p000eSgT9tf1AuzAaaAMG47GihGrk5YggAh2zYxKvJMoiRRwIwd7tFfp7RZlEEXlG/6wKXDMMNoDsfxRWpPkoejOOHQ5KOEerbdTBHSlOHDJoDEt9A9FIjp1DOt+yc94RGJIO/DZjkg+Wf9xvie9MMfHGpfTFij99yOUBIgrAmtcTed3vOWbUXfYiX6zhSnJ6defzt03Tm4esGHzrSvyr84DlQ/NYSgjsd+B4wlYLIrtKaqmw5r7GNtU97kTE2caiSB0pwUU8nghxtgSf/dzYDqHa8kpfFf7l3vMIcQ68IIPxBr+NBQuRh3QlVe8E7C4OEyxUpTD+dK/+s2YPEJWgyYneqoRKK3dfjuuFuzw/SLbCqk4/dmHdEemZnDHWscRy4n5G9LBoVVIPUUpxe0cgzTsiYq6X803iPskC6pCsBYLB37rmkwS5llCfipj1XqfUNT01XmRmvQikJWPE7CK+TC2YUt5PZEYh99MRC+TyyJodNzTB2auL8FGFJ51Hg1Zicz6VVMhCi+G04JfRlAVFYclhD8d4dBboDWT8dzI/LnwcqmuS4OTdlAWTqLPTg9hizAfxtHp4tJFi57rHJCupmkdEVpLFttRd9iJfrOFG+wihoEHfiJ2yooR3rR3bFjBfVosytm4w+w5CPuIzPya9CKQlY8TsIr5MLZhS3k9v2s1D2kyMWnMdwO7xcwqNuLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhROuWzVkkYHV3wSA0ahigD6Tzr/ZBmu0bANol77WNAY2/J6/nou/PGxoQzo+xFDDesOgH3CGeeYPqWiXs4VWi+d0aejMJk+S1xKGKeBDxXybhKar2s4P+7y1fJdfYoxciEMn0t4TEvvZPGLGDSF+CVNEYGX9ylO4vk6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcrZk9I4Ew831nM+f3x4X/14tUf2Bkgs2RzokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyfnj9i0dWGvi9/93mZ2TR9HPxd0F7ZZU05oyoIXeJbFuwNu9pJr5KepciTUmVl2NyLaph3YSB0q0NBQUlLIPgxU2EM6jlg+dX8wvcQ79a/M2OHAgZShzLsag18ZZFxsrf1uhkf50lBKTUe4+pr40+z8BYLB37rmkwNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOkqBrVh6zEKD2dlkuVjPjlcBYLB37rmkw+xl4LFtVes5RCWbeSOoaDeYkZzDDBaT7wFgsHfuuaTATGOzkkr8idiYO8dPPbfEqHrSBiMTQxNm7cHGcmccaLbdTi1x3mcIYkNEPMoCb13pUQ5qLWeLe44XVa5kVzYX2wFgsHfuuaTD2qgcg2eo1NMOTyNLgcNdkQIaAy+tSTHGq/E96ZInMfqg18ZZFxsrfBsrdFIRoGlM5IPln/cb4ntXoFLuUIVmGNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOElqjsKdbEtkXlG/6wKXDMA7Mara6L1S++xl4LFtVes5RCWbeSOoaDeYkZzDDBaT7wFgsHfuuaTAzoX/kY9emE0fanTTR5KBPMRky4G1yPMi7cHGcmccaLau89FjbHlF3E9c1gpRGLR+OL9z0IaBXzIL1NfmwBjAaQsq0SxPkXVwLHF+E65zkFG/yOlKCkRXXJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfBsrdFIRoGlM5IPln/cb4nls95sBH4O1QNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOElqjsKdbEtkXlG/6wKXDMCwsHchF7Onh+xl4LFtVes5RCWbeSOoaDeYkZzDDBaT7wFgsHfuuaTAzoX/kY9emE0fanTTR5KBPmyy7R5vu+py7cHGcmccaLau89FjbHlF3E9c1gpRGLR+OL9z0IaBXzIL1NfmwBjAaQsq0SxPkXVwLHF+E65zkFJGLKma6UlxOJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfBsrdFIRoGlM5IPln/cb4nlKCotR+OcP/NJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOElqjsKdbEtkXlG/6wKXDMDgwUsXUH9ob+xl4LFtVes5RCWbeSOoaDbtwcZyZxxott1OLXHeZwhizpuBjY2VybSH7L/kpD1/cxglGv1riOPEfC1kBC0aVm21MTiQgElzkbPz/c6/JJ/2iPRAJAhOGHoL1NfmwBjAaQsq0SxPkXVwxZZG42AAG+LEl5Si1z+ZzJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfBsrdFIRoGlM5IPln/cb4niXwcmFu+eV0NJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOElqjsKdbEtkXlG/6wKXDMBIB0oPclnJv+xl4LFtVes5RCWbeSOoaDbtwcZyZxxott1OLXHeZwhizpuBjY2VybSH7L/kpD1/cxglGv1riOPF5BkrfCQut5G1MTiQgElzkbPz/c6/JJ/2iPRAJAhOGHoL1NfmwBjAaQsq0SxPkXVwxZZG42AAG+BCdq8S7YMFyJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfBsrdFIRoGlM5IPln/cb4noWUEJUMQrqcNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOElqjsKdbEtkXlG/6wKXDMGyB5lyBFdVj+xl4LFtVes5RCWbeSOoaDeYkZzDDBaT7wFgsHfuuaTAzoX/kY9emE0fanTTR5KBPVlyt5qtbmIK7cHGcmccaLbdTi1x3mcIYkNEPMoCb13prVatREbv36IyoYtFp7GgKRuhrsJReP7T2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTKRx6G6Y3CZNTzAnJNrY57r8W32jf1Y5gMvydDPl7I1qECGgMvrUkxxN+zZPe2/uq4Ya77f8vmAHVoMmJ3qqESit3X47rhbs8MykFBdRlxZwTQ68/3TNPUeGmM340wuvpGzpuBjY2VybSH7L/kpD1/czYDqHa8kpfFf7l3vMIcQ621MTiQgElzkbPz/c6/JJ/2iPRAJAhOGHoL1NfmwBjAaObh6wYfOtK9lxPJECl51eBCdq8S7YMFyJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfx/Qis4Up03Ejw4o2he+6PsBYLB37rmkwNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOxmoGyhcGGitN2UBZOos9OL0prYqxmTzK+xl4LFtVes5RCWbeSOoaDeYkZzDDBaT7wFgsHfuuaTDy58HKprkuDk3ZQFk6iz04R7f/Z43QsIi7cHGcmccaLbdTi1x3mcIYkNEPMoCb13oiEFgcKS80jKWdRgA3CYSvMpBQXUZcWcE0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm0xnN5zg1hvpm8nfbON8CfGwFgsHfuuaTA0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek7xhA+nGH43aDa5c70WeNYpk8rBnyA2a2eY2Nk+uxLPvcuT6SxIGKL0s8TuxAbbviixSLbK2nsPGFAkSuU96ebilpwAZIX2MBvYrqEx1I9NHJGMZSUNb0n0ElhgOkSxvx2wsiM+ceaaCsxBPmd3IyJnOyxQZ13Y28ciwNAP34iStikJuMch/Os1uWDl+4FOsmihKlCAG3SxEkb4H8hrATh4fPBntcazikktwnqTq6NAuxhrvt/y+YAdN+plWTQJSyyCSKAiy43mJhUEU0INUM9QuKPqxC7RtK+DKkvY++ZbwdP1wyS/3aSrGGu+3/L5gB22iW8nonK7EzLqI6u0j+FXaG/2ofzXiiywb5BE4LPl1sMfPBlsntgLplJeHDglFh+OHAgZShzLsag18ZZFxsrfMZzec4NYb6b40muXOoOHZ5JIJff7NywdC15MEywTNkDsZ+HD2URmm/4Fh0Qr5vNq/1U4QQ+VIc/9FHc1iKADHEmpY1EOJIl0ZbE/A46UybqoNfGWRcbK32o5HDNB0yTFAoHnaArgPt3V6kmAJ4eDlgwoAcRhnygGsgQYUFr9YowYa77f8vmAHR36V+tUnb18zg2xdgp8no0d+lfrVJ29fAs1LPn6HgQx8Q3aPXoTFS2u6fnFt336nDjgq5bS0R06HfpX61SdvXx3k9A5MdWTCIQReu5uH1PuYxK9uLmj5jcCgedoCuA+3ZGMZSUNb0n0N4SUY7lQA7K16i0mUQtXQ6f24hpCv4lMfNdZqQwejkCOeAt1ewM0/sBYLB37rmkwM6F/5GPXphNH2p000eSgT7f5COxpDxYeImj7vy7rUifxDdo9ehMVLYkTUVibScnLlidT7bPQijPAWCwd+65pMMBYLB37rmkwRIoLn9egg/BH/aTihIVCKrQojrs1fywOGGu+3/L5gB3AWCwd+65pMMBYLB37rmkwwFgsHfuuaTBUQ5qLWeLe413so7/7iF17O6dZqM3gPAKRx6G6Y3CZNTzAnJNrY57rM/2kRNgvXw/6mKU2THl66+BogNuogAOMGW00sQPhj2EzoX/kY9emE0fanTTR5KBP6ONzp+7hXDGHPXlibT90mZGMZSUNb0n0EizaPfb3cbrNuixhPog1YIL1NfmwBjAaQsq0SxPkXVwxZZG42AAG+GKvNqPuoqOLFJsutPhWnAUXlG/6wKXDMMpYEYyxiFvVEffU5rv2DP/AWCwd+65pMMBYLB37rmkwRN7coAtNOaSL2Y7OhP68ULwwAh8cTZElwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTAGyt0UhGgaUzkg+Wf9xvienaIh30sE96LAWCwd+65pMDOhf+Rj16YTR9qdNNHkoE/4N8T7k72rpmexTkzDK04OOSD5Z/3G+J4FBPbvxVaVh8BYLB37rmkwwFgsHfuuaTDAWCwd+65pMESKC5/XoIPwEQ5TdQq6YFm0KI67NX8sDhhrvt/y+YAdwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwlr+ygDqvd8xCyrRLE+RdXDFlkbjYAAb4bKGaAV46YCvj5RcgwgjQhQ8PxmQ971X9emN0zedPSLS7vihb8ZETmgnSstrzOjdxkcehumNwmTU8wJyTa2Oe6+LCHDRBA7JhLirM+NHltlQEw2W9SYdJ0InXxmFhT0za8vW25wxRx1GOymG4mwLpAF3so7/7iF17yyZEpp3jEryRjGUlDW9J9P6yxc7Et6q1zbosYT6INWCC9TX5sAYwGkLKtEsT5F1cCxxfhOuc5BShHe2vw3ELfxaJiTslwsXZGW00sQPhj2EzoX/kY9emE0fanTTR5KBPB1dvVDZvlRBhG1YDzFw/vkTe3KALTTmk2t5JCjnSzRu8MAIfHE2RJcBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwBsrdFIRoGlM5IPln/cb4nly3AX5roWG1wFgsHfuuaTBvGmZYvZ6Rpjkg+Wf9xvieae2MJgG5lf9nsU5MwytODjkg+Wf9xvieesjA98mAqWJqdAZaq+1S7ymeB61MDrynLDrxri4gVNTsvs13HGK2qjzAnJNrY57r8W32jf1Y5gMm/FsGqxUtHjzAnJNrY57rLTqW1K22MmjU+0JrU4Wj4tL4tUjYqPlgeYlKCdCnI5OoNfGWRcbK30hktkF8Zqu5SspUvMPS3DGU1YyGTrnjE5lBTmlRMXB7GGu+3/L5gB2h1DrW9vEsE4nXxmFhT0zaFm44zKYzgwIpuYy5eMZGUOmQnyJT2hswh6gGBmPEJ+/2Mtq573DaJvEN2j16ExUt6UKy6HtG6CrAWCwd+65pMIwPJOfwW7QeMD0ktcLH7SqoNfGWRcbK3wbK3RSEaBpTOSD5Z/3G+J5oXFkLyIYs6BnJEViV2WJBmT3jF9rhCmPAvQf9U4/chYyoYtFp7GgKZOFmhAL8IsKaadZBAWn6fq0vB7aGVL+n+DaldfTwJjRFecCozoQv+4m81zCsbjdDwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwElqjsKdbEtkXlG/6wKXDMF2vGOFFzwj9v+BI22dOZAuRx6G6Y3CZNTzAnJNrY57rLTqW1K22MmhbX0FxEDOBmKiao9ZS5E+V3K0BMX5li8NCyrRLE+RdXEYH0QCtiGDpR9vSXKfqf47dfQ2eJPzG5ZGMZSUNb0n0NQzLe6b5AxHNuixhPog1YMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwodQ61vbxLBOJ18ZhYU9M2jW6aToNP7rugvU1+bAGMBpCyrRLE+RdXBJRhXxUBWUrnrQMNNogG98WiYk7JcLF2RltNLED4Y9hM6F/5GPXphNH2p000eSgT2WDQKEUUAU0AyxGFtzVFvtoiFvadXdngS1AYxVX/WNzvDACHxxNkSXAWCwd+65pMMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMAbK3RSEaBpTOSD5Z/3G+J6+LEv4cXmyx6g18ZZFxsrfvWonbqyIlKW2f69x6ZFzBcBUbemBPy35DxSybk4EmijAWCwd+65pMDOhf+Rj16YTR9qdNNHkoE9ujC37r/G82iJo+78u61In8Q3aPXoTFS1hw6npbjMOemyntUQhEu87scySv1+2J/gcTrv6tkFuN0SKC5/XoIPwR/2k4oSFQiq0KI67NX8sDhhrvt/y+YAdodQ61vbxLBOJ18ZhYU9M2p9OwdCmkAEb1/rylGn9XFGuwkNDcJGIqMIypRx1QSEFOSD5Z/3G+J46vkVT48948eWcBDOJsKPIFOPV/94X/vq9xLR5NNK4ADA9JLXCx+0qqDXxlkXGyt/AWCwd+65pMMBYLB37rmkwwFgsHfuuaTBRbaECQSOEDZk94xfa4QpjwL0H/VOP3IWMqGLRaexoCiiKfvWE7COHmmnWQQFp+n4nI4HlVbgl2xJao7CnWxLZF5Rv+sClwzD5y+9P+EBA6Che5TH98v4d4OcO8boaHfeQUmWM+w322zzAnJNrY57r4sIcNEEDsmGknQM3Gmmxs8gb2V3YicvpBD5rApKkucSB3Y5Qs5wnn3A9braIZnlTwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTAzoX/kY9emE0fanTTR5KBP0c27w92zFd9E3tygC005pDOhf+Rj16YTR9qdNNHkoE/TsWw6PlYF6DOhf+Rj16YTR9qdNNHkoE+3VJH78NDE6lSBZIgI35Rgbs37l3tbKUHj5RcgwgjQhQ8PxmQ971X9Tk0wwOfr5mg6P4C/QXl80tru3h4LMjmqhBJMQjlhdgiC9TX5sAYwGkLKtEsT5F1cRgfRAK2IYOkWSWrOjCwtXSLMSFB9p6vVscySv1+2J/hJ8A8pbn8qSGkkkiw4KT96idfGYWFPTNqySGBBht/JVkTe3KALTTmkkDHd5DolrDG8MAIfHE2RJcBYLB37rmkwM6F/5GPXphNH2p000eSgT1TPaSqv6T7LUHk7KWmEpPux7Lu2DuBUvMQB+NFEmBdPidfGYWFPTNqB1Vcf9unqxnzHzDCQWp80Ng1uyzYlp0EX7b9stNUTSbQojrs1fywOGGu+3/L5gB3AWCwd+65pMMBYLB37rmkwwFgsHfuuaTC1/rmJlpZgcK7CQ0NwkYiowjKlHHVBIQU5IPln/cb4ngNVWnXmXRSP3//8L+0A/42zpuBjY2VybSH7L/kpD1/cxglGv1riOPE2EeL1XVzlxCtFEuYojIBWAFp8iw/NHFvnQleYRn8KcxeUb/rApcMwODBSxdQf2hugHWHK2OqaEHrn4dNdXxf+H9X2vrh0Pbkwse1ueKHTmuwYQmRDouy9wFgsHfuuaTDAWCwd+65pMMBYLB37rmkwgvU1+bAGMBpCyrRLE+RdXAscX4TrnOQUMH+LEnvKnQASWqOwp1sS2ReUb/rApcMwoHtwGCLmljUoXuUx/fL+HeDnDvG6Gh33kFJljPsN9ts8wJyTa2Oe6+LCHDRBA7JhTyyhTOlsc8N3eyRu+y5XFQQ+awKSpLnEyPpm/aCFLcxwPW62iGZ5U8BYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwM6F/5GPXphNH2p000eSgTz2kveNzFTWGwFgsHfuuaTDqKfJtv+Q6dsMOagnZakaQvIloYzi3xYxFxUH3xE4WlRhrvt/y+YAdodQ61vbxLBOJ18ZhYU9M2ksDIE38PTknKbmMuXjGRlDpkJ8iU9obMIc19A5g5jGXTOBPw9xnBRDpkJ8iU9obMD77SfHGUr2QwFgsHfuuaTCMDyTn8Fu0HjA9JLXCx+0qqDXxlkXGyt8Gyt0UhGgaUzkg+Wf9xviezUX1vwI14aYZyRFYldliQZk94xfa4QpjwL0H/VOP3IWMqGLRaexoCud5BARb0+1FmmnWQQFp+n51oPI+kxv529YECjH0+TckRXnAqM6EL/uJvNcwrG43Q8BYLB37rmkwwFgsHfuuaTDAWCwd+65pMD4MYUc/RHM1GZJOpVn06og6iAskkn/YSsYJRr9a4jjxNA9unhEzZJhJnmz4KwcZ/jQPU4ruUfy7kcehumNwmTU8wJyTa2Oe6y06ltSttjJoPPMO1YhK5PqomqPWUuRPldytATF+ZYvDQsq0SxPkXVxGB9EArYhg6S+h8/+3fDf6NWXTWSR9he6RjGUlDW9J9EBtUrMA9/6hzbosYT6INWDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMKHUOtb28SwTidfGYWFPTNoLK7y92zrZZYL1NfmwBjAaQsq0SxPkXVwSUYV8VAVlKx46uWwrHngJFomJOyXCxdkZbTSxA+GPYTOhf+Rj16YTR9qdNNHkoE8/fVjt4b4+UvFyUWHJsVl1huGB4EQ2mQt4plZLtn54pLwwAh8cTZElwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTAGyt0UhGgaUzkg+Wf9xvieTEPGIHKmNtGoNfGWRcbK30asS5s0ZU2JqABxiMA7tjS7KDkxR4EMUiFSL396+9SJgkUsdCB0GeLAWCwd+65pMOiPvJJ+NIbiaTDIcH+vkJUykFBdRlxZweGYAskJ+MSZPMCck2tjnuvxbfaN/VjmA/jupxcsQCulodQ61vbxLBOJ18ZhYU9M2lzPw1/cCJZMs2gh8uecdEm0KI67NX8sDhhrvt/y+YAdWgyYneqoRKLnZfjdr8eWA8BYLB37rmkwz95BZ7YqC7lCyrRLE+RdXBJRhXxUBWUrjsrC2bolm4m2LvgKmInRkzkg+Wf9xvieANMisYrSaCpGfJRfHgOL1zA9JLXCx+0qqDXxlkXGyt/YQMsg2YSFRV2AmpsGeZs/RMYRhORWz638Ug8BLyqKN82A6h2vJKXxQOLYBBrowD6LB3MAU+nGqUyEDGhlCheCwFgsHfuuaTDAWCwd+65pMNqo0Ae5JUh+RXnAqM6EL/sFEBYxyXz1YPz1a6e87zLTMI3DWUUS8YSu/IZ0pdubmvCm+DhBNHfx7hvpiF9PRvTyPGvPnkDfx8jXTyvILzO2WBdYkXdJQ9jyIAb/6P9JEjm4esGHzrSvZcTyRApedXh49/7CPZG1+Kg18ZZFxsrf6omUlvf51h2t7POW0dfaMT/VJTEmSSzWPlbuxWje9MW6NMakaRBDLMu9jmdGv5feGGu+3/L5gB3ZBliDJCuKeP2CrOx6AZNuOYahnWFEIlx19gRVcWBVwa3s85bR19oxfNl5SS+okjxEiguf16CD8EkzR4dI11lEtHU+MvysWv5s8jOyjwnVpBySiUbXia6OqaB7yhk1J4BC9k6h5Y71X5TK09xkZJv1Zdg9HJi/Q9XhhQd5G/Xq5OYiqiWWtCZqkqBrVh6zEKDG13tPUhWWZKfiqBihguvhXeyjv/uIXXsu6l9D6gyxUcBYLB37rmkwDB2TZHWspj1JqWNRDiSJdPEN2j16ExUt2XeX8ktiuY8Ya77f8vmAHb23f9HiueSywFgsHfuuaTAuxPUN2+8SQg2WXzfm1gjjbVY5+BLn0ZXkZZKVsZGPZDBPsFxd3p2GwFgsHfuuaTBgrcIThxdfF53j9Df7gZDz4SEjjhM6QQJQ4zJDkwRGqJDRDzKAm9d6EPQTFGz2CFvS7BO0G2nPRETe3KALTTmkhdVrmRXNhfYOP4w+tHXso6oJPrd1Rgqz5UaCTKMoCzQh+y/5KQ9f3MYJRr9a4jjxXRJiKZ4+jS71girRWgAdKWPuNpNzh/xkQsq0SxPkXVxGB9EArYhg6Qwrr1D1wJHY4cMmgMS30D0Ya77f8vmAHaHUOtb28SwTidfGYWFPTNpXltGWD4p/POI0EhXVLVmzjKhi0WnsaAooin71hOwjh7Om4GNjZXJtIfsv+SkPX9zGCUa/WuI48faE8A6S0ZZo9YIq0VoAHSlj7jaTc4f8ZELKtEsT5F1cRgfRAK2IYOn0kXct+otyDuHDJoDEt9A9GGu+3/L5gB2h1DrW9vEsE4nXxmFhT0zaTLKvmTiOgv+3BrWU01tJZvxSDwEvKoo3xglGv1riOPE0D26eETNkmDjgq5bS0R06bUXfYiX6zhS9qwVKBkKzMON2FWO++CkhYWaM3bdub3AzUgudAoIV8+aMqCF3iWxbPs1XzEObJXP1h2+Z+wg/MUynDVY9Smyv8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLfc9CSVHsOFPheU73Klzgb9JsavxjE8f2s4yHKOV+vAh437qMTokd4LHnvN3f51aJEuxPUN2+8SQqr3neLkrrD6OiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHJR/tlyZ6V5A6A+HhePZxTkn2tbnjiZkgG3rM51h07VHlkeW9vGFC/iWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFlyy7PpeE6MgOhOQdnuEaIsM2ev42Ezam8FY5PTEMo3z5OT24kS10JBx7sPzAhhk/bilcidqhM5mEW+PLWHJwcdsoKmVcgLNIxSykisypGmm3zrogeifzvRR8jRLnCqHAbsCUIkFv5qe3PHrYr99U5d+ZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4hMY7OSSvyJ22N71FU5195hWOT0xDKN8+Tk9uJEtdCQce7D8wIYZP263OQSZ56IRu1vjy1hycHHbKCplXICzSMUspIrMqRppt866IHon870UfI0S5wqhwG7AlCJBb+ant4GMXMmDet/smWM7sg7m9pItp3y7fmTZdcVSVVRNYpozshsyfOCZT+LQGI+luyLZumDkt/4rqvxDVjk9MQyjfPk5PbiRLXQkHHuw/MCGGT9uPo25JUioSDJb48tYcnBx2ygqZVyAs0jFLKSKzKkaabfOuiB6J/O9FHyNEucKocBuLsT1DdvvEkKiRgj03pBs15ljO7IO5vaSLad8u35k2XXFUlVUTWKaM4uF5rQDhiQ11IybwRAazvML1TEereSyJuJwLZK3pRcbsZObORxDgNDMB79ko66rEToalT2jA9ioCQ2AdkZql9BwfFE3jEDu6x+Xvs0mPLDR6dGM3GzqJngwHeFlQlDk6Qwdk2R1rKY9IRDs3+pJdXmjwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+zsi8kDgweUqWel5v1mcFYLrh9/sx4J4ZcNuo+KvlQHfBxuLSKOWBKb/Teo4jMnl3Ty/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR2pu4hMG3CBrDXz/9QgbnfFKhsSCkbvUz3C6TA2VzpP6H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Ld4IyBLZpBiVJ/yVU3ZlmB+jEIUzLcAFCu3L1ItaP0xqENUeFFIS2pdJ1GxjPklkEyea9cc3w1wpQvkfclH6CdBm/GHvZjoUD5U+fKgA4J2sm2utZi+wc2dqpZSkKI9QQlLgB9YwaOIMsulkJz9NFOhtweqD1MqXb9n+UYSQNlGadnWUc0rmwGbEh4ZYMZnP+J8INnicMgBu/nfIMm83p+HzHdP6daf35EzYWBrk4CmlNmcjidK2GUszmkN4NvJP45rBaSix9SEwMZWQ/t+vjg24S7MtAeUHgua9hF2AWlHqMjXUlPGluXsHdA6JnAJKc4JppTCIZXB2xAc0k8FOSJeOJzN1aWbkWul13NcfrtCt6CFTH9NElHHLKVEcAzrpp14gOZlIYAvylVI5U9r6HGuzaskJ0t8DF4Y14cu4wOOWOFXZPAKpZADnkspgM9yDOLWdTihq5fNsUfyNj3fdwuL0LKP82o7u7JyuEjckbVktW5TwB2gV6RRNJu74PkAwaW3cu57R+r0QAyrlX0gor6kt07wCLvaFL0sjHjPOUb0zcUECgwZXCjE1yGHQHFsp1jMdMjFP6oCH0KWvjiqZu2f4QQY2ggkjI+4Thz2RZWraXcjdROOYkivQpa+OKpm7Zu3wi7RwaKz2XPav8BEGLU3YAdZrAqa9Mwg+SFO4YWYS4sHs5YKNom+QJ2hHn9a8aVS7MXWCJPL8lG/wQo8u2TW+pbmcnCDUJaRJEXOL5s/3my8G10yS4nHEx4kZVvK4LPmzJjv0jbyHoEixDSOaunbw8yrBlALsZk/l92SRuPTl836aGJ6c8Fb/5eWNM29TOkggVfaYiee2LGLbTW5DQLQ9f5MSqbLD8CMnlLxQHHMfA9nJ+iH6Y1aG92mvSKuyJRPASFTGAlbGHJE0BCHjrbBmxANNNUZAyw+X/Plo19sJ5Tb+spHGP86Optg1IoOK/UAnTvq7uXQhPh+vqqcWlNP2r8TIH2uO0kn3sgcdrMwsNz4rRwjBiQZE14vDqwgyyR6R2Io1Apt6iQ6J/V1vTdYgGMQTaPjz4XKMWHy5Xllwm2utZi+wc2RRPYn3R5zTRnGuANZTsWW6wKiLOWMEK+Rph5S9PiMfC+R9U44PrDq7mlwjuN09KXnMTnspNe37kjDz18Ia764Xp3v9OgOxUf8gX+lOdzu8wQW6A1k/HcyM0PjlidWHKnzdCSRiEUsATFKZjcaqZgVuRWJoAkfDaqblrCFXfVz7+ZNChmFOPz7M81+yMnQp2Nyo5ozFHJQV3+4yNGfFXJqycFmUMNY9FzR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/X0mFXQGDwUBfxxgLW/DpkietI52dApanS0ZwazF+DSia1Dv3sAhvWmfnNRqgv4UiYRGFaybmRCQWc02j3u+2kOy44C5ZqFQCn5vz96kpWbarmDIzkr822b6s8qwQE970EPDmeXSehv1knBXlhDPOgjbPf3JibGS9KAiuTcO6Px1knBXlhDPOidKCAKe7ioPLBQFOQvZ3yiVjW1fM47WbtJi8mo3u4XzqNUbehcOlfX6pOtkR5QI7rnkyOhxNuHYvuKiazyQ07CygDEbahTo5m18mOKd8EkIcL8CR+13B7XkmbmMQAYscojA4Ul7SfdWts7gbstDN5asFAU5C9nfKKmCrQtaJvfTpSneC5GunO6sZObORxDgNCTgqIdp7VhNdJCZTW10xy+0kpBS5r4LY4+/8gGLek9mp3E3uavtjBHa6sMkM+revdIECM44M6zSyTns76LF6di+5w6DyHzunJHqlF7ubtva1h5E0gkpomTYDx0oL8iJkpmAmFR3LKaecIKQH9xapKWm5wIy7VEbo3tIPi8/JGwoF4JAwcpRs2wpWqh0Oh2IWULQ66nxKXucTrs7IZ1ypQh3Jw9PGjYEhWUzsVX+qjJ2cFhRLHtr5z2lMrT3GRkm/U3VEkFOPxs0V4JAwcpRs2wpWqh0Oh2IWUcyI5pET4IalzGchwav//MHqUIOpiz3xD4GKLMDrjCPkWFOUwRSz7Ap3F2/KZDZS25G6XRReeG2It9mDkl+tWoKNKs5jPsTZHsY21T3uRMTZ+gA4ucyggfPwGopGN5FQ7sSi8p14YFtKqQD3q+pGjRHEcuJ+RvSwZzysUlAo8iA2xHoMmoJRXKqOnyOzoOHz81Zicz6VVMhCgnI8G7oo/IVFYclhD8d4eVd4cjsjZBW+zpQddyRRcRHdtxg6oOGCPveW98boqideHDJoDEt9A9akY/FF8AzWhRx8k0NEWRjFCCcmaBVJKejfuoxOiR3guycuDfKaqf+rkOsWPaq9s573lvfG6KonXhwyaAxLfQPfj10qKusZM2nA6cAXe2AmJCFBodbJdoT6qQD3q+pGjRHEcuJ+RvSwZzysUlAo8iA437qMTokd4LG3ox6OkpsUe5DrFj2qvbOe95b3xuiqJ14cMmgMS30D349dKirrGTNmepWlV3h5bLQhQaHWyXaE+qkA96vqRo0RxHLifkb0sGhWOg6iIp1UbuDmirbUrVEvcp/eEZRPWUoA1fRcFMeMBv1BljVnPz/q4Ga14AP/SQcyP8LAktKTHyA8Y33xR/3r3/3eZnZNH02VAHAPePKsOCEmw+NwTtK9Bmk/RnodzdrZ+y1R+IOdIAKmSo8Nxy/ZGV/HFcSs5eZdsjXDviZ5w0g+b0azBmc8Mqoq3XbdxqWfoJvbUlc1mP3CT8+Dul5Yk9A6Vhmag7l0eY3Tq5s88KvCL+HSA6aIE+jOBsGK0KE/34Z3y6pISUytPcZGSb9TdUSQU4/GzRQW6A1k/HcyPsvccCkeJVeV4ruVEFfBRDaUCqUsoSsGlJ25ku1+CC14tJFi57rHJCCa1xN53e85ZtRd9iJfrOFG+wihoEHfiJyTlMu5OxK3HCCD8Qa/jQUOZW32EHlUV1wuDhMsVKUw/nSv/rNmDxCcCUIkFv5qe3o6Fxp5dO7pUpim5dgZrhdGvQikJWPE7CK+TC2YUt5PaH/7UNU58jTvHeW8nb43dkFLE6gy+KXP1YggAh2zYxKvJMoiRRwIwdnjTu2O+dB5RcDU+ErvoJgItJFi57rHJCCa1xN53e85ZtRd9iJfrOFG+wihoEHfiJJ+K7bVNLNKjX5NnXYXS47aP33I5QEiCsHEcuJ+RvSwaFVSD1FKcXtE9CnTVxY3vYPwGopGN5FQ4lmrhao9NqsZ64K/wQvn7OD3Vtl8iFR/xUVhyWEPx3h0FugNZPx3Mjd/LzmrCWut7V3amXOXEZSrgzMGFy6BD4Hmu720KXEVwNu9GXfU3btedK/+s2YPEJodQ61vbxLBOJ18ZhYU9M2rJ2lf7LOhOaqpAPer6kaNEcRy4n5G9LBoVVIPUUpxe0xvZrfAFJ45w8wJyTa2Oe6zP9pETYL18Po6Fxp5dO7pUYGXhDpCZo02vQikJWPE7CK+TC2YUt5PYaBqWUz3QgT4yoYtFp7GgKht7ZsYjD8fR7td2RznPfJEYLxxdtWkL34cMmgMS30D0UiOnUM637Jz3hEYkg78NmOSD5Z/3G+J6LOzTU/SEynItJFi57rHJCAnGtjK+v0BVtRd9iJfrOFKcnp15/O3TdQsq0SxPkXVwxZZG42AAG+GaYQhqPazlY3rZtq8XFOj3sY21T3uRMTZxqJIHSnBRTyeCHG2BJ/93GCUa/WuI48TO5hFXrrKRowgg/EGv40FDOq35Y6l2k/8Lg4TLFSlMP50r/6zZg8Qmh1DrW9vEsE4nXxmFhT0zadG53MZeqtq24MzBhcugQ+ObV9EPoBEz3VFYclhD8d4dBboDWT8dzIzOhf+Rj16YTR9qdNNHkoE/sU2Z71Tky1t9NOFo/gkIUWIIAIds2MSryTKIkUcCMHe7RX6e0WZRBF5Rv+sClwzD5y+9P+EBA6JKHozjh0OSjQuZhsD7PaVLhwyaAxLfQPRSI6dQzrfsnPeERiSDvw2Y5IPln/cb4nnB0sKTpK3byxMUzSIq7Wq7H8YPSoAnQYMLg4TLFSlMP50r/6zZg8Qmh1DrW9vEsE4nXxmFhT0zafW1pqfczPjk4LDrX5pCNrxxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnDzAnJNrY57rLTqW1K22MmjPpffILJP9yx7wLlbrB15Ha9CKQlY8TsIr5MLZhS3k9hoGpZTPdCBPjKhi0WnsaAreJqV/niaV7DVmJzPpVUyEKr+CAO2uy01UVhyWEPx3h0FugNZPx3MjM6F/5GPXphNH2p000eSgT9B/ek/RaITV9Dyfl9n8vc/1girRWgAdKW1F32Il+s4UpyenXn87dN1CyrRLE+RdXAscX4TrnOQUDysPxsmjpWg+youHJ0sXU+xjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3cYJRr9a4jjxd+M3Bws3M3nCCD8Qa/jQULe+KiDarvwvwuDhMsVKUw/nSv/rNmDxCaHUOtb28SwTidfGYWFPTNrvpVQOQUqSLnSAJKXVVxU9HEcuJ+RvSwaFVSD1FKcXtMb2a3wBSeOcPMCck2tjnuviwhw0QQOyYZ1/qcGxeC8OKYpuXYGa4XRr0IpCVjxOwivkwtmFLeT2GgallM90IE+MqGLRaexoCoXgkpKH6TlpNWYnM+lVTISepapIUmNOAVRWHJYQ/HeHQW6A1k/HcyMzoX/kY9emE0fanTTR5KBPnZO/8FBOclChOq9sRsET/liCACHbNjEq8kyiJFHAjB3u0V+ntFmUQReUb/rApcMwXFoKZw2tfBOSh6M44dDko22EMoS8Ahib4cMmgMS30D0UiOnUM637J2LT9QW2XVLTXYCamwZ5mz9dOs0IYu1Ci6P33I5QEiCsgcZdMvisFLttRd9iJfrOFKcnp15/O3TdObh6wYfOtK8sDFMPqFVMSqCOx34HjCVgG89wpqN26FXsY21T3uRMTZxqJIHSnBRTyeCHG2BJ/93NgOodrySl8YKNuRJmdBRXwgg/EGv40FC5GHdCVV7wTsLg4TLFSlMP50r/6zZg8QkLmLkS6L2UIQup2fdyAurZSxfzUhAFD7dS0pd/SoDbqxxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnP2CrOx6AZNuOdM3OLYTtuZLmWUJ+KmPVSmKbl2BmuF0a9CKQlY8TsIr5MLZhS3k9kRiH30xEL5PubMUiPEHCqdhujk21+NMk3u13ZHOc98kRgvHF21aQvfhwyaAxLfQPRSI6dQzrfsn3b+3M0b5yi+vux6JMIhErRSxOoMvilz9WIIAIds2MSryTKIkUcCMHWlAqlLKErBpGl6aGdzskH41Zicz6VVMhCgnI8G7oo/IVFYclhD8d4dBboDWT8dzIwwdk2R1rKY9o6Fxp5dO7pUpim5dgZrhdGvQikJWPE7CK+TC2YUt5Pb9rNQ9pMjFp9Ijj35PgicaqpAPer6kaNEcRy4n5G9LBsjzVMb2Werg+VqsHKyV31Sht71Lx03BVTDDPOxma7izDoB9whnnmD7ZDNSSn5ftIfhaLaESChLI7bBBw/qXKbomgIOXbwqvbemQnyJT2hswXa47ZGoVCtPFX/ozmn9HsBMVqPovgrpw4/7CDGWMONIBLmdLVRh/xFvVIAgx1sm4aDcb8kPEFtZTA+jtY2bE9m3gjXOEok0StlY9qxRdVGrRKV9HBqAm1LSR3mCRd2pm54NARHvgdqrC5B7hjBvB1ges1r3OeJy5x7oTl03mhREEEyoZAjAoDNEUaFVzusiyCg082Ol+YzQ6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcu+ViV8SzXCDVq4lp3Q3E4tgoGYRI7CS9JdDD6unk4J+tP/8iyWTRROXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZq7yBPxzHmKG2W/fuVNNz/ImEqpsA+sej/xScREvltrsHDZMRgFfe1OrGISi5pGmyy8V8b58GG7aywKTkKJerd+XIk1JlZdjcvlb6sRvxeiu4SSlnUTC2QgxnN5zg1hvpj7jts9D9Vf69qoHINnqNTQT1zWClEYtH4XLjiOTjsUyMZzec4NYb6YDRpGjFGzDGiVfbovfMR6DMMIMVCYg7BmoNfGWRcbK30qiFeKDhAZk9qoHINnqNTQT1zWClEYtH4XLjiOTjsUyMZzec4NYb6YO7nzba2P/xyVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3wKlnV9VTt8z9qoHINnqNTQT1zWClEYtH4XLjiOTjsUy9xovJ2mxAzRLvnX2Duhfj3UWKJQ6R9GzprfkM6pnQKu/EUKWXiWm56g18ZZFxsrff600u7C6i61wMz/WqplQkXyA/Cw3lzwqR8iPFqfBHPU67OyGdcqUISYj5WNFHWMZcQr3mv20Raxi7mYxX0WepLFItsraew8YU4sSWeE4EReWnABkhfYwG9iuoTHUj00c/1U4QQ+VIc8n4rttU0s0qE1T/XKuGrakQIaAy+tSTHE37Nk97b+6rhhrvt/y+YAdvbd/0eK55LLAWCwd+65pMMCUIkFv5qe3lfxdCVK0plLAlCJBb+ant0quPrqKexhDfituwZjT2jy9qwVKBkKzMF1o37kFIzi3RIoLn9egg/DX8AjISKtMcDhszRjqw8t8fSMyXoLumZf8DWxmzGd+ycBYLB37rmkwkZH2/nXjRmPRhWLP1OR+C4hOdYUHwfkX4SSlnUTC2QjAWCwd+65pMJ5R1LlXox2Zax/eKhbB3Vxw7Ea2f5QtARhrvt/y+YAdN+plWTQJSyz/dmxyum6USj8BqKRjeRUOfituwZjT2jyhKlCAG3SxEhJrdWXyxuQTjK6BxsmUurV/NShQVMzpIcBYLB37rmkwwJQiQW/mp7f4O43a0O1PgooJ2edU1i1iqDXxlkXGyt/WLm3eKt4OT8BYLB37rmkw1uhkf50lBKRJ6shrRPWUp8smgqJhmepjGGu+3/L5gB036mVZNAlLLH3vzCCnNr0Tntym+tHv+zaoNfGWRcbK3zGc3nODWG+mDu5822tj/8cCpZ1fVU7fM5DRDzKAm9d6kqBrVh6zEKD+ePzjN8nMzbtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXehD0ExRs9ghbdwwqZv6zyy5qORwzQdMkxQRM5a3QoG6cNv1C5IcM1159+qWmlydBZquwSwszM3a5nb5JfkbWY532vCk8ezaIWDokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyHh5H/kQeq4iz8hPZk9AeGZ3eQ9NTAuFhcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJN9Y9kCMWWVDNumJ9zDsK75UygcE7sJiDRwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk6P7+01uBmdkjA+OnBq18uLGfZ/DmqPyQ4V/WU3qpupr7Z36IFzy/QUfILcYi00x4udtI/0UeRgdZFdkSnhQ3bdyErauFowuZk/kMqEp6+Cp4YUHeRv16uTmIqollrQmalRDmotZ4t7jhdVrmRXNhfbAWCwd+65pMPaqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+qDXxlkXGyt8Gyt0UhGgaUzkg+Wf9xvie1egUu5QhWYY0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4SWqOwp1sS2ReUb/rApcMwDsxqtrovVL77GXgsW1V6zlEJZt5I6hoN5iRnMMMFpPvAWCwd+65pMDOhf+Rj16YTR9qdNNHkoE8xGTLgbXI8yLtwcZyZxxotq7z0WNseUXcT1zWClEYtH44v3PQhoFfMgvU1+bAGMBpCyrRLE+RdXAscX4TrnOQUb/I6UoKRFdclX26L3zEegzDCDFQmIOwZqDXxlkXGyt8Gyt0UhGgaUzkg+Wf9xvieWz3mwEfg7VA0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4SWqOwp1sS2ReUb/rApcMwLCwdyEXs6eH7GXgsW1V6zlEJZt5I6hoN5iRnMMMFpPvAWCwd+65pMDOhf+Rj16YTR9qdNNHkoE+bLLtHm+76nLtwcZyZxxotq7z0WNseUXcT1zWClEYtH44v3PQhoFfMgvU1+bAGMBpCyrRLE+RdXAscX4TrnOQUkYsqZrpSXE4lX26L3zEegzDCDFQmIOwZqDXxlkXGyt8Gyt0UhGgaUzkg+Wf9xvieUoKi1H45w/80nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4SWqOwp1sS2ReUb/rApcMwODBSxdQf2hv7GXgsW1V6zlEJZt5I6hoNu3BxnJnHGi23U4tcd5nCGLOm4GNjZXJtIfsv+SkPX9zGCUa/WuI48R8LWQELRpWbbUxOJCASXORs/P9zr8kn/aI9EAkCE4YegvU1+bAGMBpCyrRLE+RdXDFlkbjYAAb4sSXlKLXP5nMlX26L3zEegzDCDFQmIOwZqDXxlkXGyt8Gyt0UhGgaUzkg+Wf9xvieJfByYW755XQ0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4SWqOwp1sS2ReUb/rApcMwEgHSg9yWcm/7GXgsW1V6zlEJZt5I6hoNu3BxnJnHGi23U4tcd5nCGLOm4GNjZXJtIfsv+SkPX9zGCUa/WuI48XkGSt8JC63kbUxOJCASXORs/P9zr8kn/aI9EAkCE4YegvU1+bAGMBpCyrRLE+RdXDFlkbjYAAb4EJ2rxLtgwXIlX26L3zEegzDCDFQmIOwZqDXxlkXGyt8Gyt0UhGgaUzkg+Wf9xviehZQQlQxCupw0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4SWqOwp1sS2ReUb/rApcMwbIHmXIEV1WP7GXgsW1V6zlEJZt5I6hoN5iRnMMMFpPvAWCwd+65pMDOhf+Rj16YTR9qdNNHkoE9WXK3mq1uYgrtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXemtVq1ERu/fojKhi0WnsaApG6GuwlF4/tPaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMpHHobpjcJk1PMCck2tjnuvxbfaN/VjmAy/J0M+XsjWoQIaAy+tSTHE37Nk97b+6rhhrvt/y+YAdWgyYneqoRKK3dfjuuFuzwzKQUF1GXFnBNDrz/dM09R4aYzfjTC6+kbOm4GNjZXJtIfsv+SkPX9zNgOodrySl8V/uXe8whxDrbUxOJCASXORs/P9zr8kn/aI9EAkCE4YegvU1+bAGMBo5uHrBh860r2XE8kQKXnV4EJ2rxLtgwXIlX26L3zEegzDCDFQmIOwZqDXxlkXGyt/H9CKzhSnTcSPDijaF77o+wFgsHfuuaTA0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek7GagbKFwYaK03ZQFk6iz04rPpCrRID6Nv7GXgsW1V6zlEJZt5I6hoN5iRnMMMFpPvAWCwd+65pMAwdk2R1rKY9xP174gDGwo8etIGIxNDE2btwcZyZxxott1OLXHeZwhiQ0Q8ygJvXeiIQWBwpLzSMb9SjuyaHp2TAWCwd+65pMPaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMqEqUIAbdLESImsZrxj6swPAWCwd+65pMIL4r2VJ/f/JQIaAy+tSTHE37Nk97b+6rhhrvt/y+YAdLsT1DdvvEkKspjmAQ+WM6zKQUF1GXFnBNDrz/dM09R4aYzfjTC6+kbOm4GNjZXJt1ltRIiC3WqEn4rttU0s0qMHKfGlhZjJmbUxOJCASXORs/P9zr8kn/aI9EAkCE4YeDCuNVCU7v0plzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZqR8iPFqfBHPU67OyGdcqUISYj5WNFHWMZcQr3mv20RaxEiguf16CD8FkZQfsOmazj0mYsgD7uX+0rJgj0vjeWlFRDmotZ4t7jhdVrmRXNhfan4qgYoYLr4V3so7/7iF17d/LzmrCWut4L142YVxSj9DafoqSRYJzvgjipf+V29wGEelDZxKY0tJQx43UyoUIdCVaiK2Kix+dEiguf16CD8Nq6gnw/xVmhZcjgIoSriUqYOYcdscO6cJQ3hIX2RJDecQKHQC7AFJeoNfGWRcbK3wbK3RSEaBpTOSD5Z/3G+J5lQGNtXQicj6x3W73WWWwNd/LzmrCWut5crRe/j/NFEHWVa4W6Yn4OwFgsHfuuaTDAWCwd+65pMMBYLB37rmkw1v73wpaYW/0wse1ueKHTmuwYQmRDouy9wFgsHfuuaTDAWCwd+65pMMBYLB37rmkw/1U4QQ+VIc/pkJ8iU9obMExCYiTvrzNes6bgY2Nlcm0h+y/5KQ9f3MYJRr9a4jjxD9RQIvAhGoyW4qSiO3qj3+DnDvG6Gh33kFJljPsN9ts8wJyTa2Oe6+LCHDRBA7Jhe4AEvgqHKXIt1hWhhI8E4tDsxVBsgkPTMLHtbnih05rsGEJkQ6LsvRJao7CnWxLZF5Rv+sClwzDDaA7H8UVqT40AgtPQ4RQzwL0H/VOP3IWMqGLRaexoCmOH6UWvbqlfeseThdMUJvzAWCwd+65pMMBYLB37rmkwBD5rApKkucSDMC97q/CYU3A9braIZnlTwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTAzoX/kY9emE0fanTTR5KBPpi/QQ3QAU/GRx6G6Y3CZNTzAnJNrY57r8W32jf1Y5gP6mKU2THl66zOhf+Rj16YTR9qdNNHkoE9WRmc3I1j5WcBYLB37rmkwwFgsHfuuaTDAWCwd+65pMJGMZSUNb0n0QG1SswD3/qHNuixhPog1YMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwFJsutPhWnAUXlG/6wKXDMPnL70/4QEDo6Bk8CTARz3yoNfGWRcbK33Vv8dmQgalVsT40ok7+2lAl2EOZyiVQ+TU+PtULq1mZIfsv+SkPX9zGCUa/WuI48cP7JM61hW5CepLoJLvA5Fc7/6lGH2ZmzUoC1u7PX7hJYm+edmtI3b2OymG4mwLpAF3so7/7iF17DzcIhqGMLQZEiguf16CD8Ef9pOKEhUIqtCiOuzV/LA4Ya77f8vmAHaHUOtb28SwTidfGYWFPTNq7IDVYZOvF+Nf68pRp/VxRrsJDQ3CRiKjCMqUcdUEhBTkg+Wf9xvieBZZ8Z/Vi35iSWV0SSxDYDsBYLB37rmkwvcS0eTTSuAAwPSS1wsftKqg18ZZFxsrfwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwIfsv+SkPX9zGCUa/WuI48bqPTo1ovmtlqDXxlkXGyt+zpfNKPqguCMYJRr9a4jjxu3QvpD8Laur8Ug8BLyqKN8YJRr9a4jjxx2nul6v+n4niaLXwDYlDoHq74vYNDVBSSBljzD6HSXpE3tygC005pDOhf+Rj16YTR9qdNNHkoE/4MOc6UfiqaTOhf+Rj16YTR9qdNNHkoE+vTb/K3ch6oFSBZIgI35Rgbs37l3tbKUHj5RcgwgjQhQ8PxmQ971X954R8ww9UdCf8CyejKSfcq9MOEg5Kmw8L6F+0TU7SlHNrVatREbv36IyoYtFp7GgKZOFmhAL8IsJy+5nx1JzUfFG71n0QjkmsQVJx+DTr+3Jrvxpl2yBkDg9kl0t7I5W6SgLW7s9fuElzWp6/L+DmbkTe3KALTTmkkDHd5DolrDG8MAIfHE2RJcBYLB37rmkwM6F/5GPXphNH2p000eSgT7SNbHLYVtHtUHk7KWmEpPux7Lu2DuBUvMQB+NFEmBdPidfGYWFPTNrKl0ASdoesmH9s7v6Rh/xlNg1uyzYlp0HCtytBf/n+KbQojrs1fywOGGu+3/L5gB3AWCwd+65pMMBYLB37rmkwwFgsHfuuaTBrVatREbv36IyoYtFp7GgKZOFmhAL8IsKzpuBjY2VybSH7L/kpD1/cxglGv1riOPHZPbL0NbZsyStFEuYojIBWAFp8iw/NHFvnQleYRn8KcxeUb/rApcMwXa8Y4UXPCP1cFoDmkkq8WlVSrfydKQA2ZfrJxuQcP1gwse1ueKHTmuwYQmRDouy9wFgsHfuuaTDAWCwd+65pMMBYLB37rmkwgvU1+bAGMBpCyrRLE+RdXAscX4TrnOQU4f8pwwKG1T0SWqOwp1sS2ReUb/rApcMwLCwdyEXs6eEoXuUx/fL+HeDnDvG6Gh33kFJljPsN9ts8wJyTa2Oe6+LCHDRBA7JhlHhcsLe8CONCFshD+MKNkAQ+awKSpLnE8DfdRW84p5VwPW62iGZ5U8BYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwM6F/5GPXphNH2p000eSgTzR2a+mV9uguwFgsHfuuaTDMmLAuFeHUq9IWZyRNlzQG8O9daMoxy/IczBNUAZSJKZHHobpjcJk1PMCck2tjnuviwhw0QQOyYXE06YPwylW4BMNlvUmHSdCJ18ZhYU9M2j6/8VZz3SBibKe1RCES7zuxzJK/X7Yn+EWDREuSGLipwFgsHfuuaTBqE1QcA6aRlEV5wKjOhC/7ibzXMKxuN0NrVatREbv36IyoYtFp7GgKnSun8r5JRK1eMUppIQnshhmSTqVZ9OqIOogLJJJ/2ErGCUa/WuI48dZxaMp1DURtSurNT19gaRz1hRx9HzAnCjZEuQmNlq1ZvRzyiucKSmrAY9hMEVNowcBYLB37rmkwwFgsHfuuaTDAWCwd+65pMLfxIr8u7o7LAFp8iw/NHFvnQleYRn8KcxeUb/rApcMwJC9RKyns6UGmuXXfCLpGAl3UkXiCZPwNgvU1+bAGMBpCyrRLE+RdXDFlkbjYAAb4I7qjzGYNMwoWiYk7JcLF2RltNLED4Y9hM6F/5GPXphNH2p000eSgTy/rbOln0OJc6oGRy8U0dYRbmdcWHQPF4D2uRqRD9lfGvDACHxxNkSXAWCwd+65pMMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMAbK3RSEaBpTOSD5Z/3G+J558aUJngmAnMBYLB37rmkwbxpmWL2ekaY5IPln/cb4npEoeNptTdpDZ7FOTMMrTg45IPln/cb4nts7r/SbThDaanQGWqvtUu8pngetTA68p0gidVlk9IH4RN7coAtNOaRka1OHephHjOz4Fc2e0X1d2+1kpzkJkZrF4Z9KOnTL5Rhrvt/y+YAdodQ61vbxLBOJ18ZhYU9M2pOpaizKHemRKbmMuXjGRlDpkJ8iU9obMJBs9CVRsYQLovwwPQ17bBN38vOasJa63lytF7+P80UQ/AnPdtIKD2YNJ3jH8EHgV8j6Zv2ghS3McD1utohmeVORx6G6Y3CZNTzAnJNrY57rM/2kRNgvXw+e3ckpOSqm3qiao9ZS5E+V3K0BMX5li8NCyrRLE+RdXEYH0QCtiGDp1wKB4iWa1CqSWV0SSxDYDpGMZSUNb0n0tO6P2Jsu6kjNuixhPog1YMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwFomJOyXCxdkZbTSxA+GPYTOhf+Rj16YTR9qdNNHkoE/qKr/0LvHA/NWDsvwNdcAuqDXxlkXGyt8Gyt0UhGgaUzkg+Wf9xviek2PDFW7dGF0ZyRFYldliQZk94xfa4QpjwL0H/VOP3IWMqGLRaexoCooRJKV5vHKKWpyTSXtAQwWWJ1Pts9CKMz1NNttoK7+1RXnAqM6EL/uJvNcwrG43Q8BYLB37rmkwwFgsHfuuaTDAWCwd+65pMBJao7CnWxLZF5Rv+sClwzDWAdhLH9wLIJDRDzKAm9d6a1WrURG79+iMqGLRaexoCpZ1yBBP9kehXjFKaSEJ7IYZkk6lWfTqiDqICySSf9hKxglGv1riOPH2hPAOktGWaMY7xD5B4tMmVRb9ucwOXndYHcceC3bt8L0c8ornCkpqwGPYTBFTaMHAWCwd+65pMMBYLB37rmkwwFgsHfuuaTCRx6G6Y3CZNTzAnJNrY57rLTqW1K22MmgQooj+XTH/pUTe3KALTTmkq4axkiVew5pJsbxTgx2xTnOEdIhM+5oQ3mh+MdrdPHuC9TX5sAYwGkLKtEsT5F1cRgfRAK2IYOm3yRNRAF9ZhSLMSFB9p6vVscySv1+2J/ivLtwfF9+TzEzgT8PcZwUQ6ZCfIlPaGzD1avesNVM4IezC7kCnMi5Q1c4I1gKMyQm9HPKK5wpKasBj2EwRU2jBIfsv+SkPX9zGCUa/WuI48XkGSt8JC63kK0US5iiMgFYAWnyLD80cW+dCV5hGfwpzF5Rv+sClwzASAdKD3JZyb6a5dd8IukYCeHk1KFd3gKK4V1J5A3Af8TCx7W54odOa7BhCZEOi7L3AWCwd+65pMMBYLB37rmkwwFgsHfuuaTCRu3fB9AtaM+DnDvG6Gh33kFJljPsN9ts8wJyTa2Oe6+LCHDRBA7JhIDekynISIlI/jrHiIaKYbcBYLB37rmkwM6F/5GPXphNH2p000eSgT9qtlQbJK2NbUHk7KWmEpPux7Lu2DuBUvMQB+NFEmBdPidfGYWFPTNowcR8KHJN5hRDrDNdBi0vINg1uyzYlp0ERDlN1CrpgWbQojrs1fywOGGu+3/L5gB3AWCwd+65pMMBYLB37rmkwwFgsHfuuaTBrVatREbv36IyoYtFp7GgKhgRhdyfWkwUYa77f8vmAHaHUOtb28SwTidfGYWFPTNr3rUk9OI8MgNf68pRp/VxRrsJDQ3CRiKjCMqUcdUEhBTkg+Wf9xvie0YjX0B28Z1JvYc43mJDana0vB7aGVL+nWiGFct8+LIUwPSS1wsftKqg18ZZFxsrfwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwIfsv+SkPX9zGCUa/WuI48VyrraijZYOn4+UXIMII0IUfwldyFtbWW0DgKakAXNf0JstPjDBPaOCu9qLHVD0aFuBtSgGxG0pAqDXxlkXGyt/YQMsg2YSFRV2AmpsGeZs/8sWSENY3+22sd1u91llsDTOhf+Rj16YTR9qdNNHkoE+xCJDuu7SW7AgtNr+icS9ajKhi0WnsaAr7noL/O6vQyB1/Y1qVnlIzRXnAqM6EL/uJvNcwrG43Q5OYFEBJfSIYnJWN2CoNMljLnjvKRySunC+kiTE2ksC9xAH40USYF0+J18ZhYU9M2mWLzE26sPNtSk6Q9mKICGrGCUa/WuI48cj1GLDWfTcHYXFtq2LTFzG9HPKK5wpKasBj2EwRU2jBIfsv+SkPX9zNgOodrySl8YKNuRJmdBRXGkP0uvMTnYWLB3MAU+nGqQ352ruhypEw6I+8kn40huKBM78zXkGVC8BYLB37rmkwwFgsHfuuaTDlPU2piCym8zCx7W54odOajFIo0AQQWSREiguf16CD8CaMiRZuGXn4UHNt0Z0aS3WFxxUK63QlUdHgE6Z29mzTqWopDhWrLUWhG37csGjubujqSFmk3zYp5RwB2j+JUvV64c4tVCczmbd1+O64W7PDePC9WQS2+5+zpuBjY2VybQD16ny9fmk7uPNtE1N6OPVYjyLSXV5MUrSkkB3ZsLwyT6Eu2xBENNS8S4xcFwaTxgKB52gK4D7dkYxlJQ1vSfSZBQcV0y5PD9ZrtGVbf/q3wFgsHfuuaTDZW9Tc6xei2yRKXyckhTIizkyQmBmQ0jrzKeD8chZTSHqD0cdP7ibjB/0N7qXtgUuCFfgvXHzSEYhG4yiXNnPTiky4eUIJ2/h82XlJL6iSPIL1NfmwBjAaH7mUaPtluaoEA5MlnbvkHmBscT8ZbRQBqKAR8vN2ScAYa77f8vmAHYfTI81FpnVHJ+K7bVNLNKgZ5V+uIEEK7+EkpZ1EwtkIwFgsHfuuaTCI0PYO4nCkHmjBahxDGarMeujSh4bHHPcI9LbUH5bZsy7OEyCMGDLsmibMoEx3LXhXN19zG3yZ/cBYLB37rmkwYK3CE4cXXxeslEAzcwzIV+mQnyJT2hsw6EBIT5eD8Z+zpuBjY2VybaEqUIAbdLESq+yikjuA+Lqn4qgYoYLr4V3so7/7iF1705ppnroUMtDAWCwd+65pMGCtwhOHF18XcfY1xzdEc8bpkJ8iU9obMCi6SR3bv1/Bs6bgY2Nlcm2hKlCAG3SxEux6tfF0RwGJp+KoGKGC6+Fd7KO/+4hde9lexNhGeYmwwFgsHfuuaTDGkK0gp48bmD8BqKRjeRUOua6FTEyXtZM8aap62hUdQcBYLB37rmkwYK3CE4cXXxdJHC45IMqSTc5MkJgZkNI6fP1aoJraG7HAWCwd+65pMGCtwhOHF18XwBWjihVXPhnOTJCYGZDSOqX3WF2Y3rQ1wFgsHfuuaTBgrcIThxdfF4dIbzpDUcTwzkyQmBmQ0joK3NJesgeaM8BYLB37rmkwYK3CE4cXXxeh6gHmwahysnLF9nXsbQ9vbiZYGAQw3lOoNfGWRcbK32o5HDNB0yTFAoHnaArgPt3V6kmAJ4eDlixxeV5qTehQfzJ/5MKN2KyoKTJI3aJglCsmCPS+N5aUa1WrURG79+iMqGLRaexoCh1VaNo7Z/F6HEcuJ+RvSwbUjQSoiA5mQjzAnJNrY57r4sIcNEEDsmGnJ3lxfxKwZMLg4TLFSlMPwFgsHfuuaTAzoX/kY9emE0fanTTR5KBPHr7TzVVAUitnsU5MwytODjkg+Wf9xvieOr5FU+PPePGQ0Q8ygJvXemtVq1ERu/fojKhi0WnsaArGogDVmQ8JoRxHLifkb0sG1I0EqIgOZkI8wJyTa2Oe6+LCHDRBA7JhHSa25ZxUIyLC4OEyxUpTD8BYLB37rmkwM6F/5GPXphNH2p000eSgTx8XqBOH8J65IVAmq+H+WJbiNBIV1S1Zs4yoYtFp7GgK5ZvcISo7WdQcRy4n5G9LBnPKxSUCjyIDEPQTFGz2CFt3DCpm/rPLLq0yD9MfwDAwm7Cl/JGm4dRMzOo1oB5ATYcwxAzjdp4XoA1fRcFMeMBQbYN8kK6rh/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4Ull/LbH3nTjfuoxOiR3gtHoVpcdwyZrAwdk2R1rKY9Bslab2P8omcMHZNkdaymPR0/XhGDCcxKeppZo8RsuOzTmYJPsMg+Q6bFeBOZiXGcJsavxjE8f2u0vHvd+5v00/4ndrcguBFspnhPA16MAjVnqVpVd4eWy6xxATWFVpDn8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/FUFF0KLvkcR5ELwYuCrySacRvD4lXwsnO8H3QNHdsh00gEgh5rwTB4l2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZRpjNvcV01fPgH6mKA8iOZTzr/ZBmu0bBLB5ndRVGHnYcwxAzjdp4XoA1fRcFMeMBd/eezngX2H8owH89/P7+CsOW9w8BUFblrS1TXObGJTlOqZzn61y5rtlY9qxRdVGr6XH3k8uFaYyrNd65etilFWDiA6bJiA7/4aIi/A+pRzjGWibpKknJBy/BJV9UtiIl8aWSUg45QJwNTo9MmY6L+yXH6M6sq4/6CvRW48IRHZRI26MsU3OoLPQuqIONPkd2UTAApspO4z2XmK7xcbFXj52NFPl31wE3Vky97a5W3s6EM6PsRQw3r8DhOAb9OTiBDsZ+t3i1dSCd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+FQRTQg1Qz1D9aDJodEP4LuRq8whmI13Pvf/d5mdk0fTZUAcA948qw+ooThGF5bBxVnOhCGoXArhwEU0yBqKU7RmOYgTRnNP30iQ/6mZ9pEFTfNmEUmqMgcFqtQFTH7C9FkYtbPg8Yg+ZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4qvV8ZIoYFr4C9UxHq3ksibicC2St6UXG7GTmzkcQ4DQTM5VhMW6nM06GpU9owPYqAkNgHZGapfQcHxRN4xA7usfl77NJjyw0enRjNxs6iZ4MB3hZUJQ5OkCpZ1fVU7fM8fLpL/P9hSAPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuvmNJa65VppwBMloxPdDN7kLT9KQ3pbn9GhzDEDON2nhegDV9FwUx4wF3957OeBfYfRJvI/8fpSgqw5b3DwFQVuWtLVNc5sYlOU6pnOfrXLmu2Vj2rFF1UavpcfeTy4Vpjh90imrnfcKmH860fPQD/v/hoiL8D6lHOMZaJukqSckHL8ElX1S2IidvqxD2AqzaTGutIgRi3ZDX3A9iPSC2exowPjpwatfLik3woVAL15GWjg/EhHtVuttqqgvbqIhfPpH+iYXN2p5ZQyvkqv1zB7Ah8gkp9XXDmoi1Hn//j9/BCkjmt314ynziILP11PrKfD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDwSZka4SgeV+cDpwBd7YCYgvVMR6t5LIm4nAtkrelFxuxk5s5HEOA0EzOVYTFupzN3dNMSYyqYosJDYB2RmqX0HB8UTeMQO7rH5e+zSY8sNHp0YzcbOomeDAd4WVCUOTpDB2TZHWspj2EsIoIFO5TJj7fBSngAeVpmkFWFrOe10MVdf0sP8GLr3nOzk9EhQmWXbkwgwVzovW4ugDXg6fOP5Jm5jEAGLHKIwOFJe0n3VqlfgKZxfTm7DgGxpVeYde9LEXGmfgOzLPKX3++GkmMpJx2QQ8NPRzdWn1fZW0i5InteD0WCGyQkm/2NXYf/YzeQZl+0QKwT4iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUgvhzZ/roxehwzLic26TZGFv6uQ1bQ+V1P5g+3VUkwsBNEUaFVzusiycCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPavvlersphWFrgSNBvfq0O8iUoVEULW/wAyrlX0gor6h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC5phREvPgpvHBpIYeA2rj5kBghSAkob+RtcYPplyneb5FgMEVi6IXblsFshSxqvZfeXR15LUBDW8Q9t/s4jiy19tVJMf5fqF0qOH/tgCkP0SSPXFdmWcYdt4ARkxInittcjDCGziKbjMv35wrSemaxXEncUfC4oj29m0sv7LJtanH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LvOELWtFYaJAxkL91+oXh1AAHKLhj4L3RjWp4X/fEthWNsdqxvyc0pvvhO+I7b9wou5ATpgb+4aq6ErXIdZ7wR5yW6ej+suMWMlqR6Ss0rWpS39lrM0Fjh+0bWTRss2SZ7boMQ9kCHfld5S7zHloRbUxnruitJTU5fo7z4kSyXGiUjiULvKTmuR2NmUzZZGl6r2nM1TdOPxpIPYjjdDk1OnCoBis/Sfzy5For6NVNWKf7+Rd6RVecWt4CB2+x1dCck3zbSoOQRx3nR5uG9nhR7eaC4KLgH1HIl3ZD3COIklUNHcpaKnhBw/6v3udftxxal/X7Vgwpq1m/3bzWigGMNu5v4tY598oSxE0hI8hd/EjxOCWQOf9lxKeGWg1fXWs47Otr8I6qXgGhV61CriVOEh1Y0sTZ2JVscAnADdIoyLp6mtXJ04t5ye/kCaG/Cips5R6rCXSgUSRgc6Vj+6CkAiEPrBEBknua9NxLPlGB5uCHZR4Z3+uu+vf4N/Me3q2agSiDi/n/D6umI6XsR1CKHGvDAd9udy7/RMyaiOE3wmFrkWU1DDwtGUA+shqDm5LRcQovbn0UBCek01yr933bI3rnzuleuJhvIQ+sEQGSe5qPTkVUE8JgL+5oythSdMPw/5ZEpvnnCbeHi01zgwg6osjTDan1LY/bEZAC3bvJxP5meILWUKgVMGuRZTUMPC0Z5zv/wJGiTbL8SvJXScv/ZXeMgv3oRcDnJvEZO9mKBpshD6wRAZJ7mjuO7n0C1r4WTwo92JO+lNOYbhkpwC4T/9JeSNvONVLyibe6J08G1E4zC7wQK4TzmIypvzpPlRBwhCHFYzNkpjRT4A85W96WwMNJMecpme9JPxeVHY2ukRH8AB54KP2dtSEPrBEBknuaIHJ+u4OHV5jmVQgcWasZb/sj43xyIb4eusfdNB/IdZxcYAomaEwmZIQOXtDU5u889qQ5v7YHwpWJwEzYb4hXIW+Y0dg3b+F80PHPcHSInAdUx6MurK0KvAGPwkw2U4rIIQ+sEQGSe5qGipHRm0sXuJAuzK6wbsDqctJkFf8ZfvbiwIK8U41mvnCznftZbQGvM8L00CbT6wY/sqjk+k9SposZMhxvkGHbHSatHr5It4DFvcgvmb80lTtpxcGpQbshyTVheLnKFqUhD6wRAZJ7mmnGWJ+fzudCLG9cd+T+HoQwJ1eCSwCIfeWuZc9aJE4AcLOd+1ltAa8Drb9s7cm2wvw3vXiN4TaoQ0yc6HjW9tpbrZZ5iiCZDdCHlB2vCDHXgU+XL9pinxJNc+1jOjQNgCEPrBEBknuaI6rvJVVs8srol4gFzMlsFaawhz4FPe1LktIgbfynmZFws537WW0Br3+YgywUPINFKL+0xOIS6BRDTJzoeNb22pOVhTXHK3UQ0IeUHa8IMdeBT5cv2mKfEpFMtcg5h2HKIQ+sEQGSe5q98s1PqbkGsciuJ1vYj11amlE62q4H78TlrmXPWiROAHCznftZbQGvmRtgKQvxGIAj0kHpIYKDgonATNhviFchUOwu5X+nlCbFvcgvmb80lTtpxcGpQbshFKCOCWH8bBwhD6wRAZJ7mgknJXF6FDyfveyCH8xBFnbl/lMG4EAUquLAgrxTjWa+XGAKJmhMJmSl7r/l8mHptbfQ4cVtAgihcAnADdIoyLqAR5IctJYlo9Dxz3B0iJwHVMejLqytCrx3EPxnSZ1p6CEPrBEBknua9uNazyGYieZyHXf7GYdcBK9NeIOhCnx/usfdNB/IdZxcYAomaEwmZB7bTh8KXRU6otOqXZeJO0CEIcVjM2SmNGUzihLU9H1Sw0kx5ymZ70k/F5Udja6REQvQwdh199lHIQ+sEQGSe5qcAir8rvOatkg6WJaGjhW882nCLk2rkijSXkjbzjVS8om3uidPBtROFFhsDsXhTtpuBWiL0HuiQ/8C2SZVmDNdaCpNmYWFotr8SvJXScv/ZXeMgv3oRcDn9W5PCuoKIQYhD6wRAZJ7mqX2OKRWT8TXyMW3xiZ69ToUIy4Z1cIdQIeLTXODCDqiyNMNqfUtj9vHupnIqnGSrn42VhiMLM0RicBM2G+IVyFGcq2QeZUzenEKL259FAQnpNNcq/d92yM8G47iTSfwNCEPrBEBknuaerkFeqhhROz002Riix/MNtf9NgLi2KrHgSiDi/n/D6umI6XsR1CKHFY9CrR8sc6DVP2ytLPYwZPoOI/l4KNd8ZDN2fyyNG4X7+QJob8KKmzlHqsJdKBRJJZMuIx4Gai0IQ+sEQGSe5pcYc5JF1GcMf5jxIIwenTUW9yfZxjxmx6nhloNX11rOOzra/COql4BlJXT/1SmazfSiOOniWREO+aC4KLgH1HInklgbTjURxMNHcpaKnhBw/6v3udftxxaPp/nZsYtffG/3bzWigGMNho0bmLTcIruNV3pNOhM8SA5rErLfUGP6/v5F3pFV5xaZMXpaMfGrGKTfNtKg5BHHTeOYR8p3goC5oLgouAfUchTT3ZYhximWKg+0cbVI0KI/q/e51+3HFrwd8QvOvqfHr/dvNaKAYw2vT0wsN4LwH9ZfXe8LoxOrfE4JZA5/2XECoy6wKFWQsFFEde3ZxAAVKFXrUKuJU4SxOC7gTSKuN1wCcAN0ijIumSkD5mog/nvua20TykTKW7lHqsJdKBRJPGJaYh+6I/+uYeHg3QpABL03Es+UYHm4HVoKyJwGrrB9/g38x7erZqZnXKC21cYBEqq5hzqTqJUa8MB3253Lv8OwvBssuGCOWuRZTUMPC0ZAN5EPRILQnirBfYRnJT/PKTTXKv3fdsjMh2mmPF9OD65h4eDdCkAEo9ORVQTwmAv29wkxMp1hED/lkSm+ecJt6av25hibhltSvDmWDgh1+gRkALdu8nE/lyUWm5V6c8pa5FlNQw8LRl5CKeVaj4YZBeVIxxCJM1/d4yC/ehFwOcc338tO+Ojg7mHh4N0KQASO47ufQLWvhbtBGlZxGho4JhuGSnALhP/myq6TgNFCPOpKfz6XsqAqzMLvBArhPOYafv6gndPMeqEIcVjM2SmNKzczXOESz00sALoOg6Ow/I/F5Udja6REVhVvtJrCnNyuYeHg3QpABIgcn67g4dXmK0GeMJlV3nm+yPjfHIhvh5tnDga7h4e0mwCydbQ5eYohA5e0NTm7zzkRCVZFvzcXYnATNhviFchAs7iqUfiASJsKKfQqLU90lTHoy6srQq8ucUhPvL1ZXa5h4eDdCkAEoaKkdGbSxe4x95n7l1B7HJy0mQV/xl+9rYeGN5DTz2kdO41lfCW3CUzwvTQJtPrBsvVhVtecDA8ixkyHG+QYdvLNhocnH8B3FXfvz6Hn1IJO2nFwalBuyHeV3nk+mUu57mHh4N0KQASacZYn5/O50IS+AgU4u1kNjAnV4JLAIh9kLTjdD5o6nt07jWV8JbcJQOtv2ztybbCVkKIg2mTtoZDTJzoeNb22n5nErH3kgJR5LZvwy6Rt3mBT5cv2mKfEoI5K9vSc2jSuYeHg3QpABIjqu8lVWzyyvlJsCkR2H7AprCHPgU97Uu31h1GQ8SZEnTuNZXwltwlf5iDLBQ8g0Wg5sMqtsLs9UNMnOh41vba7MUyVqJ6gPXktm/DLpG3eYFPly/aYp8SDeWmNqKs5Me5h4eDdCkAEr3yzU+puQax+J2RHekLYJqaUTrargfvxJC043Q+aOp7dO41lfCW3CWZG2ApC/EYgEEvujMjvMuKicBM2G+IVyFuGyupup3illXfvz6Hn1IJO2nFwalBuyEjy1Bokzk1j7mHh4N0KQASCSclcXoUPJ8cqJvGgupYH+X+UwbgQBSqth4Y3kNPPaRsAsnW0OXmKKXuv+XyYem1PxLCciJ8i+NwCcAN0ijIurGhAtdoZut0bCin0Ki1PdJUx6MurK0KvOqpSPzleLKVuYeHg3QpABL241rPIZiJ5rZE4NeIDE6+r014g6EKfH9tnDga7h4e0mwCydbQ5eYoHttOHwpdFTr8zzSvpYX+v4QhxWMzZKY022xV5qNoe2awAug6Do7D8j8XlR2NrpER0IP+bBPZ3oi5h4eDdCkAEpwCKvyu85q286tjQTq4WfHzacIuTauSKJsquk4DRQjzqSn8+l7KgKsUWGwOxeFO2kZotewlp9ZE/wLZJlWYM10DPU+xyyynyBeVIxxCJM1/d4yC/ehFwOcRQzpnHqrnjrmHh4N0KQASpfY4pFZPxNd26d4mM3vXtRQjLhnVwh1Apq/bmGJuGW1K8OZYOCHX6Me6mciqcZKuZn5AeGihWuSJwEzYb4hXITYk1GfyHPxhqwX2EZyU/zyk01yr933bI3gwjzTzyFOmuYeHg3QpABJ6uQV6qGFE7PhWaJ7e93p31/02AuLYqseZnXKC21cYBEqq5hzqTqJUVj0KtHyxzoMAwmCRzxlGSug4j+Xgo13xkSwZA0FErhq5rbRPKRMpbuUeqwl0oFEk4ig3pcBR38G5h4eDdCkAElxhzkkXUZwxYlDX+6nWOmpb3J9nGPGbHgqMusChVkLBRRHXt2cQAFSUldP/VKZrNzwaflW2p/865oLgouAfUcg0/MitnYoY/Kg+0cbVI0KI/q/e51+3HFqXK2eQGAai/L/dvNaKAYw2zCa/bhNMUhOm26qLvQyifYJJvbdxS96ROMKA1BJV2ZOY2sBIU160RIJrvo36wB1+pmH7SyfPW5XouUwLdVD4znbHIi3kdRDOcLOd+1ltAa/tyRxTCew0adtbpwbGUdZo5oLgouAfUcj/W4Qtf+OPl9CHlB2vCDHXgi2Bbl1JsG1pnb4+bN9piCEPrBEBknuayrowlNjg55hZU5jk7QuxatxpACsWd+h/27dqUGjYXypws537WW0Br8R5UTINsWCHBWvEr5xzlXdwCcAN0ijIugmcVWaYVkeCbN3gKdTpp6yZC1PtrPWOOiwBhf1bym2MIQ+sEQGSe5rFsLrrE7m/y7iRw+BG0Jigi0ZvLnB9+wiY5XC4M6wzTnCznftZbQGvD/Xe78B73XcQdufLkr7vwXAJwA3SKMi6LNQgGT1eRLgTd1pAT9xUTu59oK9n9cckTnjbADMlkCchD6wRAZJ7mnrnoVTk5qICbDi6dn53kM2uVy24x2hFCf5dO7jhULAIXGAKJmhMJmRNvJtWZbWYVt3ot96Yqd3c/wLZJlWYM13N2oP9M5yF0RjRfT9W3GmoKotHhtD9VModrsXzaL0V+iEPrBEBknuasz/zA05H38xM9uG33/7HMVvcn2cY8ZsenlNtHCGV7JSJt7onTwbUTrnzHJ7DoowY0Dk/lVIngM1rkWU1DDwtGXCKN66Hifr84Fcp/wDvyx/adQMEFm7KCWxFFnxb/D0HIQ+sEQGSe5ppbGSW3qoZLSqhzdXrMu9a2uvRE6wBfZ/Q/KEka7FrJMjTDan1LY/bAZl2IwTnMp/I1Di5r8cE8YnATNhviFchAOFK2RNW09Gk+RWUOrCRIe/Y+iZAf4HBQjg5dCdHJz4hD6wRAZJ7mmFcv5ZUu0I98rGGWWRjqIblFBqrrLEEjIexyVEQ9Ul0piOl7EdQihw8qW2NM2Ca2yu5Drc11vdC5oLgouAfUcjbQ1hf6/sDoJMcgGIxLsPCCk7QPmljLUaZilziUFKR2yEPrBEBknuaGXxVQvJ/IBbkcc+tUU8Yxlieewh70aIa1+kLox4HyMfs62vwjqpeAQmD42Ga+TYIrvi1Ru/bfqdwCcAN0ijIunswvoXijCXvZVRog99tUC8M4FzmHpcse9Hdy3vUqEc1v9281ooBjDbFnm8bH25dpnanVXz3QgowprCHPgU97Uu7YO7F+IrCJKg18ZZFxsrfoOnJ35NqY8YNp0AGygJ+1eg4j+Xgo13xxvdjSm/7XnRyLsaH48FjiuvwwEk+muBoErmCahRFRzy/3bzWigGMNgp+QdVc8JxRQCaTFIyA7uamsIc+BT3tS3j8oe6N0aToRRHXt2cQAFQJg+Nhmvk2CFMjUfxttUYHhCHFYzNkpjTOkJeHLiTY6LkUInUSLxfjdrSs/+hsjXnXg0jiwlNda7mHh4N0KQASQr9Eb+F4mVzSiu2ttxxdPqLBFVg1NSGXI9gc0/oYpWZKquYc6k6iVDypbY0zYJrbkosr/qu3NDHoOI/l4KNd8dBmhEZ9rOeU5jLXNv2NJnUDxSRolJs0QtWP5B/C+41VuYeHg3QpABLtGr/FxDe7Okln8DHjmNDzm3iYmZPLdYhNAvGTGeHNr0rw5lg4IdfoAZl2IwTnMp8HJIPWgLc0IeaC4KLgH1HIUgsltFmSqwg1n6NfvXMRIn/9zzow/yknG4s4e8gG4Mm5h4eDdCkAEu9NFmf2568OQ3Q1w0X0b0w8niBbeUChi06+ywEyiw2xqSn8+l7KgKu58xyew6KMGAkbc9joz4tncAnADdIoyLpAI0fZ8y0AnYP5zZCdRSElWRYnF1fHkDdRJWM0mYTHIbmHh4N0KQASJ3/NyB/1QoyLVqEEcRd8bc02TRyV9LkiTzbWGioskbdsAsnW0OXmKE28m1ZltZhWgLDR7uktF/HoOI/l4KNd8UIS8jByShWxbCin0Ki1PdIM4FzmHpcsewTRRR1mvX3PuYeHg3QpABLy0MjFZ+oR4RDKbf/pDTz4MCdXgksAiH3x+3juSi4pRnTuNZXwltwlD/Xe78B73XdnVuM862WZJ4sZMhxvkGHb5U+izjLHkQ1V378+h59SCSZhO/W05NS6nWaKA+qi/9O5h4eDdCkAElHEU9eu/xSYCr5oiyIcerjZr5pdGhkLS2wXZoUXjxKJdO41lfCW3CXEeVEyDbFgh9FOtHKjuFdz/wLZJlWYM11zZijc6tw6ZOS2b8Mukbd5cHv4EM2dWRr3PDqLPphGxLmHh4N0KQASKSzbQtOYNI/yB7up3I8vFIRwMi+5L7VmnvFYOKw+U0t07jWV8JbcJe3JHFMJ7DRpwOgC+pWkf5DmguCi4B9RyJjfHQIHzfdn5LZvwy6Rt3mCLYFuXUmwbfc8Oos+mEbEuYeHg3QpABLKujCU2ODnmA5OB0V8h5Vb3GkAKxZ36H/mr2PhPU8zhHTuNZXwltwlxHlRMg2xYIfRlQ4BvXrmwXAJwA3SKMi62GBrlu0g/n+wgxjdf6gG7JkLU+2s9Y46nWaKA+qi/9O5h4eDdCkAEsWwuusTub/LxsX/FPumLdGLRm8ucH37COVgaBkON9l+dO41lfCW3CUP9d7vwHvdd0YmOsSFBUVGcAnADdIoyLpZrZtxfJxb9+J4EuxpMgIj7n2gr2f1xyQE0UUdZr19z7mHh4N0KQASeuehVOTmogL4gGoW9p3Pe65XLbjHaEUJ6rasPFbPGkNsAsnW0OXmKE28m1ZltZhWPaHJOBy8RN//AtkmVZgzXZ2Rkmpcdj8DiXKSUTM5p08qi0eG0P1UylElYzSZhMchuYeHg3QpABKzP/MDTkffzN85aG65qN7eW9yfZxjxmx5PEwaPwE8NOakp/PpeyoCrufMcnsOijBh1tjX+G5nNSWuRZTUMPC0Z8fYKkxarmSkcuCgX1JANq9p1AwQWbsoJG4s4e8gG4Mm5h4eDdCkAEmlsZJbeqhkt4XncQ5yKj6fa69ETrAF9n5uGJItctMgmSvDmWDgh1+gBmXYjBOcyn0kUILI6C+FpicBM2G+IVyE+VXMfrRu6EQyAbVbZPJEJ79j6JkB/gcHVj+QfwvuNVbmHh4N0KQASYVy/llS7Qj1ad97KbXS8o+UUGqussQSM5O4AyNbvs6BKquYc6k6iVDypbY0zYJrbuMDb+5YGYQ/mguCi4B9RyNiJheDS93Vj8V9urnRrVwQKTtA+aWMtRteDSOLCU11ruYeHg3QpABIZfFVC8n8gFsuts9AF9rgvWJ57CHvRohrwHB4L9LfMr0UR17dnEABUCYPjYZr5NggQRnU30TKfKXAJwA3SKMi6O367zJl2y82NtKSn6oHBFwzgXOYelyx7ErmCahRFRzy/3bzWigGMNpZyQmZDQjZriEFHedsM3fqmsIc+BT3tS7zqY0Vv7nnbqDXxlkXGyt+g6cnfk2pjxmKZ9lRvvHFW6DiP5eCjXfF7iUoUDrPkXDvpUsUMN47E6/DAST6a4GjR3ct71KhHNb/dvNaKAYw2NYYH/VFqT1nmMC1JclDc06awhz4FPe1LNlC5M6GoWwHs62vwjqpeAQmD42Ga+TYI59rPlqTkdMOEIcVjM2SmNC239gbavXJbhN3zwFwsOwh2tKz/6GyNeZmKXOJQUpHbIQ+sEQGSe5pCv0Rv4XiZXH5VXX1Qmot0osEVWDU1IZfGbGpZXYbsg6YjpexHUIocPKltjTNgmtvBC0ud0n29yOg4j+Xgo13xb38SaZDx3yy+GdLknoyCyQPFJGiUmzRCQjg5dCdHJz4hD6wRAZJ7mu0av8XEN7s6hFyVlM3wIx6beJiZk8t1iG++rhWmjSxdyNMNqfUtj9sBmXYjBOcynwffCVCKW+U05oLgouAfUciswqZwiflE217r+PZNVZx4f/3POjD/KSdsRRZ8W/w9ByEPrBEBknua700WZ/bnrw4g7jUBaDdwMjyeIFt5QKGLbiZYYmTOLGyJt7onTwbUTrnzHJ7DoowYMogXB0XCVppwCcAN0ijIuiP2faVRDuq32UPAztLtTmpZFicXV8eQNx2uxfNovRX6IQ+sEQGSe5onf83IH/VCjEr+lJYP56OgzTZNHJX0uSLwTAxvn2HXM1xgCiZoTCZkTbybVmW1mFZjRsqc2JHa1eg4j+Xgo13x2iQsjeFRrJ/Q8c9wdIicBwzgXOYelyx7TnjbADMlkCchD6wRAZJ7mvLQyMVn6hHhtvky23maCnMwJ1eCSwCIfd42/BlqqNCIcLOd+1ltAa8P9d7vwHvdd06HRF8e2o1HixkyHG+QYdtpgGFXn8Q7QsW9yC+ZvzSVJmE79bTk1LosAYX9W8ptjCEPrBEBknuaUcRT167/FJhzNTrg4CLh19mvml0aGQtLKx5o61xTZSlws537WW0Br8R5UTINsWCHgldcmqEXe1T/AtkmVZgzXZV57QTphx8i0IeUHa8IMddwe/gQzZ1ZGmmdvj5s32mIIQ+sEQGSe5opLNtC05g0jycycrvZ9Z05hHAyL7kvtWbQ5GFWrTQQzHtGVKQ7oCj/beCNc4SiTRLmbFK7/HUvHIgbGbHfZNlDkMABQU0zL8vx3YAxNXoX5OeViVMdq//ldR9OXVDwvGK/3bzWigGMNiCvWPBMpx/ngqatO6IboJG/3bzWigGMNiCP9qd3hq8Si++SkKr1CXS/3bzWigGMNobEa9xB4lwh3h/AUyMzKHu/3bzWigGMNi0K7wMWsEU+nUiIMtve0ve/3bzWigGMNjxtYM5t1qQaM9kGsLNoNCm/3bzWigGMNjfOB3h5FVLnQR6C3jk98KG/3bzWigGMNhGFdRZnphLKWDVqAHPa7by/3bzWigGMNmjVYdo+Vxv1F3wRWU1Tc1e/3bzWigGMNujiOCGGiqEwmloH4ml7qau/3bzWigGMNjpqFW8wFpNA5UBa6FTJHHW/3bzWigGMNpIpZ8LFkOmZF4/iidHK+B2/3bzWigGMNsdzzjyr40VREhAhJFT8BKK/3bzWigGMNkVh2CTTj7Jxgh5jVicR9BG/3bzWigGMNlqkgG3mrBqnqCylWFDutm+/3bzWigGMNm0f1yA5GfkY0I50Iols50+/3bzWigGMNkwLyRKj7KuuWKp8boJAKeW/3bzWigGMNp0bp52Di3KHJ4qeJxyde66/3bzWigGMNgBARs4ONDnhByO/BzEFTXe/3bzWigGMNtqaccdkiIT0gPbQpobktDG/3bzWigGMNsVodNteGJ4BbtxWzFBvVyK/3bzWigGMNlrI8uA0l53/HQhd/gOsqry/3bzWigGMNr2QNfjhza4ESU0GGXwm356/3bzWigGMNlqfmJorMq0nFCzpAA4983C/3bzWigGMNqvPTsbv/j4E/l8Q/0qFAsG/3bzWigGMNhCj3FOhSnAx6sRMWG1Sqpm/3bzWigGMNhy3QUftfavDPh4uP4SquJG/3bzWigGMNv3BnV4JNxk/WALHfaS/6uO/3bzWigGMNqGiXRY3Aj4OQvlghDdGh+2/3bzWigGMNpe9M443RO/wlUjNPSzzpEi/3bzWigGMNkyCuaJ7g4mXyMW3xiZ69Tq/3bzWigGMNqAuBx2gfOvPKqHN1esy71q/3bzWigGMNs6kj3tyB6hk9HE6s1KOwH6/3bzWigGMNnUbfaOp0iG/QGrte0GihUW/3bzWigGMNk5QkkqcVbM7EobwtsVxu4+/3bzWigGMNmqLbz2uuLBSIO41AWg3cDK/3bzWigGMNnPdQufnNvSXsAwy6zANxwu/3bzWigGMNpRaeXgkCa00kg/b+E93xWi/3bzWigGMNklxgB12k0ZZVCyP7/ealgm/3bzWigGMNvsjcbggxu4ridrDytpv01e/3bzWigGMNgdUqgGvcKirxgvSIVAf2zi/3bzWigGMNtnl1lLqoqNEMqi3sFSmujm/3bzWigGMNrao7+9S8aGd1eIZaHfswH6/3bzWigGMNoufyEkpZi+IBpZmUhRyTOG/3bzWigGMNhXaQhlf0Vqcch13+xmHXAS/3bzWigGMNn/hQaDm0QwgG5j9XqZ6Rsy/3bzWigGMNn2jmQQbnR4sxYLi9RT/qt6/3bzWigGMNsneAU+V27EwvPL5fVlGryC/3bzWigGMNgL7HeR4p5VR9rX2oojpnUK/3bzWigGMNiNPg2VcGo53Yffh7lSwrj2/3bzWigGMNp88iVLEh2HI2Y99n8nmnVS/3bzWigGMNkq/YFq6XRmckzE3O1ucmUq/3bzWigGMNj+nfDopYk9pJPbtM08KQkS/3bzWigGMNsXg3CT/aoucF+YnPoLEy7a/3bzWigGMNrptykQpCf7vc6HRvERjdTC/3bzWigGMNi/C/3lCBzqfvtYYln4l7/G/3bzWigGMNhmjHMQQRqiYi1M1R306lDy/3bzWigGMNsBnLGm8zE/vqBUtnyByA6q/3bzWigGMNm4eMUqsMuLiWSuHbUbCKYu/3bzWigGMNgkEcVsxcMAWUft5RbHMsWi/3bzWigGMNmARTp6EDFA0evqBBkIp2B+/3bzWigGMNnVRL0lHewKg4lhPJE2ogdq/3bzWigGMNjbiKPKLL+NNvVwgFpkjlre/3bzWigGMNoP9O5zPl9Kqui5/JkSHSGK/3bzWigGMNqBHQUsJOfs7B7kBgYzgui2/3bzWigGMNuW+2YtRaFnutWYY0A+iTF+/3bzWigGMNuglQAa1S4w24ZHO0/ICCJ6/3bzWigGMNp7pO7nBgeOe4Xk8+dJXWWK/3bzWigGMNjWiHlf+JB79967bLb2K8/m/3bzWigGMNmHQuN1e0vSPoigxv1Sk04K/3bzWigGMNsrf9oha9bKLvsSOfd5ugfC/3bzWigGMNnRqQKwu2U26nMrlsWam1Yi/3bzWigGMNmDW15ZZDCKqHEKgePOCbfS/3bzWigGMNuzQTpu2BYvkSlVkaoAtUiW/3bzWigGMNtd8q+35uajbxYkgNOk80lm/3bzWigGMNn4Ru7Xuhc6MrUBfsfTRHG+/3bzWigGMNhM0IrdEFXb3dL0tSrdIf52/3bzWigGMNp20l+ObS89vLN3TIZf9gw+/3bzWigGMNnph/wWPZ87A+VxgRDQ9ywu/3bzWigGMNqQOv137JpdrF7zZF9VjrwC/3bzWigGMNlJfM+gqXnQoNZn2MPNrwU4hD6wRAZJ7ms0zoynRYXMhPN0Cl8OvGyghD6wRAZJ7mr3bPn77j4QLl3bXNWmn7OMhD6wRAZJ7mhLCDTnClTPSnvSQQW7UbRghD6wRAZJ7mpxIlWkWJXvszCtXgSSXdwEhD6wRAZJ7mnKthAu0BlH9XJAqxt/A+1chD6wRAZJ7miJMXnKrXPMhMfRWbmIbP18hD6wRAZJ7mljdHDj4GmB3YOH8ilFvbMMhD6wRAZJ7mvzunp1YH77pDhY/fSk+5vghD6wRAZJ7mh9ZUXWcamPKEPaPwApekSQhD6wRAZJ7mvPOhOx5YMZQMN7db0Gj94YhD6wRAZJ7mlN86itW+5AVoBhefcypId4hD6wRAZJ7mq0hSfOrMRcUZpZ4uFstFZ4hD6wRAZJ7mkXhXwC/YnbMsJlUZCrd0ZAhD6wRAZJ7mleRuMo8IcRo/K/xnSf2SGwhD6wRAZJ7mqTswrBfw0Pm6D7IGJewNF4hD6wRAZJ7mlCv1JW+BeAt0dz6brN7aq4hD6wRAZJ7mnTBqVAjRXaXRXXfwSqseBQhD6wRAZJ7mq5xI2eu6p5h/D4jLeb+88EhD6wRAZJ7moTA6gp+za4wcf4nhgkgLachD6wRAZJ7mlseSEBwrMVueLO23HdK93chD6wRAZJ7mhLN8fXIaoSHXhNdNPF8G0EhD6wRAZJ7msI1Q4puL8WEzO78aTAIw8ohD6wRAZJ7mtqasNOs9FBh7rpdjUL9ZdohD6wRAZJ7mi77esJ4TjoAYIPYgsIFs2QhD6wRAZJ7movoTHIa9/7SXuXmQ7yeJSMhD6wRAZJ7mvkmGk1QTW95zBzRIDEkICwhD6wRAZJ7msspYlPKuA9Gh9jpQD26Js4hD6wRAZJ7mi/jUaYwS7vzpnDiULBcxZAhD6wRAZJ7mhDPRi4RKVeem0AaSahmhv0hD6wRAZJ7mncMerNh9MdlvWpe1aWalMAhD6wRAZJ7ml4HpSpEu+HgdsdNVha+uf8hD6wRAZJ7mph/IffJmDLQ74sAi99ZogkhD6wRAZJ7mnLI3hDrN2lvE88GqQcYWtQhD6wRAZJ7muPCtPMgTlBtA6Y4UVKiBHwhD6wRAZJ7mp+94yENyMh7wlKb3qoTtUIhD6wRAZJ7mqnFuBBCJlXgtiiR2j+B3A8hD6wRAZJ7mp+l/J4kBs+jnE2tlRQYdbYhD6wRAZJ7mvFs+kkRiEuSDCDftjKsrVshD6wRAZJ7mrYycYS/XmgweWrOsRGpwlghD6wRAZJ7mkqwWrllEGGNJL+k4EiE70khD6wRAZJ7mjY7GDOI6LFmb3Q5HJn3HTMhD6wRAZJ7mutEd8erVCZhSzfBGN1qn/8hD6wRAZJ7mu1tjkQ5yCmy4QMr+0DihOQhD6wRAZJ7ml6P8hCgYnEGlE9LmF0CLZMhD6wRAZJ7mtikvbPXpIAD6IHjwtNi7nQhD6wRAZJ7mhNJrUeL3WSwRf4VclqrwhchD6wRAZJ7mjYbQwx9Jd4OoMcrJQ/RQKYhD6wRAZJ7mk/rL84vNybYjMPfC77s2Y90ehU8dWq+uSvU6lSnQCeoYmABKohTdQLxaBuWUrhj6m5EUEFx0rygaDHA85r5sJmgZVy++TWyOdCHlB2vCDHXldzse6NiQBeN9nOlPo+AaSEPrBEBknua9Wzp+SMPf3Hol4gFzMlsFRQjLhnVwh1AktIgbfynmZFws537WW0Br+3JHFMJ7DRprvdMvneY+ljmguCi4B9RyKBlXL75NbI50IeUHa8IMdeV3Ox7o2JAF432c6U+j4BpIQ+sEQGSe5r1bOn5Iw9/ceiXiAXMyWwVFCMuGdXCHUCS0iBt/KeZkXCznftZbQGv7ckcUwnsNGmu90y+d5j6WOaC4KLgH1HIoGVcvvk1sjnQh5Qdrwgx15Xc7HujYkAXjfZzpT6PgGkhD6wRAZJ7mvVs6fkjD39x6JeIBczJbBUUIy4Z1cIdQJLSIG38p5mRcLOd+1ltAa/tyRxTCew0aa73TL53mPpY5oLgouAfUcigZVy++TWyOdCHlB2vCDHXldzse6NiQBeN9nOlPo+AaSEPrBEBknua9Wzp+SMPf3Hol4gFzMlsFRQjLhnVwh1AktIgbfynmZFws537WW0Br+3JHFMJ7DRprvdMvneY+ljmguCi4B9RyKBlXL75NbI50IeUHa8IMdeV3Ox7o2JAF432c6U+j4BpIQ+sEQGSe5r1bOn5Iw9/ceiXiAXMyWwVFCMuGdXCHUCS0iBt/KeZkXCznftZbQGv7ckcUwnsNGmu90y+d5j6WOaC4KLgH1HIoGVcvvk1sjnQh5Qdrwgx135pivyILuXTa5mH6RgyVREhD6wRAZJ7mo7dCAZ0A/pR6JeIBczJbBVihw1tijCQfIG+quVOWQpjcLOd+1ltAa+pwbnWmLiplK73TL53mPpYixkyHG+QYds3jrHyQe+Yh9CHlB2vCDHXfmmK/Igu5dNrmYfpGDJVESEPrBEBknuajt0IBnQD+lHol4gFzMlsFWKHDW2KMJB8gb6q5U5ZCmNws537WW0Br6nBudaYuKmUrvdMvneY+liLGTIcb5Bh2zeOsfJB75iH0IeUHa8IMdd+aYr8iC7l02uZh+kYMlURIQ+sEQGSe5qO3QgGdAP6UeiXiAXMyWwVYocNbYowkHyBvqrlTlkKY3CznftZbQGvqcG51pi4qZSu90y+d5j6WIsZMhxvkGHbN46x8kHvmIfQh5Qdrwgx135pivyILuXTa5mH6RgyVREhD6wRAZJ7mo7dCAZ0A/pR6JeIBczJbBVihw1tijCQfIG+quVOWQpjcLOd+1ltAa+pwbnWmLiplK73TL53mPpYcAnADdIoyLrjKP87N5hhPNCHlB2vCDHXaLZpG3LhexgGd2/X8w6XySEPrBEBknuad27tRNVvGFzol4gFzMlsFfjH8kgwMRj/yHHDZiuayzhws537WW0Br57HQ/9cWCZMrvdMvneY+lhwCcAN0ijIuuMo/zs3mGE80IeUHa8IMddotmkbcuF7GAZ3b9fzDpfJIQ+sEQGSe5p3bu1E1W8YXOiXiAXMyWwV+MfySDAxGP/IccNmK5rLOHCznftZbQGvnsdD/1xYJkyu90y+d5j6WHAJwA3SKMi64yj/OzeYYTzQh5Qdrwgx12i2aRty4XsYBndv1/MOl8khD6wRAZJ7mndu7UTVbxhc6JeIBczJbBVCJSJQ8JmgiU5xosr6WW2YcLOd+1ltAa8H1MgAUYzoOK73TL53mPpYVjDFFn+2SgScO0bStFiJG9CHlB2vCDHXbsT+phbpGyECH7QqVoxcISEPrBEBknuaIzB/9eJZ+6Tol4gFzMlsFUIlIlDwmaCJTnGiyvpZbZhws537WW0BrwfUyABRjOg4rvdMvneY+lhWMMUWf7ZKBJw7RtK0WIkb0IeUHa8IMdduxP6mFukbIQIftCpWjFwhIQ+sEQGSe5ojMH/14ln7pOiXiAXMyWwVmMEu+JWkoYB+amxH3jG973CznftZbQGvCYyESxSEGPiu90y+d5j6WInATNhviFchlC51k5PUZ0PQh5Qdrwgx13B7y5T3RPq0WA4ue+TQSiIhD6wRAZJ7mmeTN+vlz+T46JeIBczJbBWYwS74laShgH5qbEfeMb3vcLOd+1ltAa8JjIRLFIQY+K73TL53mPpYicBM2G+IVyGULnWTk9RnQ9CHlB2vCDHXcHvLlPdE+rRYDi575NBKIiEPrBEBknua/maR4s+D39nol4gFzMlsFUI8QhDRs5vIKsoVg6eHDShws537WW0Brx7os/XNCsrLrvdMvneY+lj/AtkmVZgzXX+4GsTIRoGk0IeUHa8IMdfqgIGvqQQnRWs3aDDNmg2yIQ+sEQGSe5r+ZpHiz4Pf2eiXiAXMyWwVQjxCENGzm8gqyhWDp4cNKHCznftZbQGvHuiz9c0Kysuu90y+d5j6WP8C2SZVmDNd2fjv5jX4apHQh5Qdrwgx19pUocIq6zxe9nx2gHG187shD6wRAZJ7mqGNX8Bkkql96JeIBczJbBVBMkmZvxLRjziHdv7jHnDzcLOd+1ltAa9kHTFvKESG5673TL53mPpYa5FlNQw8LRnZ+O/mNfhqkdCHlB2vCDHX2lShwirrPF72fHaAcbXzuyEPrBEBknua5lW4ilKzuz7ol4gFzMlsFd/ktAaaR/xkYZanZRJkLfVws537WW0Brymhmx8Q67gc5vMvmaTaGJWEIcVjM2SmNHSVKCWus/Iy0IeUHa8IMdcwUSSYaTP+Tpt7fV/hgrI5IQ+sEQGSe5rmVbiKUrO7PuiXiAXMyWwV3+S0BppH/GRhlqdlEmQt9XCznftZbQGvxJLs4F+ArQLm8y+ZpNoYleg4j+Xgo13xXHfAY4+o9iPQh5Qdrwgx18c3b/ZTBaX2MafOxlb4T/4hD6wRAZJ7mipT6yK3uiyg6JeIBczJbBVsoQZyXj6g6fAZU3po3gZvcLOd+1ltAa/EkuzgX4CtAubzL5mk2hiV6DiP5eCjXfE3x3580t4xvdCHlB2vCDHXvMSiGrmydcjlN9JiBGoVuyEPrBEBknuapQSim0dLldXol4gFzMlsFdxpACsWd+h/25R4klbiemxws537WW0Br2VfSuEwf7nW5vMvmaTaGJVDTJzoeNb22jfHfnzS3jG90IeUHa8IMde8xKIaubJ1yOFV9mmYDz3SIQ+sEQGSe5rPwGSgX4E3I+iXiAXMyWwVNIpP2sfz5OSe0ll+5h08AnCznftZbQGviI/mhTgvhuLm8y+ZpNoYleaC4KLgH1HIBi+rrBUXpnvQh5Qdrwgx1+7+7/eRj+si4VX2aZgPPdIhD6wRAZJ7mmD8t0Jn5Xui6JeIBczJbBUrooGX81rsjLO/65Nfmq8jcLOd+1ltAa/WGouOT1rAq+bzL5mk2hiVixkyHG+QYdsrF//VyKIgddCHlB2vCDHXYg8gz0Cp2TkzTu2q2+JQ0CEPrBEBknuaYPy3Qmfle6Lol4gFzMlsFVieewh70aIa5ep4/IQj27Nws537WW0Br7SvQkCqPPue5vMvmaTaGJVwCcAN0ijIuouVyutkftVS0IeUHa8IMde4YTo1jtIAqFPPtY5o/i1hIQ+sEQGSe5r3oKtKF+SG2+iXiAXMyWwVh9rATNG1pu4bCF6NnZ4ZdHCznftZbQGvsYEK3wC4tPDm8y+ZpNoYlVYwxRZ/tkoEpx6LP5vbX1PQh5Qdrwgx12TD6UN6kcwU2AY+DwX8Ol0hD6wRAZJ7muwat/7Ib3Rw6JeIBczJbBU8HVd7vWAgfOKCJTsKr4FHcLOd+1ltAa8uoXjUzkBCwubzL5mk2hiVicBM2G+IVyGoRjq3ByLhH9CHlB2vCDHXQtrfnAsueuOQq0VrD5tgdyEPrBEBknua0PjuB1mZhWzol4gFzMlsFTnqLpES0sCm52E7HB/+3KFws537WW0Br0KKK+FCes2A5vMvmaTaGJX/AtkmVZgzXWuNIirURLVC0IeUHa8IMdfxQ2J6/6GnVA+aa/dBTyMnIQ+sEQGSe5q0P51+vEeb5OiXiAXMyWwV5RQaq6yxBIyxl/I0avveE3CznftZbQGvIeQV4Z+ppWvm8y+ZpNoYlWuRZTUMPC0ZJ1IA4kgWs4bQh5Qdrwgx1zlgH+K3uJWNK2WizVml68UhD6wRAZJ7mtdXIlKtMCc26JeIBczJbBVlOcFn5ufXktBHYFJRF/bRcLOd+1ltAa+FnXh7Y47tk9tbpwbGUdZohCHFYzNkpjSBixSH3ND03tCHlB2vCDHX7l7t0yvkyq9JmxAxv2KFkiEPrBEBknua+n0ScDwkr9Dol4gFzMlsFUMM+Edcab/ctG0cCHOzvepws537WW0BryYngUFNV2ND21unBsZR1mjoOI/l4KNd8ayLE2NSDATa0IeUHa8IMddHFFJtTSuLpIpLz3+PbS84IQ+sEQGSe5p5Bb6afthBRuiXiAXMyWwV33r5ce1KypPoO9eV1w7NbHCznftZbQGvn189neZelNHbW6cGxlHWaLxrTRMnRJOkDsMHTjZeXWPDxZ60dJOq58gAE2ekCjgsAMq5V9IKK+ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwuaYURLz4KbxwaSGHgNq4+ZAYIUgJKG/kbXGD6Zcp3m+RYDBFYuiF25bBbIUsar2X3l0deS1AQ1vEPbf7OI4stfbVSTH+X6hdKjh/7YApD9Ekj1xXZlnGHbeAEZMSJ4rbVQRM3Gc+S9egGtkf1mj3HKliZFPd+JzvjvtQTrroWfUQDKuVfSCivq03NQQFCgtDwfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctPT/IbYgO2uVnwg/IMu6/6X3GFc3FY3ZPv+ggUqaEPvXOGXMNJvXM3NonL3dWzRS56qn3s1umVquYMjOSvzbZvqzyrBAT3vQQ8OZ5dJ6G/WScFeWEM86CNs9/cmJsZL0oCK5Nw7o/HWScFeWEM86Ns7gbstDN5asFAU5C9nfKLolAfj4G6tkBC4FyK6L/AUHEvd2ySFhq/KAMRtqFOjmeiNuPW/CDp0x7oTl03mhREEEyoZAjAoDKP6KF+0082mK+TC2YUt5PYsIxenHftXO+xNtcbkLGLjp1WBz+fQys9ceXkISJnAR+dK/+s2YPEJYgC8UwPsxZTXrMEQnCbaDyJ7st+o4ixz/JyRd77vY9tvsIoaBB34iQePKFnQHK2Y9iri0bUW3lRGDR4XXyl3Afl5GWqPsztuXIigbRpCe1ePuFEQpJW7QTCRl2xo1KzWeIEWMn685D4r5MLZhS3k9lOcgM1yvyiUR6IvRtsBNB8OEt53KmNdrRSI6dQzrfsnpTdHK4QUqaZB84UJBNDhoFx5eQhImcBH50r/6zZg8QlgjcDJo9n9bZNysM0H/beDDKv9ENpWIf9BboDWT8dzIxUW+myAUVjrKqyDWSNA+o38nJF3vu9j22+wihoEHfiJagpUwam8thzoSNNC4bGfFXLBbzwYjMF7LTGR1s2MiycftDjtC/XPqm+wihoEHfiJagpUwam8thyHT7+7+DXSRFXFdmfLZSgZSD2I43Q5NTryX1Fjn5Ez7AEuZ0tVGH/EW9UgCDHWybhoNxvyQ8QW1lSVdNvXF73h7boMQ9kCHfld5S7zHloRbZcuiL3kkrXAPSX+5s87cFdwukwNlc6T+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3eCMgS2aQYlSf8lVN2ZZgfoxCFMy3ABQrty9SLWj9MahDVHhRSEtqXSdRsYz5JZBMnmvXHN8NcKUL5H3JR+gnQZvxh72Y6FA+VPnyoAOCdrJtrrWYvsHNnuoeOzclB8GBz+GzdbA8ObbmNcw6kzQbxjhI6oKFdIyvt/5Fw87SHagCvMDmp2o5MfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvGsVqECQ9P1fMK16swBak6aDrV0SaupysaHlTmKsmfKgFg0CdygaSDdwS7MS5Y9KycDP+1jQ0/h7dx6Orf8695LKBmmOe67LI7T6JQ+hpNEaI0UfY20Pp+SJTlKIewzw5uGqxOMXTsGOkOdenP1NYvWsxs9IP0pnBPCIRv2FGzuAX1AASdlQAAEImZiMR65mYoQ+5TvnXRb50aJuwOjnKObmNcw6kzQbxSApTvk90uZxuofeqqBDYt7hrgqqBwcKPB0ccR9Vzx+RzrYuMgECcZwFgsHfuuaTBKYijmPzIIkYlZunU3QS6KOiONu6+bwfrKhw221tyLQozD3wu+7NmPgbd5esuM2q0cAJOOq9NkjSZvCCGiKac6wFgsHfuuaTDAWCwd+65pMHYbNu+Fr0Eyhu9aeTRVvOydqFMDJi9aoPoCSGYvHeNHOMKA1BJV2ZMT6WuC0VzVyqI4QKHmoIxJ60aQLEfXaN1SnllT1OJZtcBYLB37rmkwq+9yLK/bVb9tiIMdLAg5rKU/hvYt1n+EpgZPCiXftU5Nz7Ynn829T6mQRsCW0lNd5pNyqlkQKKfhwEYlgJb7LHrocQZzasscXA1PhK76CYC/dP79Ds9NObQtn3CtrIhnFhn+9MKSpcr7dQJDr86z2huofeqqBDYt7hrgqqBwcKM5ITC48ak19Q3mfW5gzSZ9FPKVr8xhesRKYijmPzIIkYlZunU3QS6K5dEl9DCehMRqD2j1XTd1p4zD3wu+7NmPgbd5esuM2q0cAJOOq9Nkjf/Ja8bBSafimJxIw1OSzVWvpHauJwoRp3YbNu+Fr0Eyhu9aeTRVvOwmDhfaPCP9I/oCSGYvHeNHOMKA1BJV2ZMT6WuC0VzVyqI4QKHmoIxJ60aQLEfXaN2eceORd2EjlsBYLB37rmkwq+9yLK/bVb9tiIMdLAg5rP+m/qXdPk1DpgZPCiXftU5Nz7Ynn829T6mQRsCW0lNd5pNyqlkQKKfVBRUrA6q0OHrocQZzasscXA1PhK76CYC/dP79Ds9NOfgEO8eC8wxdFhn+9MKSpcr7dQJDr86z2huofeqqBDYt7hrgqqBwcKM5ITC48ak19ZE1UvcYM7BXFPKVr8xhesRKYijmPzIIkYlZunU3QS6K6fIVdifx5rFqD2j1XTd1p4zD3wu+7NmPgbd5esuM2q0cAJOOq9Nkjf/Ja8bBSafi7vmOgFb8V5CvpHauJwoRp3YbNu+Fr0Eyhu9aeTRVvOwB3etOUjP5QfoCSGYvHeNH2v01L/YnV47EHR0jURoJ3C7GKcYkY3bf9P2w1qjfMOTpDnXpz9TWL3XlaFtbYtPeH5vL4yVciF1y6VrBZqP2W/GwAIE0kyRpdyvNX5JepqHOgMYqSUM+Q2gZM1la6Pu45w4ejLjiCSUcu92WgJjSbGCwvJtFTmNtOSEwuPGpNfXnGTYGKRPSm1B9Yd2pZFfQSpFTj9M4F4rWNvD+U/2X0pAEB4y5lxQjZhXzxArgHaCNk0KoTqVA4Ry73ZaAmNJs1lrf3MAW+LBUjSEEMa6eRm+MPjUmAcNOYEZ1rj4dO3bWmH0QnDKBioTGSR7/wOaPOB129t1fowXsfegtNRsNtu7mlytUNHbRfpgikR+ILxdGpjsL3U4MpayECM1hQM845mw8QDXyQrEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvDvs4X13is5a+X2U2Sr4h2tfpPQ2kXFtYhzzdEPSJT5a+7grw2Uuih50Nrz9FNAQEPr2LbsPFQc/85hXRHi13qvfqYTuVYKVl0u4Abt8zT7TWUWgnEYxS+SkDw5m5NjMoLYT91JalH4CMgHRiT624YyqKLF5ZhqmfZtLL+yybWpx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7zhC1rRWGiQMZC/dfqF4dQAByi4Y+C90Y1qeF/3xLYVjbHasb8nNKb74TviO2/cKLXyY4p3wSQhQun+fadIqyRtOCB1pVP/YIVe74nJ6edzid0R9SwaTlvBBQDkg8Q3rOQ9zsKk8AIidXQoFv1vZWB532mKjRs8AuQ9zsKk8AIilgAHyd0stRO66YATYoWs0DNis1qs5hxN7RtZNGyzZJnymAz34CM8TekOdenP1NYvWO0HZMQy281p35Zthlj87WgxwPOa+bCZuX3CwhwA79owICxouRz2wyCL0/lDTkTEO95IiZfXcDT5dLolfq/xY8EfppvqcUz6AavDmDTROJFI+ewdy3Rna4aELzFZeL6+QHV5xeL4xickIDeNs7bqVjAgLGi5HPbDIIvT+UNORMQ9sRnqdohw/rInvCB4XJTTAWDQJ3KBpIOfoAOLnMoIH62LiTlmATyVMCAsaLkc9sMCLmfIM/UTQBwoQZER5Qwea9CKQlY8TsIdg1suZ9E6/+FUC5JyaHrvXgkDBylGzbDVmaIohTeKh69QIF4Myn71WIIAIds2MSqzpuBjY2VybUj2QowWZ18NQhQaHWyXaE8BYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h4oak6uU6IRXG+n1s+QzRGCUzsVX+qjJ2cFhRLHtr5z2AY7DohsgeLJbslkf323799Xhyp5wRBnnlrD/BzgDbunDz5/Wn/KoAGJu0vDWy4qIlM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw+pd036qvfaAzkhMLjxqTX1Kf/V7ycg6kNxX2xf0wa4os3NonL3dWzRF/O8s64DUvK6maR0RWksW21F32Il+s4UTWToPteyKxE4Fz2wTKAvWmnCcfykCW93XgkDBylGzbDVmaIohTeKhxVrctsH/OmEWIIAIds2MSqzpuBjY2VybSXbC0NoZwHP60aQLEfXaN0is88qvK7zdsEfppvqcUz6rR508ZTGndGpcg1sRIlPCWvQikJWPE7CHYNbLmfROv/mk3KqWRAop9UFFSsDqrQ4tprO255FFziUzsVX+qjJ2SOL0yshwRnP7EthwE8LM8XC4OEyxUpTD4eiwO9xP+5his56PQm0umWY3JjE6+3cOPWqEdoGn7o3Bj1IlHszAVRPxOboHLSP5CvpaDe6pRF9Jeg+iExCMrmtHnTxlMad0RKYACBo8PvF4cMmgMS30D11ZMnUofCOemHAPT7xp+aotGwLZityvxOKIOYTGdbNXiBkf8+t9vrD1ZmiKIU3ioevUCBeDMp+9ViCACHbNjEqs6bgY2Nlcm3rOASvJyBn0DkhMLjxqTX19MpFthW8Fe1CFBodbJdoTwFg0CdygaSDksVqJxdxStwOGp1msVUhnVRWHJYQ/HeHBj1IlHszAVRKkVOP0zgXigfHKEpWtWA3/qi9tma2Ui4l6D6ITEIyuQGrw5g00TiRXBfVVxFmFh/mk3KqWRAop9UFFSsDqrQ4WGMfX5IfxBasPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPXVkydSh8I56YcA9PvGn5qi0bAtmK3K/E62EIDuudjQfIGR/z632+sPVmaIohTeKhxVrctsH/OmEWIIAIds2MSqzpuBjY2Vybes4BK8nIGfQOSEwuPGpNfX8WktWje8BUkIUGh1sl2hPAWDQJ3KBpIPhQdEXYU/SbPKYDPfgIzxN6Q516c/U1i+LxqgEbQGiQuSOCFwaOINhKN+o8Y3BzwugGYbnhsuuELnQQQixnI7IERS6cvX3J4AUiOnUM637J+dceKXRUJo8xj2xuG2LhpacaiSB0pwUU007V+j040uDhauMtfc3NEsBYNAncoGkg5LFaicXcUrcOB129t1fowVtRd9iJfrOFOjjhCoiburJGOc+HiWwXb2UzsVX+qjJ2SOL0yshwRnPTkGSJu/s69jC4OEyxUpTD+dK/+s2YPEJ8V7vSBv/Nd8BYNAncoGkg5xqJIHSnBRTmm20Jd5iXPesPWg6FSenyHeAIBdpfm+x/0ImPkJmWxowO89C+dp7ip/UvLitUeOwFIjp1DOt+yfWS5qOPsKoa+3EeOPoqNzDMDvPQvnae4oCLmfIM/UTQNqTlZfCjsNca9CKQlY8TsI4MCPTRacQbHK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiYrwj6/ble3V20GmV5DU87zvQ25D4d2Paby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMTsglqTDpbG9sS5LPshKV/6vbpM1DWlPc/G8MS9PnKJHV0KBb9b2VgaN3SXsBwel7LRhPgGFlt59Crq+9aP37oqDXxlkXGyt9Yt+40/kUJWGf52OwzgI9ts8TuxAbbvigaeSEc5Yud19epfUFxPX1+l5VLDx54rUFE3tygC005pDTkS24pPPLGsKC38YHLOwovufeYUOXH4uiD5Y6BVN2PyRClOEIV4iy8qkyybZPDJhuI6d4fCdOI3GlKF/MfOq4vufeYUOXH4nvqzdifKM1tAMI/ezIQEtyzxO7EBtu+KKWqYVWBnUw+mBdAEbtIgEAUcHXO09MXFFWb87ctC+RSiU5xkatEkaTM6GC9NLPeIJGMZSUNb0n0zasixnaPUTKGhC8xWXi+vkB1ecXi+MYnlDYYvbSvdRqAE7TNzfAu5YNWBUbEQksWrmXAkBhazfSoNfGWRcbK366vse09xFj3BiOD7Cu0vs4CN0nQxNKM1osRvXKU+PMJW2Nsp2cpbugX4gsx3pBAj3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4uljxQy0PgHiVynIiZoshFJTuU3JkJFIp6ZsnxGchEBsqIRi0VMcAPCWGbSapYwqcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMjmJGmnDlH5ffTv7ig9fqTuvCep1L35Qxqjc1IscbNw5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm9cU6E4LOfuh6/71/BcnnXOaMqCF3iWxbsDbvaSa+SnqXIk1JlZdjci2qYd2EgdKtDQUFJSyD4MVNhDOo5YPnV/ML3EO/WvzNjhwIGUocy7GoNfGWRcbK36F2IlEkBcGdwH2wOq/fkXM0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm1cF9VXEWYWH+aTcqpZECin4cBGJYCW+yzpfGNFm6ZkuVEJZt5I6hoN5iRnMMMFpPtmPJKZ4to+yqF2IlEkBcGdOBc9sEygL1qtMRfD4H29qDQ68/3TNPUeGmM340wuvpGzpuBjY2VybVwX1VcRZhYf5pNyqlkQKKfhwEYlgJb7LJZWH16/+TeYenPTtAYOt1ZcF9VXEWYWH+aTcqpZECin1QUVKwOqtDjpfGNFm6ZkuVEJZt5I6hoN5iRnMMMFpPtmPJKZ4to+yqF2IlEkBcGdOBc9sEygL1pGnIbMNLh/CzQ68/3TNPUeGmM340wuvpGzpuBjY2VybVwX1VcRZhYf5pNyqlkQKKfVBRUrA6q0OJZWH16/+TeYenPTtAYOt1bzqGF3/y/2hqcZNCgGlPXmbglCZfq9SqOvnYUlb1kWV1eYB5ioJUYgZjySmeLaPsqhdiJRJAXBnTgXPbBMoC9aNB+Jl5TV3RF2qGJ/T63OOGY8kpni2j7KoXYiUSQFwZ04Fz2wTKAvWo6LZStoIP8ydqhif0+tzjjMQT5ndyMiZ8xkVW9vDPYGV5gHmKglRiDAWCwd+65pMGUmuIEf6izZHylZdJlKPU7AWCwd+65pMOeZUFsfq5UAMKVufBmMpuTAWCwd+65pMP9YOIVlvcdJHACTjqvTZI0mbwghoimnOkv8MthD2qTcwFgsHfuuaTChdiJRJAXBncB9sDqv35FzVbujO5Wg4siIil5J5hTKsaWoJuy1vbXJGGu+3/L5gB14Oyl8S5kmyhq/Qzj08fGxKhYlwlva71cKN/W0WpqKosqJ+k5q9hXVwFgsHfuuaTBcF9VXEWYWH+aTcqpZECin4cBGJYCW+ywrn3ZFGlK59lfgGehlBGJjKhYlwlva71fDZBJb1raC65DRDzKAm9d6pAc/hVAOtpjJUu6i4j6R0UqRU4/TOBeKB8coSla1YDcgaJXbcfIaIcBYLB37rmkwsUJYN6b3gXv9odWZ/Pd0wutGkCxH12jdb5Alwbg/16pgpYxBgkNjhUqRU4/TOBeK0V4Tx5FIIGp3fNfKtXeOasBYLB37rmkw0TtSsmzc9o4qFiXCW9rvV2GQTlOpCr5UBXWszM5IXVeQ0Q8ygJvXeqQHP4VQDraYyVLuouI+kdFKkVOP0zgXipTnmDH7+vkS854vOQaLL0vAWCwd+65pMLFCWDem94F7/aHVmfz3dMLrRpAsR9do3ckktFNyXochYKWMQYJDY4VKkVOP0zgXitY28P5T/ZfSd3zXyrV3jmoeZa/KEJx66PS8G0PpPuB9abPF51YYnoO0bAtmK3K/E26509W9q/53qDXxlkXGyt9mPJKZ4to+yqF2IlEkBcGdOBc9sEygL1pGnIbMNLh/C1W7ozuVoOLI9zvVG0uYXoi0bAtmK3K/E2kWABr1bcQgwFgsHfuuaTAGPUiUezMBVEqRU4/TOBeKlOeYMfv6+RI16IvKftbJJXD3jZufTTGBHmWvyhCceuj2wBYjwj/QGuzf2+SW3Kh8wFgsHfuuaTDdiU2I7GLQGKg18ZZFxsrfnyMGKRvnXNUtmJaBJcfH6hD0ExRs9ghbdwwqZv6zyy6tMg/TH8AwMJuwpfyRpuHUTMzqNaAeQE0LLXl/6S7X0VK+LNInXRCt8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWXsHhv35Z6JyYPnDJ/QYHRSmqNzUixxs3Dl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGb1xToTgs5+6Bu/Lsybc3KEIPEEOOs5sYJFhs+T6mvC3Bp5IRzli53X5CRqz7/gFKofUxVuCXS5Y32Pkite4rtGKQ9XKZKOL02NVcWq422EsmDUy0bAGUzIwtYC11BuhLU0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek7xhA+nGH43aDa5c70WeNYpk8rBnyA2a2eY2Nk+uxLPvcuT6SxIGKL0YNTLRsAZTMjC1gLXUG6EtTSc3R/HQ5ndZL+814w1rJaAnC2OPa2fiuxAJYl05q/fDug+TuqWkX/ruAsn4JNJFag18ZZFxsrfj82zPk7UNQ+/EUKWXiWm56g18ZZFxsrfKap2DOjhkd3+7du2loyvwMBYLB37rmkwoUe3BxAoiF5hG/Dvi8gsq8BYLB37rmkwRfOp6ip8MKHuGuCqoHBwo8HRxxH1XPH5CAkvP3UcHknAWCwd+65pMHvZzLAQalyc04oKQ+o6teoLT3Bzvh6oZhxNtEOd6XfNwFgsHfuuaTD/WDiFZb3HSRwAk46r02SNJm8IIaIppzpL/DLYQ9qk3MBYLB37rmkwSPZCjBZnXw2Iil5J5hTKsbtZK8yRV0MzPFxh3NDvXjbtxHjj6Kjcw5DRDzKAm9d6pAc/hVAOtpjJUu6i4j6R0UqRU4/TOBeKB8coSla1YDfzni85BosvS8BYLB37rmkwf0h/5H1vCppX4BnoZQRiYyoWJcJb2u9Xw2QSW9a2guuudS5Pr3/gXDkhMLjxqTX1Kf/V7ycg6kOQ0Q8ygJvXeqQHP4VQDraYyVLuouI+kdFKkVOP0zgXigfHKEpWtWA3IGiV23HyGiHAWCwd+65pMH9If+R9bwqaV+AZ6GUEYmMqFiXCW9rvV9FUcAzFf15drnUuT69/4Fw5ITC48ak19fTKRbYVvBXtkNEPMoCb13qkBz+FUA62mMlS7qLiPpHRSpFTj9M4F4qU55gx+/r5EvOeLzkGiy9LwFgsHfuuaTB/SH/kfW8KmlfgGehlBGJjKhYlwlva71fDZBJb1raC6651Lk+vf+BcOSEwuPGpNfVG1iRz8J27qpDRDzKAm9d6pAc/hVAOtpjJUu6i4j6R0UqRU4/TOBeKlOeYMfv6+RIgaJXbcfIaIcBYLB37rmkwf0h/5H1vCppX4BnoZQRiYyoWJcJb2u9X0VRwDMV/Xl2udS5Pr3/gXDkhMLjxqTX1A2GjIfMR/uGQ0Q8ygJvXeqQHP4VQDraYlxFofANwh+ZoVOelkqJIZ8BYLB37rmkwRNZGJa2HJb/AWCwd+65pMJYTnZDwGLlXkNEPMoCb13phZozdt25vcB+pBQUd/IzhvoiGCRllu1SRftjjGWJHTS9udGlOlsAWEd9TOS5JxzRZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3PaQRqM/EDxFb919yWa4zkk4Feq0u3fyx3Mf7t/Frf+I+yxT25U6A77bbkld5sbnJxz38vshk4xKN+o8Y3BzwtEVRlw+CYWvdcB9u/qWYJQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LuByd/PverQFaqS53zBtL8hnLXdIfXO1vNpQQWf5HvYU+eoa6rFNJu/QSH2YZFW3xFeE6ZypoaFfbWmxzHlS9XPhY+xAPB4d3kggVfaYiee0Hir08408efyDyVW5fvLJZWeKdmTkEiU0K2xFvcFFIVwDKuVfSCivq03NQQFCgtDwfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctPT/IbYgO2uVnwg/IMu6/6X3GFc3FY3ZPv+ggUqaEPvXOGXMNJvXM3NonL3dWzRS56qn3s1umWY9BCSCKyXy1gWv4xlzFUdpfSZQ1rylVvtG1k0bLNkmZ5RRDns/Z1n8DwKRTyX3NLC/Akftdwe10azJJLiCUOBtfJjinfBJCHC/Akftdwe113lLvMeWhFtzf48rPx8NWywUBTkL2d8oqYKtC1om99O8p7aAH4eqChGpjsL3U4Mpe1r32W9EobICqD4nUayamL3FBVXLnrdhYLkAzBtEkvpXgkDBylGzbClaqHQ6HYhZSqiwbt8jjHaOLU5nnUugAcwICxouRz2wyCL0/lDTkTEGB6jBl007Ic8OcUvtKIUaMtTNNKBXsMOsfEoSEIM7uVeCQMHKUbNsKVqodDodiFlyvZhKluyThkfcsHapQOQ0JTOxVf6qMnZwWFEse2vnPZYXgyXk/raPV4JAwcpRs2w1ZmiKIU3ioclBrYPaT/VkOxjbVPe5ExNn6ADi5zKCB+lqmFVgZ1MPmYCYVHcspp5nRpRErudjt6lr9eQQZ3jNxxHLifkb0sGc8rFJQKPIgPYMn+n/hOve2aUWvu4AhcMlM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw9Vm/O3LQvkUuPqFpjzn2ScrD1oOhUnp8hO7JRb/x7EOE1H72YelCd04d25Ov43oRL9fWYL+PrUhR2DWy5n0Tr/C09wc74eqGa5Dxmmqoeuzaw9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9akY/FF8AzWjk7vOH1LLGLR72ncro64s3bFg2Or5Tn2CxQlg3pveBe7Uw8m9dq1DWJFFahibdzyJxztYHphKvOAIuZ8gz9RNA2pOVl8KOw1xr0IpCVjxOwjpKB/H5OuK2oXYiUSQFwZ04Fz2wTKAvWraSExDNWfYfSeCdmyU1jT/P4IOPj2rD7GvQikJWPE7COkoH8fk64rahdiJRJAXBnTgXPbBMoC9aRWpniozq7B5J4J2bJTWNP8/gg4+PasPsroTqTSgJi7T4SW4WqIeN7/ql0b95iYOXudBBCLGcjsjAV/O7+mBoupwX0GRKw5bQvt0W25erGIQD9tcnMj9RLm0x5H/lly5vjFEgqd1+mTahIXdDSvqLtivkwtmFLeT2EhfxS9iprzW0bAtmK3K/E4og5hMZ1s1elM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCVnM1cGH7eekB8coSla1YDcL/crejE9lKs3NonL3dWzRF/O8s64DUvI4HXb23V+jBW1F32Il+s4UC8g1E4M0/TYqFiXCW9rvV2i5rzxk0Nib0+q/glx2ZgvVmaIohTeKh69QIF4Myn71WIIAIds2MSryTKIkUcCMHXNszWGG6djIb4w+NSYBw04g2hSnxXHovK+HjxaB4B74rR508ZTGndHwthhZvKXBo2vQikJWPE7CK+TC2YUt5Pbl1Zp261EHWiPssU9uVOgOPc0I368GozjVmaIohTeKh9cmIYqSm9q57GNtU97kTE2caiSB0pwUU8nghxtgSf/d5pNyqlkQKKfhwEYlgJb7LP2etmX0678cnRpRErudjt6lr9eQQZ3jNxxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnP2h1Zn893TC60aQLEfXaN3EjcMxCv+bMgFg0CdygaSDksVqJxdxStwOGp1msVUhnVRWHJYQ/HeHQW6A1k/HcyOhdiJRJAXBnTgXPbBMoC9aKl0Z8puAdIOsPWg6FSenyHeAIBdpfm+xxvZrfAFJ45z9odWZ/Pd0wutGkCxH12jdmTY7f6kcrckBYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h0FugNZPx3MjoXYiUSQFwZ04Fz2wTKAvWjWK/7yXhm8DrD1oOhUnp8jqbdmcoQYqPFgZNuL2sSDi4cMmgMS30D0UiOnUM637J9ZLmo4+wqhrOSEwuPGpNfX8WktWje8BUjA7z0L52nuKAh7GJdVdRXcRgZf3KU7i+Q2k7OKvdEGVjFEgqd1+mTYLInudpCvlYqwllGw4+2H7LtIzPkI1jT+iOE5XnmHnvQrc4luuChwCI/Bt3qO0PQqzxO7EBtu+KOOjsLeQ0/cg0uQfh0LiyLUvufeYUOXH4puhHwoq8y0TrGWufpBe56aJxx1WK5LYoJGMZSUNb0n0yMokQ8Xzmo/R8jzVqDLOsT0WfHBgXkxdQG4QiHntQdTsiWL5M7qTAMr2YSpbsk4Z+hGhqX5cvLANULrWKsJVwe6+0ZjaPn9Bb3XN+LvwPDptxbng338D5C+595hQ5cfilVUL9qNGJFcnlvZGpiniSFTszs8iePtfjZpRn0I8htYK/0QP5j9MMbZmjHDNp2DBqDXxlkXGyt/NVaB58sH37Se1DLEygSLqv9281ooBjDZNR+9mHpQndOHduTr+N6ES/X1mC/j61IWoNfGWRcbK34VTxHkWmBnXfHWjXjdtXbsH+7JZe9gI3npWtUmfjM5zs8TuxAbbvihKkVOP0zgXigfHKEpWtWA3w8alrUQHJV4qFiXCW9rvVwo39bRamoqigEqH4O9/vb9NZOg+17IrETgXPbBMoC9a3Cz20f/neMFLsOcyU709DetGkCxH12jdUSVeyZa4Joz6fgaOMo9KuioWJcJb2u9XaLmvPGTQ2JvbnYP/owPYhW+MPjUmAcNOzdy+6tPm5P2oNfGWRcbK3yXbC0NoZwHP60aQLEfXaN2PqZ3uwiHxwuaTcqpZECin1QUVKwOqtDhPs5nBXQ7LOMJ051v7yRlxPjDLnEtHk9ibxtFos46qE+I3sv05ME8NsUJYN6b3gXu1MPJvXatQ1s8ISqMdJlEC6zgErycgZ9DtxHjj6Kjcw7/dvNaKAYw20TtSsmzc9o4qFiXCW9rvVwo39bRamoqijkGiclllg6JKkVOP0zgXigfHKEpWtWA3gLBW88bFphmxQlg3pveBe/2h1Zn893TC60aQLEfXaN0W/ru0ZOKHVaF2IlEkBcGdOBc9sEygL1qGSh6bgqv4AmDUy0bAGUzIFb919yWa4zlvjD41JgHDTiimEGmqLZu336fLQW943BgqFiXCW9rvV2GQTlOpCr5UNyB9cSD20sRcF9VXEWYWH+aTcqpZECin1QUVKwOqtDjU+kUR+qnOyP2h1Zn893TC60aQLEfXaN3rsKOrJeaVAYNWBUbEQksWYcA9PvGn5qi0bAtmK3K/E26509W9q/53OUb99pwMO7pvjD41JgHDTlf3sBC6UUi8qDXxlkXGyt/rOASvJyBn0DkhMLjxqTX1/FpLVo3vAVKbvgjOrX4mneaTcqpZECin1QUVKwOqtDhVDUsmMpH18jokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyt5JVmvTzF7rqi4g5nKdTjZ+E8U2gV8rJOBc9sEygL1qbYDmy63yFvKasjIyYzneg8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTIGEjBijipE1KkVOP0zgXimjQ9PcbIOOVhX9ZTeqm6mvtnfogXPL9BR8gtxiLTTHi520j/RR5GB1kV2RKeFDdt3IStq4WjC5mT+QyoSnr4KnhhQd5G/Xq5OYiqiWWtCZqWczVwYft56QHxyhKVrVgN0YBtSUAOeeaQIaAy+tSTHE37Nk97b+6rp7WNoaMRI3YKhYlwlva71eaGGgmy74fKsNwP71HnkU4bPz/c6/JJ/2iPRAJAhOGHlo1LtHNujgmb4w+NSYBw05Qs5TED4fZ7zSc3R/HQ5ndZL+814w1rJYvxMuc4I56TqgxK8NU4X2xtGwLZityvxMhM0qVZ/PNsLtwcZyZxxott1OLXHeZwhgETOWt0KBunJJ3ezUKUQNvZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYcQr3mv20RaxC9k6h5Y71X6F2IlEkBcGdOBc9sEygL1r6Afunv0u1DxE7nNp8sszc5iKqJZa0JmqoMSvDVOF9sbRsC2Yrcr8TcWpboDb4ci05Rv32nAw7um+MPjUmAcNO2ZGfUYU51f+oNfGWRcbK386FAbo9HW2L60aQLEfXaN1vkCXBuD/XqqF2IlEkBcGdOBc9sEygL1pMnazpShb/KpflSbQ/7r+gNv1C5IcM117MQT5ndyMiZzlG/facDDu6b4w+NSYBw04t9eqo+YceYykJuMch/Os1uWDl+4FOsmiJRkkmMiKGuDgXPbBMoC9ahE8I+GjfVBQ8XGHc0O9eNjkhMLjxqTX1RtYkc/Cdu6qQ0Q8ygJvXeqgxK8NU4X2xtGwLZityvxMhM0qVZ/PNsDlG/facDDu6b4w+NSYBw07YWAuy43ftn6g18ZZFxsrfrTIP0x/AMDCDPmhAtpi4ZmsezOrWWHiu9orqZYAgHpsdWsUzXETiNzkhMLjxqTX1I6uWZM4WiPDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+XJ3oG7RzGOQSpFTj9M4F4oHxyhKVrVgNzV7zIVb1C5ZYdrvGZRgZ1BvjD41JgHDTrPEKKh2QiyNe7zqVFgic2tyzBRZimRsFTgXPbBMoC9a/VUeKNysqlvszYnLau54Rv2h1Zn893TC60aQLEfXaN00d3mb64F3741bY5YhZOjlOSEwuPGpNfUDYaMh8xH+4XujoQl/csKl7P9PFRuz6r5vjD41JgHDTl4pqn/CERX0QzAT0rgnVAh2bHqbKgtnFHMj/CwJLSkxQofVGkA14n9Qxzx4BSYyoB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCwDKuVfSCivq1Uq2Dto8OhUHcHIYr9UE6eIrdrTIszmZFBAObT4XJblwKtGsbPg3isU/BOF/jE73fkpwVdcZXA0sU3rguAfkIwDKuVfSCivq5UPY8o2c6sP87xs4Igtz+ft/5Fw87SHagCvMDmp2o5MfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvGsVqECQ9P1fMK16swBak6aDrV0SaupysaHlTmKsmfKgFg0CdygaSDdwS7MS5Y9KzSgIrk3Duj8Y+YStKhYVkrvWyKpZe+sEzXqdpuCbaDKLCOjqeEmbrfNg0ZOIlCNdkv94TlSlGhCUZ6CCfYNpaWND5/1YD7AQ8v94TlSlGhCXjazt+6rrfB+Ko8VlHmIOiCeBlNilgh9jJakekrNK1qQkb41xZ0+zJ532mKjRs8AuQ9zsKk8AIidXQoFv1vZWCiB9WB76XcZLBQFOQvZ3yiVjW1fM47WbuugXT7eLWvflucMDlUgErFND5/1YD7AQ8v94TlSlGhCS7SMz5CNY0/93jaDoJOdeiCeBlNilgh9kVxXVWyCsBA6Q516c/U1i/bO4G7LQzeWrBQFOQvZ3yipgq0LWib307yntoAfh6oKEeVRRrIbJxinwOmAujGGLoiTYgnaEY9ipwtqEPKcLSowR+mm+pxTPoBq8OYNNE4kdKDEt0ZXQvCabaYySE8y06sPWg6FSenyE7slFv/HsQ4OyxQZ13Y28c34Nvk7H7rocEfppvqcUz6AavDmDTROJFklm0yLGFEkHLkwrR+v8SSp3F2/KZDZS3sxsfasFm1PlKUnG7T12N5i0kWLnusckK6maR0RWksW21F32Il+s4UEtRfj9IyqtVcV9VAj7OHu4t9mDkl+tWoMZPML60V2LXsY21T3uRMTZ+gA4ucyggfPwGopGN5FQ59toKzMgaeL57z2bM2B/fLTkGSJu/s69jC4OEyxUpTDwH9bAy+mJtKg5WcJPKVWHNyfFt1tmECVnVgpvDe2lFKHEcuJ+RvSwZzysUlAo8iA3wIO8c5E+3g+N086PV5FEsrKQvEtQJT6s/gg4+PasPsa9CKQlY8TsI24X1LNvxtz9Xhyp5wRBnnJWtTBfHE+fTDz5/Wn/KoAPfIsUQ0jlrJrD1oOhUnp8jqbdmcoQYqPHPT6yNUvnsS4cMmgMS30D1qRj8UXwDNaFHHyTQ0RZGMUIJyZoFUkp6N+6jE6JHeCzQ7e1k80QpnH0km0H4E0GIpim5dgZrhdGvQikJWPE7COkoH8fk64rYMHZNkdaymPSsoshgLutmaNWYnM+lVTIQoJyPBu6KPyEx7gBn3LDygw1IMUJ5zDzvyntoAfh6oKPhm3//nFZf+rZk23b3pB/JUBKPN3GUEFodcDF+PIeNo6Q516c/U1i/RMgNHSLmAHm3gjXOEok0SFaxWXSQHf9Gev1XJ64vHB4bvWnk0VbzsKcFDnmYTcQFH7YX+0q2tls/fgeW7+hConrgr/BC+fs6IhdTrbbAMB1RWHJYQ/HeHQW6A1k/HcyNUVB/nV0W7J0HI9aDL4/wTg3EgxiHOanvhwyaAxLfQPRSI6dQzrfsnEjbJKiHgK4VH4j/NjnSpDzA7z0L52nuKAi5nyDP1E0C+H3zUE+AHXrcGtZTTW0lmnGokgdKcFFNC17pbbRwO+JkLg62wnfIEMDvPQvnae4ogi9P5Q05ExEFugNZPx3MjNKeerljP17mI7fwuiHXfkQFg0CdygaSDnGokgdKcFFP4MMNVGwB+ioG3GviY1gpyMDvPQvnae4ogi9P5Q05ExEFugNZPx3MjvAxOxpSNoEDKr5wcIRQebFMzMTd2VbLAK+TC2YUt5PZV2JP4bUIOyVuWK92u6/4CPc0I368GozilaqHQ6HYhZedK/+s2YPEJSpKqD9UHtEFIvXN9qra2Y4jt/C6Idd+RAWDQJ3KBpIOcaiSB0pwUU4C+XPtIrJshuwWlpXTkn4OsPWg6FSenyHeAIBdpfm+xzDLAEHanyPOxbQFtYIvNeT3NCN+vBqM4pWqh0Oh2IWXnSv/rNmDxCZIHAVMsU3P9yq+cHCEUHmxTMzE3dlWywCvkwtmFLeT2tABR3yk+d/+ZC4OtsJ3yBDA7z0L52nuKIIvT+UNORMRBboDWT8dzI7e3hHkj6OA7Dles2xfXwOkRaygtE5naOViCACHbNjEq8kyiJFHAjB1pQKpSyhKwabASKP3W8lapkoejOOHQ5KMomfIY+Y3JZuHDJoDEt9A9FIjp1DOt+yeysXhkHKmrsDK32yL1KO64i0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+Il2Uvsf3ICB5f3QKvhcCLHPMZPML60V2LXsY21T3uRMTZxqJIHSnBRTzM3XQzV7lJmQa5o65mLcbp64K/wQvn7OuRh3QlVe8E7C4OEyxUpTD+dK/+s2YPEJogDrY8w0JEg5NouTrV/Nc1TM/LO5RPzdJ97wqLFSjbNUVhyWEPx3h0FugNZPx3Mj2vJWBwm3MZTYg8PKAP8lIBwzO7OLXCoB7GNtU97kTE2caiSB0pwUU4C+XPtIrJshahmfDTGjj9OeuCv8EL5+zj7t8wpOtE3LVFYclhD8d4dBboDWT8dzI15pOM2U1ORYjUonnWknetJmfPrlWAGhChxHLifkb0sGRVxgon0onxx5v5RzOTsGdDfRPHCarIS0Qcj1oMvj/BPnkjRpdXAmkuHDJoDEt9A9FIjp1DOt+yd5D2rB2KwTxupzYTLIoYhdytYQDdKpC4RIYQ4pQCMNLSK9zEzIsSkd2wPHIWOU7dznR+tQd3WcZavvciyv21W/UlBsfAG9u8PhqrQcXYw6hpxqJIHSnBRTX5dT1uFDwVD52yY94aShO4+ECzyoDEkO7GNtU97kTE2caiSB0pwUUxJ4SPDkCA54Qn6cdsG0uo6PhAs8qAxJDuxjbVPe5ExNnGokgdKcFFPbsntuFnlMp/nbJj3hpKE7j4QLPKgMSQ7sY21T3uRMTZxqJIHSnBRTpp/8oKj5YIhCfpx2wbS6jo+ECzyoDEkO7GNtU97kTE2caiSB0pwUU5+SuzlDLH2bq6HeRI058bqCNw2vYZ1NRI+ECzyoDEkO7GNtU97kTE2caiSB0pwUU5+SuzlDLH2bq6HeRI058boYf+TYwVS4kI+ECzyoDEkO7GNtU97kTE2caiSB0pwUU5+SuzlDLH2bTbl/EUOT3V2CNw2vYZ1NRI+ECzyoDEkO7GNtU97kTE2caiSB0pwUU5+SuzlDLH2bTbl/EUOT3V0Yf+TYwVS4kI+ECzyoDEkO7GNtU97kTE2caiSB0pwUUzsbvkIC2oOYgTQrGf59Sxdce6gJfrhvWotJFi57rHJCgcZdMvisFLttRd9iJfrOFKcnp15/O3TdSZPOCZaguuN8FyHxX8VRCJKHozjh0OSjyJask47xBrjhwyaAxLfQPRSI6dQzrfsnQ6E/cqmx8G6AT1ueVk2HLhNKpC45fGJah4jRU0S74lhYggAh2zYxKvJMoiRRwIwdxU3M2T/kMpB9BDX0RjbgsM6Emqho75RJNWYnM+lVTITu+49+N5j8NVRWHJYQ/HeHQW6A1k/HcyN9BDX0RjbgsPyFDQea6P7Hj3F5vxN4vEbsY21T3uRMTZxqJIHSnBRTn5K7OUMsfZutV3RFUpvZ3TVmJzPpVUyEq4yOERp1nZJUVhyWEPx3h0FugNZPx3MjfQQ19EY24LDjRkmphqfq+n6BQePAhrS5a9CKQlY8TsIr5MLZhS3k9gwVVKVZChi47E21xuQsYuO33De77oBSSIeI0VNEu+JYWIIAIds2MSryTKIkUcCMHTO6wNMXY2pO0+yOMqqMIvXXrMEQnCbaD7W5VQZO52ca6n1DU9NV5kZr0IpCVjxOwivkwtmFLeT2ysSmPrK5fjBUHJ01rNlq0txTPL7s1Vxvj4QLPKgMSQ7sY21T3uRMTZxqJIHSnBRTABKLJIyCVUTkXbfrnrGzqhl8kz+spx1yg3EgxiHOanvhwyaAxLfQPRSI6dQzrfsnYE7NNkWoR49tPVM7sSVoAcIIPxBr+NBQb/dQ2czp4u3C4OEyxUpTD+dK/+s2YPEJp9mOyCf3RrSK2GiDW7KhizERImOBVL5e7GNtU97kTE2caiSB0pwUUwASiySMglVE2lsipotIURSSh6M44dDkozaG3MIh2AzVwuDhMsVKUw/nSv/rNmDxCWsVH2Gwy/qzq3h3LJ68A/S1uVUGTudnGup9Q1PTVeZGa9CKQlY8TsIr5MLZhS3k9g2EcLWlm5nRgdyAXHv78ZN/rmlOCs+pkSjSrOYz7E2R7GNtU97kTE2caiSB0pwUUzjqIP3K9HgnIo4O+YMlIBA9LaGidc4WLxSxOoMvilz9WIIAIds2MSryTKIkUcCMHebMkZ2fEVkD0TJg68Pxohyym6TZ+4ZAL8TFM0iKu1quZ7v/Kw4/e5ANu9GXfU3btedK/+s2YPEJxsUzRLntQIEW72BR20ZnxLBiobIKCIsckOFC3nBXjR+j9a4NkQvW6fJMoiRRwIwdc2zNYYbp2Mirod5EjTnxuoI3Da9hnU1Ej4QLPKgMSQ7sY21T3uRMTZxqJIHSnBRTBNa77cixzGvSYzw1lBVSfIaYHTMW8JqPKYpuXYGa4XRr0IpCVjxOwivkwtmFLeT2AAEp26K0QYZYSuqVtH+R9pKHozjh0OSjyJask47xBrjhwyaAxLfQPRSI6dQzrfsnoaHdRVajFyyOY/Zz5BTbEsIIPxBr+NBQ5lbfYQeVRXXC4OEyxUpTD+dK/+s2YPEJoeuA5Mirn0be1qNZioQyIAsyjBhW1qfXHEcuJ+RvSwaFVSD1FKcXtKcLd6wnWbHqE+0qe10QYTRjuqaY4wcJjhwpgDUH9R9fa9CKQlY8TsIr5MLZhS3k9rQAUd8pPnf/B7Oxmcvj1hpjBfVosytm4xwpgDUH9R9fa9CKQlY8TsIr5MLZhS3k9rQAUd8pPnf/E+0qe10QYTRjuqaY4wcJjhwpgDUH9R9fa9CKQlY8TsIr5MLZhS3k9rJsJpzbWmJ4IkKR3IvQI8iZJoS14FBVjvUYK9rKqt/ywuDhMsVKUw/nSv/rNmDxCfHmz+BvnaU8uZpoX5z1OOspfoWQz0YWbrqZpHRFaSxbbUXfYiX6zhRvsIoaBB34idsqKEd60d2xYwX1aLMrZuMpim5dgZrhdGvQikJWPE7CK+TC2YUt5Pb9rNQ9pMjFpzHcDu8XMKjbi0kWLnusckIJrXE3nd7zlraJ8/lTY3NynAnqRY0tzpmXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZmkeZDENNQiLjQTiMFQj5Fijq1iJ2SgVkpdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmTyWwC/bRyxBlh1+mBHY9E564K/wQvn7OfO3i5SZEQvnwiwWgJ+7QozM1NjMSpFCDjrzbpUr/iWCU9XczSMtPKPszmn3y2/0NBSV51MktsHakUv84M1SLLCCEhntrBV+cE+h1JLLPn+qUzsVX+qjJ2SOL0yshwRnPo7T1pRQ63F7L7To5FoCCydWZoiiFN4qHmp16fspb4dnx/NWum6aNbjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyMj1EomkBOXDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8ZP9vSwZxnYAOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHLlYlQlOkI9vzaMWyOJnvaYpmRSLqrDyOGA61zq5LyRKADNFTHDXYzP5v3z4BoloQOwb5BE4LPl1hp5IRzli53XmFInidWHoGXYrqEx1I9NHIHyuUN/TYhgir1AJXJarU4lX26L3zEegzDCDFQmIOwZqDXxlkXGyt+glhNV8qicNbLHdE6hK3m2QIaAy+tSTHE37Nk97b+6rujMteNf9cfp/uoMRIZf43L2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTLwQFJvaXTD8+RpYN5qRry4DY1iAzS0/iJWWZ0DjHaUEHbMOhvMOjthqDXxlkXGyt9Z+gm9tSVzWb1tbidPYvITNDrz/dM09R4aYzfjTC6+kbOm4GNjZXJt86hhd/8v9oanGTQoBpT15m4JQmX6vUqjr52FJW9ZFldXmAeYqCVGIMxBPmd3IyJnOyxQZ13Y28eB8SJ0Eoctp8uT6SxIGKL0GGu+3/L5gB1DUfp2UPpHMcm+zkrrBdbdLYW4B002kb1exiS1n92oFmkcaxGusi5nsCB20QNKFLQdB0Al9P1lUx7wKoR3+QP1nvIw9bSbQXyoNfGWRcbK35uA+xX6r6MrntpxF5Xd9SgdB0Al9P1lU/9lZ436iW/ZqDXxlkXGyt+Qmd/cNiaCSlHp7xYKUAciaRxrEa6yLmeTo3e2umQ5q7EXavObQprQkNEPMoCb13rC2pgAuKXPY8TJ94F7L83+y/BJV9UtiIni6NijPWSXfSCT8V7G3NBEHEcuJ+RvSwYQvkdla5p3Cwo87QNhWHJ850frUHd1nGXCbYKEuMHqNO2N5ot3ufNuHQdAJfT9ZVNF+jyPXqXgzaee5spar6GAkNEPMoCb13phZozdt25vcKg18ZZFxsrftjgv6aFjGp5fBFRjSASZefGU7Yaa/ltVjHkTuid8rq/45IRa06TYebRsC2Yrcr8TP7Ma1XYBKh0Y6KXCSDj5F+PlFyDCCNCFilVRhs+0ObpH4j/NjnSpD9AHpDVKFDk05tCyWgEiKXtlWchJ70S7PvfvvZGFwKPyrDVmeF0AhpUcRy4n5G9LBvHw0l8WzOdVmQuDrbCd8gQETOWt0KBunDb9QuSHDNdeffqlppcnQWarsEsLMzN2uV4eBkldpXel8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3Z/sInISWfn1UPnPI3akLZs1xOkrv9mo2+GOKrqhBY73772RhcCj8isfCkcVtcnhcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMNKfTS1aPKqZJH7Dr7SBOurqgselVXw2ny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8bs+d2pFfQrbrGUcTp8V9i6Ff1lN6qbqa+2d+iBc8v0FHyC3GItNMeLnbSP9FHkYHWRXZEp4UN23chK2rhaMLmZP5DKhKevgqeGFB3kb9erk5iKqJZa0Jmp0kToM5jgJRzSc3R/HQ5ndZL+814w1rJYvxMuc4I56TuGu/GBSs/BGw3A/vUeeRThs/P9zr8kn/aI9EAkCE4Ye4e9Dh8lxhBUA0CsrL1TEzUCGgMvrUkxxN+zZPe2/uq7jqS2b4yIpdqnQtyZxDfebu3BxnJnHGi23U4tcd5nCGARM5a3QoG6cknd7NQpRA29mzfnCvpTk9bhdDjKl/Ez7cEVQvmZs4ZhxCvea/bRFrEL2TqHljvVfNKeerljP17mB8SJ0Eoctp8uT6SxIGKL0GGu+3/L5gB10kToM5jgJR/TzsTrIT/0QyD7Psl+asFt/WCNz4K/0/HWBGAt0vX4Foan+dLQcY7MYa77f8vmAHQih5UzjWkOq9POxOshP/RDIPs+yX5qwWyKAhcK4f6qPdYEYC3S9fgWhqf50tBxjsxhrvt/y+YAdLG2KyO1nrRf087E6yE/9ECYqdB9zl8frf1gjc+Cv9PzgWZgmZ0ccTaGp/nS0HGOzGGu+3/L5gB1lm7+N33q6mPTzsTrIT/0QJip0H3OXx+sigIXCuH+qj+BZmCZnRxxNoan+dLQcY7MYa77f8vmAHYGA51/eN3IYegQEcfOW8epHaRTsYmwPn6g18ZZFxsrfrTIP0x/AMDCDPmhAtpi4ZmsezOrWWHiu9orqZYAgHpt8qC7wYSWXdUMThgOCryD2BLHXILXug7by/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPFpbEnY3Ckt2M3TyG6JpEQpIT3ce60XvKcwUhrOHwTVkfiP82OdKkPpJTzZpExTfo6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUci5uZGGoe8WQOgaEDoJHRzeJdxYUiParVk/6zjsel3ed8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTsrNWYQz+pTB9BDX0RjbgsDBhAG9cJcbnJl5pP+/w5LVg8M/XPHF9qOQkas+/4BSqH1MVbgl0uWOXt14nAyWWX0NaRZr5dtq7lcwbKRQEQlmWnABkhfYwG9iuoTHUj00cGEQXuDjAvKNdy8CtVyGrD0JgWLIeqDPpcQr3mv20RawKPO0DYVhyfIE0Kxn+fUsXY69bQ3K9J0CIZqMNe2dGd6g18ZZFxsrfND+gw4XgwxtYSuqVtH+R9uzNWXIR7349svZocreqjFVZ7jm7Ur1mMIBPW55WTYculpOZ+n1K42xx2+R8PZCp4Bac4htHVSbngyg1kDodHEcl75f+1G19Y6uh3kSNOfG6xtH52OG0xKznzHgVog13GAo87QNhWHJ8gTQrGf59Sxf8hTjvWNjdA4hmow17Z0Z3qDXxlkXGyt80P6DDheDDG3Ayk+IiB0GE9PmvC//CR55JgvW095XUsr2rBUoGQrMw43YVY774KSGEV/5uS3r+fNJjPDWUFVJ8QQ9eyk4W732wQhh0pcAK0Wo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa2wULyPbYaeuqQ7Jo9aE8RX9QLeJ0Ku6wPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8WlsSdjcKS3w24ojaO+Xb6rod5EjTnxusbR+djhtMSszcRjlSAArIdqaIwjnVb6nn6PNq8dQEb/p/toiHwXQ2KnCZoSaiIUUZCqxpLATr7/gTQrGf59Sxf8hTjvWNjdAwih5UzjWkOqpOLexdwWs1qgbimBuFce4RF0CZnA1o4s+2yJBPCihQ8jYa8N06d/3zQ/oMOF4MMbcDKT4iIHQYRXMVxEKZuZHCXVMBWtR9g7oDQNxTANHbCB8SJ0Eoctp/aF54fL6y7Lll4RdywoIIzn1D4PvyxBtNQFXSg/+Y/DBJkRRSsPqcKWrZ5ZKcPlTar3Uf148eWiuJMq7VCULOU6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZW5BCAWusjPebZkuCtnFqVHAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTuvFlDLeVAgzYhpwO952DPqO9b/CSYJy6IPEEOOs5sYKI6I2xjDEQ3C8V8b58GG7aywKTkKJerd9LvnX2Duhfj3UWKJQ6R9GzprfkM6pnQKu/EUKWXiWm56g18ZZFxsrftjgv6aFjGp4nu3HfAAlZQqg18ZZFxsrfJmzaQoAueoDSYzw1lBVSfOvf3QJG+4FVgE9bnlZNhy6FFzBmfV8+hVeRs+988DR/gTQrGf59SxdFS2m0Rhxp0UqSqg/VB7RBRdUPMe7YwCSoNfGWRcbK3yZs2kKALnqAXUrkOzw4JZDr390CRvuBVYBPW55WTYcufOoONLnRFEpXkbPvfPA0f4E0Kxn+fUsXa7JBGmZ8Dl5KkqoP1Qe0QaExFltfGT2sqDXxlkXGyt977N95KPgA/Ver61Mz6ccbfID8LDeXPCpKkqoP1Qe0QblmHjFw+jP+SZPOCZaguuMkVp5M0JkVg/7uLr4i1X3J1AVdKD/5j8Pj5yT0H1ER4FnuObtSvWYwaHGmnSlmR8uIc/9sx4RXmNQFXSg/+Y/DM5K+elT6eANJk84JlqC643Ayk+IiB0GEkNEPMoCb13pJABgwKu/lQI9HL9fBaD3ov5YvryNWNrQl75f+1G19Y0vpv8GSFMOISpKqD9UHtEF4CQuQ51KPK5XRbIfXsO7oBEzlrdCgbpw2/ULkhwzXXn36paaXJ0Fmq7BLCzMzdrnQjS9Y30whPhkVy0JPbV8hcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNyukvJ0+dhsJmo1m768rOu+6KP0OZGTDsTCwOKYR7CtX5dkcyguCL99+IiKSVI2SrdHNoKxKXwQLwMTsaUjaBAF03/mTVO1RaZC4OtsJ3yBBrnUAqt0p/IrHEBNYVWkOeaWK6kom03KoDXnCgBbXhAFAgfy5oikWemg2a6thA6og+wjudaZdNLMevofOtLahN6IfOpWQZiMJRbcYTh6GFXrcT8eyl/0y4hTjj57LvU90C8OIornqDi8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEfv2RztNZnVWCx2tiJQLxVJWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJO+mx+WMZOI2Wd8Z4UpbHw0uNSd7jJV/9wmf0g7T8uikTmdjCz+epvdf0N2LXKhc58DXHDjv1yxOgAg8H/eMiiuF4iEljlli5BByPWgy+P8E+eSNGl1cCaS4cMmgMS30D0npv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWs1XPzOFWEX+vnECxWJ+ZR2PaqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+gGwFmQkytbgP1ziX8hdVw2N7AhKNvBXLfCf1a1PYXmtrLsSh2Hw2xeEkpZ1EwtkI/0+nXrAtOe6t1Us1yOUS3vlBN2g//N548SmTLoMMx8CoNfGWRcbK3/R+7e50mN32JwNf9wGtoGSBgOdf3jdyGIRweIGYy0fZSvXkPabCstaA8+8fyuFjDFB5OylphKT7sey7tg7gVLwRjnHMJPFmDqIKIf16unyHu/+ELO4kdpEs8GueonihwlAadsLr1qYpwFgsHfuuaTC38SK/Lu6OywBafIsPzRxb5Uu+2svBKxz+pNzirPND8f0JPsPRESoNtJelJ2P/PoESJICPeT2raZ8A84lnmGTMnqFJ1wn/hzwx5ryufnuHSAvxdtMQ3+XX6My141/1x+l8O9/lmpDJyQ5/7HavQMhIEd89j/BZuIM14+ko1WhanRa7zoMzwU8uQYrSQJBv7P4m4Cs6NtgPEf7EyRNyHfiq8IMB0jorXOitMg/TH8AwMJuwpfyRpuHUTMzqNaAeQE2oQhcuO4+bqlLw+bLG0tqNOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHLBjnWyfSULUyqFVeARFJVo446nnlC6Jml+WDN1P4BA6oaphD75swo+O6WJZXM/p+z+JYZOh8gdAI0nk+Bh9+WJI7YmO/Juo5XmjKghd4lsW/1xkVp2NLD9NMZY/k2FuejfD2SbpJ8WsSO2JjvybqOVp+WKE9AG629rnuPQR7bsgZ9PWYNc42vk3M0i2UsHFFDbPyHo3ZO5owcc3ogdkqWwcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Jgb1e9FaeuJQqUP47Zts2kKg4ZEwM3vRL3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTuvFlDLeVAgxxFwkNSjx8R7Uda/Df4hrj5oyoIXeJbFssqisAKpLZ9Cem/tdTojcxABpLkx4DeSBlzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZqtolvJ6JyuxOzkZ5XLSI2Dag18ZZFxsrfqXfoT0uSK9QTk9xFozd/EjVmJzPpVUyECKTogwhiX3akj0qk1xQxGJDRDzKAm9d6p9mOyCf3RrQVTnOQGWevRjXjrdZ2biuXbXyK9WL38YScKTuURxbQ/O0nUfNDFyrJcRcJDUo8fEdB6b+5wfP5ft+DlieiQjQwxAV5snqf4dqrXW/Lngz1XTXftv/gwZeS42B5hyENdIdi11TfDsEnIB+pBQUd/IzhvoiGCRllu1SRftjjGWJHTVyT4dfEL/inQiVAWBgw1HBOvcYwCjMniXAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JovMoZgNf4RBJ6BAASQm2UoG0Y/tGaX5TMXNhc1TVpiuLICuKpniw7IKadvTV2Cv94mtPmXKriGrVACtDY6oJrN4GEzOpq6cHNZTjuwSoh6Uq9LBbPu84Eb5Qpu39MOATjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRy6NnIV7qdz1/T7I4yqowi9deswRCcJtoPiFN34nXB0lH8UnERL5ba7Bw2TEYBX3tTqxiEouaRpssvFfG+fBhu2ssCk5CiXq3flyJNSZWXY3L5W+rEb8XoruEkpZ1EwtkI753r7z1uKWsZUqcucZyzIgAzkJCJoBMZQIaAy+tSTHE37Nk97b+6rmFcV6pKQIgY0xppYqyutR8ZUqcucZyzIgAzkJCJoBMZQIaAy+tSTHE37Nk97b+6rlVbcOIpGTPC/QGttesYKYDNinA5JzIHRy9nAOXMoiDEDCuNVCU7v0plzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZq8qVePvYVwa2bNcTpK7/ZqCkJuMch/Os1uWDl+4FOsmjvnevvPW4paxlSpy5xnLMiNbhL5G5GLNwPsI7nWmXTS8uDSGpSh1alqDXxlkXGyt+tMg/TH8AwMLPE7sQG274oCE+KhaIWDMrxOUvVKUGSD5acAGSF9jAb2K6hMdSPTRw7hw+8jMcJvtPsjjKqjCL116zBEJwm2g9uQcKSvvB8RDLYve3nwTNoUIejvdUmFwMWnOIbR1Um54MoNZA6HRxHxZBydf5r6zWeMjyWMYBdYwHSysqpY4h1ouJoANjKSdsZUqcucZyzIr+Z7XH2HrV6vasFSgZCszDjdhVjvvgpIfJhNjB2HOn/W5Yr3a7r/gI0TqWNKWaeePE5S9UpQZIPBEzlrdCgbpw2/ULkhwzXXn36paaXJ0Fmq7BLCzMzdrkluoVrZUgurKt/6obduUPpWyQ6rG9bTZuXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZqNtVn0GSBMFmzXE6Su/2ajb4Y4quqEFjvfvvZGFwKPyhSmClL5kJWen2Y7IJ/dGtHfiq9uADSO9BrqqWjh33U15WPQGbvn42fNvrw/EzzjiWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFlzJgvaaFBapWcRcJDUo8fEdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk76bH5Yxk4jZ07HhY7BFg8qlG8KO+O2lmiZeaT/v8OS1YPDP1zxxfagzfIcJGnly/Xp5MwVrdLSb0kfhGIVJ+sp4LB8SnYnkWJuhHwoq8y0TY59MtPd72sG5YOX7gU6yaAD1dGCILjYtYpS2VcoJdBssGaW6ielPxFEJZt5I6hoN5iRnMMMFpPv3GKSbJQo2s/eBG8KWa740kKxaDasfPpti/QZxTA2ygikJuMch/Os1uWDl+4FOsmjkgw4hj87NG+N/Fi4B0FwXlpwAZIX2MBvYrqEx1I9NHJGMZSUNb0n0ynkdVxrpQSOimCUn4MQS/MlkgnfFIyU3ykgMr9iKesZN/xGCJWsccGohSSi0mKWlcVrIoVc6ZeH9s+Z7SxRm5KfZjsgn90a0x8Rln0b/RmYWnOIbR1Um54MoNZA6HRxHgsX2cBltbUx6CKPxjjRCIXXUXy0wb/1SAoSEas/7EsKPuFEQpJW7QdcKS2PyV/OHaj9JfMVzGs3/rdqFdmhrd+/MiU0EfcK0qXfoT0uSK9SBGrP+kd/5qABKVBuglOW+ax7M6tZYeK5qORwzQdMkxaICI0ezhqA3hX9ZTeqm6mv1CiDMyziG/InLUojYFv+//NqCpndR1dPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+fy9XVZwkl1dzYpwOScyB0cCQZtiLovMJYRjIpqXdgryhZegRHAfelaXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZozlgiUSSlJPn4AaHQvH1b7NReFosymZhDokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyymkKrPAXuCTttcR8WpyGg90A30UpVmtaoWFgEdetSo1nauqvuIr+zGpQqLKO6hlOG5ijMvAwQDKo1fNd3oasbSKODvmDJSAQDles2xfXwOkUsTqDL4pc/ViCACHbNjEqs6bgY2Nlcm0gotVE/6BHkK4Jk1m5wAEigI+jAtt4bO01Zicz6VVMhCgnI8G7oo/IVFYclhD8d4fm/fPgGiWhA7BvkETgs+XWGnkhHOWLndeYUieJ1YegZdiuoTHUj00cN+plWTQJSyxJb3vtfaweaTQ68/3TNPUeGmM340wuvpGzpuBjY2VybdboZH+dJQSkDi7bRPfSArK7cHGcmccaLbdTi1x3mcIYkNEPMoCb13rAlCJBb+ant8gGZMNnOJAmJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfeygR1a92YwMfrh1j7P7yEkCGgMvrUkxxN+zZPe2/uq5VW3DiKRkzwkt823SW/R2iJ15JUQF1w9ovB2RBqE8Qg/GED6cYfjdoNrlzvRZ41imTysGfIDZrZ5jY2T67Es+9y5PpLEgYovSzxO7EBtu+KLFItsraew8YikQAyWKXI4K/EUKWXiWm56g18ZZFxsrf1uhkf50lBKSrJshmE1ZfTWxHoMmoJRXKsvummJ6cYLwYa77f8vmAHcCUIkFv5qe3gnI6ZltxUmIVBFNCDVDPUNQA6jzimz0WwFgsHfuuaTB7KBHVr3ZjA1G5mylj9mW/PwGopGN5FQ7zMTThNfQr8/9VOEEPlSHPdlL7H9yAgeVJWgIGkfD1HHsoEdWvdmMDuKPqxC7RtK+9qwVKBkKzMON2FWO++CkhNiM/3IusMSybNcTpK7/ZqJ0Jsfa36wdxhvCMT6MdX9OfAPOJZ5hkzOOv2o7NCN8yWvq0tzIfbEGpv2qnHTf9g7T//Islk0UTQvZOoeWO9V+9Oslpscp+fIHxInQShy2ny5PpLEgYovQYa77f8vmAHa4Jk1m5wAEirm8GEJCzh9IiaPu/LutSJ/b0ZVcbjQTSW5FZH+ZGdxzAlCJBb+ant/MxNOE19CvztY2ChAhRVj9ztHZMAPMdzZyfzgHf513mBMNlvUmHSdB1hxOPGSuxJkzgT8PcZwUQdlL7H9yAgeWyNcfwmy5SoZvhQT+f1furGGu+3/L5gB2uCZNZucABIq5vBhCQs4fSImj7vy7rUieDlZwk8pVYc2ZBWAsg+pKjwJQiQW/mp7fVe1ooB9wnMbWNgoQIUVY/c7R2TADzHc2cn84B3+dd5gTDZb1Jh0nQsMdWVVIHobzuzk/UUKvbj3ZS+x/cgIHln5pkv+29tQAQ9BMUbPYIW3cMKmb+s8su0jiJ1b77BtzRMmDrw/GiHEHRmpIQ7tIkKvz/8yBkR601JD5J2pzGV5Oc+HX4RSdW2c64Cr8Xadbqa9p+s51GzkZrApfLiXT1DFMtBFY3sZqB3IBce/vxk2mF9NC7O+C6QPVHMmkNW9O3BrWU01tJZrtdDpSOynH30TJg68PxohyQ0Q8ygJvXesbFM0S57UCBFu9gUdtGZ8Q1atilW5y4K2E88nbISAJHyPeJqedH2Vr7lb+MngCU+BgHK07y28LVB/0N7qXtgUshUCar4f5YlnOvYDcCdEcznPKByz5hZQ4fqQUFHfyM4b6IhgkZZbtUkX7Y4xliR00OgHp18yZGfXIVGuvHLOGqQtLc4hcd0haXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnkDEh4cK+avIo4O+YMlIBCzGnDL6qMecIHcgFx7+/GTWuHzQuAYPLxS5R9byV2hR0HtWYjlWU/S8uUUFTosjZYcYkg3lk+Yb1aS6I1Th7GcANJsFoQX1LJZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWXYezyHFFaWl99kHlmR50LyfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxfGpeaTsz15ytmiXGHs8cQ+aMqCF3iWxbLKorACqS2fQnpv7XU6I3MQAaS5MeA3kgZcxmz9AAC0ynxG91hzMy4FFj5+cursX8ETuc2nyyzNzmIqollrQmaraJbyeicrsTs5GeVy0iNg2oNfGWRcbK34s37kzPB+IhY69bQ3K9J0BrFR9hsMv6s6t4dyyevAP0uHkcmlnxQWAXobiViRArXDIdbayeN9KhqrlQHW6bvlaB3IBce/vxk5+aZL/tvbUAIpc30DAikYVYSuqVtH+R9n+CkJ1/R0P5av0Cps8hBu2+EjR0npuqLlo1LtHNujgmTbl/EUOT3V0oAV/uiNJ7uYNHXGeH2LC0RXoTiWnhAYRE3tygC005pJ2PjdxlApxGre8A8KaCEouJRkkmMiKGuFeoiPowlP6r+hWb3LoWbbwkVp5M0JkVg4KapVqiRmGifBch8V/FUQiQ0Q8ygJvXeqHrgOTIq59GneP0N/uBkPOLN+5MzwfiIbUCk9u5djIbizfuTM8H4iHiIXogJzL+u72rBUoGQrMwvnE5wKNaMBRiCjv/vpJYcPPDrTfYYTjKa57j0Ee27IH/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyPXyMGM0AOBbyXAZ9o/vsM2B/p4Vpoz/Drs7IZ1ypQhpnbfE/C2mMCscQE1hVaQ5/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx7Gsb06a6vcxJ84SfQL8uXkBEPjeRLrhKcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPACRbAxUqn6wqOJ/8fex68lhXjuJgudJM2jFsjiZ72mKZkUi6qw8jhgOtc6uS8kSgAzRUxw12Mz+b98+AaJaEDsG+QROCz5dYaeSEc5Yud15hSJ4nVh6Bl2K6hMdSPTRwkwZIjBcGCGBr6LiX5vnG2NDrz/dM09R4aYzfjTC6+kbOm4GNjZXJtEOl/aQLOm96XkYrNcNg/4btwcZyZxxott1OLXHeZwhiQ0Q8ygJvXemPKonJwCA9HV6iI+jCU/qs0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4BuEW2SpeduhPtKntdEGE0fvOR2XnFrlVs/P9zr8kn/aI9EAkCE4YeX4CHGxF1gxNvJcBn2j++w/TnBVw5PkIIenPTtAYOt1bzqGF3/y/2hqcZNCgGlPXmbglCZfq9SqOvnYUlb1kWV1eYB5ioJUYgRN7coAtNOaSF/yc7SCzNRecpI1FuFZpa/4RPiruSzIEUJzSMEUKMwQOk7IQVzJHiYlp83Az1u0SjJSv4Ka0sWKVmuzIYksrLNpsE1zwo/C+jhG4beAcEch6f2/rGKUm6CJvvwm5Ml1aLN+5MzwfiIReAIzzXgm7Z/auuQkqIl6gAf03y83Mqy5Xsr229kkEcE+0qe10QYTRMpVL58MJBQoGAnvueMkLemzXE6Su/2ai6g3AJ2dqPgzudpJy86nmIzEE+Z3cjImdjyqJycAgPR36PNq8dQEb/ETuc2nyyzNzmIqollrQmaiTBkiMFwYIYGvouJfm+cbasuRwhskqGjIGJj2Qh3IiJljiIpZs9yIQAf03y83Mqy43LOJGYrv79qDXxlkXGyt8Q6X9pAs6b3peRis1w2D/hY8qicnAID0fE91vB7WqOp7V9K+vyG9GCE+0qe10QYTTlfRNP3a/oxpflSbQ/7r+gNv1C5IcM1169qwVKBkKzML5xOcCjWjAUYgo7/76SWHDzw6032GE4yuL26A76c5IbmiHaSj0fmrVZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk0MSw/dqK9HHl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGb8AHUmsrXqV0bGd7ABmna7Vzdfcxt8mf06JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcp4Tl0cp2WclDqDsw3GBFyav8a9H81GpKKFhYBHXrUqNZ2rqr7iK/sxqUKiyjuoZTiem/tdTojcxABpLkx4DeSAfILcYi00x4sYtchMc4mmUcQr3mv20RaySoGtWHrMQoMbXe09SFZZkNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOIhBYHCkvNIwee83d/nVokbtwcZyZxxott1OLXHeZwhgETOWt0KBunJJ3ezUKUQNvZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYcQr3mv20RaxC9k6h5Y71X5TK09xkZJv1GaKbeJvuZdVXmAeYqCVGIMBYLB37rmkwDB2TZHWspj10B9jT4Fn4OAMJfh4Q4NFonDKHD3t4wrBD06ZKOxjpTHKVSDuBUUILDgiDJbz5BY6hKlCAG3SxEhzWEKD2PpNXdg+mmYluNhyZAvZJHgRkvfL3UeuSfCGgYQjH0WBFruMLiUET6cS6kbOm4GNjZXJtajkcM0HTJMUETOWt0KBunDb9QuSHDNdeffqlppcnQWarsEsLMzN2udosEuxiz72pnZ6hdWFNOl86JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUclqc3dGkLbiP2yooR3rR3bGj1LPZE6uc4sLGR8ZjESG20Oe6Y2oFJJEc1hCg9j6TV7PyE9mT0B4ZtF4E6dtJ6DI6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZJxySuyuWh3uG2wQmryA5pfaoV1U/wv+YeQNK+vHa1FwL39q2OrdvMfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxTrls1ZJGB1d8EgNGoYoA+k86/2QZrtGwvkPST7jLNQPiDA7VOaQ+AiDxBDjrObGCiOiNsYwxENwvFfG+fBhu2ssCk5CiXq3fS7519g7oX491FiiUOkfRszjpyXrOGgoLV5gHmKglRiDMQT5ndyMiZ4RVz/N5tm+MgfEidBKHLafLk+ksSBii9Bhrvt/y+YAdYgC8UwPsxZTXrMEQnCbaD2WHX6YEdj0TL0NCG4eImb6ZsjU/M7eLPgHSysqpY4h1s6bgY2Nlcm3WLm3eKt4OT8BYLB37rmkwQPdBX//cRrcB0srKqWOIdSE2/WqAu5XREiBKXmipad4PsI7nWmXTS9/eDlBQWb2ikNEPMoCb13phZozdt25vcKg18ZZFxsrfEn0RGm3rB0SKRADJYpcjgr8RQpZeJabnqDXxlkXGyt8TxCRFdTZu1RRH6g+4YcPzbHRUnNvOTNBSU7lNyZCRSGhTwpKQqniXq3h3LJ68A/QZ/C4f1hSg0cnWxrCCADH9iC2SXKNBKbWa/sbTdmm9xTYv1yiOX8cUc7R2TADzHc1WwqLOPfeSacBYLB37rmkw/W0qT3FpEXaP4G9/8qtgnC9DQhuHiJm+loYTYXP7ZuuaFHHSvsBMv5DRDzKAm9d6vbd/0eK55LL/VThBD5Uhz+dxfhcQh13L9iri0bUW3lTCbYKEuMHqNL8yIR2yBElvykgMr9iKesa+of7UZ4UUWKg18ZZFxsrf+UY2dcl8nIaene9YsPK4t8vwSVfVLYiJ8C3urU+V8bD7lb+MngCU+Gb7dfJYiVXHydbGsIIAMf2BVMhkQY5kVpr+xtN2ab3FNi/XKI5fxxRztHZMAPMdzVbCos4995JpgypL2PvmW8G+iIYJGWW7VBD0ExRs9ghbLNKtkJNGg+W4EkG4xCRtzIhBemq8LWWMpUm29/YKOmlLUyznmsp5qY58TgH9jycGCQ2AdkZql9BwfFE3jEDu69CfBfrEEOqbARO2FI0qUBw9NbvLVSRh08vJyVyAn9P4q4j0S+aVfp5Lek8xFmzmIlJTuU3JkJFITtQr8I3+EpwK3i/ynA4SUrT9KQ3pbn9G4++p9PuNtvdPKdBsNUvW7SxFxpn4Dsyz9rmT0ugJIkAaGVCbZOT3hsCUIkFv5qe3Qhj5/ds432uZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4re3hHkj6OA750bbJiIZC3e0byk0i9kWazPIGY4aVIbeVnOhCGoXArhwEU0yBqKU7ZAntCuCluV+iEQPT9/I9pShjpELf/aCKUqe2oMdKD1yKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTyNOGBYR8d3lMgAR/8oyPRSgvVMR6t5LImagpUwam8thwIyMY/vV7Tn14eOBK7vhtvwxXRPxIwFahA95t9lk2aNTudyJIkz+VJCQDErCrJjjonenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvhUEU0INUM9QM4Wm5eVjRrO4ugDXg6fOP13lLvMeWhFt6Pd4OdMbLSVl5iu8XGxV4z2TQ1QOCohiC4j2MM04Y1HV25U9Uq4lMvuLTEYhdwuUD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDAqplN3cVEzU/AaikY3kVDsN1GxF8bVtarA4cDybZAivpDnXpz9TWL9qqgvbqIhfPpH+iYXN2p5akPIN6OlF1sbK2EmmuheO85xwP35XTd6rzIdIlMUJc4ZljO7IO5vaSLad8u35k2XXFUlVUTWKaM7IbMnzgmU/it7eEeSPo4DvnRtsmIhkLd7RvKTSL2RZrM8gZjhpUht5AMig+TYo8W3ARTTIGopTtkCe0K4KW5X61LAK7MCLqZMZcSLb94zxG86VtEiHnpQqjwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+yerg4Gueif9HZS+x/cgIHl3gy+nTaA/69L4v38+snsvd5or/D1mwhGW+PLWHJwcdsoKmVcgLNIxdFBzzIvZu6EbEOj5C+YdsxdAqKbN5zmlErU1VCxcQ8jPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuvmNJa65VppwCDlZwk8pVYc2Dkt/4rqvxDS1Ms55rKealE1yn/4DsSygkNgHZGapfQcHxRN4xA7uvQnwX6xBDqm4a8Uq5yqTerjAHVhPDekxjLyclcgJ/T+KuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSMPPBDcBy1gpCFJ8W5xmekysDhwPJtkCK+kOdenP1NYv+lfEbkbVJpOkf6Jhc3anlqQ8g3o6UXWx6lc2YFG6Gzu0bAtmK3K/E7wPLueC2ZXK+GiIvwPqUc4xlom6SpJyQcvwSVfVLYiJx/mGnXcyWIjLb/+4WYqS27i6ANeDp84/XeUu8x5aEW3JBnkp7WtTJ2XmK7xcbFXjPZNDVA4KiGILiPYwzThjUTSnnq5Yz9e5olnDTr2SABCZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjPtjeaLd7nzboSgGQJusI1+fm07Jj+SqtNL4v38+snsvR+xB9XjAweb4rn6MKGc2hMoKmVcgLNIxdFBzzIvZu6EEmne35LIf33Ed+yAS0DMXaPA8XIE0tuMKaIn7NYNLGIL5ZgXVjx77Dwm/Oxmv/Ln3tqXZ0AkX2u0byk0i9kWazPIGY4aVIbepGiSv363aRlwEU0yBqKU7ZAntCuCluV+TPrbn2WH7eny5osjpT6EQZljO7IO5vaSLad8u35k2XXFUlVUTWKaM5DZsbNvEjC2GB+Qg0r3LE6sDhwPJtkCK+kOdenP1NYv9amjwIgKLhSkf6Jhc3anlqQ8g3o6UXWxKuyHgyoF7/Wvf7ic5DhLBw/IYWiIqjyhXlB9PcWZIklyA8lDag+GgwKotuQtH8+glDMnpLGc+Ze4ugDXg6fOP13lLvMeWhFtyjug6FVLIrtl5iu8XGxV4z2TQ1QOCohiC4j2MM04Y1GojPSwEcqobCd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+EiyUqT/eAKq0/SkN6W5/RuPvqfT7jbb3+arq2Sh2UhgsRcaZ+A7Ms/a5k9LoCSJAGhlQm2Tk94aBgOdf3jdyGG/3Az9mqEJIPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuv4XjR4xtY9fiitg/iIcX3Jri6ANeDp84/XeUu8x5aEW1czZfT91SAb2XmK7xcbFXjPZNDVA4KiGILiPYwzThjUaA0DcUwDR2wolnDTr2SABCZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOWcVEDmcTkfl3LwK1XIasPfm07Jj+SqtNL4v38+snsvR+xB9XjAweb7ru/9ZjM+U8oKmVcgLNIxdFBzzIvZu6EEdmj9azFT33XrMEQnCbaD7i6/LGWU6AbKVF6ecgnJ+Z0gwoF2P6DULU43JJavBLSAdLKyqljiHXDFR0jIQgdxKpNS6+zNLwMPcMSjj9uY2yw5b3DwFQVuWtLVNc5sYlOMW1BDnS8vOGfbV8LENMHnNvHnyRR2QhLJ3p6Q0i4QRB3IGxObWMORRKby4maNfc8Mti97efBM2iIGSgXJT5yfKwOHA8m2QIr6Q516c/U1i+dnTpLGZ8G36R/omFzdqeWpDyDejpRdbFpk16XGVhxQK3VSzXI5RLevA8u54LZlcr4aIi/A+pRzjGWibpKknJBy/BJV9UtiIkXaU5ZoCi+JDZuUPrgWB3wtG8pNIvZFmszyBmOGlSG3mVw2ZfJfIRwcBFNMgailO2QJ7QrgpblfpwKRDU3TqT8W5Yr3a7r/gJKntqDHSg9cilRennIJyfmdIMKBdj+g1C7ZNdaujmE8p23ifjuZvPzEm/7NCMCMO+0/SkN6W5/RuPvqfT7jbb3gqqRull2UYosRcaZ+A7Ms/a5k9LoCSJAGhlQm2Tk94ZQiFhm5PpcuevCkWcx1kIlD8hhaIiqPKFeUH09xZkiSbb8RmN0mlx6av0Cps8hBu16pW3YA+enM7RvKTSL2RZrM8gZjhpUht5ri1+w5FZjlHARTTIGopTtkCe0K4KW5X6cCkQ1N06k/BRH6g+4YcPzL822C5Gep9o+3wUp4AHlaZpBVhazntdDF5JNeqzxZVKreHcsnrwD9FpDd51og9sbagpUwam8thz5YN2Labsty14eOBK7vhtvwxXRPxIwFahA95t9lk2aNeyrCYVQJYGrvA8u54LZlcr4aIi/A+pRzn7e4xvVnKJTw4tTa6h2OqXDFR0jIQgdxKpNS6+zNLwMuygSZ/jWHjqw5b3DwFQVuWtLVNc5sYlOMW1BDnS8vOH3fsKPXehUMMvJyVyAn9P4q4j0S+aVfp64PvMfONWqcAnDUfOHSA2AtP0pDeluf0bj76n0+42290O2ltKwEvjoLEXGmfgOzLP2uZPS6AkiQBoZUJtk5PeGsGkGdB5JKgInenpDSLhBEHcgbE5tYw5FEpvLiZo19zyBUV36z0rilLi6ANeDp84/XeUu8x5aEW11xOsmwjwOsWXmK7xcbFXjPZNDVA4KiGILiPYwzThjUatf0y2WNVsLD8hhaIiqPKFeUH09xZkiSbb8RmN0mlx6aohEu0KiVP2sDhwPJtkCK+kOdenP1NYvsTMTBjF5sSOkf6Jhc3anlqQ8g3o6UXWxaZNelxlYcUCTY9Q5WJEAIkqe2oMdKD1yKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTy6kwPYLzYAqH5KWFgRmyG17i6ANeDp84/XeUu8x5aEW25HKF5TRk9BGXmK7xcbFXjPZNDVA4KiGILiPYwzThjUQwdk2R1rKY9e9DNL0JiEfk+3wUp4AHlaZpBVhazntdDFXX9LD/Bi695zs5PRIUJliwfVEDW7E8KtP0pDeluf0bj76n0+42295mOowEtaVTrLEXGmfgOzLP2uZPS6AkiQBoZUJtk5PeGLsT1DdvvEkK9qh1he6jlAKPA8XIE0tuMKaIn7NYNLGIL5ZgXVjx77OyLyQODB5SpZ6Xm/WZwVgtAvDiKK56g4k65bNWSRgdXfBIDRqGKAPqogwm4UoeHslnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTXde6LA/loEVa4EjQb36tDvIlKFRFC1v8QNfkIgbM1NhQxzx4BSYyoB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCwDKuVfSCivq1Uq2Dto8OhUHcHIYr9UE6eIrdrTIszmZFBAObT4XJblwKtGsbPg3isU/BOF/jE73fkpwVdcZXA0sU3rguAfkIwDKuVfSCivq5UPY8o2c6sP87xs4Igtz+ft/5Fw87SHagCvMDmp2o5MfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvGsVqECQ9P1fMK16swBak6aDrV0SaupysaHlTmKsmfKgFg0CdygaSDdwS7MS5Y9KzSgIrk3Duj8Y+YStKhYVkrvWyKpZe+sEzXqdpuCbaDKLCOjqeEmbrfNg0ZOIlCNdkv94TlSlGhCUZ6CCfYNpaWND5/1YD7AQ8v94TlSlGhCXjazt+6rrfB+Ko8VlHmIOiCeBlNilgh9jJakekrNK1qQkb41xZ0+zJ532mKjRs8AuQ9zsKk8AIidXQoFv1vZWCiB9WB76XcZLBQFOQvZ3yiVjW1fM47WbuugXT7eLWvflucMDlUgErFND5/1YD7AQ8v94TlSlGhCS7SMz5CNY0/93jaDoJOdeiCeBlNilgh9kVxXVWyCsBA6Q516c/U1i/bO4G7LQzeWrBQFOQvZ3yipgq0LWib307yntoAfh6oKGga1gz5GvAbCqD4nUayamL3FBVXLnrdhYLkAzBtEkvpXgkDBylGzbClaqHQ6HYhZSqiwbt8jjHaOLU5nnUugAcwICxouRz2wyCL0/lDTkTEpdntYsoL4Pu7BaWldOSfg14JAwcpRs2wpWqh0Oh2IWUcyI5pET4IalzGchwav//MwV5kUMSlBLg/AaikY3kVDpfLoXhFCw66nvPZszYH98vmVt9hB5VFdcLg4TLFSlMPAf1sDL6Ym0pa+hqimJ2X8nJ8W3W2YQJWqpAPer6kaNEcRy4n5G9LBnPKxSUCjyIDbEegyaglFcosfCRz2v5wfslQhwwd/5HsKYpuXYGa4XRr0IpCVjxOwh2DWy5n0Tr/eygR1a92YwPO2tIEHj2/xDVmJzPpVUyEKCcjwbuij8hUVhyWEPx3h5V3hyOyNkFbvHc7g4cZMrv/N2MTaHVG9xSxOoMvilz9WIIAIds2MSqzpuBjY2VybRUEU0INUM9QplmD20//tk4d23GDqg4YI+95b3xuiqJ14cMmgMS30D2ncXb8pkNlLbIzZIlGboVyUpScbtPXY3mLSRYue6xyQgmtcTed3vOWbUXfYiX6zhQS1F+P0jKq1fho39ocamqTi32YOSX61ago0qzmM+xNkexjbVPe5ExNn6ADi5zKCB9vjD41JgHDTtzqtxk1FboUKykLxLUCU+rP4IOPj2rD7GvQikJWPE7CHYNbLmfROv84Fz2wTKAvWu3RjnCbT5ZXUzZu75YUdPUpOZdZQhNYheHDJoDEt9A9akY/FF8AzWgLsYsz9m1HAZucCMu1RG6NkTl0OxTClGmfAo4nHH+TJzAgLGi5HPbDAi5nyDP1E0Dak5WXwo7DXGvQikJWPE7CNuF9Szb8bc/V4cqecEQZ5yVrUwXxxPn0w8+f1p/yqAD3yLFENI5ayaw9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9akY/FF8AzWhRx8k0NEWRjFCCcmaBVJKejfuoxOiR3gs0O3tZPNEKZx9JJtB+BNBi6n1DU9NV5kZr0IpCVjxOwjpKB/H5OuK2DB2TZHWspj0rKLIYC7rZmjVmJzPpVUyE7vuPfjeY/DVMe4AZ9yw8oMNSDFCecw878p7aAH4eqCh2IatuiP3BOfO5LdK+3b+OS3cdS8o8J0QWF+uipddfz8PFnrR0k6rnq8SgVy+zu84wJ4EETcBLLA+KJYYrPZrPZx8t+nfC0Ey/dP79Ds9NObI5MhPxLR7eFIjp1DOt+ycQNRCftE4V/94QhPwzwbP2tzdiLT7PbX7sY21T3uRMTZxqJIHSnBRTzK4p5Lzi4SX/FGkkN2jrQJi3nmW7jCeRHEcuJ+RvSwaFVSD1FKcXtL1iAFT9aMIUOuzshnXKlCE5TwY8yyMYUQFg0CdygaSDksVqJxdxStz8ChqcrOjAqoJ4fh36Dqz5QW6A1k/HcyO9Oslpscp+fIjt/C6Idd+RAWDQJ3KBpIOcaiSB0pwUU8zN10M1e5SZgbca+JjWCnIwO89C+dp7iiCL0/lDTkTEQW6A1k/HcyOgNA3FMA0dsIjt/C6Idd+RAWDQJ3KBpIOcaiSB0pwUU5+SuzlDLH2bmzXE6Su/2aivh48WgeAe+AGrw5g00TiRpyenXn87dN39Aa216xgpgOImk+vwn70GlM7FV/qoydmdE8lMvwJei4zRM3BMuGLvgE9bnlZNhy5BMikM6wATmDA7z0L52nuKIIvT+UNORMRBboDWT8dzI9UdmtwVO0PMW3kjooUhSQTCCkB/cWqSlhSI6dQzrfsn1CU7K2tVmUTiJpPr8J+9BpTOxVf6qMnZnRPJTL8CXotzbM1hhunYyJs1xOkrv9mor4ePFoHgHvgBq8OYNNE4kacnp15/O3Td3V/w6VymHZCI7fwuiHXfkQFg0CdygaSDnGokgdKcFFMEqBWW0JLx7qv563jy/A5Swgg/EGv40FDmVt9hB5VFdcLg4TLFSlMP50r/6zZg8QnAlCJBb+ant+kwTowJRidXqpAPer6kaNEcRy4n5G9LBoVVIPUUpxe0BLRI3+DyLvmhjpELf/aCKWMF9WizK2bjKYpuXYGa4XRr0IpCVjxOwivkwtmFLeT2h/+1DVOfI06RR2zVUAzA8jVmJzPpVUyEKCcjwbuij8hUVhyWEPx3h0FugNZPx3Mj5/jRE8SyBFAOV6zbF9fA6RSxOoMvilz9WIIAIds2MSryTKIkUcCMHWlAqlLKErBpIpuHBpG5C2SSh6M44dDko+95b3xuiqJ14cMmgMS30D0UiOnUM637J7KxeGQcqauwd4iQbWx/SUiLSRYue6xyQgmtcTed3vOWbUXfYiX6zhRvsIoaBB34ibIzZIlGboVy/dAq+FwIsc8o0qzmM+xNkexjbVPe5ExNnGokgdKcFFPMzddDNXuUmdM3+t8ynYkOQcj1oMvj/BPP4IOPj2rD7GvQikJWPE7CK+TC2YUt5PYOg5gcINTo7nywa0RFid4cUzZu75YUdPUpOZdZQhNYheHDJoDEt9A9FIjp1DOt+yfyinADNDfiGTlldVhPPkI+Qcj1oMvj/BPP4IOPj2rD7GvQikJWPE7CK+TC2YUt5PYOg5gcINTo7iVNvb6LcPpV46FnwlZdCSgbz3Cmo3boVexjbVPe5ExNnGokgdKcFFOAvlz7SKybIXS8Z7sV3QKfnrgr/BC+fs4+7fMKTrRNy1RWHJYQ/HeHQW6A1k/HcyM9KJubS1PxJklBGq0NZ6EPHDM7s4tcKgHsY21T3uRMTZxqJIHSnBRTaG/Uv/vY6DOM+V+dOjIKw+OhZ8JWXQko5SlBBdGQPdNr0IpCVjxOwivkwtmFLeT2Ef/gKQa4BuUFR3aqwJTIx9IJYVZDMZbwKHKNfOIaCSwNu9GXfU3btedK/+s2YPEJyH2yugjmPZ1kGo8zBIu9yzlmsLGCk0KdWIIAIds2MSryTKIkUcCMHf8h5LLpZRdhdLxnuxXdAp+/dP79Ds9NOXCuVTJSltfSXag9LGFh998UiOnUM637J1wD88tylpEK6nNhMsihiF3K1hAN0qkLhEhhDilAIw0tIr3MTMixKR3bA8chY5Tt3M3gWMhyfR+Mi0kWLnusckKBxl0y+KwUu21F32Il+s4U2wPHIWOU7dwrZq1/nSg9wotJFi57rHJCgcZdMvisFLttRd9iJfrOFMjbiI4yTVEYzeBYyHJ9H4yLSRYue6xyQoHGXTL4rBS7bUXfYiX6zhTI24iOMk1RGCtmrX+dKD3Ci0kWLnusckKBxl0y+KwUu21F32Il+s4UpyenXn87dN3cTTNx7Jxvy5KHozjh0OSjyJask47xBrjhwyaAxLfQPRSI6dQzrfsnXfNYji9oG1j4Ce28IabRf4eI0VNEu+JYWIIAIds2MSryTKIkUcCMHcVNzNk/5DKQyPbkAJYLEsk1Zicz6VVMhO77j343mPw1VFYclhD8d4dBboDWT8dzI5aw7BlOiBHqrPRz0IwRjerqfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7NJjPDWUFVJ8GXyTP6ynHXLqfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7NJjPDWUFVJ8hpgdMxbwmo/qfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7F1K5Ds8OCWQGXyTP6ynHXLqfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7F1K5Ds8OCWQhpgdMxbwmo/qfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7FAYurdfid1pGXyTP6ynHXLqfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7FAYurdfid1phpgdMxbwmo/qfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7HfQBJMFZG1JGXyTP6ynHXLqfUNT01XmRmvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7HfQBJMFZG1JhpgdMxbwmo/qfUNT01XmRmvQikJWPE7CK+TC2YUt5PZV2JP4bUIOydQFXSg/+Y/Dayn+ngB8GIlS0pd/SoDbqxxHLifkb0sGhVUg9RSnF7RPQp01cWN72JEWaU5oIUtyMh1trJ430qHCCD8Qa/jQUG/3UNnM6eLtwuDhMsVKUw/nSv/rNmDxCfkmO47DGbmeTbl/EUOT3V2CNw2vYZ1NRI+ECzyoDEkO7GNtU97kTE2caiSB0pwUUzsbvkIC2oOYgTQrGf59SxcMZw6zxP+1SItJFi57rHJCgcZdMvisFLttRd9iJfrOFNsDxyFjlO3cgTQrGf59Sxedf6nBsXgvDn6BQePAhrS5a9CKQlY8TsIr5MLZhS3k9izRkTMzGcrsYRaoiSTcFSUpfoWQz0YWbrqZpHRFaSxbbUXfYiX6zhTbA8chY5Tt3IE0Kxn+fUsXBcsOI3TA2xl+gUHjwIa0uWvQikJWPE7CK+TC2YUt5PYs0ZEzMxnK7J4c1F7f0gw0KX6FkM9GFm66maR0RWksW21F32Il+s4UyNuIjjJNURis5t926S4NqQHSysqpY4h1koejOOHQ5KMsK+jXre5gqOHDJoDEt9A9FIjp1DOt+yeHgbP8kp4oYuxNtcbkLGLjt9w3u+6AUkhATI9K6TW/dliCACHbNjEq8kyiJFHAjB3xv0zWEMki4teswRCcJtoPtblVBk7nZxrqfUNT01XmRmvQikJWPE7CK+TC2YUt5PYoIk3/ccJlRDHr6HzrS2oTwgg/EGv40FBv91DZzOni7cLg4TLFSlMP50r/6zZg8QmFJV3FR4VTsUO5yz0DaC9CiDb5dVcOsGITCaQLmHTSSxxHLifkb0sGRVxgon0onxzMMsAQdqfI8218ivVi9/GEb2UQtFxHUvOtZUUNxhjnkvgAhU0hdZFD8Rp7kdD9W9cr5MLZhS3k9h5vftVx1b/p0mM8NZQVUnwZfJM/rKcdcoNxIMYhzmp74cMmgMS30D0UiOnUM637J2BOzTZFqEePfBch8V/FUQiSh6M44dDko8iWrJOO8Qa44cMmgMS30D0UiOnUM637J2BOzTZFqEePWErqlbR/kfaSh6M44dDko/4yfXr78HOawuDhMsVKUw/nSv/rNmDxCafZjsgn90a0jmP2c+QU2xLCCD8Qa/jQUG/3UNnM6eLtwuDhMsVKUw/nSv/rNmDxCafZjsgn90a0shZVy0qMOFxSbsE9Q+MK/ViCACHbNjEq8kyiJFHAjB3kIw7O/EbQUWzsgR+/54LWwgg/EGv40FDdiz5sAoFbqcLg4TLFSlMP50r/6zZg8Qmn2Y7IJ/dGtL/n5c40/HouJ+lEkYsDOQYcRy4n5G9LBoVVIPUUpxe06w8Ifk+Bes8MYggcGWYrj4tJFi57rHJCgcZdMvisFLttRd9iJfrOFNsDxyFjlO3cGxCMksGIlTY1Zicz6VVMhO77j343mPw1VFYclhD8d4dBboDWT8dzI2r9AqbPIQbtVdiCjiSqy7pS0pd/SoDbqxxHLifkb0sGhVUg9RSnF7TMMsAQdqfI8xRH6g+4YcPz3FM8vuzVXG+PhAs8qAxJDuxjbVPe5ExNnGokgdKcFFM46iD9yvR4J3uOBRbQo7WPNWYnM+lVTITu+49+N5j8NVRWHJYQ/HeHQW6A1k/HcyOWhhNhc/tm6/3QKvhcCLHPj4QLPKgMSQ7sY21T3uRMTZxqJIHSnBRTOOog/cr0eCeugnYA7ZxAZsIIPxBr+NBQb/dQ2czp4u3C4OEyxUpTD+dK/+s2YPEJDShEp3DmBhj25WSigQZFN1LSl39KgNurHEcuJ+RvSwaFVSD1FKcXtKVhm+/DsKKisXNaftNNASSwYqGyCgiLHAT+IgNtG1ooHEcuJ+RvSwZFXGCifSifHKVhm+/DsKKinG53X3/V1luwYqGyCgiLHAT+IgNtG1ooHEcuJ+RvSwZFXGCifSifHNvjoDHADN6c2c64Cr8XadaINvl1Vw6wYt8wKDiXsdoYCa1xN53e85Z7eGoQHY5J32+wihoEHfiJALbMopyIA7KNSiedaSd60obblYwMskv6KCcjwbuij8iCeH4d+g6s+UFugNZPx3MjizfuTM8H4iFce6gJfrhvWotJFi57rHJCgcZdMvisFLttRd9iJfrOFAvINRODNP02eyNjLtaVpdPBlFKzfwtBkFLSl39KgNurHEcuJ+RvSwaFVSD1FKcXtKcLd6wnWbHq9BFWe6f/sJITSqQuOXxiWoeI0VNEu+JYWIIAIds2MSryTKIkUcCMHXNszWGG6djITbl/EUOT3V0Yf+TYwVS4kI+ECzyoDEkO7GNtU97kTE2caiSB0pwUUwTWu+3IscxrUBi6t1+J3WkZfJM/rKcdcup9Q1PTVeZGa9CKQlY8TsIr5MLZhS3k9gABKduitEGGtYICTu0jmJeSh6M44dDko8iWrJOO8Qa44cMmgMS30D0UiOnUM637J6Gh3UVWoxcsJqpeike1brDCCD8Qa/jQUG/3UNnM6eLtwuDhMsVKUw/nSv/rNmDxCaHrgOTIq59GZqhUe+mBnjM1Zicz6VVMhO77j343mPw1VFYclhD8d4dBboDWT8dzI4s37kzPB+IhnX+pwbF4Lw5+gUHjwIa0uWvQikJWPE7CK+TC2YUt5PYAASnborRBhuaTooksoI785UPoysWHMRgcRy4n5G9LBoVVIPUUpxe0pwt3rCdZsepIoTKdzhpiG8IIPxBr+NBQ9Rgr2sqq3/LC4OEyxUpTD+dK/+s2YPEJoeuA5Mirn0YYpXq4jKQpyo9xeb8TeLxG7GNtU97kTE2caiSB0pwUUwTWu+3Iscxr//5CLNN4ngTKr5wcIRQebFMzMTd2VbLAK+TC2YUt5Pa0AFHfKT53/z3o+EmYPp9Bwgg/EGv40FD1GCvayqrf8sLg4TLFSlMP50r/6zZg8QljyqJycAgPR2EWqIkk3BUlKX6FkM9GFm66maR0RWksW21F32Il+s4UpyenXn87dN1dvVjznlk1jxuYXwitwQHjQEyPSuk1v3ZYggAh2zYxKvJMoiRRwIwdxU3M2T/kMpCLN+5MzwfiIbdpvtuCo9TYfoFB48CGtLlr0IpCVjxOwivkwtmFLeT2smwmnNtaYngiQpHci9AjyDVmJzPpVUyEm7JnuSs5/oVUVhyWEPx3h0FugNZPx3MjsExDDgvDqPc9LaGidc4WL8wp1kpdMEDcWIIAIds2MSryTKIkUcCMHXNszWGG6djIGOlRK8S506GI7fwuiHXfkQFg0CdygaSDnGokgdKcFFNjVw15zPf/9w4SmoRsz5QcuwWlpXTkn4OsPWg6FSenyHeAIBdpfm+xT0KdNXFje9j9zxObilZJy8xt7tWekkK/Pc0I368GozilaqHQ6HYhZedK/+s2YPEJkqal3AnGOSH+TKikSQkkQjVmJzPpVUyEKCcjwbuij8hUVhyWEPx3h0FugNZPx3MjewAGHEttSo9STO1s8R4om4tJFi57rHJCCa1xN53e85ZtRd9iJfrOFAvINRODNP02aW7rsgznvxKYVjWGVBK0ZKqQD3q+pGjRHEcuJ+RvSwaFVSD1FKcXtKcLd6wnWbHqM1bvZ+IR89E9LaGidc4WLxSxOoMvilz9WIIAIds2MSryTKIkUcCMHTpbX7ibJJn8P/b4Y7Q9hp81Zicz6VVMhO77j343mPw1VFYclhD8d4dBboDWT8dzI+EhI44TOkECY7qmmOMHCY7qfUNT01XmRmvQikJWPE7CK+TC2YUt5Pb9rNQ9pMjFpzQ7e1k80Qpni0kWLnusckKBxl0y+KwUu21F32Il+s4Ub7CKGgQd+ImVhqsillAnUmO6ppjjBwmO6n1DU9NV5kZr0IpCVjxOwqExlKxSUW3tOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2R+JOhZGjs2qfBzt+PhrTzkgFxsc7HdT9fL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk6xambyK5ZxNCQ3bmdTTHwSU9XczSMtPKNmon17on6hJWKagsUyzNiV40l1lb1OXtEisFUyYgp+4QZMeFQwgW5KeuCv8EL5+znckWoY56cgvX/VuTF7etTfBA2zjeKRdg+6gnuh/ZnB5q0SLj91Ue6/VmaIohTeKhzh9A8064LSKe1TYiCbn8biUzsVX+qjJ2SOL0yshwRnPQnjH9mQ9QSGuH3+zHgnhl/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk2wB+7h+Ops6cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPLFTffQ8Vjhg/cS70TOfxv8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTIGEjBijipE36BwFmlAXzTSDxBDjrObGCRYbPk+prwtwaeSEc5Yud1+Qkas+/4BSqH1MVbgl0uWN9j5IrXuK7RikPVymSji9NjVXFquNthLL45IRa06TYebRsC2Yrcr8TytzgvjvoHUVRCWbeSOoaDeYkZzDDBaT7mX4CuzABKAbrRpAsR9do3aOQsokbvxIJbPz/c6/JJ/2iPRAJAhOGHjxLClSgbNjYMHmt5YWbIR/K3OC+O+gdRVEJZt5I6hoN5iRnMMMFpPuZfgK7MAEoBh0HQCX0/WVTy2bpv2tbObpAhoDL61JMcTfs2T3tv7qu6My141/1x+n+6gxEhl/jcvaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMvBAUm9pdMPz5Glg3mpGvLgNjWIDNLT+IlZZnQOMdpQQdsw6G8w6O2GoNfGWRcbK31n6Cb21JXNZvW1uJ09i8hM0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm3zqGF3/y/2hqcZNCgGlPXmbglCZfq9SqOvnYUlb1kWV1eYB5ioJUYgzEE+Z3cjImc7LFBnXdjbx4HxInQShy2ny5PpLEgYovQYa77f8vmAHUNR+nZQ+kcxyb7OSusF1t0thbgHTTaRvWLuZjFfRZ6k1mfzUC43/Fd3K81fkl6moX7CWyVyXUgBvxFCll4lpueoNfGWRcbK34eankdbrxdvdWmDUGkabyyfis3C105LtDB5reWFmyEflhHj5R0eum2U55gx+/r5EpDRDzKAm9d6m+FBP5/V+6sYa77f8vmAHYHyuUN/TYhgNCu50u+mZD32qgcg2eo1NBPXNYKURi0fhcuOI5OOxTKDKkvY++Zbwb6IhgkZZbtUYu5mMV9FnqTWZ/NQLjf8V3crzV+SXqahSzsc7kDwkmu/EUKWXiWm56g18ZZFxsrfh5qeR1uvF291aYNQaRpvLBzcV/u2s/MqMHmt5YWbIR9k420gPMzwli6E8nLwjXFLkNEPMoCb13qb4UE/n9X7qxhrvt/y+YAdgfK5Q39NiGAlTb2+i3D6VfaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMoMqS9j75lvBvoiGCRllu1QASlQboJTlvsmhdMzPTwDOzEE+Z3cjImcCQZtiLovMJYRjIpqXdgry0dTODdBGb49xCvea/bRFrESKC5/XoIPwn5X61vvONpmfz+rM9N6t83NIoH30Y/1TpgUsNqHpUHniRElPR3NRSv7qDESGX+NyBhrrVfbC2BJ1aYNQaRpvLDf+GbhgpLcQDq3FKZ22cDWoNfGWRcbK3/nIPgN1sFPdk/viCEKra9VSU7lNyZCRSMPPBDcBy1gpYkpOYQqBvWc44KuW0tEdOvjwgmfs3gFhwFgsHfuuaTB1gRgLdL1+BSE2/WqAu5XR5hk53ZMwrsZpHGsRrrIuZ5XzRZzhb/NMC091b+oWTTHJWr97XimORG+ZYXaK5+VoqDXxlkXGyt+bgPsV+q+jK57acReV3fUoHQdAJfT9ZVP/ZWeN+olv2ag18ZZFxsrfkJnf3DYmgkpR6e8WClAHImkcaxGusi5n+FW5X3rK/qGj9a4NkQvW6XPKxSUCjyID4e9Dh8lxhBVriwKdAZkr2hV1/Sw/wYuv6/TSGMYmkCd1aYNQaRpvLJHLX41lHrivlsksW/e/RJaQ0Q8ygJvXegtOodBjAsd8xMn3gXsvzf7L8ElX1S2IieLo2KM9ZJd9u8is7ymztxQn3vCosVKNsxHIGztG3D59l+VJtD/uv6A2/ULkhwzXXqg18ZZFxsrftjgv6aFjGp5fBFRjSASZefGU7Yaa/ltVjHkTuid8rq/45IRa06TYebRsC2Yrcr8TlVceTXqIAKg4Fz2wTKAvWlZCe9Kqf+Obh5qeR1uvF288S/+qybeRrjPnogiOyLI4LoTycvCNcUsCgedoCuA+3Q4r3iaUp86T9++9kYXAo/KWrZ5ZKcPlTar3Uf148eWi+A2Q9roXEgnm0LJaASIpe2xIXvOJu4IsOOCrltLRHTp+mnOnSKRQEFn6Cb21JXNZUQDEX4lGWKytMg/TH8AwMJuwpfyRpuHUTMzqNaAeQE3HF9S0XUQIvJdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmcKCqXitt0N6Btxr4mNYKctAHpDVKFDk05tCyWgEiKXt8/VqgmtobsVnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZdLZvM0qnBXIiWVPnLuOv5i8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEf1CiDMyziG/IPNzaDvCFIaJl5pP+/w5LVg8M/XPHF9qDN8hwkaeXL9enkzBWt0tJvSR+EYhUn6yngsHxKdieRYm6EfCirzLRNjn0y093vawblg5fuBTrJou1+rpQQR+Jr2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTKYf5Ka5/GWqF1Y+ITbQJudUQlm3kjqGg3mJGcwwwWk+3TElC9B8dfJ/NCiX9/UY7UlX26L3zEegzDCDFQmIOwZqDXxlkXGyt9eREAmXnDwtjQ68/3TNPUeGmM340wuvpGzpuBjY2VybRGAB4d3kht7ANArKy9UxM1AhoDL61JMcTfs2T3tv7quVVtw4ikZM8KmnLdBGvECu/aqByDZ6jU0E9c1gpRGLR+Fy44jk47FMrdioAahW9MfuAif+5RWQnq7cHGcmccaLbdTi1x3mcIYkNEPMoCb13qgttppKKgo0l1Y+ITbQJudUQlm3kjqGg3mJGcwwwWk+/cYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaLtfq6UEEfiabTBt9inE+0XI2kGhH7Do5h2NmUzZZGl68I7wplOQWXeN2Kc840t3yqg18ZZFxsrfkDMKGytpghA5DvZFJtWwPVZtjBO6mc1dtQOf/kCuU5Hu2cXNH2ENcTqaIbAMJIYidMSUL0Hx18n80KJf39RjtUHDfgQTDHM+s3tuhVgWpeWhN/ZkCh8PGpTLzgBCqrCe1xM6IgAtBYCbyNJo9XB7TYi//KVA67Yp78bAujZ95cr0IHpdFep4nL4Bg1TWUJjZLLfyZ5DREnSzpuBjY2VybfrdlCN08jk03wQsbQn+yHH+6gxEhl/jcgKB52gK4D7de5Jwaop+SgX80KJf39RjtZZyfE+45JLdVVtw4ikZM8KmnLdBGvECu+zNWXIR7349svZocreqjFWWrpKnmLHyTfzQol/f1GO1U5kwTVsOpVJVW3DiKRkzwlIBGKdgzAnsgFD+rULB/nSy9mhyt6qMVeDL1Go9tUpeioJv280BYJR4Vr0xScR7MUVijJJDGkeqEPQTFGz2CFss0q2Qk0aD5bgSQbjEJG3MtDp30dyAqvO1NlDNPhOvtv+o6hWtmGM88v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTI9fIwYzQA4GgNA3FMA0dsHqvOorn9k/PWfoJvbUlc1kuyoBCnecoakC8OIornqDi8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEevRTlP7GPsob+7O8JtvNsEpqyMjJjOd6Dy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTdeswRCcJtoP/+r7mHvH0IImXmk/7/DktWDwz9c8cX2o5CRqz7/gFKofUxVuCXS5Y5e3XicDJZZfQ1pFmvl22ruVzBspFARCWZacAGSF9jAb2K6hMdSPTRyyImF4gLRZAeLoelQsoS2rdZW6GV6T+u2EV/5uS3r+fNJjPDWUFVJ8syQFQwHsB8uWcnxPuOSS3Rt8p0X0CdD2gTQrGf59SxdFS2m0Rhxp0aC22mkoqCjSsvZocreqjFWEV/5uS3r+fF1K5Ds8OCWQsyQFQwHsB8vb/PP8Oh3FIBt8p0X0CdD2gTQrGf59SxdrskEaZnwOXqxdYru6EBsCWsxoLAaN8uiEV/5uS3r+fFAYurdfid1psyQFQwHsB8vb/PP8Oh3FIBt8p0X0CdD2gTQrGf59SxenTLSfFhOuFaC22mkoqCjSsvZocreqjFWEV/5uS3r+fHfQBJMFZG1JsyQFQwHsB8uWcnxPuOSS3Rt8p0X0CdD2gTQrGf59SxfNgiPRdbyekqxdYru6EBsCWsxoLAaN8ujtJ1HzQxcqyeBpNHE6AO1ure8A8KaCEosl75f+1G19Yy2a8VzUKxdPm6vlv538ueskVp5M0JkVg6ZlWgsvFSgf0mM8NZQVUny3AuAs/L/6LDQ/oMOF4MMbW2z3zrfD5s59BDX0RjbgsDuIYx+sMCpeSpKqD9UHtEGhMRZbXxk9rKg18ZZFxsrffQQ19EY24LBSVAvyGLNP7dQFXSg/+Y/DGlqDXon/BIWBNCsZ/n1LF+P2Tm9llXVZyWSCd8UjJTcOocV65N45nYhXBDOhBH1FKeQPCOwHc30Xzw7EV/WenoBPW55WTYcurF5UEaGE8BBc4sUPyiMvv4iNPLs1jxwFQEQ+N5EuuErjqS2b4yIpdqzm33bpLg2pAdLKyqljiHWIVwQzoQR9RbdVdc/6vWrbSpKqD9UHtEFKXBKO9XCukH0E/+qieaVTMti97efBM2gmjOcw44iM30qSqg/VB7RBcgSHKsJX9UIOocV65N45nQRM5a3QoG6cNv1C5IcM1159+qWmlydBZquwSwszM3a50I0vWN9MIT4ZFctCT21fIXAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTXiu5UQV8FENUHJ01rNlq0ri8y1dJoq9dNBS2whqH9mEHMocwcz6EblQcnTWs2WrSg2UaAsx1tH5/5/InIEaeQ1JJV5ASN217JoznMOOIjN9312Ws+pWq16+ANuIaJlP7Mti97efBM2j+mc0j4BRwi69nm6T95JrFcrpLydPnYbCZqNZu+vKzrvuij9DmRkw7EwsDimEewrV+XZHMoLgi/ffiIiklSNkq3RzaCsSl8EC8DE7GlI2gQBdN/5k1TtUWmQuDrbCd8gQa51AKrdKfyKxxATWFVpDn8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/H97zWiwGO4gPTpcLDwCAwEcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPzpqcbuHqpfkUiFX6ucTVQhs1ODzxVU26hYWAR161KjWdq6q+4iv7MalCoso7qGU4bmKMy8DBAMqjV813ehqxtgPPvH8rhYwxTNm7vlhR09bmYpk9pEF9gwuDhMsVKUw8vFfG+fBhu2ssCk5CiXq3flyJNSZWXY3L5W+rEb8XoruEkpZ1EwtkI0PjHSkdNmghAuqEmiSrMnDSc3R/HQ5ndOSHV1ZqHYJlRCWbeSOoaDbQLbwE2vp5paLqzJmflsPSXt14nAyWWX0NaRZr5dtq7lcwbKRQEQlmWnABkhfYwG9iuoTHUj00cUDPDrcroLQg30TxwmqyEtDyysjm0YoAWqWHocdWP2uifAPOJZ5hkzM1ezGbHNKH/XRgIlQNYHRw9KJubS1PxJkMwhzoXyEYq19g6lp1V+7GiuSxudVJCDRaJiTslwsXZGW00sQPhj2HLgs+B63nnzqCjVRLdaXwd66Iair6YAZJ0gwoF2P6DULZHfpHkei6vwFgsHfuuaTDAWCwd+65pMKiao9ZS5E+V3K0BMX5li8MBwBPDHhdUeqxeuD6shnAJn5PxXDoT3t1pXZsUodBpfEC8OIornqDi/0+nXrAtOe50WCl5tquQpORGAqNNDZF8cfLXy3xyXq3Q+MdKR02aCEC6oSaJKsycC9ZMPlT/XfDdZyxSv4Zf/Xw73+WakMnJbEhe84m7giw44KuW0tEdOoPAwalWIkWMHXasYX9cU6KDPmhAtpi4ZmsezOrWWHiu9orqZYAgHpvNQ9JN+x23ikUiFX6ucTVQ8CiSttW2UI7y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPFpbEnY3CktyVOMdBkfdnjQ7016U0+K/3IfbK6COY9nchpSuQmq6TBe26IMgzJNWlKkqoP1Qe0Qd4LveOj/NI2I7YmO/Juo5Wn5YoT0Abrb2ue49BHtuyBvWBA5bsASShMIKaHK0YKEl1ul6GEKswzybh0OcInYcCscQE1hVaQ5/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxPE9t4zk7Q4eAc0DG94l4sKGoL2EFUF5oWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJO0+9OeXqeBZEIlQFgYMNRw/Ex7qZTK5HWFf1lN6qbqawiZh+PEFdAj1/PJ4sblFSDJNH5QjMIPaPeBG8KWa740kKxaDasfPpti/QZxTA2ygikJuMch/Os1uWDl+4FOsmhklm0yLGFEkG+kvUXQ7VbvsR10XrjdKUSn2Y7IJ/dGtIyl9TPv9aQY8Akk+MZCkjxQa9NPTh61csaBMYSGv4d94vTbZ33JAvgHAEEBNnDrw9JjPDWUFVJ8ovChepCyRuHXrMEQnCbaD7h5HJpZ8UFg8T58fugMkrRYSuqVtH+R9sQB2b/uFxUshXVn8uxRcdTIfbK6COY9ncwvVJ4HZdpmW/XOQYwY44NNuX8RQ5PdXWWLZ9yzgwesbXyK9WL38YScKTuURxbQ/O0nUfNDFyrJcRcJDUo8fEdB6b+5wfP5ft+DlieiQjQwjB4lYwrh6+oSBbque5PdCNJjPDWUFVJ86t8wuTNiFPSrod5EjTnxuslMZq/nPC1mBwBBATZw68NJeu9TPMn5UqfZjsgn90a0Ot2vJvzuloPjYHmHIQ10h3Ayk+IiB0GEBEzlrdCgbpw2/ULkhwzXXn36paaXJ0Fmq7BLCzMzdrnB3fJ3X1lv+lijxMpjjZ4ZWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNpYBh0eiRuF+9AMCS2HM0oNgf6eFaaM/w67OyGdcqUIUScDcCKHI1bcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Jgb1e9FaeuJQqUP47Zts2kImyODlNNZJBvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyBhIwYo4qRNIIEuW/bgSsdCJUBYGDDUcCYSqmwD6x6P/FJxES+W2uwcNkxGAV97U6sYhKLmkabLLxXxvnwYbtrLApOQol6t35ciTUmVl2Ny+VvqxG/F6K7hJKWdRMLZCAVgSqTJ69V1Y64/DcGpme1AhoDL61JMcTfs2T3tv7quG3ynRfQJ0PbH/Tuy6YXF1jQ68/3TNPUeGmM340wuvpGzpuBjY2VybY7ZnRJu8d57Tf8RgiVrHHA0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm1aZTVtdcidZk3/EYIlaxxwNDrz/dM09R4aYzfjTC6+kbOm4GNjZXJt/IfhQIZsaT2RB/VAmrYbaJXZg+ub6CpKQIaAy+tSTHHkQK/WNyYU+xpjN+NMLr6R6NLvPlfAjkbII4eyFRziJQ247Akmt7VKyLp3vGdAsWslX26L3zEeg4h4BdF8CI0lZL+814w1rJaskPxLL+8gffcaLydpsQM0S7519g7oX491FiiUOkfRs6a35DOqZ0CrvxFCll4lpueoNfGWRcbK35w5rfimeDIdUHh6yh593qrXrMEQnCbaD3ESIhp2mBn38n2qUKCbsXpAxDl9RRXHVCUWghz150BsE0aZheK3Y6vAY9hMEVNowfyH4UCGbGk9kQf1QJq2G2guROT6lfVa/RlSpy5xnLMiAgT227uRo+UIloowW2NqfEO5yz0DaC9CbEhe84m7giw44KuW0tEdOiCfPNFuEz5DGVKnLnGcsyK/me1x9h61el9C9Fa8In6vAdLKyqljiHVSQiTI9fxSylJJV5ASN217Q7nLPQNoL0JiqNKeR+wbkA247Akmt7VK3KjZPqsRiGA2n6KkkWCc76kKusz0wYsiUklXkBI3bXtQh6O91SYXA6g18ZZFxsrfs3Loq3+daHh6IfOpWQZiMKt/6obduUPpLy6osqpOnWtxzX8IzbCgTrESjECqoTOlE2vz5fSFcLHLf7OcpqTG3LOm4GNjZXJtWmU1bXXInWbo6D1NqqC2u77ri61RX9XzkQf1QJq2G2h5NVr6G45QSAa6qlo4d91NeVj0Bm75+Nmu/BBmSMNhoNcTOiIALQWABWBKpMnr1XX1MasXt3Je5z1MWKLPPEQJ3wRV2REAOwNfQvRWvCJ+r/Uxqxe3cl7nf4KQnX9HQ/nfBFXZEQA7A2o5HDNB0yTFogIjR7OGoDeFf1lN6qbqa/UKIMzLOIb8ictSiNgW/7/82oKmd1HV0/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln5/L1dVnCSXV3NinA5JzIHRwJBm2Iui8wlhGMimpd2CvKWBNo/t02XSXK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiYb4NjkZHww2bP3znU/tfvrxRI1cnD8VOzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8dME68gBnvurfdvJ74Vf+IcmXmk/7/DktWDwz9c8cX2oM3yHCRp5cv16eTMFa3S0myHtmpgoIVG9Gqu0gl7pG4oOV6zbF9fA6YeI0VNEu+JYWIIAIds2MSqzpuBjY2VybSCi1UT/oEeQbEoVhd0E5R9juqaY4wcJjup9Q1PTVeZGa9CKQlY8TsIDXHDjv1yxOgAg8H/eMiiu0TJg68PxohySh6M44dDko8iWrJOO8Qa44cMmgMS30D0bmKMy8DBAMqjV813ehqxtnYSSf8uMLUzCCD8Qa/jQUG/3UNnM6eLtwuDhMsVKUw8vFfG+fBhu2ssCk5CiXq3flyJNSZWXY3L5W+rEb8XoruEkpZ1EwtkIMZzec4NYb6ar+et48vwOUjSc3R/HQ5ndZL+814w1rJYvxMuc4I56TjfqZVk0CUssvXcglnBhkDU0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm3W6GR/nSUEpCz8Jbk9XpVdu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6wJQiQW/mp7eI3HDwKglicSVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3706yWmxyn58eq86iuf2T89Jz5ieEfkatPcaLydpsQM0S7519g7oX491FiiUOkfRs6a35DOqZ0CrvxFCll4lpueoNfGWRcbK35GR9v5140Zjfo82rx1ARv8RO5zafLLM3OYiqiWWtCZqN+plWTQJSyxJb3vtfaweaYyugcbJlLq11B/hnW2VFgKoNfGWRcbK39boZH+dJQSkDi7bRPfSArJsR6DJqCUVyqJrhHCVEGtbGGu+3/L5gB3AlCJBb+ant8gGZMNnOJAmFQRTQg1Qz1CoZdbSBAJ1D8BYLB37rmkweygR1a92YwMnUW7njO3Sez8BqKRjeRUOt+MY7xhd1OP/VThBD5Uhz9YPVpt3iCD57pGVIJuZfk/n+NETxLIEUBeAIzzXgm7ZoSpQgBt0sRIpuQHGbGDppiF0aihglkmU1g9Wm3eIIPmyNcfwmy5SoZKga1YesxCgtpJDG80CZhhrH94qFsHdXOBrhOuzEZKSUQDEX4lGWKwxnN5zg1hvpvho39ocamqTfPBntcaziknsGlVUz7L5yZDRDzKAm9d6rTIP0x/AMDBVW3DiKRkzwkt823SW/R2iCXNkpSkyQv7DHzwZbJ7YCykxBOVOb0E2dAZGmnX1qCi7b1/bmJ4Tra6YaK6MHNtgXMZyHBq//8yKPVGY51VV1kVbZy8pJ/RImQuDrbCd8gSWnABkhfYwG9pF9h3bz9HOtY2ChAhRVj8Jl1NFOe4kqtLo+YNVEj9S7MbH2rBZtT5MNaotUtg8tLsAWh//fc5aqGXW0gQCdQ/rr3MUWOscivflsg/0WVC5k/oV+KvNGVm1b9voaeofh1/440+5RR7TPV4hxirwMUplTF2+N3xKiydod/Ond8KrCz4/agvEWoOubwYQkLOH0iJo+78u61In9vRlVxuNBNKtSBpYKGglSsCUIkFv5qe3V0cMx+Kv2f3c1RXu+ASqfoAA7FXlHWIfk/oV+KvNGVm1b9voaeofh6dkxe0PHbEs05WlmcxWU5mwEij91vJWqZDRDzKAm9d6G9mMN0D2P/ak3QePlbRsxiLMSFB9p6vVPgVXQMWUer0Cvn9oRv44mnsoEdWvdmMDF4AjPNeCbtmj3iIBMOu2QzVVmlW4swPlrHdbvdZZbA23t4R5I+jgOxpTyVI+0Rbog20tG8A6fN827xr4UtD2lRhrvt/y+YAdDShEp3DmBhjvfucLnmY7zwTDZb1Jh0nQsMdWVVIHobzwTbDAWmmQL3ZS+x/cgIHln5pkv+29tQA7hw+8jMcJvmE88nbISAJHrHdbvdZZbA17KBHVr3ZjAxpTyVI+0Rbo8VFulHs7TBGia4RwlRBrW5flSbQ/7r+gD1fnJnzCLtq1jYKECFFWPwmXU0U57iSq0uj5g1USP1LWD1abd4gg+Uw1qi1S2Dy0uwBaH/99zlpBAULY/Z3PHeuvcxRY6xyK9+WyD/RZULmT+hX4q80ZWbVv2+hp6h+H6hYCVnK6tyw9XiHGKvAxSuwaVVTPsvnJJ2h386d3wqsLPj9qC8Rag65vBhCQs4fSImj7vy7rUifGLAPFSbSS461IGlgoaCVKwJQiQW/mp7c1F6qgSOWLOdzVFe74BKp+gADsVeUdYh+T+hX4q80ZWbVv2+hp6h+HkxzJjwVNYWbTlaWZzFZTmSKbhwaRuQtkkNEPMoCb13ob2Yw3QPY/9qTdB4+VtGzGIsxIUH2nq9W8dzuDhxkyuwK+f2hG/jia7akzeH9Wt1EXgCM814Ju2aPeIgEw67ZDNVWaVbizA+Wsd1u91llsDef40RPEsgRQGlPJUj7RFuiDbS0bwDp832TaldLgfTclGGu+3/L5gB0NKESncOYGGO9+5wueZjvPBMNlvUmHSdBkZLXtljtbkPBNsMBaaZAvsjNkiUZuhXKfmmS/7b21ADuHD7yMxwm+YTzydshIAkesd1u91llsDe2pM3h/VrdRGlPJUj7RFujxUW6UeztMEXc2LLIQUSV4l+VJtD/uv6A2/ULkhwzXXkTe3KALTTmkxsUzRLntQIFIqjQdmY20w2MScYILr8nKiZjvtPUD3cSpw0Y6nHfIOLFzWn7TTQEkNWrYpVucuCtMNkpqivOHwhnKVJ5kbyk23KjZPqsRiGA2n6KkkWCc76kKusz0wYsi0N+JEZC++Y6Q0Q8ygJvXekmfK2kzO7tiyLp3vGdAsWtXAcLtp0uZbesj33dP6cGqDQgoGk+LoghA9UcyaQ1b07cGtZTTW0lmu10OlI7Kcfe4o+rELtG0r2CaTrEplOv9TDZKaorzh8IGbvZiXsyjpkw2SmqK84fCOisph8/gxawWu86DM8FPLkGK0kCQb+z+JuArOjbYDxGAAOxV5R1iH5+aZL/tvbUADGbasUVKklEQasdgistmE1MAfNQn7pi183CpvSddyU+ZYiVWx1lcYdyo2T6rEYhgNp+ipJFgnO+pCrrM9MGLIn2OSVadm6r+TKVS+fDCQUKtMg/TH8AwMJuwpfyRpuHUTMzqNaAeQE2hnIvEqGgKSNXYbEBvMxW1cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNEqlxRRwUCgJaGE2Fz+2brKQ5uRK95glexc1p+000BJP6czgXuboJkdCLs2mCxTVNatqTBUlyP2dx7kaiycy2ZdLDqCJsjzKEi/IPGWCoHNtj7Q3h6NJ7Yra9aAEFD8ODOzyb4WaSBlv1+Afw4xpmdH/Rcg2T4nO/JYaCE0WWwV6O6FjFNPKKIFu9gUdtGZ8T+nM4F7m6CZFnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZdh7PIcUVpaX32QeWZHnQvJ8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/F8al5pOzPXnK2aJcYezxxD5oyoIXeJbFssqisAKpLZ9Cem/tdTojcxABpLkx4DeSBlzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZqtolvJ6JyuxOzkZ5XLSI2Dag18ZZFxsrfizfuTM8H4iFjr1tDcr0nQOrzCup29yc4JEnllLjIiqigH8j97JF7ZPQRVnun/7CSSTPx7JpBH3nc8I5nhc3JFFEAxF+JRlisF6G4lYkQK1w63a8m/O6WgzyPrhAZoHsommuxJZ9+SSmoNfGWRcbK34s37kzPB+Iha7JBGmZ8Dl4NKESncOYGGGiltrHRijybWjUu0c26OCZ248PcNP/fQDYhvoxpF4ftFEfqD7hhw/OcKTuURxbQ/CKXN9AwIpGFtYICTu0jmJfT2MYMpUPXkfPQgrWiPALPntY2hoxEjdh7I2Mu1pWl0yw31CEDEPpmav0Cps8hBu2+EjR0npuqLlo1LtHNujgmKeQPCOwHc30oAV/uiNJ7uWQPlj3JDLZCUQDEX4lGWKzIrYnIgvY8cII3GJU310hIqDXxlkXGyt+LN+5MzwfiISRXZeEO95njq6HeRI058brbKT5m8Xzrfauh3kSNOfG6yUxmr+c8LWYilzfQMCKRhVts9863w+bOizfuTM8H4iG1ApPbuXYyG4s37kzPB+Ih4iF6ICcy/rugH8j97JF7ZEihMp3OGmIb+hWb3LoWbbwVoI9zVSo3v4KapVqiRmGitYICTu0jmJeQ0Q8ygJvXeqHrgOTIq59GJmGb4TafsQv0EVZ7p/+wkve7dY5Hmwcd9BFWe6f/sJKsXlQRoYTwEGo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa5mi5I5hfW+zGRXLQk9tXyFwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3WRBYbZjfDBCo4n/x97HrzNinA5JzIHRwJBm2Iui8wlhGMimpd2CvLW8genp3nEPjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyvnnKX1cBwe8AyqRUp3Gnve3yLki3bibXJsjg5TTWSQby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTR6f2/rGKUm6zdqaoR8Vowbo4qykUuU1hyZ/SDtPy6KROZ2MLP56m91/Q3YtcqFzn9fzyeLG5RUgyTR+UIzCD2jV1nSmtbA90OzKeOakhOUTV5gHmKglRiCjhG4beAcEch6f2/rGKUm6BBmLc/DklrVRCWbeSOoaDeYkZzDDBaT7o4RuG3gHBHIen9v6xilJulbFwslpr0+NUQlm3kjqGg3mJGcwwwWk+6OEbht4BwRyHp/b+sYpSbrGHvhbWhrIW1EJZt5I6hoN5iRnMMMFpPujhG4beAcEch6f2/rGKUm68rTEx555MqNRCWbeSOoaDeYkZzDDBaT7oB/I/eyRe2RD06ZKOxjpTPHq5bfbk4rSbPz/c6/JJ/2iPRAJAhOGHlo1LtHNujgmwh/4DHdrSAL2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTL3Gi8nabEDNEu+dfYO6F+PdRYolDpH0bOmt+QzqmdAq78RQpZeJabnqDXxlkXGyt9kcx/p4foiFBPnedAgbGM0izfuTM8H4iF+K27BmNPaPIGAnvueMkLeB+aQ/+cVPEacXqvRwOhsL0pcEo71cK6Q/auuQkqIl6iZc+dqyDmN6DQKBcmLoXUzps6jUsIsxoOjhG4beAcEch6f2/rGKUm6JmGb4TafsQtDZT1zmdUdsag18ZZFxsrfsExDDgvDqPcuea/JZVNP2V29WPOeWTWPrHV3yM1I7DUxoSRAcePrbHg+hS0ejj4YwcesO5ZsEqeJRkkmMiKGuL/upSyKfvPZxTiGUmZ6kCVIoTKdzhpiG6nvgA4oVJBkHp/b+sYpSbopoTcoCFi+Lh+pBQUd/IzhvoiGCRllu1SRftjjGWJHTTrwQPJBxam4AH9N8vNzKsuaCXfrnlSWcnG90bLZRE848v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCThSWX8tsfedPx5s/gb52lPP9SGguZxlVw0AekNUoUOTTm0LJaASIpew6zfVlYV37XOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2QHGoib4C6luzOMNiTSfs4EmgWrNl8ART5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmN/vNvNnELELRkJneEdv3rnaPBZ/13BeeNoxbI4me9pimZFIuqsPI4YDrXOrkvJEoAM0VMcNdjM/m/fPgGiWhA7BvkETgs+XWGnkhHOWLndeYUieJ1YegZdiuoTHUj00cqDErw1ThfbGU7VrDN8NfmPaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMolGSSYyIoa49GTRF6zpt2h+85HZecWuVWz8/3OvySf9oj0QCQIThh5aNS7Rzbo4JmivXTTcnB78X85afUIPTVlRCWbeSOoaDeYkZzDDBaT7oB/I/eyRe2QzVu9n4hHz0R+uHWPs/vISQIaAy+tSTHE37Nk97b+6rlVbcOIpGTPCgb5omef4MLL2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTIA9ep8vX5pOx1G+6PPF8Eiu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6Y8qicnAID0ePQYbkacjSXCdeSVEBdcPaLwdkQahPEIOBo8aI3e2NZA4SmoRsz5QcpIT3ce60XvJ2qGJ/T63OOPcYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaJYHVFCkyjKo2jSfulCZUF3v6Lme4o3Ymwo7RsYlkEXyWKfcPMjclXh8aP5VfZylvKe41mqWIQm6kNEPMoCb13qSpqXcCcY5IfrNx2ec/K5PEubNgLUCnDE9TbRnjQLkYw08zc6vAj5WKLm1tWbhqqpW67dAVN7b/ag18ZZFxsrfewAGHEttSo/9cxCU8JqaDJKmpdwJxjkhJ7o2QGsj9Cie1jaGjESN2Glu67IM578SQHEBG9CbUyd7AAYcS21Kj/HqFE7O5cHsqDXxlkXGyt9t2rMcl8Fer7Q4A9Ut2sTHltgzb/UQpAHY0ncO/huVADudpJy86nmIo4RuG3gHBHL9zxObilZJy8xt7tWekkK//6YNQLRwHeywTEMOC8Oo99A9MX1yFb7bqDXxlkXGyt+HhJINuPA8+w4SmoRsz5Qcfo82rx1ARv8RO5zafLLM3OYiqiWWtCZqvw2+/GkjeP0Im+/CbkyXVqipKfrZ4oariog76M1gpCesSCpEIzenkpKmpdwJxjkh9+qP3omDG7MYa77f8vmAHd7b4gHqNbarZQqJeaycKAnvTbB6rYie9K/ieSfkGwQtYLI8guliKJNpbuuyDOe/En29qKkoTGZVAEpUG6CU5b5rHszq1lh4rmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa1E8SHrrD8e1ajDRsE795I9VaEqJdyTGF1nKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTNyQ3dT7+qhvy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8W6vjSPm5YQc3eCsK/0mfbvC7kl74s55mnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTJOt9hnGoEMpdoavfMvuAaGfxJQcoKRy75oyoIXeJbFuwNu9pJr5KepciTUmVl2NyLaph3YSB0q0NBQUlLIPgxU2EM6jlg+dX8wvcQ79a/M2OHAgZShzLsag18ZZFxsrfDB2TZHWspj1fzlp9Qg9NWVEJZt5I6hoN5iRnMMMFpPuhKlCAG3SxEhzWEKD2PpNX9qoHINnqNTQT1zWClEYtH4XLjiOTjsUy9xovJ2mxAzRLvnX2Duhfj3UWKJQ6R9GzprfkM6pnQKu/EUKWXiWm56g18ZZFxsrfkZH2/nXjRmN+jzavHUBG/xE7nNp8sszc5iKqJZa0JmoiEFgcKS80jJCGwyPdZ4tc3tviAeo1tqufmmS/7b21AJKga1YesxCgTFc+ZFbYaF+OvGyENI5RRdDGO9kj+CC/AEpUG6CU5b5rHszq1lh4rmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa+EzWJzjtpJnVZYjAhYqgUglU23QLyr3EPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8WlsSdjcKS33PQklR7DhT4XlO9ypc4G/SbGr8YxPH9rOMhyjlfrwIeN+6jE6JHeCx57zd3+dWiRLsT1DdvvEkKq953i5K6w+jokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyUf7ZcmeleQOgPh4Xj2cU5J9rW544mZIBt6zOdYdO1R5ZHlvbxhQv4lnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZfV8l19ijFyIQyfS3hMS+9kw+ZeNpnwdkS0byk0i9kWa7nQQQixnI7IVBi0BQyCqiVl5iu8XGxV4z2TQ1QOCohiC4j2MM04Y1G3t4R5I+jgO+DvNscTmwbco8DxcgTS24wpoifs1g0sYgvlmBdWPHvsnq4OBrnon/TsxsfasFm1Pt4Mvp02gP+vS+L9/PrJ7L3bgdhqyGFu6YyBQjaes1fNpH+iYXN2p5akPIN6OlF1sbK2EmmuheO87MbH2rBZtT6O00zWO5v4Fz7fBSngAeVpmkFWFrOe10MVdf0sP8GLr5jSWuuVaacAWvoaopidl/Jg5Lf+K6r8Q0tTLOeaynmp4CiHdOOQTLlWc6EIahcCuHARTTIGopTtkCe0K4KW5X6IRA9P38j2lKGOkQt/9oIpSp7agx0oPXIpUXp5yCcn5nSDCgXY/oNQu2TXWro5hPI04YFhHx3eUyABH/yjI9FKC9UxHq3ksiZqClTBqby2HMcIh/gOQ6jVW+PLWHJwcdsoKmVcgLNIxdFBzzIvZu6EsIv8frgmXJJlTF2+N3xKi7wPLueC2ZXK+GiIvwPqUc4xlom6SpJyQcvwSVfVLYiJfGlklIOOUCd0uP3scM9aVcMVHSMhCB3Eqk1Lr7M0vAw3pOvMiZf9UgkNgHZGapfQcHxRN4xA7uvQnwX6xBDqmwETthSNKlAc1zMViyFVrlHLyclcgJ/T+KuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSE7UK/CN/hKc2MftVaX1jbS0/SkN6W5/RuPvqfT7jbb3fAg7dd8A4oBeHjgSu74bb8MV0T8SMBWoQPebfZZNmjU7nciSJM/lScpaSeInzJC1J3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb4VBFNCDVDPUAF+9KDaJKdluLoA14Onzj9d5S7zHloRbZf0NAqtoDd7sOW9w8BUFblrS1TXObGJTjFtQQ50vLzhd1vEdc79Hexo/rRCPEaO2Q/IYWiIqjyhXlB9PcWZIklyA8lDag+GgwKqZTd3FRM1PwGopGN5FQ4UHpW4r5KymqwOHA8m2QIr6Q516c/U1i+Oa4G0vYE4WCxFxpn4Dsyz9rmT0ugJIkAaGVCbZOT3hsCUIkFv5qe3lPGe/JeCeh2ZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4u2pM3h/VrdR50bbJiIZC3e0byk0i9kWa7nQQQixnI7IT7duLr1b6xtl5iu8XGxV4z2TQ1QOCohiC4j2MM04Y1HV25U9Uq4lMvuLTEYhdwuUD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDAqplN3cVEzU/AaikY3kVDsN1GxF8bVtarA4cDybZAivpDnXpz9TWL8BiL2AI2jGTLEXGmfgOzLP2uZPS6AkiQBoZUJtk5PeGxors/i7NUfZOCM34lF8GUyd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+FQRTQg1Qz1AsJW2OIXB1B7i6ANeDp84/XeUu8x5aEW0EH5Izf2RPqV4eOBK7vhtvwxXRPxIwFahA95t9lk2aNTFKywb/ZbsY0fk+KBarJZy8Dy7ngtmVyvhoiL8D6lHOMZaJukqSckHL8ElX1S2IiXxpZJSDjlAnJljlkQz5247DFR0jIQgdxKpNS6+zNLwMlTJW2tuWBBpb48tYcnBx2ygqZVyAs0jF0UHPMi9m7oRsQ6PkL5h2zF0Cops3nOaUStTVULFxDyM+3wUp4AHlaZpBVhazntdDFXX9LD/Bi6+Y0lrrlWmnAIOVnCTylVhzYOS3/iuq/ENLUyznmsp5qeAoh3TjkEy5AgayiJy279Okf6Jhc3anlqQ8g3o6UXWxsrYSaa6F47xO8hukoSimAs6ADuCH/t1YmWM7sg7m9pItp3y7fmTZdcVSVVRNYpozshsyfOCZT+Ln+NETxLIEUBiU/p0DOgMLtG8pNIvZFmu50EEIsZyOyIplkdhOUHyOLEXGmfgOzLP2uZPS6AkiQBoZUJtk5PeGxors/i7NUfYi1UmvxCq2Ayd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+FQRTQg1Qz1ABfvSg2iSnZbi6ANeDp84/XeUu8x5aEW2KOvrmQrsyv14eOBK7vhtvwxXRPxIwFahA95t9lk2aNTFKywb/ZbsYgflouSyzQ7e8Dy7ngtmVyvhoiL8D6lHOMZaJukqSckHL8ElX1S2IiXxpZJSDjlAna/mcyvVdsqzDFR0jIQgdxKpNS6+zNLwM6179c57c6tdb48tYcnBx2ygqZVyAs0jF0UHPMi9m7oRsQ6PkL5h2zF0Cops3nOaUIfo+LNS+G2Q+3wUp4AHlaZpBVhazntdDFXX9LD/Bi6+Y0lrrlWmnAL8r3pApf+vIYOS3/iuq/ENLUyznmsp5qeAoh3TjkEy506KWkBwNGU2kf6Jhc3anlqQ8g3o6UXWx6lc2YFG6GztpHGsRrrIuZ6VMzWpAWqw3mWM7sg7m9pItp3y7fmTZdcVSVVRNYpoz7Y3mi3e5824dB0Al9P1lU1EPOqDVn3NCtG8pNIvZFmu50EEIsZyOyPbyvIjEXLmZLEXGmfgOzLP2uZPS6AkiQBoZUJtk5PeGogDrY8w0JEjDTcC/whQl7yd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+oJYTVfKonDWX5xFdfKFrG7i6ANeDp84/XeUu8x5aEW0/bgZIaf5BR14eOBK7vhtvwxXRPxIwFahA95t9lk2aNaFtpeZyOIqcKDmlhXEIPcEnenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvhTy5ECdSP9vD0CRkVZQ1Cu4ugDXg6fOP13lLvMeWhFtuq0ux7PeRANeHjgSu74bb8MV0T8SMBWoQPebfZZNmjWhbaXmcjiKnE8Lnbawo0HHJ3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb4U8uRAnUj/bwWq/DRK8wSnuLoA14Onzj9d5S7zHloRbdpr+ZC4yq0JsOW9w8BUFblrS1TXObGJTjFtQQ50vLzhw+r2cJXreqH561IRAzEqwCd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+NKeerljP17muE6JTDfvrb6wOHA8m2QIr6Q516c/U1i/y1IEAX0f7sCxFxpn4Dsyz9rmT0ugJIkAaGVCbZOT3hpaFXVriTBzXy8nJXICf0/iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUi6/DQ+ZOYvbcMVHSMhCB3Eqk1Lr7M0vAwWMRMuNkrGzQAIENq7GEAzcHxRN4xA7uvQnwX6xBDqm1ATX2nhzMFdC6RJeCfkY9Q+3wUp4AHlaZpBVhazntdDFXX9LD/Bi693CqaFP+lbtDOfWRtly443S+L9/PrJ7L3bgdhqyGFu6RSppcJyXocTpH+iYXN2p5akPIN6OlF1sSrsh4MqBe/1r3+4nOQ4SwcPyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoMCqLbkLR/PoJQzJ6SxnPmXuLoA14Onzj9d5S7zHloRba1VT/kIUyL6sOW9w8BUFblrS1TXObGJTjFtQQ50vLzhOjAHB5VUJi68Dy7ngtmVyvhoiL8D6lHOMZaJukqSckHL8ElX1S2IiSAz0BU+sVVVC9UxHq3ksiZqClTBqby2HK78NVxnZNe1O+s8ug+1q8YoKmVcgLNIxdFBzzIvZu6EYpeHW65Q7ClLc6Z6890kLid6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+PSibm0tT8SZf9wWEKqdZBEtTLOeaynmp4CiHdOOQTLm/sfa9jALcjnARTTIGopTtkCe0K4KW5X7ah3mwK5S6Gl3LwK1XIasPpI1CoiH+uAY+3wUp4AHlaZpBVhazntdDFXX9LD/Bi68B3A2T3qpozIG3GviY1gpyC9UxHq3ksiZqClTBqby2HK78NVxnZNe17ru/9ZjM+U8oKmVcgLNIxdFBzzIvZu6EEdmj9azFT33XrMEQnCbaD7i6/LGWU6AbKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTyy233oHX1+xTf3g5QUFm9osMVHSMhCB3Eqk1Lr7M0vAx55QNr85CZMAAIENq7GEAzcHxRN4xA7uvQnwX6xBDqm1MvRQL67+kiAdLKyqljiHW8Dy7ngtmVyvhoiL8D6lHOMZaJukqSckHL8ElX1S2IibeiksmvUX4myfXj6NVyhlC0/SkN6W5/RuPvqfT7jbb3hKzKYCAiqhheHjgSu74bb8MV0T8SMBWoQPebfZZNmjUKJeHv8RHe2Zc9sUYd/sqMmWM7sg7m9pItp3y7fmTZdcVSVVRNYpozTni2OUN2i8Wkj0qk1xQxGMMVHSMhCB3Eqk1Lr7M0vAwxGveDghcw7QAIENq7GEAzcHxRN4xA7uvQnwX6xBDqm6rGWlM4VTEBo6qqHj5lJ4XLyclcgJ/T+KuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSLxsAvDc1eDHrhOiUw3762+sDhwPJtkCK+kOdenP1NYvC/6Akex4GGMsRcaZ+A7Ms/a5k9LoCSJAGhlQm2Tk94ZQiFhm5PpcuevCkWcx1kIlD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDEiBKXmipad56CKPxjjRCIc6g1O9nq0TwtG8pNIvZFmu50EEIsZyOyMwXOrNR3vS/ZeYrvFxsVeM9k0NUDgqIYguI9jDNOGNRynkdVxrpQSPuaBI0PEgyg5ljO7IO5vaSLad8u35k2XXFUlVUTWKaM78yIR2yBElvFEfqD7hhw/MKAkXFLbbX0Uvi/fz6yey924HYashhbukWP9HXts+1cKR/omFzdqeWpDyDejpRdbHbVHsQQE1htJXnWNF/r/F9mWM7sg7m9pItp3y7fmTZdcVSVVRNYpozHSIcacghCjhy68JNIwXdMgvVMR6t5LImagpUwam8thzHCIf4DkOo1eCajVB9GseUKCplXICzSMXRQc8yL2buhAunTJOC3k0uu9zhK/3OZSE+3wUp4AHlaZpBVhazntdDFXX9LD/Bi68/ryOAX0ooXZmR0kHlni5swxUdIyEIHcSqTUuvszS8DMW9si9Dm7obAAgQ2rsYQDNwfFE3jEDu69CfBfrEEOqbZVEdPVLE+FNn/QYuNLPkKSlRennIJyfmdIMKBdj+g1C7ZNdaujmE8tyb491uwysZ79S84+xtvvm4ugDXg6fOP13lLvMeWhFtpw4U83KVte6w5b3DwFQVuWtLVNc5sYlOMW1BDnS8vOFCFrkZy+1OvMvJyVyAn9P4q4j0S+aVfp5Lek8xFmzmIlJTuU3JkJFIPXaWy+/uEFi0SlBB0iY8I6wOHA8m2QIr6Q516c/U1i8zlnNsGy/dmSxFxpn4Dsyz9rmT0ugJIkAaGVCbZOT3hrvJEchibIzb0h6FQ/som+ajwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+wTNAErLQx12YJj7cJSeNuawxUdIyEIHcSqTUuvszS8DBW+8rKv1iNxAAgQ2rsYQDNwfFE3jEDu69CfBfrEEOqbARO2FI0qUBwvuopUtWZLuyd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+DB2TZHWspj3eDL6dNoD/r0vi/fz6yey924HYashhbul6tvGsUUp/A6R/omFzdqeWpDyDejpRdbGythJproXjvJWGqyKWUCdSP5yt0sHrkJwpUXp5yCcn5nSDCgXY/oNQu2TXWro5hPLjIdMxbSJaruDhEHI21dy0/7jVhqh8NgZ+b0ESL3prLxxuLSKOWBKb/Teo4jMnl3Ty/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOOr9b8OdjuH+rdgUVHazgAVASjzdxlBBYHYu2cbBVC27SCXgofxdjQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Ltx5v2R/2i7QW6cR3ugt84yOSikUR84Jm6vt7lh6NPTEyIl9tcDvIrKwQFMBrptmFt2FocRTvBr2+YkbIMZ8A+du/y3mwoDlqvnujeI7UaGwAyrlX0gor6uFtH4CBmEku99O/uKD1+pOawKYBavthoH2q801yQRY6YZnynTrgorqLBsEY5rCh9x+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCxOkt2vc9ZNFnlFEOez9nWfw9MlWEq9WakLp/n2nSKsklM7FV/qoydlVr5987fmvr+erqih1M4/juhK1yHWe8Eecluno/rLjFjJakekrNK1qUt/ZazNBY4ftG1k0bLNkme26DEPZAh35ER/L5RBJnizlDeT6t1fqC+Td+E65KKgBnRom7A6Oco5uY1zDqTNBvADqgENC9mCx0CLpsTroN4suFJk9qIBqt23gjXOEok0Svg4z4i8XZ5/O1vv0WSUjnGKokewPSrr+wFgsHfuuaTC/V+HK7PruUXsDzbt9n/3hkUF8SM2bHqoV0obUMXT9Anih+5YDBrMY8nr+ei788bEm5qj0sPQYIBI26MsU3OoLJm8IIaIppzrAWCwd+65pMCR64g5RIKvAmo59SWkrRX6BVQJc9viB46HSBYNLJWQtMCeBBE3ASyzziCaTcQUoHHqOk6a1qF+lFCNaiJ5DIyxW18zeCoGwTCScuw28rHqINrBKvbSWGziDk0+X1bOhZpOy+UhRy3RuvCbxyBk0EuXET/gv9cMW9aU36m9F1OXaA0RlPktigXsbXdvOLveqRW3kfBhmCLGRYbo5NtfjTJPGPbG4bYuGlpvRR6m0pbhSa61hnB7UJsyQt1DnHGtR+23gjXOEok0Svg4z4i8XZ5+IJ+VFi0eGOpoguXkotD1GwFgsHfuuaTC/V+HK7PruUXsDzbt9n/3hr4NXqWw7OA8V0obUMXT9AiaCF2hswYBm1thYfaJ+QITI24DrHhlRZk3Ptiefzb1PqZBGwJbSU11zUTVDaWp20aAjxHiaRbJUwFgsHfuuaTBcDU+ErvoJgL90/v0Oz005BI3JdyDdQVEWGf70wpKlyoYzsSsNWFJ0G6h96qoENi14sER4MYVG7l5ujH7GFmkHKVP553NK9K4etuq7YO628EpiKOY/MgiRiVm6dTdBLoo8c55Lao1U+sqHDbbW3ItCjMPfC77s2Y+Bt3l6y4zarcj8E2OMD64IdjhLaH2iFg7bzi48hZGtVVdHdts/DWOPdhs274WvQTKG71p5NFW87EVevCI8GMK8buknetUlFrQ4woDUElXZkxPpa4LRXNXKKI1sG+05K7PwSyN8YfBDhRuk0ZDeP3PXwFgsHfuuaTCr73Isr9tVv22Igx0sCDms59c/arLlPPSmBk8KJd+1Tk3Ptiefzb1PqZBGwJbSU13ETDykGosMFlzon9+dkVuOV0d22z8NY49cDU+ErvoJgL90/v0Oz005Ac5k/CLrjLYWGf70wpKlyvt1AkOvzrPaG6h96qoENi14sER4MYVG7mHTdqcStfnQnPvrzUAkMW1LBoCyTaf/g0piKOY/MgiRiVm6dTdBLoog2jOC4V9ficqHDbbW3ItCjMPfC77s2Y+Bt3l6y4zarcj8E2OMD64I4m/RGRXCtaZafD/+ALxcOgQTfNBnHK/9dhs274WvQTKG71p5NFW87OhMeW5tgSm2+gJIZi8d40c4woDUElXZkxPpa4LRXNXK6wVaUP9dt9ApU/nnc0r0rqPBMYH68KDQKWG/7xJRim6r73Isr9tVv22Igx0sCDmswn6sV8B+j7zCX3TpPARXBQwr236jwPR1xkgkULL5AvswJ4EETcBLLPOIJpNxBSgcTAlx2aeLfB8krfxm4sTn+8BYLB37rmkwwFgsHfuuaTA2sEq9tJYbOIOTT5fVs6FmPi2JqhGkBE/NttVaLPBczsRP+C/1wxb1pTfqb0XU5dpwdEvRp/kjAajekj7PLyzl8qtBmK7Vxhdhujk21+NMk8Y9sbhti4aWd4C/rFdtJPeNbMoYuP62oJCy0+ORsx9DbeCNc4SiTRK+DjPiLxdnn10t3pJwKv8bbesCLgYotUMsgmFctB+RL79X4crs+u5RewPNu32f/eFWvCc3tR+FwRXShtQxdP0CeKH7lgMGsxjyev56LvzxsSbmqPSw9BggOnQHfseN1W1yX0LWnL5dmMBYLB37rmkwJHriDlEgq8Cajn1JaStFfp20c1L0keWjodIFg0slZC0wJ4EETcBLLPOIJpNxBSgcRxBMyE748g6e/noWG6oc5gu8FWz+jCVowFgsHfuuaTA2sEq9tJYbOIOTT5fVs6FmuurTE2YqxrlXq23rZrzOw8RP+C/1wxb1pTfqb0XU5dpwdEvRp/kjAVRUYYV/VM7FOZdUF8riElm6a1gZMsAzDMY9sbhti4aWd4C/rFdtJPcDWyxE7GeNVZCy0+ORsx9DbeCNc4SiTRK+DjPiLxdnn10t3pJwKv8bauayXcdn5O5Zb/h0F1jGIqPvn/94l6eXewPNu32f/eH+xdMIF2IPahXShtQxdP0CFVx6xUxL6WLyev56LvzxsSbmqPSw9BggqN6SPs8vLOUh1Yef+0iajacB+idEPRV+JHriDlEgq8Cajn1JaStFfud6Ol02C4gTodIFg0slZC3BjnWyfSULU3NRNUNpanbR7nH6SILg7/AbqH3qqgQ2LXiwRHgxhUbuXR0jtwLGTLDOldSBr0GXkcBYLB37rmkwSmIo5j8yCJGJWbp1N0Euis3DenaJbTEkyocNttbci0KMw98LvuzZj4G3eXrLjNqtyPwTY4wPrgjRoNlryl3GkKD6vHWL1wQ48E0Y7HTDO+V2Gzbvha9BMobvWnk0Vbzsre40+b/MNUJu6Sd61SUWtDjCgNQSVdmTE+lrgtFc1crrBVpQ/1230PjigiH2ZjOYj+fVYC3WCMLAWCwd+65pMKvvciyv21W/bYiDHSwIOayTOmi3OtgZdmbQFTYqvlIwTc+2J5/NvU+pkEbAltJTXdWYYYKPNgs1PHs+R7GWvOt48J/v6skEC1wNT4Su+gmAv3T+/Q7PTTlX2D6IDAZ5GRYZ/vTCkqXK+3UCQ6/Os9obqH3qqgQ2LXiwRHgxhUbuFtoNCfe/cTeB4H05I6QIyMBYLB37rmkwSmIo5j8yCJGJWbp1N0EuispIxYYsbAUCag9o9V03daeMw98LvuzZj4G3eXrLjNqtyPwTY4wPrggisSVjG7T/iuIOlwCGjPIYFro93WK9Tpd2Gzbvha9BMobvWnk0VbzsIOplzsorDExu6Sd61SUWtDjCgNQSVdmTE+lrgtFc1crrBVpQ/1230ClT+edzSvSuo8ExgfrwoNCJ709CpHQmiavvciyv21W/bYiDHSwIOazlXVDp/7cALaYGTwol37VOTc+2J5/NvU+pkEbAltJTXcjsdcB259qXEjboyxTc6guruDnuKlgiyT2cC5KCVzZov3T+/Q7PTTn6mnAfDr9bvBYZ/vTCkqXKJqQPqEz95bTnmVBbH6uVADClbnwZjKbkTc+2J5/NvU+pkEbAltJTXQtPcHO+HqhmcGFqrX5nWBDAWCwd+65pMFwNT4Su+gmAv3T+/Q7PTTkd1sSG19NTFBYZ/vTCkqXKhjOxKw1YUnQbqH3qqgQ2Le4a4KqgcHCj1Kh2dBfoHzMxjHhxXS1Mv8BYLB37rmkwSmIo5j8yCJGJWbp1N0Euiqw+nOOnWLAsag9o9V03daeMw98LvuzZj4G3eXrLjNqtHACTjqvTZI04Fz2wTKAvWg3EgB4kcemWwFgsHfuuaTB2Gzbvha9BMobvWnk0VbzsXrC/Y8nYV376AkhmLx3jRzjCgNQSVdmTE+lrgtFc1cqiOECh5qCMSetGkCxH12jdbdBtjhEDk97AWCwd+65pMKvvciyv21W/bYiDHSwIOawyevBJuJtTUqYGTwol37VOTc+2J5/NvU+pkEbAltJTXeaTcqpZECinJkNifELz+tUYxlHvSQBSZlwNT4Su+gmAv3T+/Q7PTTmhCf5T1PzJ8xYZ/vTCkqXK+3UCQ6/Os9obqH3qqgQ2Le4a4KqgcHCjOSEwuPGpNfUN5n1uYM0mfeQY4ctLCg/WSmIo5j8yCJGJWbp1N0EuisNn4muq/50vag9o9V03daeMw98LvuzZj4G3eXrLjNqtHACTjqvTZI04Fz2wTKAvWnzIl9piDpgtwFgsHfuuaTB2Gzbvha9BMobvWnk0VbzseJI3sQqZe9T6AkhmLx3jRzjCgNQSVdmTE+lrgtFc1cqiOECh5qCMSetGkCxH12jdZDEoYbsCdwzAWCwd+65pMKvvciyv21W/bYiDHSwIOayGNPdbLt/UTqYGTwol37VOTc+2J5/NvU+pkEbAltJTXeaTcqpZECinJkNifELz+tWOhG3mMm0lvVwNT4Su+gmAv3T+/Q7PTTnx5bynw5fwNRYZ/vTCkqXK+3UCQ6/Os9obqH3qqgQ2Le4a4KqgcHCjOSEwuPGpNfWRNVL3GDOwV+QY4ctLCg/WSmIo5j8yCJGJWbp1N0Euik7wuCbKyq7tag9o9V03dadyukvJ0+dhsAa7uYpL5T0mbmNcw6kzQbwA6oBDQvZgsdAi6bE66DeL3z1d3inx7vwqVmtebrbNeVA+qUgeAqkYBf3g5Th79ziZtOaV3rbA45OWF8KnLZwBUD6pSB4CqRhREutXY27C0H0UQNyGAT5px9QUA4n2k7Q/m4zwAVWJRxFguxXMgMsXYsacUWhCF6CjlvYZ+HpI7pnPGMX0SF8DnI+PlatupIlYnxsFlxAQE/iiwGl157iWfPyipdPqDuabhlmvWfHeKcBYLB37rmkwqhwPFfueNRUQxkdRtXHGGHOxgWow/G6LkvlBHiy3LejVy0TFImojNkbPQKB5piy2G+MOqean6icdt59ZyKqN42WsdLKWHhR9G13bzi73qkVzCnp+ua6ixkmgX40HHjm4bKDOXxvAme2WhJoEOKDjb0odg7Lws3CNS+NUGOoRoh/JeV/VJ1seV+WKUQGTYMurDCvbfqPA9HW2Wc5osDyA81aL8oOAfFS548GcdeSei/nO0Sga0ocbDwwdk2R1rKY9YrLI1Ow0ElbWmH0QnDKBioTGSR7/wOaPupmkdEVpLFvqHHI1yiAGK82Su4OGpqX+9EV/ZVHeofgVcmAJ52QFaOZqm+7wZO0V4m/RGRXCtabiN7L9OTBPDZm05pXetsDjINI/05OX1ov50STVWBusOeEyOT6Jg5gwBb40+j9JBClzT2WEQwLY8QmtcTed3vOWBzF0cu6U6b2tc9O5lUpeTPjigiH2ZjOYXAUL4wWgKHLjwZx15J6L+c7RKBrShxsPdjhLaH2iFg7bzi48hZGtVVCtKGqLmpTaWPCrRU0PtFqsJxgRh210YKjlKiOs0gRlDCvbfqPA9HU6dAd+x43VbeTWdIsLxu3YmbTmld62wONkiyOTbSu4w/BLI3xh8EOFVoncAGm6YKpmFfPECuAdoI2TQqhOpUDhHLvdloCY0mxB2HI455bXqRbaDQn3v3E3VhbouAeKK6/jwZx15J6L+c7RKBrShxsPCmSzK+vxonL0CZHEz0EvamHW9k/xEsA/HB9mT1rH5CwcRy4n5G9LBgNM9J4T6Hm6YLkXeRIMPlVUVGGFf1TOxarkM8V49Rbn1lrf3MAW+LDT7hLSAvyDIMCTsqSLk1SmXslGlDKq0rb25cUiCOkQlcfUFAOJ9pO0Om5cZBqGn8kRYLsVzIDLF9RipjlsWqciMlkMGSopX0EB0rdEwIGjwTToHlm2V76QcLGGvjlbJ3XWmH0QnDKBioTGSR7/wOaPAYCZgsLQ7uZjrlimj3MII23gjXOEok0SZ8uMTcoUeKzZ0wVTcQ9wy18S7ejBSGb4HgAv45hvKaOajn1JaStFfvicPyAERY7grXPTuZVKXkwpU/nnc0r0rrltu64zkjsb1lrf3MAW+LDT7hLSAvyDIKjekj7PLyzlIdWHn/tImo1iMk/Dg6PNKWgZM1la6Pu4LT3FN64V7B4RYLsVzIDLF3K6S8nT52Gww8WetHSTquemrIyMmM53oIKmHB1ENW07Bf3g5Th79ziZtOaV3rbA48UCWtKJ2eUIVG1UeuuDwd9h1vZP8RLAP5vBSCgTR+xFWIIAIds2MSoSmq9rOD/u8uaTcqpZECinB7ccNGtUQ0ozbXroVfCi1jN2f/DBhJMLtGwLZityvxMDj+ey6aTLrcfUFAOJ9pO01CdIBMgddrpYggAh2zYxKjB5A2Omnc40KOVxHZHvWGwqFiXCW9rvVwXzyuO1cQKjSh2DsvCzcI1L41QY6hGiH7oR2TMvCqiEq80xvBvfgqtG8h0UlviqMDD5G33ufRzxWsxs9IP0pnAwyhm+u5mfsdcB9u/qWYJQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LuByd/PverQFaqS53zBtL8hnLXdIfXO1vNpQQWf5HvYU+eoa6rFNJu/QSH2YZFW3xFeE6ZypoaFfbWmxzHlS9XPhY+xAPB4d3kggVfaYiee0Hir08408efyDyVW5fvLJZWeKdmTkEiU0K2xFvcFFIVwDKuVfSCivq03NQQFCgtDwfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctPT/IbYgO2uVnwg/IMu6/6X3GFc3FY3ZPv+ggUqaEPvXOGXMNJvXM3NonL3dWzRS56qn3s1umWY9BCSCKyXy1gWv4xlzFUdpfSZQ1rylVvtG1k0bLNkmZ5RRDns/Z1n8DwKRTyX3NLC/Akftdwe10azJJLiCUOBtfJjinfBJCHC/Akftdwe1xEfy+UQSZ4sI2z39yYmxkvvCv6L7me0zRSDh87mOL7fWO0HZMQy281p35Zthlj87WgxwPOa+bCZuX3CwhwA79owICxouRz2wyCL0/lDTkTEO95IiZfXcDT5dLolfq/xY8EfppvqcUz6AavDmDTROJFI+ewdy3Rna4aELzFZeL6+QHV5xeL4xickIDeNs7bqVjAgLGi5HPbDIIvT+UNORMQ9sRnqdohw/rInvCB4XJTTAWDQJ3KBpIOfoAOLnMoIH62LiTlmATyVMCAsaLkc9sMCLmfIM/UTQFRbFgavAZiva9CKQlY8TsIdg1suZ9E6/+FUC5JyaHrvXgkDBylGzbDVmaIohTeKh69QIF4Myn71WIIAIds2MSqzpuBjY2VybUj2QowWZ18NQhQaHWyXaE8BYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3hxTocKi3omLwhpxmZtCvVSVaX9ZvoJe6cvhqXJzaLMaODCIWhhTCDVYjbDmrSNx7SWYCYVHcspp5nRpRErudjt6lr9eQQZ3jNxxHLifkb0sGc8rFJQKPIgNF1pLizt+ffhS2UoimbAzEsmIfj2FrPeDMxV44XkACLfWCKtFaAB0pbUXfYiX6zhRNZOg+17IrEdNERnB9b9x1ZgJhUdyymnmdGlESu52O3qWv15BBneM3HEcuJ+RvSwZzysUlAo8iA+1GgG/AnejDBH5d5Nb5sfkd2Ig3SMjFLVe6bBKRjbs1DtMs5EUaUZBYggAh2zYxKrOm4GNjZXJtnGqV60+sEsT44oIh9mYzmMYIuX+MRwG2Uc8EGIRRT08PJo5BvLOJdliCACHbNjEqs6bgY2Nlcm2capXrT6wSxNA83omXDZzLn7Mk+3l1IY0zFssQVwf33y+QHRyogQoLHEcuJ+RvSwZzysUlAo8iAx2uj9gT5waOTQbM7YMtlDbiDpcAhozyGO3YYSLvZJDyTCZg+YTqmpoPdW2XyIVH/FRWHJYQ/HeHfroUhiOicc46Tj/7B21oNlrRF5rgcU0J20plasIhJg4wICxouRz2wwIuZ8gz9RNAlZnKzUlpyj5r0IpCVjxOwh2DWy5n0Tr/5pNyqlkQKKfhwEYlgJb7LBs068yiHao0nrgr/BC+fs5OQZIm7+zr2MLg4TLFSlMPqXdN+qr32gM5ITC48ak19fTKRbYVvBXtEFxjJGuPLY+LSRYue6xyQjgddvbdX6MFbUXfYiX6zhRNZOg+17IrETgXPbBMoC9a6972h+nDsDcGCB+gdLSrKRFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybSXbC0NoZwHP60aQLEfXaN3oPGdfu84ZIispC8S1AlPq+oTU3PJ5KN9r0IpCVjxOwjbhfUs2/G3P+eN/hBVIbTMnDRel4faEa3CAjfd7xQL2dWTJ1KHwjnrCHTnGJiwHXcTZrR9MdAnrJFFahibdzyJxztYHphKvOAIuZ8gz9RNAlZnKzUlpyj5r0IpCVjxOwjpKB/H5OuK2wSRpLZa1rDsYpvJFpyu2Qkzv77OQ7L2nlNYBnFeoylz4AIVNIXWRQ2vQikJWPE7COkoH8fk64rbBJGktlrWsOwpksyvr8aJyrrNgBgSLhZq6fle4Myn11YNHAzIEMAyd7GNtU97kTE1HZ9WYTKq9U4jwWvntcuJiqN6SPs8vLOUh1Yef+0iajY5FsGDdYBkE4XWtGD/Rq6kPJo5BvLOJdliCACHbNjEqs6bgY2Nlcm2VrUDlzL3COQGAQX2IpawmpKFk2NHyLDnmwLkSqPVwnqKvaI5Zmr6glM7FV/qoydkji9MrIcEZzw91bZfIhUf8VFYclhD8d4cGPUiUezMBVPj2we/Xwe+zhByivyDfY+EqEHNKcJDhm5OIIHKIWQir9KM91k9syYvH8YPSoAnQYMLg4TLFSlMPsUJYN6b3gXvzkgYjmawpSilT+edzSvSuo8ExgfrwoNCUUggCRWdzyiBkf8+t9vrD1ZmiKIU3iocEUr80Y7LPoOxjbVPe5ExNR2fVmEyqvVOI8Fr57XLiYm5jMyU+AnNu/nLahDZxASjnhJ6iW2E7I3HO1gemEq84Ai5nyDP1E0CVmcrNSWnKPmvQikJWPE7COkoH8fk64rbBJGktlrWsOxojBQdksktf4hRkqU2sgD6MxXhNV2oUijGTzC+tFdi17GNtU97kTE1HZ9WYTKq9U4jwWvntcuJitlnOaLA8gPOin7d3Husz3h1ULW2AWLCOdWCm8N7aUUocRy4n5G9LBnPKxSUCjyID0TtSsmzc9o4j7LFPblToDhvp9bPkM0RglM7FV/qoydkji9MrIcEZz+bV9EPoBEz3VFYclhD8d4cGPUiUezMBVEqRU4/TOBeKB8coSla1YDeQi5O8bQYGf0ngnZslNY0/D7DkI+4jM/Jr0IpCVjxOwjpKB/H5OuK2oXYiUSQFwZ04Fz2wTKAvWmnCcfykCW93HVQtbYBYsI71zdBAlwTmSxxHLifkb0sGc8rFJQKPIgPRO1KybNz2jioWJcJb2u9XYZBOU6kKvlSir2iOWZq+oJTOxVf6qMnZwWFEse2vnPbrOASvJyBn0DkhMLjxqTX1RtYkc/Cdu6pe8gHhuo5/I1TM/LO5RPzdKL4bTgl9GUBUVhyWEPx3hwY9SJR7MwFUSpFTj9M4F4qU55gx+/r5Euy+CFWbAgfCSeCdmyU1jT/6hNTc8nko32vQikJWPE7COkoH8fk64rahdiJRJAXBnTgXPbBMoC9ac8CebNyyCTpipQ3jNDYXS9DMZffV+OpzxF5kW0MLn8kUg4fO5ji+34vGqARtAaJC5I4IXBo4g2Eo36jxjcHPCwmjeAwihDl36UBzba09Q7BhEABmpbOO19fXI7Nh9lUtNrBKvbSWGzj85jILoHNoPqZI+Qiu6A4wiU5qh9cbfcRQkaz+Fo8ShJxqJIHSnBRTgp7dEfopuCc8Hfe4JT2CyZ0aURK7nY7epa/XkEGd4zccRy4n5G9LBoVVIPUUpxe0EwXPrxhxdLM0YRGHlQeoH6VqodDodiFl50r/6zZg8QkLhoIxd52G3lMzMTd2VbLAK+TC2YUt5PYwsdeXQDWrkJTOxVf6qMnZnRPJTL8CXovu0V+ntFmUQSSJw00xaEzAZd/yTly2zIKhjc+n+qcPo50aURK7nY7euEyNknZEVqhYggAh2zYxKvJMoiRRwIwd7tFfp7RZlEFEYxRziOLSXPiY6kXZLM45a7ik3ABrJWmDRwMyBDAMnexjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3cRMPKQaiwwWXOif352RW45ruKTcAGslaYNHAzIEMAyd7GNtU97kTE2caiSB0pwUU8nghxtgSf/dyOx1wHbn2pcSNujLFNzqC5YlHfB/zqZzDWSX1+HDlqSDRwMyBDAMnexjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3cjsdcB259qXEjboyxTc6guruDnuKlgiyQ1kl9fhw5akg0cDMgQwDJ3sY21T3uRMTZxqJIHSnBRTyeCHG2BJ/93IAIyXWxsyLm8Oxz8TxEyn46FnwlZdCSgxk8wvrRXYtexjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3cgAjJdbGzIuWJ7/LE7Dk+ghc9PbYqAbFhFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHe7RX6e0WZRBT8Tm6By0j+SFooqTaar4ls3NonL3dWzRF/O8s64DUvIcRy4n5G9LBli+KRiVnTXVnAnqRY0tzpmXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZt7lATO+fQUOvnb+3Ba03evx8+ho+XTVupzN/l4anUH+OiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHKx1f1+XtgrToR+KHV4rtaleh7vTtA6Y2z8UnERL5ba7Bw2TEYBX3tTqxiEouaRpssvFfG+fBhu2ssCk5CiXq3flyJNSZWXY3L5W+rEb8XoruEkpZ1EwtkIzMkqBzwJG4Pg2YerELivI7XwTXmaZPyNsHkkgh1IqBUlX26L3zEegzDCDFQmIOwZqDXxlkXGyt9HnrOJuwmGUi8HZEGoTxCDV0yH7pXjXLcvZwDlzKIgxEeskJCHxHLFZDpqtZrfo5tourMmZ+Ww9Je3XicDJZZfQ1pFmvl22ruVzBspFARCWZacAGSF9jAb2K6hMdSPTRwoqTFCFnhtH8JtgoS4weo0CEXZx67/VYaqw6hbRq2ZocvdpbV7OJGSqDXxlkXGyt+k/f5AuYfucgQYimGjnqelqo+/6VQ2n/aD6pd7T4wICCDkaXfatq4nqDXxlkXGyt/0l4nob285ilY+I3KRG/XjPWKN83VYbStVW3DiKRkzwlqGBdlZwtkjgMpAlEzTVMPQnS2lYR1pzhUjqW31aQvzrTIP0x/AMDCbsKX8kabh1EzM6jWgHkBNGflyiQPJklWh4ZO8WllMNTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyMj1EomkBOXDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8QGOw6IbIHiyvDwW3zPXFw8TMRllKl4+FmzaUnbp7B7W8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTsrNWYQz+pTD9x/2wXHAq7Hoe707QOmNs/FJxES+W2uwcNkxGAV97U6sYhKLmkabLLxXxvnwYbtrLApOQol6t35ciTUmVl2Ny+VvqxG/F6K7hJKWdRMLZCCH7L/kpD1/cJw9YlomiUp8JXZAhY8A6K/Hq5bfbk4rSbPz/c6/JJ/2iPRAJAhOGHhJao7CnWxLZRGMUc4ji0lz4mOpF2SzOOfaqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+qDXxlkXGyt/BJGktlrWsOwpksyvr8aJyiOBKVzxmGVUlX26L3zEeg4h4BdF8CI0lZL+814w1rJaskPxLL+8gfSH7L/kpD1/cyOx1wHbn2pcSNujLFNzqC5YlHfB/zqZz9qoHINnqNTTDk8jS4HDXZECGgMvrUkxxqvxPemSJzH6oNfGWRcbK35WtQOXMvcI5AYBBfYilrCakoWTY0fIsOebAuRKo9XCePj7SyAJdO89s/P9zr8kn/aI9EAkCE4YeElqjsKdbEtn49sHv18Hvs4Qcor8g32PhKhBzSnCQ4Zt+85HZecWuVWz8/3OvySf9JV9ui98xHoMJmtXG2aPKGZDRDzKAm9d67OW8m3j208NdLd6ScCr/G2rmsl3HZ+Tu+jci+PTO5rqECi/rk7guZlEJZt5I6hoN5iRnMMMFpPtmPJKZ4to+ysEkaS2Wtaw7ftncQJK48aeBg57WamN5zOyvfg8iGk0+QIaAy+tSTHE37Nk97b+6rlVbcOIpGTPCm6GX1On6ntn3U4yioDBJC7EVN8+GDJBiyLNO9bmKzQ1mlj87A5FHjBpjN+NMLr6Rs6bgY2Nlcm0EWaoAMA0T8qjkWIc3LYL+xBsWOBf1OjogbaRGBa63erCipxj3is3EUQlm3kjqGg3mJGcwwwWk+5HHobpjcJk1tTDyb12rUNYxMlr698GshCVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3+s4BK8nIGfQOSEwuPGpNfUp/9XvJyDqQ/aqByDZ6jU0E9c1gpRGLR+Fy44jk47FMrFCWDem94F7/aHVmfz3dMLrRpAsR9do3W+QJcG4P9eqJV9ui98xHoMwwgxUJiDsGag18ZZFxsrf6zgErycgZ9A5ITC48ak19Yag663Wr0fXjRBmQQXz8GWoNfGWRcbK3+s4BK8nIGfQOSEwuPGpNfVG1iRz8J27qvaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMrFCWDem94F7/aHVmfz3dMLrRpAsR9do3aqfhyI4IdU/JV9ui98xHoMwwgxUJiDsGag18ZZFxsrf6zgErycgZ9A5ITC48ak19fxaS1aN7wFSjRBmQQXz8GWAbAWZCTK1uA/XOJfyF1XDY3sCEo28Fct8J/VrU9hea2suxKHYfDbF4SSlnUTC2QixQlg3pveBe7aOQZwLKZ7xMA6OixUw6rRBUf+h5bl0QsNwP71HnkU4bPz/c6/JJ/1P+uEQL8hFMHUt0LNTvpDLYOXiu5r1A9YP2rrHdb1eRgY9SJR7MwFU+PbB79fB77OEHKK/IN9j4TK4kLrElPLVDAko/mYmeUUlX26L3zEegzDCDFQmIOwZqDXxlkXGyt+VrUDlzL3COQGAQX2IpawmpKFk2NHyLDliI0tlVN5G8z4+0sgCXTvPbPz/c6/JJ/2iPRAJAhOGHoNWBUbEQksWYcA9PvGn5qi0bAtmK3K/E0lMbGpMLalIL2cA5cyiIMSDVgVGxEJLFmHAPT7xp+aotGwLZityvxN+4gQPL1DzMi9nAOXMoiDEQvZOoeWO9V+RX2BSyKrCs3EK95r9tEWsCjztA2FYcnwqgHrgP0Ys0NjTutw/wzMvRIoLn9egg/AqVmtebrbNeTBOxsWdPiRLwFgsHfuuaTD/WDiFZb3HScj8E2OMD64IauayXcdn5O4BgwWK04qNgEjBpGmAhK5EgvU1+bAGMBrCHTnGJiwHXcTZrR9MdAnrMTJa+vfBrIRgpYxBgkNjhSSJw00xaEzAdDNUb3ycDXtLZd1ieTRwWLgWCEjsdZ8lwFgsHfuuaTD/WDiFZb3HScj8E2OMD64IftncQJK48aeBg57WamN5zAZ0/x117MyJwFgsHfuuaTCxQlg3pveBe7aOQZwLKZ7xMA6OixUw6rRBUf+h5bl0QsNwP71HnkU4bPz/c6/JJ/2SQsgUWCpujcBYLB37rmkw35uVDSA9htMm5qj0sPQYID8BqKRjeRUOcLN2H2dvqf2oNfGWRcbK35HHobpjcJk1xDOnbRINvwN8q3Yc1Z3rs7miAasUKv6TrbQbr0Wc1efUUVSQ6WhdvsgAjJdbGzIubw7HPxPETKfo0u8+V8CORh5lr8oQnHro9LwbQ+k+4H1NPyGslk1x0eUo8iDNXpzHy1/0mkD5lMAYa77f8vmAHRJao7CnWxLZA0RlPktigXvsHJ6m4HEG7LmiAasUKv6TrbQbr0Wc1efUUVSQ6WhdvsgAjJdbGzIuWJ7/LE7Dk+gwscktoq3WFsBYLB37rmkwDCvbfqPA9HUaTV1KG5vCDRhrvt/y+YAdeDspfEuZJsq+DjPiLxdnn3AbcsFcxHrhwJEVuN6gT0FoVOelkqJIZ8BYLB37rmkwqelc3ICaMs86dAd+x43VbSM11Dv7cr6DFu7lHgQvYkzSFpE9iGhjyODXEbg5AnphOnQHfseN1W30LsRL+XZTYxhrvt/y+YAdeDspfEuZJsq+DjPiLxdnnzktmzEVy2n4iJmaDkV14LHte3qWuRx69MBYLB37rmkwBFmqADANE/IW2g0J979xNxHdkgd81/Bh7zexPibMk63QW8ISDeu3BqzkHOTCS30lOS2bMRXLafix91ggRJwKhrOm4GNjZXJtWsvbF38YWeRrZ+Gtr7w0eusFWlD/XbfQ0DzeiZcNnMufsyT7eXUhjV4gg1k7kjBXwFgsHfuuaTAGPUiUezMBVADnBcUjTELbBLo4purMT196IyjIK4Jm/Fd5WV8gU76CcPeNm59NMYEeZa/KEJx66PS8G0PpPuB9U/CeJIgVd11aaAG/u9P6rTwUXoSBXj+QmDHBrdsEygeoNfGWRcbK32Y8kpni2j7KwSRpLZa1rDvib9EZFcK1plp8P/4AvFw6WOShFsK1eb2GS0bEBp88iXpz07QGDrdWwFgsHfuuaTDBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDryH6zaN8puUfAJJPjGQpI8qTTBWlHyLSSB/JGDlqdOXlpoAb+70/qtPBRehIFeP5Do0u8+V8CORh5lr8oQnHro9LwbQ+k+4H1T8J4kiBV3XVpoAb+70/qtPBRehIFeP5Ak96MM5hLRSqg18ZZFxsrfZjySmeLaPsrBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDrg8MxZ7cKwooZLRsQGnzyJenPTtAYOt1bAWCwd+65pMMEkaS2Wtaw74m/RGRXCtaZafD/+ALxcOg0CDPmJpTJ88Akk+MZCkjypNMFaUfItJIH8kYOWp05eWmgBv7vT+q08FF6EgV4/kN+3BFUyRUa0wFgsHfuuaTDNkruDhqal/qHbIOVVkhdDwFgsHfuuaTBF86nqKnwwoXiwRHgxhUbu0PpIV6W3I+AW4UzD/Lz2a0v8MthD2qTcwFgsHfuuaTDBJGktlrWsOxim8kWnK7ZCp6EZaAJxX+WYxYB6PUv8lg4ldsB3gKsrkez6ymeMObwYpvJFpyu2QvBLaZvQ8UKGwFgsHfuuaTBF86nqKnwwoXiwRHgxhUbuFtoNCfe/cTdO/KKaXL7gi2hU56WSokhnwFgsHfuuaTCp6VzcgJoyzy8jKhI7hEwpOvnqAzq55s41e8yFW9QuWcQiqV/8gaQqWoAfbmEZUToW2g0J979xN0YBavpdlFWjkNEPMoCb13qkBz+FUA62mMlS7qLiPpHRcHRL0af5IwFUVGGFf1TOxTmXVBfK4hJZpxMO70QHN//AWCwd+65pMFwX1VcRZhYfhr/7NekDA/okWLnzM+eAUtVumz2A9tWGNkn/94itCst6c9O0Bg63VlrL2xd/GFnka2fhra+8NHrrBVpQ/1230ClT+edzSvSuo8ExgfrwoNBRbOPR3LlP5hhrvt/y+YAdg1YFRsRCSxbMU4UVpv+iFFpoAb+70/qtPBRehIFeP5APAtSrS/jN9A4/6C2GHvfpkNEPMoCb13qC9TX5sAYwGsxThRWm/6IUWmgBv7vT+q08FF6EgV4/kPC0s2De/udNtNd3+Ny1F6z4hMiC1gWTDyDSP9OTl9aLKVP553NK9K5OCSomSQ12P7Om4GNjZXJtWsvbF38YWeRrZ+Gtr7w0eusFWlD/XbfQKVP553NK9K6jwTGB+vCg0EFlPVRfR4xHGGu+3/L5gB2DVgVGxEJLFsxThRWm/6IUWmgBv7vT+q08FF6EgV4/kHgrJanED3+jDj/oLYYe9+mQ0Q8ygJvXeoL1NfmwBjAazFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QyFlmPrTnC+W013f43LUXrPiEyILWBZMPINI/05OX1ospU/nnc0r0rk4JKiZJDXY/QLw4iiueoOLAWCwd+65pMGuiOljGxGW0NFO/NoUYFKbAWCwd+65pMN+blQ0gPYbTJuao9LD0GCA6dAd+x43VbWMlVwJEAHW5SMGkaYCErkSC9TX5sAYwGhmkhUZruG54fpRLPm1xe9x9bM6EFqs+eFM2bu+WFHT1qTTBWlHyLSR3ljnjqNbx+X6USz5tcXvcMIXRUjR+vcXAWCwd+65pMN+blQ0gPYbTJuao9LD0GCAvIyoSO4RMKVZurVyHEK9cS/wy2EPapNzAWCwd+65pMMEkaS2Wtaw7CmSzK+vxonLnXQh1cHIHWRbu5R4EL2JM0haRPYhoY8jg1xG4OQJ6YS8jKhI7hEwpZWPmHBCXX86oNfGWRcbK33mI+vqzK689qZBGwJbSU13mapvu8GTtFb3DQeqZhZgzYFGpEEAiKOFoVOelkqJIZ8BYLB37rmkw7OW8m3j208OjlvYZ+HpI7pnPGMX0SF8DJ6/XdsslDegOP+gthh736ZDRDzKAm9d6pAc/hVAOtpjJUu6i4j6R0fj2we/Xwe+zhByivyDfY+EyuJC6xJTy1YK8JXE08oaRwFgsHfuuaTCxQlg3pveBe/OSBiOZrClKKVP553NK9K6jwTGB+vCg0J64Fa3BVLwhNaQ+/yt3IYuoNfGWRcbK35HHobpjcJk185IGI5msKUopU/nnc0r0rqPBMYH68KDQR4AnUVgr+S01Zicz6VVMhGCljEGCQ2OF+PbB79fB77OEHKK/IN9j4Qwx8+Gz2w+KkNEPMoCb13qkBz+FUA62mMlS7qLiPpHR+PbB79fB77OEHKK/IN9j4SoQc0pwkOGbKGHwLihVpzzAWCwd+65pMLFCWDem94F785IGI5msKUopU/nnc0r0rqPBMYH68KDQio1N7wGOgC81pD7/K3chi6g18ZZFxsrfkcehumNwmTXzkgYjmawpSilT+edzSvSuo8ExgfrwoNBJPQwzh1FLnjVmJzPpVUyEYKWMQYJDY4X49sHv18Hvs4Qcor8g32PhDDHz4bPbD4oCgedoCuA+3USKC5/XoIPw+G3ThEbqJl/LGIGtbraLex5lr8oQnHro9LwbQ+k+4H1U/ra7yV2SsQGDBYrTio2ASMGkaYCErkSC9TX5sAYwGpE5dDsUwpRp5xA0oF7DLRduL6S/eYL/s8UCWtKJ2eUI7whiIHij6dbAWCwd+65pMEXzqeoqfDCh7hrgqqBwcKM5ITC48ak19Sn/1e8nIOpDaFTnpZKiSGfAWCwd+65pMNE7UrJs3PaOKhYlwlva71cKN/W0WpqKonsigqtHOVe20FvCEg3rtwZX4BnoZQRiYyoWJcJb2u9Xw2QSW9a2guuzpuBjY2VybVrL2xd/GFnka2fhra+8NHqiOECh5qCMSetGkCxH12jd0s6pjFM+9QoYa77f8vmAHYNWBUbEQksWYcA9PvGn5qi0bAtmK3K/E2mLuqmjv3qpUzZu75YUdPWpNMFaUfItJPc71RtLmF6ItGwLZityvxOfCJxtsOnNSMBYLB37rmkwsUJYN6b3gXv9odWZ/Pd0wutGkCxH12jd1MI3MmnKoMjRtVyF7/T9TcBYLB37rmkw/1g4hWW9x0kcAJOOq9NkjTgXPbBMoC9aUgW2JZuK+B1IwaRpgISuRDr85uOqE8NxFb919yWa4zlvjD41JgHDTlCzlMQPh9nvFu7lHgQvYkzSFpE9iGhjyFwM2C47wN8ib4w+NSYBw04v2SAfuBCHvqg18ZZFxsrfeYj6+rMrrz2pkEbAltJTXeaTcqpZECin1QUVKwOqtDjS1jvHBWk/j8BYLB37rmkwBj1IlHszAVRKkVOP0zgXipTnmDH7+vkSHq2CWF0RLWhUzPyzuUT83WCljEGCQ2OFSpFTj9M4F4rRXhPHkUggalRyCw+1qvISwFgsHfuuaTBcF9VXEWYWH+aTcqpZECin1QUVKwOqtDgcp4hvhbTsNuIv8vZq+ewAwFgsHfuuaTDnh+dvDcAIMg8eoX8wDqdowFgsHfuuaTClgpZlbNijNpDRDzKAm9d678dX2DDyHREIQ8qf4uyP172rBUoGQrMw43YVY774KSFhZozdt25vcDNSC50CghXz5oyoIXeJbFvGgQMzhW4dwqvRAO/RtUdE8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3Z/sInISWfk6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZWeKdmTkEiU0TMczVmxwA6NHGil1XtixJOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHLBSay3l6556Ko6S20Gke3I5oyoIXeJbFuwNu9pJr5KepciTUmVl2NyLaph3YSB0q0NBQUlLIPgxU2EM6jlg+dX8wvcQ79a/M2OHAgZShzLsag18ZZFxsrfSPZCjBZnXw32qgcg2eo1NBPXNYKURi0fhcuOI5OOxTL3Gi8nabEDNEu+dfYO6F+PdRYolDpH0bOmt+QzqmdAq78RQpZeJabnqDXxlkXGyt9I9kKMFmdfDfaqByDZ6jU0E9c1gpRGLR8Pkewz8hTS5eQnfxo58a0PwNSgROhYtQu+6dBkYMzRxIm81zCsbjdDJGt93FLnFxYRO5zafLLM3OYiqiWWtCZqnLeundAyWWpvbEeOIXIN/Bhrvt/y+YAdUGGnNXOa/EjR768ZeCgbj6g18ZZFxsrfeYj6+rMrrz2pkEbAltJTXScPWJaJolKf3xP5p7A5hlmoNfGWRcbK32Y8kpni2j7K3OXkGArzLsPlwA+e7vpE+EQZs2Apd9RcuHkcmlnxQWBay9sXfxhZ5Gtn4a2vvDR6V68Rit0cPmJQPqlIHgKpGCr/TOL9TExIGGu+3/L5gB2DVgVGxEJLFqmXs2T5MYpVJw9YlomiUp9NOMIRwaIAjsWz+BjCIGE8KfOysdJt4XYAQnJ+BiGA7qKg6ef+jn55GCAa+dPV1zrAWCwd+65pMP9YOIVlvcdJyPwTY4wPrggaIwUHZLJLX8tf9JpA+ZTAGGu+3/L5gB2DVgVGxEJLFqmXs2T5MYpVyACMl1sbMi5vDsc/E8RMpwQR3LGsnLGJnRpRErudjt6QmayYsXTbfsQzp20SDb8DfKt2HNWd67O4FghI7HWfJcBYLB37rmkw/1g4hWW9x0nI/BNjjA+uCAwdk2R1rKY9cLN2H2dvqf2oNfGWRcbK32Y8kpni2j7KNmcKzFr+wOcDRGU+S2KBe+wcnqbgcQbsCrFEFU3DiuABYNAncoGkg5LFaicXcUrcwSRpLZa1rDsMHZNkdaymPY1SkNEqcpXgpmFERzayw5ORjGUlDW9J9HNRNUNpanbRkldJvla2lA9ay9sXfxhZ5Gtn4a2vvDR6BkU4JP+T11NgZED5XUW0vEv8MthD2qTcwFgsHfuuaTBI9kKMFmdfDfbKzPqjkHxfXR0jtwLGTLBM5A0VtvblosBYLB37rmkw35uVDSA9htMm5qj0sPQYIHIo+HkVcgLphByivyDfY+G6kKM6rsi69MBYLB37rmkwf0h/5H1vCpqs5Bzkwkt9JSEpC2QWlVtqWmgBv7vT+q0VYbUk+RlGQZTOxVf6qMnZI4vTKyHBGc9lJyf/SnjGFgR+XeTW+bH594APv36K8aa8cmJ2aAfglMBYLB37rmkw/1g4hWW9x0nI/BNjjA+uCHY4S2h9ohYO284uPIWRrVVeIINZO5IwV8BYLB37rmkwjZpRn0I8htZagB9uYRlROsLX98K6mygUD1qrowGFRhSC2sD5UBmwkAFg0CdygaSDksVqJxdxStycapXrT6wSxPjigiH2ZjOY2AtciUXIvXno0u8+V8CORh5lr8oQnHro9LwbQ+k+4H1MCXHZp4t8H36USz5tcXvctYyihw9reCUYa77f8vmAHYNWBUbEQksWqZezZPkxilXVmGGCjzYLNT0dWT5AhveRq0SLj91Ue6/VmaIohTeKh5AYdVtwThZhRGMUc4ji0lz4mOpF2SzOOXBaXHiGb44EwFgsHfuuaTDfm5UNID2G0ybmqPSw9BggLyMqEjuETCn0U+K7XkRY2kv8MthD2qTcwFgsHfuuaTBI9kKMFmdfDVWet8z1OQe6nv56FhuqHOYJCD6wYHv5F5TOxVf6qMnZI4vTKyHBGc/N4uOh+kDjVi8jKhI7hEwpDFKleI9a/u+zpuBjY2VybVrL2xd/GFnka2fhra+8NHrrBVpQ/1230NA83omXDZzLn7Mk+3l1IY1eIINZO5IwV8BYLB37rmkwjZpRn0I8htZagB9uYRlROmHTdqcStfnQnPvrzUAkMW1Qqfyq2ro4rqw9aDoVJ6fI6m3ZnKEGKjyQoEY4ar1b3iKxJWMbtP+K4g6XAIaM8hhvwPIlwyQltBhrvt/y+YAdg1YFRsRCSxapl7Nk+TGKVU57CX+OERAHVFRhhX9UzsUyfGSk/TQONqtEi4/dVHuv1ZmiKIU3iofj/vgimiURQGvu6TVpIgPAvcNB6pmFmDMAPSxBKWuLGejS7z5XwI5GwFgsHfuuaTDYMn+n/hOve2Wzkn8IqOfIuDWFmQt6wgskvkXL9ippztFFzBXMa00M9NP60c0SRhBGeTtGwlIiuddQDEsqvwiLJxNx0Um4IV8Ya77f8vmAHXg7KXxLmSbKvg4z4i8XZ59dLd6ScCr/G2rmsl3HZ+TuWW/4dBdYxiLte3qWuRx69MBYLB37rmkwe9nMsBBqXJzg1xG4OQJ6Yajekj7PLyzlIdWHn/tImo3OYUoQsWQUygFg0CdygaSDksVqJxdxStzBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDrEFQXAcv0RMJDRDzKAm9d6pAc/hVAOtpjJUu6i4j6R0fj2we/Xwe+zhByivyDfY+EqEHNKcJDhm8aVzVPzxd1SwFgsHfuuaTB/SH/kfW8KmqzkHOTCS30lXS3eknAq/xtq5rJdx2fk7oVYP8izPwbjrD1oOhUnp8jqbdmcoQYqPGeonAj/cgyPAYBBfYilrCakoWTY0fIsOcBG57Wr+0Oh37cEVTJFRrTAWCwd+65pMM2Su4OGpqX+odsg5VWSF0PAWCwd+65pMEXzqeoqfDCheLBEeDGFRu5dHSO3AsZMsLPfPmj9XUVawFgsHfuuaTB/SH/kfW8KmrB5JIIdSKgVH71nYZ2gpuIvIzaDID1+UZDRDzKAm9d6pAc/hVAOtpjJUu6i4j6R0XB0S9Gn+SMBqN6SPs8vLOXyq0GYrtXGF0v8MthD2qTcwFgsHfuuaTBI9kKMFmdfDYH8kYOWp05eBH5d5Nb5sfkLFbZouw8esatEi4/dVHuv1ZmiKIU3iofj/vgimiURQCEpC2QWlVtqWmgBv7vT+q1cum+Jd3Z/Lag18ZZFxsrfeYj6+rMrrz2pkEbAltJTXcjsdcB259qXgotjUEDptk3HnAUCV7x/vEjBpGmAhK5EOvzm46oTw3GUUHQYVZ+36CDSP9OTl9aL+OKCIfZmM5jxR0c7TiHsXhAETdKGezxdAi5nyDP1E0Di63Y6oC4qn8LX98K6mygUD1qrowGFRhSc9MSGVo5EeBhrvt/y+YAdeDspfEuZJsq+DjPiLxdnn3AbcsFcxHrhTvyimly+4ItoVOelkqJIZ8BYLB37rmkw2DJ/p/4Tr3uR7PrKZ4w5vBim8kWnK7ZCCQg+sGB7+ReUzsVX+qjJ2SOL0yshwRnPzeLjofpA41Y6dAd+x43Vbe4WfENQw4d7kNEPMoCb13qkBz+FUA62mMlS7qLiPpHR5c53VVWpRXBblxhN7uaZ/CBdQmF9fE81wFgsHfuuaTB/SH/kfW8KmqzkHOTCS30lOS2bMRXLafix91ggRJwKhqtEi4/dVHuv1ZmiKIU3ioeQGHVbcE4WYeXOd1VVqUVwW5cYTe7mmfzmtfvzyNlAgMBYLB37rmkwRfOp6ip8MKF4sER4MYVG7mHTdqcStfnQnPvrzUAkMW2UcU5/fYwwoEjBpGmAhK5EOvzm46oTw3GUUHQYVZ+36CDSP9OTl9aL0DzeiZcNnMufsyT7eXUhjQQR3LGsnLGJnRpRErudjt4GPp0kjfyJjuZqm+7wZO0VvcNB6pmFmDPBvwz4GMliPOjS7z5XwI5GwFgsHfuuaTDYMn+n/hOve5Hs+spnjDm8GP4WbMclbdleyUaUMqrSthQPBso56xSPlM7FV/qoydkji9MrIcEZzxfznETtsNccTQbM7YMtlDbiDpcAhozyGOiT4a7qoJ48GGu+3/L5gB2DVgVGxEJLFur7MnDMDSBIjmUoAoQhOLe9w0HqmYWYM0scqvz2kvPHeHcfhmRGV2d76HVCkFwS1MKRtQL/Kaal+fRVtt9AE2gnI4HlVbgl2x5lr8oQnHro9LwbQ+k+4H1T8J4kiBV3XVpoAb+70/qtPBRehIFeP5AvqBEktYUG1Kg18ZZFxsrfZjySmeLaPso2ZwrMWv7A5/j2we/Xwe+zhByivyDfY+EPOWagzpbWaBAETdKGezxdAi5nyDP1E0A4TJTxhk+Y/8jsdcB259qXEjboyxTc6guWJR3wf86mc476QwT80CFfwFgsHfuuaTDfm5UNID2G0ybmqPSw9BggqN6SPs8vLOUh1Yef+0iajacB+idEPRV+S/wy2EPapNzAWCwd+65pMEj2QowWZ18NgfyRg5anTl5aaAG/u9P6rTwUXoSBXj+QBBHcsaycsYmdGlESu52O3pCZrJixdNt+85IGI5msKUopU/nnc0r0rqPBMYH68KDQC6p3eFmTShqmYURHNrLDk5GMZSUNb0n0c1E1Q2lqdtHU7ynz82vQdVrL2xd/GFnka2fhra+8NHoGRTgk/5PXU/ADa8fsbx9WS/wy2EPapNzAWCwd+65pMEj2QowWZ18N9srM+qOQfF9dHSO3AsZMsDAOq3/jXM7BwFgsHfuuaTDfm5UNID2G0ybmqPSw9Bggcij4eRVyAumEHKK/IN9j4Rka9obXe2n2wFgsHfuuaTB/SH/kfW8KmqzkHOTCS30lISkLZBaVW2paaAG/u9P6rRVhtST5GUZBlM7FV/qoydkji9MrIcEZz2UnJ/9KeMYWBH5d5Nb5sfn3gA+/forxpslav3teKY5EwFgsHfuuaTD/WDiFZb3HScj8E2OMD64IdjhLaH2iFg7bzi48hZGtVXTnn/Q3m2GLwFgsHfuuaTCNmlGfQjyG1lqAH25hGVE6wtf3wrqbKBQPWqujAYVGFILawPlQGbCQAWDQJ3KBpIOSxWonF3FK3JxqletPrBLE+OKCIfZmM5hgluQ6tB2Q8+jS7z5XwI5GHmWvyhCceuj0vBtD6T7gfUwJcdmni3wffpRLPm1xe9welhgE7enf4hhrvt/y+YAdg1YFRsRCSxapl7Nk+TGKVdWYYYKPNgs1PR1ZPkCG95GrRIuP3VR7r9WZoiiFN4qHkBh1W3BOFmFEYxRziOLSXPiY6kXZLM45DmcHqJVUSBrAWCwd+65pMN+blQ0gPYbTJuao9LD0GCAvIyoSO4RMKVZurVyHEK9cS/wy2EPapNzAWCwd+65pMEj2QowWZ18NVZ63zPU5B7qe/noWG6oc5gkIPrBge/kXlM7FV/qoydkji9MrIcEZz83i46H6QONWLyMqEjuETCmbN/IpOSPFvrOm4GNjZXJtWsvbF38YWeRrZ+Gtr7w0eusFWlD/XbfQ0DzeiZcNnMufsyT7eXUhjXTnn/Q3m2GLwFgsHfuuaTCNmlGfQjyG1lqAH25hGVE6YdN2pxK1+dCc++vNQCQxbVCp/KraujiurD1oOhUnp8jqbdmcoQYqPJCgRjhqvVveIrElYxu0/4riDpcAhozyGGPyhEXhvResGGu+3/L5gB2DVgVGxEJLFqmXs2T5MYpVTnsJf44REAdUVGGFf1TOxTJ8ZKT9NA42q0SLj91Ue6/VmaIohTeKh+P++CKaJRFAa+7pNWkiA8C9w0HqmYWYM+zNwynoV0d66NLvPlfAjkbAWCwd+65pMNgyf6f+E697ZbOSfwio58i4NYWZC3rCCyS+Rcv2KmnO0UXMFcxrTQz00/rRzRJGEEZ5O0bCUiK511AMSyq/CIsbRK1P8MhWLRhrvt/y+YAdeDspfEuZJsq+DjPiLxdnn10t3pJwKv8bauayXcdn5O5Zb/h0F1jGIpAw1kLg9YCWwFgsHfuuaTB72cywEGpcnODXEbg5AnphqN6SPs8vLOUh1Yef+0iajc5hShCxZBTKAWDQJ3KBpIOSxWonF3FK3MEkaS2Wtaw74m/RGRXCtaZafD/+ALxcOos+NGHYh8aRkNEPMoCb13qkBz+FUA62mMlS7qLiPpHR+PbB79fB77OEHKK/IN9j4SoQc0pwkOGbKGHwLihVpzzAWCwd+65pMH9If+R9bwqarOQc5MJLfSVdLd6ScCr/G2rmsl3HZ+TuhVg/yLM/BuOsPWg6FSenyOpt2ZyhBio8Z6icCP9yDI8BgEF9iKWsJqShZNjR8iw5TzZ5bauRpRbftwRVMkVGtMBYLB37rmkwBfUABJ2VAABsp3ienJkCocBYLB37rmkw35uVDSA9htNL/SY/hOJxWe6gnuh/ZnB5aFTnpZKiSGfAWCwd+65pMNgyf6f+E697dml7fv0UTkHDz5/Wn/KoANMX9XZt2jt8HmWvyhCceuj0vBtD6T7gfVT+trvJXZKxAYMFitOKjYBIwaRpgISuRDr85uOqE8NxlFB0GFWft+jFAlrSidnlCGOCI0Z3ORy3OUb99pwMO7p10/C0a3Aixqg18ZZFxsrfeYj6+rMrrz2pkEbAltJTXeaTcqpZECin4cBGJYCW+yyNXNSQwmjP78BYLB37rmkwjZpRn0I8htYXZE2UWyd6mzkhMLjxqTX1kxtyBmu19WwQBE3Shns8XQIuZ8gz9RNAeqTX4NXeyDA5ITC48ak19Sn/1e8nIOpDs6bgY2Nlcm1ay9sXfxhZ5Gtn4a2vvDR6ojhAoeagjEnrRpAsR9do3dLOqYxTPvUKGGu+3/L5gB2DVgVGxEJLFqmXs2T5MYpV5pNyqlkQKKcu87/7MsXuowQR3LGsnLGJnRpRErudjt4GPp0kjfyJjuaTcqpZECin4cBGJYCW+ywtsoi3da+UyMBYLB37rmkw/1g4hWW9x0kcAJOOq9NkjTgXPbBMoC9aUgW2JZuK+B1IwaRpgISuRDr85uOqE8NxlFB0GFWft+jjgzOf8xiWgOtGkCxH12jdDhWQa9a3tl0BYNAncoGkg5LFaicXcUrcJdsLQ2hnAc/rRpAsR9do3ekkuHRzZ+QAwFgsHfuuaTBF86nqKnwwoe4a4KqgcHCjOSEwuPGpNfUDYaMh8xH+4WhU56WSokhnwFgsHfuuaTDYMn+n/hOve5n8KPV1dvxHOBc9sEygL1o6tWBVgXtDkKw9aDoVJ6fI6m3ZnKEGKjyuN1MGpFElgjgXPbBMoC9ameJ44+LuAP/j5RcgwgjQhVrL2xd/GFnki0LUJJpIrXXKifpOavYV1cBYLB37rmkw9Yrk216GSMEYa77f8vmAHcNmJveQkPR5UQDEX4lGWKxqORwzQdMkxQRM5a3QoG6cNv1C5IcM1159+qWmlydBZquwSwszM3a5o5ApiwLYCZD/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyPXyMGM0AOBla1A5cy9wjnR768ZeCgbjyTgV6rS7d/LrBmEj3gN/qPO1vv0WSUjnN096ji5zwFdGYSsfZpa+2kZpIVGa7hueH6USz5tcXvcjczSu8TNAe5S5qd5T4EWL/BLI3xh8EOFKJWCrVLsSynBJGktlrWsOwpksyvr8aJyiOBKVzxmGVXBJGktlrWsOwpksyvr8aJy3bOolX2jUIns5bybePbTw10t3pJwKv8bauayXcdn5O4QflWiQVdxCKwZhI94Df6jXS3eknAq/xtq5rJdx2fk7tP2As1htXkj7M2Jy2rueEbzkgYjmawpSilT+edzSvSuo8ExgfrwoNACTv6eBnWO2/OSBiOZrClKKVP553NK9K6jwTGB+vCg0IaJAM5lfzotiPBa+e1y4mI/AaikY3kVDr9GryUan92uqelc3ICaMs8/AaikY3kVDuxQILc3cqlTXBfVVxFmFh/IAIyXWxsyLlie/yxOw5Po4IjIBgwS0cgDRGU+S2KBe+wcnqbgcQbsrqtFTxYqE8cVv3X3JZrjOSTgV6rS7d/LHcx/u38Wt/4j7LFPblToDvttuSV3mxucnHPfy+yGTjEo36jxjcHPC0RVGXD4Jha91wH27+pZglAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu4HJ38+96tAVqpLnfMG0vyGctd0h9c7W82lBBZ/ke9hT56hrqsU0m79BIfZhkVbfEV4TpnKmhoV9tabHMeVL1c+Fj7EA8Hh3eSCBV9piJ57fcV7Ln6bBGwp2lhDgUDVcPpCgYVS10eezjsPT1bqW1VjaqMHLojSgksfSYnTjLdZAbdIk8JrCDetr6QPzgc5BSXmJgIALYG4gfvV2xNh8SMNRMwuztBDu64UuMI98FLMhE+/MIf2tmdbgE84d+DW3PZtLL+yybWpx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7zhC1rRWGiQMZC/dfqF4dQAByi4Y+C90Y1qeF/3xLYVjbHasb8nNKb74TviO2/cKLXyY4p3wSQhQun+fadIqyRtOCB1pVP/YIVe74nJ6edzid0R9SwaTlvBBQDkg8Q3rOQ9zsKk8AIidXQoFv1vZWB532mKjRs8Ag1fLXh+RnpyEIEpOCqB/ZTAV/O7+mBoutF2UR5TB5rHKp+MzEJ5LdcPBufqCD0fWOqodQwHie9KAWDQJ3KBpIOfoAOLnMoIH/I5P9o1JFlvcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/m6EfCirzLRNmAmFR3LKaecIKQH9xapKWm5wIy7VEbo16nDPYWVBQKxr7gmQoaTxclM7FV/qoydnBYUSx7a+c9hxd+IAGZeat6QoGFUtdHnsdg1suZ9E6/0VOThjF2eJ8rD1oOhUnp8hO7JRb/x7EOGP9xRVykDveZgJhUdyymnnCCkB/cWqSlosXUWREpEzCjuSvHYd6S3WsPWg6FSenyOpt2ZyhBio8dEL0FCtBInjC4OEyxUpTD8r2YSpbsk4ZTWxcDlor/l/BH6ab6nFM+q0edPGUxp3RqXINbESJTwlr0IpCVjxOwjpKB/H5OuK22XUHabPGTslipQ3jNDYXS50aURK7nY7epa/XkEGd4zccRy4n5G9LBnPKxSUCjyIDTUfvZh6UJ3Th3bk6/jehEv19Zgv4+tSFHYNbLmfROv8nD1iWiaJSn8Ti1pQijpegMCAsaLkc9sMCLmfIM/UTQLuZWZvb5BOW7GNtU97kTE2foAOLnMoIH9CV7yFXiMmkIzPCw2hf+8xmLz8gUkNZ/g8mjkG8s4l2WIIAIds2MSqzpuBjY2VybYVTxHkWmBnXz9+B5bv6EKgwICxouRz2wwIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTZ+gA4ucyggfcHRL0af5IwGo3pI+zy8s5cWrKszvv/rP06kW6kYzVm74AIVNIXWRQ2vQikJWPE7CHYNbLmfROv/I7HXAdufal4KLY1BA6bZNyFcFEqvNbKhz8MUNenG+KPgAhU0hdZFDa9CKQlY8TsIdg1suZ9E6/+Zqm+7wZO0VvcNB6pmFmDPtNEOHVgwN3IqNfsYn/oxSg0cDMgQwDJ3sY21T3uRMTZ+gA4ucyggfExWZul1JXMYsPDWCzFWleJ+zJPt5dSGNMxbLEFcH998vkB0cqIEKCxxHLifkb0sGc8rFJQKPIgP00/rRzRJGEEZ5O0bCUiK511AMSyq/CIvBt2t/xBQa1aw9aDoVJ6fI6m3ZnKEGKjzH8YPSoAnQYMLg4TLFSlMPh6LA73E/7mGKzno9CbS6ZZjcmMTr7dw49aoR2gafujcGPUiUezMBVCSJw00xaEzAZd/yTly2zIKznFAuVOxFiKw9aDoVJ6fI6m3ZnKEGKjzH8YPSoAnQYMLg4TLFSlMPsUJYN6b3gXtS5qd5T4EWL/BLI3xh8EOFTBfmMEiBdjqvpcCTSiWwOMfxg9KgCdBgwuDhMsVKUw+xQlg3pveBe5HseTWJFtJxy94DfxPvFWat1/Xiw9mMXymhKUrwb+quRgvHF21aQvfhwyaAxLfQPXVkydSh8I56zFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QWd+lmj5NKBs2MaPYp7K69/gAhU0hdZFDa9CKQlY8TsI6Sgfx+TritsEkaS2Wtaw74m/RGRXCtaZafD/+ALxcOv2UEWSsyzn/j2idcEsQWxrNzaJy93Vs0Woc4gm1k9npHEcuJ+RvSwZzysUlAo8iA+zlvJt49tPDXS3eknAq/xtq5rJdx2fk7iKxTx/x1+pBpAsce8A1ZdRjr71WCqHSa/WCKtFaAB0pbUXfYiX6zhRcF9VXEWYWH8jsdcB259qXEjboyxTc6guruDnuKlgiyf6ovbZmtlIuJeg+iExCMrmtHnTxlMad0XrnCnbtiaHi4cMmgMS30D11ZMnUofCOeg3SZZmoJTcfFCNaiJ5DIyxW18zeCoGwTHdNhcCP1m7KrD1oOhUnp8jqbdmcoQYqPMfxg9KgCdBgwuDhMsVKUw+xQlg3pveBe8Qzp20SDb8DfKt2HNWd67OznFAuVOxFiFM2bu+WFHT1KJnyGPmNyWbhwyaAxLfQPXVkydSh8I56m6GX1On6ntnlKPIgzV6cx+IUZKlNrIA+jMV4TVdqFIoxk8wvrRXYtexjbVPe5ExNR2fVmEyqvVMVv3X3JZrjOSTgV6rS7d/Lj2idcEsQWxrNzaJy93Vs0RfzvLOuA1LyHEcuJ+RvSwZzysUlAo8iA9E7UrJs3PaOKhYlwlva71ctcvQ+9baQxR1ULW2AWLCOHdEemZnDHWscRy4n5G9LBnPKxSUCjyID0TtSsmzc9o4qFiXCW9rvV8wiBOuPjSy4HVQtbYBYsI4d0R6ZmcMdaxxHLifkb0sGhWOg6iIp1UbuDmirbUrVEiIU7QAI0CB4JvL2HlIyp6+tmTbdvekH8lQEo83cZQQWgpvZrikp48oKxI/FfaDQceVeBx/0a7DfFIjp1DOt+yelEQYVtBkl7QGAQX2IpawmpKFk2NHyLDnmwLkSqPVwnjXCwCliMuDd1ZmiKIU3iocEUr80Y7LPoOxjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3cjsdcB259qXEjboyxTc6guruDnuKlgiySAvZetnnrzMzc2icvd1bNFqHOIJtZPZ6RxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnEnO5Tmh2rEJ0o+O65vGKt4NYzrp4FTWbcIKQH9xapKWFIjp1DOt+ycoIfJMj+PGie/5Eqm+ukWSr4ePFoHgHvitHnTxlMad0d8nmWvce47q4cMmgMS30D0UiOnUM637Jygh8kyP48aJIURZooU/2cQwO89C+dp7igIuZ8gz9RNAVFsWBq8BmK9r0IpCVjxOwivkwtmFLeT25dWadutRB1oqFiXCW9rvVwo39bRamoqip8rEBx2amh0RaygtE5naOViCACHbNjEq8kyiJFHAjB3u0V+ntFmUQUqRU4/TOBeKB8coSla1YDf5DL4JnDfRvItJFi57rHJCOB129t1fowVtRd9iJfrOFKcnp15/O3TdYcA9PvGn5qi0bAtmK3K/E8RJwUoevkHJlM7FV/qoydmdE8lMvwJei3NszWGG6djIb4w+NSYBw06nLGqSXI8EekHI9aDL4/wTD7DkI+4jM/Jr0IpCVjxOwivkwtmFLeT2EhfxS9iprzW0bAtmK3K/EzEtf4YeMykKnrgr/BC+fs7sS2HATwszxcLg4TLFSlMP50r/6zZg8Qk5Rv32nAw7um+MPjUmAcNOULOUxA+H2e9ByPWgy+P8Ew+w5CPuIzPya9CKQlY8TsIr5MLZhS3k9uXVmnbrUQdaKhYlwlva71eTOADH7kQ08KfKxAcdmpodHRAfZnbsr5pYggAh2zYxKvJMoiRRwIwd7tFfp7RZlEFKkVOP0zgXipTnmDH7+vkSIC9l62eevMxTMzE3dlWywCvkwtmFLeT2EhfxS9iprzW0bAtmK3K/E8C8zagpaakFnrgr/BC+fs5OQZIm7+zr2MLg4TLFSlMP50r/6zZg8QlZzNXBh+3npJTnmDH7+vkS+Qy+CZw30byLSRYue6xyQjgddvbdX6MFbUXfYiX6zhTzqsUZ4hmxNgH3Q7zkTtBlOBc9sEygL1oqXRnym4B0g6w9aDoVJ6fId4AgF2l+b7EwAd6g43GZAAxou1l86AvttGwLZityvxMjmefQ8sf6M5TOxVf6qMnZhPQpA70YWs8FFHdQTzdYEvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHbJ4yCCBRH8wkkY4aqKm1qbB4b9+WeicmfDlVqGPuyXOnWwuOpNw74fL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkw8panoGjgQmCsSPxX2g0HE0e8e2FRjmWI5wsN366cbVER/L5RBJnizLRhPgGFlt59Crq+9aP37oqDXxlkXGyt9Yt+40/kUJWEhPieK3qr606qm3XMv4wdY73kiJl9dwNF/sZKgIM5LBlyJNSZWXY3L+a+lqmlo52UTe3KALTTmkNORLbik88sawoLfxgcs7Ci+595hQ5cfi6IPljoFU3Y/JEKU4QhXiLLyqTLJtk8MmG4jp3h8J04jcaUoX8x86ri+595hQ5cfie+rN2J8ozW0Awj97MhAS3LPE7sQG274opaphVYGdTD6YF0ARu0iAQBRwdc7T0xcUf0h/5H1vCpqT2QQbTYkLPkj2QowWZ18Nv9281ooBjDZNR+9mHpQndOHduTr+N6ES/X1mC/j61IWoNfGWRcbK3wwiFoYUwg1WI2w5q0jce0nMAv7OgW2InRI26MsU3OoLYk+ciHfVdO5+uhSGI6Jxzu6gnuh/ZnB55NUf9KsXw/VdHSO3AsZMsJ7JkW377qQRTWToPteyKxHTREZwfW/cdfnI1rhdV9G87qCe6H9mcHm/3bzWigGMNu1GgG/AnejDBH5d5Nb5sfkd2Ig3SMjFLcwC/s6BbYidcij4eRVyAumEHKK/IN9j4YBKh+Dvf72/rU2twQqZwVZ2OEtofaIWDtvOLjyFka1V5NUf9KsXw/XC1/fCupsoFA9aq6MBhUYUfVu1bEHwO3p+uhSGI6JxzsCTsqSLk1SmXslGlDKq0rY9MdiT0cCYeHB0S9Gn+SMBVFRhhX9UzsVV7fV7Aa7Oeag18ZZFxsrfySh5PTH7gHGheTGTzEMSDxULXnWGb3lIje3TlPFyPxBr7uk1aSIDwL3DQeqZhZgzRgtjnoB2E/GzxO7EBtu+KLCXC0N1chMBVFRhhX9UzsVF1l9xS4q8fZeWqdvtSnOue+h1QpBcEtTCkbUC/ymmpWWVmqg7+gaBqDXxlkXGyt8l2wtDaGcBz+tGkCxH12jdNkfQ/WDgMETmk3KqWRAop+HARiWAlvssg1aFEXvS8w7nRfYQ6QVJOW+MPjUmAcNOk6swZ1dVcf4wys9hwcL0cLRsC2Yrcr8Tq0kfHZDJh8MvufeYUOXH4uaTcqpZECin1QUVKwOqtDjCKKZynyH/qzkhMLjxqTX1RtYkc/Cdu6q/3bzWigGMNt01OfBe54mmtGwLZityvxNuudPVvav+d1nM1cGH7eeklOeYMfv6+RKv0rC0ZJZKRIeiwO9xP+5his56PQm0umWY3JjE6+3cOPWqEdoGn7o3g1YFRsRCSxbCHTnGJiwHXcTZrR9MdAnrzwhKox0mUQKVrUDlzL3COdHvrxl4KBuP9I3FPl78GcioNfGWRcbK35WtQOXMvcI50PpIV6W3I+BMTdA565G3W+zlvJt49tPDcBtywVzEeuEmkPvW1+PXu2DUy0bAGUzIiPBa+e1y4mIvIyoSO4RMKUxN0Dnrkbdb7OW8m3j208M5LZsxFctp+ECs0j5BTIieqDXxlkXGyt+VrUDlzL3COQGAQX2IpawmpKFk2NHyLDn9EjKdxJWHoL7k/wNm3kcXyOx1wHbn2pcSNujLFNzqC5YlHfB/zqZzv9281ooBjDbs5bybePbTw10t3pJwKv8bauayXcdn5O5Zb/h0F1jGIiVgifm0v68T85IGI5msKUopU/nnc0r0rqPBMYH68KDQDrn8EXq+wzdmPJKZ4to+ysEkaS2Wtaw74m/RGRXCtaZafD/+ALxcOknNL1KMyKR2la1A5cy9wjkBgEF9iKWsJqShZNjR8iw5efN7qTiUviNg1MtGwBlMyIjwWvntcuJiqN6SPs8vLOUh1Yef+0iajeyentuaq5/lm74Izq1+Jp3I7HXAdufalxI26MsU3OoLq7g57ipYIsnAVrhE08BCVrFCWDem94F7to5BnAspnvEwDo6LFTDqtEFR/6HluXRC5dsb2UZf/n0N0mWZqCU3HxQjWoieQyMsVtfM3gqBsEw760ulS6hDBwY9SJR7MwFUA0RlPktigXsbXdvOLveqRX4/i0JUzvQQm6GX1On6ntn3U4yioDBJCxDKoUqYp/6YsUJYN6b3gXvEM6dtEg2/A45np4cZb0Z41Cnh+RIbahOI8Fr57XLiYrZZzmiwPIDzb3qcVjfDQXlg1MtGwBlMyBW/dfclmuM5JOBXqtLt38uDKJIWr5GLPE/E5ugctI/kNRjP9Z260P2xQlg3pveBe/2h1Zn893TC60aQLEfXaN02R9D9YOAwRKF2IlEkBcGdOBc9sEygL1rtPM69fvLT1WDUy0bAGUzIFb919yWa4zlvjD41JgHDTpOrMGdXVXH+36fLQW943BgqFiXCW9rvV5oYaCbLvh8qgEqH4O9/vb9cF9VXEWYWH+aTcqpZECin4cBGJYCW+ywlYIn5tL+vE/2h1Zn893TC60aQLEfXaN3iqlMtnHVpcoNWBUbEQksWYcA9PvGn5qi0bAtmK3K/E7GSiwtjHZnOOUb99pwMO7pvjD41JgHDTs3cvurT5uT9qDXxlkXGyt/rOASvJyBn0DkhMLjxqTX1A2GjIfMR/uGbvgjOrX4mneaTcqpZECin1QUVKwOqtDhPs5nBXQ7LOAY9SJR7MwFUSpFTj9M4F4qU55gx+/r5EnTF9b0wdUvcYcA9PvGn5qi0bAtmK3K/EzHsjhcX57NBcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHgFrUi5tevOEL53KpOkk63dmWdpXmEx86h7k7D1GEvvHNqyLGdo9RMlnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8w+7l25Aq3MqFiXCW9rvV8QNBqSuW6b3IPEEOOs5sYJFhs+T6mvC3Bp5IRzli53X5CRqz7/gFKofUxVuCXS5Y32Pkite4rtGKQ9XKZKOL02NVcWq422Esp7WNoaMRI3YKhYlwlva71cKN/W0WpqKosNwP71HnkU4bPz/c6/JJ/2iPRAJAhOGHlo1LtHNujgmb4w+NSYBw06TqzBnV1Vx/jSc3R/HQ5ndZL+814w1rJYvxMuc4I56TqgxK8NU4X2xtGwLZityvxMQiHeVRL+uJ7twcZyZxxott1OLXHeZwhiQ0Q8ygJvXelnM1cGH7eeklOeYMfv6+RI5jnp/dn+BTUCGgMvrUkxxN+zZPe2/uq5ourMmZ+Ww9Je3XicDJZZfQ1pFmvl22ruVzBspFARCWZacAGSF9jAb2K6hMdSPTRxu5myMb7+Ubwxou1l86AvttGwLZityvxPclTqO3gPXvr8RQpZeJabnqDXxlkXGyt/OhQG6PR1ti+tGkCxH12jdopx5R3/v3PGhdiJRJAXBnTgXPbBMoC9ay+Bh5O1IhJ4Ya77f8vmAHVnM1cGH7eekB8coSla1YDd+mOSvxVSOL2HAPT7xp+aotGwLZityvxMrUfsiE+X0TIMqS9j75lvBvoiGCRllu1RC9k6h5Y71Xz4pGS+yYrWOb4w+NSYBw04t9eqo+YceYykJuMch/Os1uWDl+4FOsmiJRkkmMiKGuDgXPbBMoC9ahE8I+GjfVBQ8XGHc0O9eNjkhMLjxqTX1RtYkc/Cdu6qQ0Q8ygJvXeqgxK8NU4X2xtGwLZityvxMhM0qVZ/PNsDlG/facDDu6b4w+NSYBw07YWAuy43ftn6g18ZZFxsrfrTIP0x/AMDCDPmhAtpi4ZmsezOrWWHiu9orqZYAgHpsdWsUzXETiNzkhMLjxqTX1I6uWZM4WiPDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+XJ3oG7RzGOQSpFTj9M4F4oHxyhKVrVgNzQKBcmLoXUzOBc9sEygL1qxf7jLkbuO1lnM1cGH7eekB8coSla1YDcdIKi4txdgBOs4BK8nIGfQOSEwuPGpNfUAKi0QDYMzvFnM1cGH7eeklOeYMfv6+RKX5p/+6Ze3JTkhMLjxqTX1RtYkc/Cdu6qscQE1hVaQ5/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxoOtkMX1nWY1IgZF8gk/1pecEU277zU0vAWVDcTjYlD0JYd7j9T2mGe9naGprhUz+8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEcs4z//HVLKAG9vfSuSvr4acedo+JueoCzJDpYeredNQgNU6sZ8BLqyUUwDM1u4gaUnsIwLE1+Myjrs7IZ1ypQh9Gheh0xg0hrRbTL2mz8el+B4LDznFf8qAYBBfYilrCakoWTY0fIsOebAuRKo9XCe3Nz1ZiHQO24O+z3TIorV+cEkaS2Wtaw74m/RGRXCtaZafD/+ALxcOljkoRbCtXm9o22LrPJSog7syy/8/9ieOvOSBiOZrClKKVP553NK9K6jwTGB+vCg0J64Fa3BVLwhf5ZqjnBY+iubvgjOrX4mncjsdcB259qXEjboyxTc6guruDnuKlgiyVb7lQsvEPggqlL50BNHhaHgeCw85xX/KgGAQX2IpawmpKFk2NHyLDliI0tlVN5G8yd5/GoddaOY0/V1T+XTxq7BJGktlrWsO+Jv0RkVwrWmWnw//gC8XDrg8MxZ7cKwomues+3EMfEYTAyg4wE5Olj9odWZ/Pd0wutGkCxH12jd4qpTLZx1aXL4hU/M2Oe/ZqF2IlEkBcGdOBc9sEygL1ohZk5QeXdfxXK6S8nT52Gw6kJFusAILs+fAxfhBIk0BL3BTyOII8sF/N6ae7tJIZPNH/ZDgVYAHmN8sXUG3n/RMO1bv9UEx+3U3SEseafKeLMgixECuy4Y9AfSPC0BZ5xlDaSwVAFb+1LqVE2RLi71WCwJTZNMBBC5cWgCyxE3TNHxZ0kVM76dxrqg5srPf0Cs6bfL0BsCGPjkhFrTpNh5Ld0RaCT/cJAD45zU2m2HryalmxDBvT6yulhRBnYeT+x4Y8XqlYotKyqiwbt8jjHafiqJ59OKOgAfILcYi00x4gezedDC0hirkYxlJQ1vSfSLQ5tkpKAu5vn7t0tzKCwwVHyeebhbnG/T1x5TqIrJNmfddM/thkk+2cboipD+QW6/3bzWigGMNkoaRYcz3zZKmzXE6Su/2agGRAiCuFlYta0zQroSE9ZxkARO2IeEWT2f5g/iCtxkFSVHGXsjrdkzXC9v2/I6sdos6dMhzFAQE6Lw7qSoagOKY027kY+hSE7qn2Nu8ODbYKepMQJ2ZS5BKKSxzQG6RNNhiXBoeiuGTOzlvJt49tPDXS3eknAq/xtq5rJdx2fk7llv+HQXWMYiMaNlgpp61l+0oqCpiNtbWc0BE0XiGAz5J6W/8c7aWJqI8Fr57XLiYqjekj7PLyzlIdWHn/tImo1m+nRDeNTOHXF7Frm+c3rWuB6/XZGBm+tWTQhnnyXMXxmErH2aWvtpzFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QsIlxtsc+EdFfWADTFbkpBDrs7IZ1ypQh/BRGDCmA/lNyd6Bu0cxjkPj2we/Xwe+zhByivyDfY+EqEHNKcJDhm/Eshj/tbNiP4jQSFdUtWbOtM0K6EhPWceqbQonxEKAT7OW8m3j208NdLd6ScCr/G2rmsl3HZ+Tu+jci+PTO5roapsBY8gKl6LSioKmI21tZzQETReIYDPkPr0i7CFTbVYjwWvntcuJiqN6SPs8vLOUh1Yef+0iajeyentuaq5/lZBz+aYFJPWi4Hr9dkYGb6/gBEy0xY0HF8OshUXtxoGV6L67qm9YqjutGkCxH12jdss3OExllqELAWCwd+65pMDefJCHSAxHTOuzshnXKlCHjAA6L8Xp1+e++cu9RckSt5pNyqlkQKKfVBRUrA6q0OBk2Hyi6fqguwFgsHfuuaTDiNBIV1S1Zs60zQroSE9ZxlSP3MtyY4Q+XYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZhmbc54Qbzm7vt0W25erGITJibuQ934z3OZsPEA18kKxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Lw77OF9d4rOWvl9lNkq+IdrX6T0NpFxbWIc83RD0iU+Wvu4K8NlLooedDa8/RTQEBD69i27DxUHP/OYV0R4td6r36mE7lWClZdLuAG7fM0+01lFoJxGMUvrE1ERmVr3ctnlDzC/UyHOcmKOTp/XSUc9AVhiGX5cAqAnUpz6IJrHphmfKdOuCiuosGwRjmsKH3H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LE6S3a9z1k0WeUUQ57P2dZ/D0yVYSr1ZqQun+fadIqySUzsVX+qjJ2VWvn3zt+a+v56uqKHUzj+O6ErXIdZ7wR5yW6ej+suMWMlqR6Ss0rWoDOFhnjRMVgSNs9/cmJsZLG6qKbKHdyHOP5V/h1cQVj8opqYJu9OzNGtjw8+7/VQTlDeT6t1fqCwFuBF7N3PvTXCCRAji/cCtoNxvyQ8QW1jqzXWRBCXLpIULKBjHbC9aWdChOLqh8I+yxO15SJPekjIrBAkhPCHm3Pox8adc/EfaUX0X95rOSIULKBjHbC9Yi5B9R1EywYtEdm4kAmD5cVcV2Z8tlKBlIPYjjdDk1OlxhWqlEb1qfFIjp1DOt+ydD9eIaXiRUpWGB2S+nN5OwJEFN2uPF39oH4hDXtDroPcvBWzzTShFhK+TC2YUt5PYpZGx5Ak1/OOSHHXMLYBB+Glgntp4CmIdywW88GIzBey0xkdbNjIsndayI23t8j5a/q5DVtD5XU/mD7dVSTCwE0RRoVXO6yLJG8h0UlviqMDD5G33ufRzxQgfeht6B/8jGIS/YfHyIGT0l/ubPO3BXcLpMDZXOk/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwt3gjIEtmkGJUn/JVTdmWYH6MQhTMtwAUK7cvUi1o/TGoQ1R4UUhLal0nUbGM+SWQTJ5r1xzfDXClC+R9yUfoJ0Gb8Ye9mOhQPlT58qADgnayba61mL7BzZ2TkZnHbsHBPxbmei8NO38d0W4BD0aFKU5lnjpedoRzAAyrlX0gor6tNzUEBQoLQ8H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3LT0/yG2IDtrlZ8IPyDLuv+l9xhXNxWN2T7/oIFKmhD71zhlzDSb1zNzaJy93Vs0Uueqp97NbplmPQQkgisl8tYFr+MZcxVHaX0mUNa8pVb7RtZNGyzZJmeUUQ57P2dZ/A8CkU8l9zSwvwJH7XcHtdGsySS4glDgbXyY4p3wSQhwvwJH7XcHtcuWTz2nKiHVApwh1Sk8uYlNGzsQ7/B5p87T6JQ+hpNEcvpGvZGvxi8I2z39yYmxkvSgIrk3Duj8dZJwV5YQzzo2zuBuy0M3lqwUBTkL2d8olY1tXzOO1m7rol5AnwLiUQAupHEAvr/j8oAxG2oU6OZtfJjinfBJCHC/Akftdwe15Jm5jEAGLHKIwOFJe0n3VrbO4G7LQzeWrBQFOQvZ3yiVjW1fM47WbsXRqUBWJNamh2xYibNt1+aIqrp3xKIxtCCeBlNilgh9g+ieKS22BvCvXHlGkjxWG2GeNe/ViWaOstjDKcKHvRArnrDy9x642jE6QHOXg5vnMgr4u3Rc6GBKtBT7RKCf92tEZK7kisEEh2DWy5n0Tr/BMlZKI/I2EqsPWg6FSenyE7slFv/HsQ4HyC3GItNMeIa+4JkKGk8XJTOxVf6qMnZwWFEse2vnPaUytPcZGSb9eY4yvlTLgmQcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/WfoJvbUlc1kiNtqSbypkwF4JAwcpRs2wpWqh0Oh2IWULQ66nxKXucTrs7IZ1ypQhc0fGqjkjIA3BH6ab6nFM+gGrw5g00TiRiDRDjyoPEdyxeSmMOxMQeSzxwGiFvskxrD1oOhUnp8hO7JRb/x7EODssUGdd2NvHElde5mwLGJQEa0I1hCAyZ5TOxVf6qMnZwWFEse2vnPbpG4jXwUtOiPEZM0BP048II8v8JpqqcQYS1F+P0jKq1f6GaqmKuq2zi32YOSX61agxk8wvrRXYtexjbVPe5ExNn6ADi5zKCB8/AaikY3kVDhCI7jomL2c5nvPZszYH98tOQZIm7+zr2MLg4TLFSlMPAf1sDL6Ym0qNMqs1LN+6SydQKgT5HtzBdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDbEegyaglFcrK5z97NvouaslQhwwd/5HsD7DkI+4jM/Jr0IpCVjxOwh2DWy5n0Tr/q9XxkihgWvgvxK0eUeOr2jVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3h5V3hyOyNkFb7sR3hygJREr/N2MTaHVG9xFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybRUEU0INUM9QU2Y1ASpUICId23GDqg4YIyiZ8hj5jclm4cMmgMS30D2ncXb8pkNlLU7a+m9o2eVLc4SNAPWFs2eLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhTq/B1JkFXPe4W02iHFTZZkcuTCtH6/xJL49dKirrGTNtsqKEd60d2xG+n1s+QzRGCLSRYue6xyQoHGXTL4rBS7bUXfYiX6zhTc9CSVHsOFPoB2QMhvPCeJBwiJMwJX0fyPhAs8qAxJDuxjbVPe5ExNCDZMI+JrJV/yaiagphboiDpKB/H5OuK2C09wc74eqGbdL4+39QNswCXoPohMQjK5rR508ZTGndGpcg1sRIlPCWvQikJWPE7CNuF9Szb8bc9geRD7LDFinycNF6Xh9oRrcICN93vFAvabnAjLtURujZE5dDsUwpRpnwKOJxx/kycwICxouRz2wwIuZ8gz9RNA2pOVl8KOw1xr0IpCVjxOwh2DWy5n0Tr/oXYiUSQFwZ04Fz2wTKAvWrZp5+hv4yrOUzZu75YUdPUpOZdZQhNYheHDJoDEt9A9m5wIy7VEbo1hwD0+8afmqLRsC2Yrcr8T3PcKCVatKGyeuCv8EL5+zrkYd0JVXvBOcdmIiNk4jAj63I2TU/dOm6+/0IL3SXd/Qgfeht6B/8hYn9y/hYl4Yr7dFtuXqxiEA/bXJzI/US6knw/ucb4G1wWJ3QAeSDW4Be6VS+6e0RtpQKpSyhKwaUnbmS7X4ILX9KM91k9syYv8BVvBnRzJscLg4TLFSlMP50r/6zZg8QnAlCJBb+ant2TWU1Lsp7f7AqDTG4YpC0BYggAh2zYxKvJMoiRRwIwdaUCqUsoSsGmlhVaSdINj+fSjPdZPbMmL/AVbwZ0cybHC4OEyxUpTD+dK/+s2YPEJwJQiQW/mp7f9lOnYojEtEQKg0xuGKQtAWIIAIds2MSryTKIkUcCMHRyesVbja0nAfLj/Ae98T6QGIjfzAKxOnD+H1ckGx1PGa9CKQlY8TsIr5MLZhS3k9ht3+qACy3G9y9Wnow4neS7ExTNIirtarvwFW8GdHMmxwuDhMsVKUw/nSv/rNmDxCddVeC51aa+hy4kEYPmGHzv0PJ+X2fy9zzjgq5bS0R06bUXfYiX6zhTbA8chY5Tt3EGUJNT4jh8n/ZTp2KIxLRGxPs6payz5TFiCACHbNjEq8kyiJFHAjB32Dzls66/2m5dD51bMdApZAhLp/oYug/muMXrqyfypnexjbVPe5ExNnGokgdKcFFM26D8CjWxi2UKcDns3JUJ3BiI38wCsTpw/h9XJBsdTxmvQikJWPE7CK+TC2YUt5PabUaApdX2MkuMScs/XMppae7Xdkc5z3yTObbBmchPkx+HDJoDEt9A9FIjp1DOt+ycV8Z0xfobCk1Ntft7E/KHzxMUzSIq7Wq78BVvBnRzJscLg4TLFSlMP50r/6zZg8QnQbM+cXhKOj2PiyCm02amHuDMwYXLoEPjm1fRD6ARM91RWHJYQ/HeHQW6A1k/HcyNjK4O4odb+ZEQTtJphwmTr9Dyfl9n8vc844KuW0tEdOm1F32Il+s4U1L4Qj+QMsx19W7fTOPwRfWGB0Nl1SZ1ScA+iQw3goQIcRy4n5G9LBoVVIPUUpxe0y5YPbm+aghb6nSv+h723Cf2U6diiMS0RsT7OqWss+UxYggAh2zYxKvJMoiRRwIwdc2zNYYbp2Mjgx/liKPdavJKHozjh0OSjyJask47xBrjhwyaAxLfQPRSI6dQzrfsn5LjWZpzfYCCCZGxSkRLzrotJFi57rHJCgcZdMvisFLttRd9iJfrOFOytpJEzauL4YRAAZqWzjteQBJXS8jpjJew2DA9K74IQWUVJ780RjuPVmaIohTeKh69QIF4Myn71WIIAIds2MSryTKIkUcCMHYoe0imlHJn9l2JIueYbPAJZRUnvzRGO49WZoiiFN4qHr1AgXgzKfvVYggAh2zYxKu0cKYY1ofMCiKbLQzHQw9fTgI+gsDxqVRF6KSzOPHtSJV9ui98xHoPTa9jgkAF3BJQ7Ubq6BOimZttLRLcDJXD2qgcg2eo1NBPXNYKURi0fW1fnvM7QjM/W6GR/nSUEpISh7aB6tUPiJj0S8EAQi+bZdrxFpecIx33RtwrgoLtUFQRTQg1Qz1B44aPP6ROqtaLAxrcu4drApRDLRDAwZjZ/l1SO89wyltMX6BQpoOXjfoXvG1eW031sR6DJqCUVynqGdqtN+uD5EbH8bXD8bq4O7nzba2P/x5Dln1fPNXkgq9XxkihgWvjGld80emDDIoZD0YxFx+drA3aCawFio+4jxo8SKEj4//54/OM3yczNK7yieirFNbM/AaikY3kVDuODuUYXZuY/FsxkDCU1BGU1G+cfhF+1AUC8OIornqDiYMizI/OU02qjfX96yewauUWAEeYJanWVBqpeThR2+Cb+JP6qpL2z5dFErYDKdudfntvjM88oDimbgd4YwAUES933zik1/D+78v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTNuF9Szb8bc/AamRELv23yFMoHBO7CYg0goWr/BMnOLby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMA/6geAhKQYfVg0Him5cM+GQudJ4tjOm0/G8MS9PnKJEFTQCciqpNfgCJkOivzq3FPkJK4xKvxsCfYmJTxiaHl/mX464GuAKflLtWFFFLAuA0tDoOZ6a/78bAQs88UG+wSNWNrcAyGzv5l+OuBrgCnL7n3mFDlx+KMyy9ofvlbCVlMoCCcErT3Yu5mMV9FnqQaeSEc5Yud19epfUFxPX1+l5VLDx54rUHAWCwd+65pMJTK09xkZJv1pfANeIcqZovDHzwZbJ7YCxCpeKsIVteVv9281ooBjDYrojOorBNgIgL0kEjdIIoXqDXxlkXGyt8S1F+P0jKq1WxLQlCoz/0vnlHUuVejHZnyMdS4CxnscS+595hQ5cfiSqIV4oOEBmQvX5QLQu0dPSKFcyjTCHX8qDXxlkXGyt8S1F+P0jKq1WLOBTMMHIWdq9XxkihgWvjyMdS4CxnscS+595hQ5cfiAqWdX1VO3zMvX5QLQu0dPXNSxNSxDBqqqDXxlkXGyt+ZQ8ZfcClobgL0kEjdIIoXqDXxlkXGyt/c9CSVHsOFPvwBWM7j/ULR11V4LnVpr6FUSwL2N+vqSBhrvt/y+YAdjfuoxOiR3gug8SmUhhzy+eFPexG1VS3coIMZfzZDR4DAWCwd+65pMP4ndrcguBFs4Qq8qes9OGxBlCTU+I4fJ0yUbN2UnoZAOvzm46oTw3G2Wc5osDyA867BGJabWD8pCbDw+IJ1H7GA7xJGOWnqZd33zik1/D+78v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCw6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcmpGPxRfAM1oTHEWGToKb366sQifaTGPokSmKLxqdSyNINHup1QjRMc6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcizDohe2/x55vf/d5mdk0fTZUAcA948qwwsie52kK+VirCWUbDj7YftnBj5okswDWqANX0XBTHjAN3nukQuP5K8YKYvSvC3NekNqfLrFo1S0A+Oc1Npth6+IQUJKyK6p0CT7q5G4g1fj+OSEWtOk2Hkt3RFoJP9wkAPjnNTabYevJqWbEMG9PrK6WFEGdh5P7HhjxeqVii0rKqLBu3yOMdp+Konn04o6AB8gtxiLTTHiB7N50MLSGKuPibpgnmJHKJkLg62wnfIEIR++j0NQlwnDHzwZbJ7YC/KT1FckFk5uqDXxlkXGyt+INEOPKg8R3FAkSuU96ebivkiE3cSYPus67OyGdcqUIWu14ZN0Jk67RIoLn9egg/Agg5X3i7JF+MfOv84W5tkyjwW6z7kL98VoVwGCkBX7dk4mo5XYWWmWAf1sDL6Ym0pUffwU56Pib+UwWAw0XygUq5HTmOMN83eoNfGWRcbK3xLUX4/SMqrVNk8nAh8ePrThT3sRtVUt3KCDGX82Q0eAwFgsHfuuaTAVBFNCDVDPUEoM1hUKn/jV5Z846Wr2vs3yMdS4CxnscS+595hQ5cfiAqWdX1VO3zNIUNHh8lhGscChmRdotHZeK+lIboRweD9c4sUPyiMvv+Asb/XcWPWF+fu3S3MoLDBhfQeIFI3IYk8OfSPAC2B3HiXY1hK7xIm+SayPXrle5CvpSG6EcHg/YX0HiBSNyGKr7KKSO4D4uh4l2NYSu8SJYLH8acWtEfYr6UhuhHB4P2F9B4gUjchiImsZrxj6swMeJdjWErvEif1C4hPnhDVdK+lIboRweD9hfQeIFI3IYux6tfF0RwGJHiXY1hK7xInAoZkXaLR2XujS7z5XwI5Gl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGbj5RcgwgjQhfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHggs0U9Q3CXdvaxYs6P9WHd6ZlZ1kXMyJD+Z1q6OOCtTdKnc/75K1rPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHsLvgEziwlwCxk5s5HEOA0Iftd2xSE13D2SQjd+5XpjLygrXTM0EsBIK9FbjwhEdlEjboyxTc6gsKTxcCKMqql9yZ5m3LYOxnSW7iwRLiwVUYa77f8vmAHY4JAYSRk1untgvkUh8wn6345IRa06TYeS3dEWgk/3CQA+Oc1Npth68mpZsQwb0+srpYUQZ2Hk/seGPF6pWKLSsqosG7fI4x2n4qiefTijoAHyC3GItNMeIHs3nQwtIYq4+JumCeYkcomQuDrbCd8gQhH76PQ1CXCcMfPBlsntgLMyNepbGO33uoNfGWRcbK34g0Q48qDxHcUCRK5T3p5uJz0uf+XOv1i+w2DA9K74IQOZHf678KxglEiguf16CD8CCDlfeLskX4x86/zhbm2TKPBbrPuQv3xWhXAYKQFft2TiajldhZaZYB/WwMvpibSlR9/BTno+JvBkSCdbsx1i7AfI0CGcsGCL/dvNaKAYw2lXeHI7I2QVvfrSm7gUc/HTvG39hDyodsh5++F3Y07N+oNfGWRcbK3xLUX4/SMqrVYs4FMwwchZ00VnrU9qUXqZdCcH00Nt6SGGu+3/L5gB1sR6DJqCUVyqZoQQMns0zM/mnqnDyu4DQ9IbBbSIoN5MBYLB37rmkwVBRdCi75HEfNReFosymZhMBYLB37rmkw/id2tyC4EWxbKJWxmn4hdH1bt9M4/BF9f0GqYj830HvAWCwd+65pMP4ndrcguBFsLfI0uWYAqiN9W7fTOPwRfaCDGX82Q0eAwFgsHfuuaTD+J3a3ILgRbI3uG4hTLmynfVu30zj8EX0stElpEoSg3cBYLB37rmkw/id2tyC4EWwSwjPtf0QyH31bt9M4/BF9OoiULZgjuwqChav8Eyc4tvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyl5bd2XULCrNdHp187/2d+Tm8NYOhjtcB6z8v+GH0Qel2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGbIrYnIgvY8cKasjIyYzneg8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTipZnrl0m6dDpDnXpz9TWLwsie52kK+VirCWUbDj7Yfsu0jM+QjWNPzg0pVXL3SacEjVja3AMhs7+Zfjrga4Apw8G5+oIPR9YNIqN+VbMSfVg9bH9EKlyyDveSImX13A0X+xkqAgzksGXIk1JlZdjcqlT71QxNftDiDRDjyoPEdx6eMGG0US47DssUGdd2NvHElde5mwLGJSJwEzYb4hXIWSWbTIsYUSQcuTCtH6/xJKzxO7EBtu+KD8BqKRjeRUO9chZ+uWFC7ZjK4O4odb+ZFKIRGvlQX5Ks8TuxAbbvig/AaikY3kVDpNFBIknP8IKYyuDuKHW/mRgNfJ+AtFEM7PE7sQG274oPwGopGN5FQ52XijdKPPJ12Mrg7ih1v5kgDhD/kl1NPKzxO7EBtu+KD8BqKRjeRUOnqG0tgT6S0ZjK4O4odb+ZLxPKmMaUTNBs8TuxAbbvig/AaikY3kVDlzrUIanGW0GYyuDuKHW/mR/o2VDPXWZN7PE7sQG274oPwGopGN5FQ4X2SAXK4uKfGMrg7ih1v5ki9ldDhgVX+WzxO7EBtu+KD8BqKRjeRUOA8i0PM2hSBhjK4O4odb+ZOXeoSx42L/Ls8TuxAbbvig/AaikY3kVDnlgyZUXiGMXYyuDuKHW/mQ4LAfg4HKCR7PE7sQG274ob4w+NSYBw06432m651I1RRr71KqWXu7/OSEwuPGpNfXVvcg86NDujS+595hQ5cfiOBc9sEygL1rGL8Fyfno8VBW/dfclmuM5b4w+NSYBw06RpAOMPTBZtJGMZSUNb0n0C7GLM/ZtRwGzxO7EBtu+KBW/dfclmuM5JOBXqtLt38sIsJMAqh2q1U/E5ugctI/kNRjP9Z260P2CxfZwGW1tTJeq9wko2zl+p+JsQGSnruDDz5/Wn/KoAKxOIZLHiZa9C09wc74eqGb2h2T0pTfGk1zixQ/KIy+/4Cxv9dxY9YX5+7dLcygsMNz0JJUew4U+X6maz8Mf8VxEf0q9KY5+N0p+eaQ/bo0WZjySmeLaPsoMHZNkdaymPUPqIEohs3X+0xZE5fRBa86QmpkzAd2XSPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8WlsSdjcKS3mUPGX3ApaG4C9JBI3SCKF9DnumNqBSSR1IybwRAazvM0CgXJi6F1M9CSS4sJ3uDo0Oe6Y2oFJJEc1hCg9j6TVzQKBcmLoXUzkE1XCQUBUWSTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHSQAYMCrv5UCV5knami9wwVVRwMjhBTMPcMdlhAEq5i2rC+8KvwcIAjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRy5elrM4Q2ayGFsfYaeB/EKeprxooDEabJJSIObhLSGyH3ru+USttpRhqonAABXb0iXh44Eru+G2/DFdE/EjAVqI/DJWHKiE741Hti/p67mk/ZdrxFpecIxzS3acJDvgW8vgL4AaErRAspUXp5yCcn5nSDCgXY/oNQu2TXWro5hPI04YFhHx3eU+3o1N5NXNK2C9UxHq3ksiZQQ2QUj3wkuZC4vBtpP5M4CQ2AdkZql9BwfFE3jEDu6zoMML3hsWFLW514rIS+wWs9R5QN+j+vQrLJB6mLJf43JMtecPzE24s+3wUp4AHlaZpBVhazntdDFXX9LD/Bi6+Y0lrrlWmnAAjlLv2k+LR0YOS3/iuq/EOe3z8Z+NJTbJlsCP0ORw3qW+PLWHJwcdsoKmVcgLNIxa1EyOt5Iwx65ynoFzf9Z5BKohXig4QGZCMrIZftmZwZq9o9aVWJm2SjwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+yerg4Gueif9NMX6BQpoOXj3gy+nTaA/6+oBVDtU0pbPWGHeXwGopL7ZXYS/bWi5dpwEU0yBqKU7bGXA4UOqbPhxYsCesoUgArAlCJBb+ant+uiprTRbSt9CjztA2FYcnyZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4kqiFeKDhAZk50bbJiIZC3fp3Xm9o85cSWGB2S+nN5OwaC6ZoYBlhyOkf6Jhc3anloUQuydf9eX6i6RLPDkLTF81UQorfXi8zuCVCIUR8otWwFgsHfuuaTAPyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoMCqmU3dxUTNT8BqKRjeRUOrjj9jzto3EnYZ0lFbE7wxQE++nePNBF98Fb6vqF5Z5dl5iu8XGxV42bR8pD1pPHUz3KYQK/+XgdgKfQ2xeWmQwgNj5V3QggYwFgsHfuuaTAnenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvhUEU0INUM9QfNZMEwKWW+W4ugDXg6fOP4vk4FH6kl8smRJ/giieFV8sRcaZ+A7MsykY9XAgGVFZ4c5mCtfmR3P0eUYOHu6/+Ddz791M+kWQQBvxHxJf6pBBmX7RArBPiKuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSE7UK/CN/hKcMcNYmiY3mmC0/SkN6W5/Rlf3MoKzgYy6T15zrifrqviw5b3DwFQVuWtLVNc5sYlOk1Q1lZpaXp51gr0IgOLLNzUb5x+EX7UB/mHQCpvWKdtYOIDpsmIDv/hoiL8D6lHOMZaJukqSckHL8ElX1S2IiXxpZJSDjlAnfo+0X2FfV8HDFR0jIQgdxPeu75RK22lGIkkZTo4MPWNeHjgSu74bb8MV0T8SMBWoj8MlYcqITvgxCL96r80dw0bnpYuXZcjIwFgsHfuuaTC+AvgBoStECylRennIJyfmdIMKBdj+g1C7ZNdaujmE8qBJP3vZnYqhnyARpKu40sahE3pMwMRX1LtyXD2M7eK7x+GxllU3P/fYZ0lFbE7wxQE++nePNBF9Grm+OxYrv7Zl5iu8XGxV42bR8pD1pPHUz3KYQK/+XgdpuOm/7DNMOv5h0Aqb1inbwFgsHfuuaTAnenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvp64K/wQvn7OCrco3HI4z+yUytPcZGSb9fBqj3YRN+QDHJ7TLaX4iiKe3z8Z+NJTbLzRxRxS5BEWM7kKG2fKh0coKmVcgLNIxa1EyOt5Iwx65ynoFzf9Z5AFfeM8YuVC/8BYLB37rmkwq9o9aVWJm2SjwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+yXhy18Cu5/VYIM+5XEPsCiIKjNnhfsJIKZC4OtsJ3yBKF4Ix21eYhDtP0pDeluf0ZX9zKCs4GMuhQAORpidNECsOW9w8BUFblrS1TXObGJTpNUNZWaWl6ePSncbD5m70AQBPDgMRNkq8BYLB37rmkwWDiA6bJiA7/4aIi/A+pRzjGWibpKknJBy/BJV9UtiIlbiYvUXNVjIoxRqGhbhr1Rr81RUQ0sYayxeSmMOxMQeR2JkK4I6MzW2GdJRWxO8MUBPvp3jzQRfQOoESseypMPZeYrvFxsVeNm0fKQ9aTx1M9ymECv/l4HAvx2yCObatv+YdAKm9Yp28BYLB37rmkwJ3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb6euCv8EL5+zgq3KNxyOM/slMrT3GRkm/XTnu2JViQJ/KPfwPl5wLvgqAVQ7VNKWz1hh3l8BqKS+wKAWdVSLp0RcBFNMgailO2xlwOFDqmz4cWLAnrKFIAKWczVwYft56QHxyhKVrVgN7Kny9Tj5a+tmWM7sg7m9pItp3y7fmTZdcVSVVRNYpozshsyfOCZT+KhdiJRJAXBnTgXPbBMoC9ahJwYO9IupbHp3Xm9o85cSWGB2S+nN5OwpnTRQjn6Oomkf6Jhc3anloUQuydf9eX6i6RLPDkLTF/ewfAsmrBwhOtGkCxH12jdnV1EDmpa2mAPyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoMCqmU3dxUTNRW/dfclmuM5b4w+NSYBw05kppt9fudVEcGOdbJ9JQtTmh+mh+WA8dAwbSyI1QUsknxNGZ5uda16A17osQw6zMZzP8KVopQKxuES9FdXCwi/nt3//eJ5+piKxVxRsyUdOQWJ3QAeSDW465Rdkf0b3L0BPvp3jzQRfXfhybcFR0Ie9WDQeKblwz7i8NIFro3BbxpcOkpH2V6WOc+MEglnTSDG7PnujmCVqNzVFe74BKp+wFgsHfuuaTDAWCwd+65pMFY5PTEMo3z5OT24kS10JBwJO9N8m1pi2K4bMLwhaiwrhzDEDON2nhegDV9FwUx4wLPy6PHnEFfDU9rzOtALlfqMD46cGrXy4pN8KFQC9eRln+uryGH3e/DicC2St6UXG7GTmzkcQ4DQ7EYIPgTc3rujAxInul5e78BYLB37rmkwwFgsHfuuaTBXaeIhBs1ltqpNS6+zNLwMAuZaNps9FxDvFxcTExeX7YDocvGCwDw4/4EhCkOfq7GoBVDtU0pbPbeRV9UujD74DF+xfZy4GZrc9ruZiEr/fwyGbs4z3x5eGl5hxdZPJpzKp+h9ynZxFaMDEie6Xl7vwFgsHfuuaTDAWCwd+65pMFdp4iEGzWW2QEl4tQOBzxL1h2+Z+wg/MWS3QgPeTtljuR79iektI/SCvRW48IRHZRI26MsU3OoLiVkb1rzZyZlWOT0xDKN8+Tk9uJEtdCQcCTvTfJtaYtgsrbAKf3b1TocwxAzjdp4XoA1fRcFMeMAhBfKX2z//SWMRYWRXjusewFgsHfuuaTDAWCwd+65pMELn3320Md3SXeUu8x5aEW0+45kjOjRlyOB7qWn4ISo450bN41F+Hcp+wYmxjDxeIcBYLB37rmkwwFgsHfuuaTDu4I7AKSoyZbngJsMhIul2mPh/pS7t/k0kEVoPbZayfgR+XeTW+bH594APv36K8abkp9bs8M+BjldM/Fl1JARPwFgsHfuuaTDAWCwd+65pMIm6r6AYR8tqMbUd0Pmm2sB7jt68uaHSWSxVFqDyYofy0aDZa8pdxpCg+rx1i9cEOFHIEqttIaW2YxFhZFeO6x7AWCwd+65pMMBYLB37rmkwQufffbQx3dJzUTVDaWp20ZwZ1ocmjguAPT8iJItjm/hyKPh5FXIC6YQcor8g32Phc80LFW5uoC/2QJjRRYiWwsBYLB37rmkwwFgsHfuuaTDJ1sawggAx/Vj5ABPnt5iWVO/qcvwCi9VWOT0xDKN8+Tk9uJEtdCQce7D8wIYZP24JyYtPBHDQSzGfUzmQkKcXDJ9LeExL72R/x+iCgxSc9pdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxmam7iEwbcIGsNfP/1CBud8UqGxIKRu9TPcLpMDZXOk/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwt3gjIEtmkGJUn/JVTdmWYH6MQhTMtwAUK7cvUi1o/TGoQ1R4UUhLal0nUbGM+SWQTJ5r1xzfDXClC+R9yUfoJ0Gb8Ye9mOhQPlT58qADgnayba61mL7BzZ2TkZnHbsHBPxbmei8NO38d0W4BD0aFKU5lnjpedoRzAAyrlX0gor6tNzUEBQoLQ8H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3LT0/yG2IDtrlZ8IPyDLuv+l9xhXNxWN2T7/oIFKmhD71zhlzDSb1zNzaJy93Vs0Uueqp97NbplmPQQkgisl8tYFr+MZcxVHaX0mUNa8pVb7RtZNGyzZJmeUUQ57P2dZ/A8CkU8l9zSwvwJH7XcHtdGsySS4glDgbXyY4p3wSQhwvwJH7XcHtcWjMJsg0T8KCNs9/cmJsZL7wr+i+5ntM0Ug4fO5ji+3/1g/k05mQJfnFRdSxayBnBSbaDc4Qlm51h5E0gkpomTYDx0oL8iJkpmAmFR3LKaecIKQH9xapKWH4XBOP/gst8kJwkoFIaeMl4JAwcpRs2wpWqh0Oh2IWUqosG7fI4x2ji1OZ51LoAHMCAsaLkc9sMgi9P5Q05ExDveSImX13A0TlFdMeLqVB9xX2xf0wa4olMzMTd2VbLAHYNbLmfROv9Z+gm9tSVzWXXXGqe/hNQ3XgkDBylGzbClaqHQ6HYhZQtDrqfEpe5xOuzshnXKlCF+KZ2cCDojUsEfppvqcUz6AavDmDTROJGINEOPKg8R3LF5KYw7ExB5hdB8abv1G8KUzsVX+qjJ2cFhRLHtr5z2lMrT3GRkm/Uudhg6xCrchw3Ja/XBIZDOAWDQJ3KBpIOfoAOLnMoIH8MfPBlsntgLEKl4qwhW15VxX2xf0wa4olMzMTd2VbLANuF9Szb8bc8riyPp1ahjhotDm2SkoC7m+fu3S3MoLDAVBFNCDVDPUJmLH3q+TbiZHdtxg6oOGCMomfIY+Y3JZuHDJoDEt9A9p3F2/KZDZS09R5QN+j+vQnOEjQD1hbNni0kWLnusckK6maR0RWksW21F32Il+s4UEtRfj9IyqtWBDWipwpEh24t9mDkl+tWoMZPML60V2LXsY21T3uRMTZ+gA4ucyggfPwGopGN5FQ6MDrbvB35M7J7z2bM2B/fLTkGSJu/s69jC4OEyxUpTDwH9bAy+mJtKaU+7FrLqupQnUCoE+R7cwXVgpvDe2lFKHEcuJ+RvSwZzysUlAo8iA2xHoMmoJRXKvKZbIPK2IYXJUIcMHf+R7A+w5CPuIzPya9CKQlY8TsIdg1suZ9E6/wKlnV9VTt8zL8StHlHjq9o1Zicz6VVMhCi+G04JfRlAVFYclhD8d4eVd4cjsjZBWzUb5x+EX7UB/zdjE2h1RvcRaygtE5naOViCACHbNjEqs6bgY2Nlcm3pG4jXwUtOiJgAg9RzrwwGtP/8iyWTRROnC3EK7+Fb/MbXe09SFZZkTCIv7ttHc26HiNFTRLviWFiCACHbNjEqs6bgY2Nlcm3+J3a3ILgRbO6hN6M8acG5uQ6xY9qr2znIlqyTjvEGuOHDJoDEt9A9akY/FF8AzWjIyiRDxfOaj9HyPNWoMs6xlmu432Q0Y6RxX2xf0wa4olMzMTd2VbLAHYNbLmfROv+u7Lc9MLOn7MEfppvqcUz6AavDmDTROJEPLQj5V8ycxnFfbF/TBriizc2icvd1bNH+BL4a1d7nnRxHLifkb0sGc8rFJQKPIgPE9j9QGxx9qNWgCIHX+u9YAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4eNmlGfQjyG1kJB9PRMhOAPJeg+iExCMrmtHnTxlMad0alyDWxEiU8Ja9CKQlY8TsI6Sgfx+TrittdFGhSV2OM9cc7WB6YSrzjrhFTlXHuZ/8NSDFCecw87tWd5+e4mmY89y/XjWEUzjGxuDd1zeOjw5I4IXBo4g2Eo36jxjcHPCwmjeAwihDl3yCvi7dFzoYHFOpZ08/IJvg2z5EyYI0PSQfXQgsgzo8iy222i2BIpcpTOxVf6qMnZI4vTKyHBGc+OMzCZJIUMn0amOwvdTgylB6zgflin7TzExfu4fqaoh5nPgLuZafO5+lFDCpo0se6APeXNQ8AQrB4FDevtDiVUFIjp1DOt+yfhBOZPNhBTGByhChvTvpUuwgpAf3FqkpYUiOnUM637J8TeLJZmqX4+sDrAXOB2kKidGlESu52O3o9ryFAi7Yx2WIIAIds2MSryTKIkUcCMHWGiJIyLcU1+paphVYGdTD6vh48WgeAe+K0edPGUxp3RqXINbESJTwlr0IpCVjxOwivkwtmFLeT24SrKfn/kqlL2DAG9vKlzX5TOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMP50r/6zZg8QlwFdadm3+LCz3NCN+vBqM4pWqh0Oh2IWUr5MLZhS3k9qA6L7eqtSNLFLZSiKZsDMSsPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPRSI6dQzrfsn1kuajj7CqGvtxHjj6KjcwzA7z0L52nuKAi5nyDP1E0Dak5WXwo7DXGvQikJWPE7CK+TC2YUt5Pbl1Zp261EHWioWJcJb2u9XLXL0PvW2kMVTNm7vlhR09Sk5l1lCE1iF4cMmgMS30D0UiOnUM637J9ZLmo4+wqhrOSEwuPGpNfVuNVFDdcWgDJ64K/wQvn7OuRh3QlVe8E7C4OEyxUpTDzLGV+OpY5jMcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPYGK9eVAshnMBqZEQu/bfIGV8705rZE15dngkk061zcZdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmhYAIjKQGxpdNcYYB1rrXDjR7x7YVGOZYjnCw3frpxtWA6HLxgsA8OF2eCSTTrXNxDqFeXIjVfUOP4r3tD8ykX0WyOTE2UwNchBdE73GNEXhycn0fczLPWCqiwbt8jjHafiqJ59OKOgAfILcYi00x4gezedDC0hirpdntYsoL4Pu7clw9jO3iu0UsXHSJTh9fwx88GWye2AtXmM/1PwQfAag18ZZFxsrflMrT3GRkm/Xwao92ETfkA75IhN3EmD7rOuzshnXKlCFEfvRNXzByUY+JumCeYkcomQuDrbCd8gSa0FkKFf/PUTssUGdd2NvHElde5mwLGJToOI/l4KNd8Yg0Q48qDxHcsXkpjDsTEHmdSONssUdyRcMfPBlsntgLSsnTb+gkzYu/3bzWigGMNjssUGdd2NvHElde5mwLGJQ6XaNLBsMOW1n6Cb21JXNZr7G/jwLhfcWoNfGWRcbK3+kbiNfBS06I8RkzQE/Tjwgjy/wmmqpxBgH9bAy+mJtK2Xa8RaXnCMf0OvMHvDYg/D1HlA36P69CUzwCUlzmNrOVd4cjsjZBW8N9WS0N3Ar0Jj0S8EAQi+YI5S79pPi0dELQhhfkIQJ6EtRfj9IyqtWBDWipwpEh2xbMZAwlNQRlNOFUfUNORDS/3bzWigGMNmxHoMmoJRXKlg4eev4gKlOGQ9GMRcfna8TV49Rk/S1FqDXxlkXGyt8VBFNCDVDPUCdWzbguOJpWbEegyaglFcpdsZsWKUWNcrPE7sQG274oPwGopGN5FQ59UmWGtPgYzhUEU0INUM9Q04AMuUKyfEYvufeYUOXH4gKlnV9VTt8zbKvuBcrZRNY/AaikY3kVDrtOYmE/873gT1nZXCU9vI1O2vpvaNnlSxSt7apcRCOKAqWdX1VO3zP/HNN5W3do95YY6aD0XR4zw4cYOmpNXIaJtYcgU9kSUIo9UZjnVVXWjfuoxOiR3gvz9TTqCcIX6o37qMTokd4LatZfxrEvPYZmPJKZ4to+ygwdk2R1rKY9fx529Q/hxwQMHZNkdaymPfBdPgDYCdLDIHo30Cu57AfeHD/Xt+YMt361ITAcx75EwdHHEfVc8flsVgFds90Qye6gnuh/ZnB5v9281ooBjDZ00pwpiy/KVzFtSD/oT5P8Bt0iTwmsIN6cttEH0AG408FOlKqDpMwodyvNX5JepqE5aSfWa6ks+7Uw8m9dq1DWP77b6RQp493TfvYTFfYPPGHAPT7xp+aotGwLZityvxOV9Q7cUMjDZf2h1Zn893TC60aQLEfXaN1rkWU1DDwtGcFOlKqDpMwo5pNyqlkQKKfTN/rfMp2JDt+ny0FveNwYKhYlwlva71cEc6Ble9y2EVnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTQxLD92or0ceXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZtFbib0IxNoKqLwSlHt4MeIG88hJpnhuTJdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmjlN8DtvWK/k8nj5HI2hxgULON7OnVU7m0fFnSRUzvp2MfiIt7lB+sEFCIQkGbbCx7biLDAQ2AyJP32Qsz4x1Zg6OyG6bnoLJ5S7VhRRSwLhnppnAJKCwxgBAaM/z24ni2T4/OyE/PSL6UUMKmjSx7oA95c1DwBCsY4a7EVtF4fPlLtWFFFLAuIV/ZdH5vFOFV3ThbjCmjuS2fZUPm+VOMLrpgBNihazQje0nSLGFZm24dN9TtPW7ZQ6hXlyI1X1Dj+K97Q/MpF9FsjkxNlMDXEHcVqgmeypWSE+J4reqvrTqqbdcy/jB1ialmxDBvT6yEZKSlycncwrS5B+HQuLItS+595hQ5cfimn3Z7mXQWQkffdSuUY3eUJHagvye4VbPYvQurHilbHUqosG7fI4x2uQ8uV/iK4s0kxGQ5DlU5Nw63KRBzNiNf58A84lnmGTMQIQAkkXI9AvOUe32hDivHrEddF643SlElMjKTBbv4Pu6qnClgm/kvfDb8ejw1EdjL7n3mFDlx+IVaVVg1Df/hPoRoal+XLywDVC61irCVcFFsjkxNlMDXEN+ruTgp9AKiOD+dc7r1Q3ASdLvMqoB3e6iqgo/5TZNsLgoSeYubrTwK1m3PL/wf5pb1tIBC0VVYNTLRsAZTMgqyzifN2olEspzTMIxSnr12DJ/p/4Tr3u+i47LNHaWl2UTyWps7apmGnxmMQCxj34ntQyxMoEi6r/dvNaKAYw21Fnqz9W3OdyV5knami9wwSuQjVJvX3zIyaBG5lFC15bSA98b+XLS7dOjr1vmDRKA7Ili+TO6kwDJoEbmUULXltSrNFnjOj4OsKnWW73hyQ7caUoX8x86rmY8kpni2j7KwCQsxpmpB15WdCXZjtZA6n7vJk4g6c34qDXxlkXGyt/jYgY1I8DT8aWqYVWBnUw+rx6WIJXkULgi+PxZxyAsvy+595hQ5cfizyX9SCyjrO/Kc0zCMUp69Y1hODlkb3GoFHB1ztPTFxTuoqoKP+U2TYgNIy7Xb5Q6e2jEewmcIsBTwfp10y41a3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR8WFYBi3y++fg8hCJk/L6jM+MMucS0eT2KokqiNWOGtA4jey/TkwTw3y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR8PFnrR0k6rngXuQoZbZBJp0tisKfj76OPBwnZcmTAaAUUsG1UV4mxH6UUMKmjSx7t4POnGkg9Q2y0YT4BhZbefQq6vvWj9+6Kg18ZZFxsrfWLfuNP5FCVhn+djsM4CPbbPE7sQG274oGnkhHOWLndfXqX1BcT19fpeVSw8eeK1BRN7coAtNOaQ05EtuKTzyxrCgt/GByzsKL7n3mFDlx+L4dxnSTBlBYCf07MPu4p6b4++p9PuNtveBe5ChltkEmkvLh2Lc3/Fc/u8GQ7ttLbw9sRnqdohw/rCp1lu94ckO3GlKF/MfOq4vufeYUOXH4nvqzdifKM1tCSIDT+JAzFO/3bzWigGMNsT2P1AbHH2o944k6CUUc4wwyEQDWnQBo6g18ZZFxsrfSPZCjBZnXw3To69b5g0SgGgtTHbsyiD7YNTLRsAZTMg9TpLdnKt3pXAV1p2bf4sLiJP9+dI2nl95apJj9XwnyKw6Vv2stUef5MenSScGPQZ8gPwsN5c8Kgf7sll72AjeeGGkxskoeYewphO9sWFUSt6vbb68OjtvRN7coAtNOaT543+EFUhtMycNF6Xh9oRrcICN93vFAvZg1MtGwBlMyBW/dfclmuM5JOBXqtLt38vfp8tBb3jcGCPssU9uVOgOiJP9+dI2nl9cF9VXEWYWH+aTcqpZECinNWgrYbbx1WLfp8tBb3jcGCoWJcJb2u9XIuZD0JykHlVg1MtGwBlMyBW/dfclmuM5b4w+NSYBw06432m651I1RaF2IlEkBcGdOBc9sEygL1o8xiSrsOp/iZdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmGZtznhBvObu+3Rbbl6sYhMmJu5D3fjPc5mw8QDXyQrEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvDvs4X13is5a+X2U2Sr4h2tfpPQ2kXFtYhzzdEPSJT5a+7grw2Uuih50Nrz9FNAQEPr2LbsPFQc/85hXRHi13qvfqYTuVYKVl0u4Abt8zT7TWUWgnEYxS+1BOE2i+qcLAtG5bhd9QY2Xvk6EmRLo0UqT/lnpuvqm3EncUfC4oj29m0sv7LJtanH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LvOELWtFYaJAxkL91+oXh1AAHKLhj4L3RjWp4X/fEthWNsdqxvyc0pvvhO+I7b9wou5ATpgb+4aq6ErXIdZ7wR5yW6ej+suMWMlqR6Ss0rWpS39lrM0Fjh+0bWTRss2SZ7boMQ9kCHfktVnK7ut7KplucMDlUgErFxD3rSogWUrZOuWzVkkYHV3wSA0ahigD6Tzr/ZBmu0bA0b9+1iilocrWbOUYtVbAK9K/J6mhZiP6saPcFSAULr69pzNU3Tj8arjF66sn8qZ3sY21T3uRMTRKar2s4P+7y1fJdfYoxciEMn0t4TEvvZI35flCh5vUV7uaXK1Q0dtFO/f05z7HQJfA0VF+rieLiPSX+5s87cFdwukwNlc6T+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3eCMgS2aQYlSf8lVN2ZZgfoxCFMy3ABQrty9SLWj9MahDVHhRSEtqXSdRsYz5JZBMnmvXHN8NcKUL5H3JR+gnQZvxh72Y6FA+VPnyoAOCdrJtrrWYvsHNmJtgJcuO1QdUcC9mrSQeEK7G3TEucUUtqd9YSz6jzRsQzthX4NBEs0AMq5V9IKK+rTc1BAUKC0PB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwty09P8htiA7a5WfCD8gy7r/pfcYVzcVjdk+/6CBSpoQ+9c4Zcw0m9czc2icvd1bNFLnqqfezW6ZZj0EJIIrJfLWBa/jGXMVR2l9JlDWvKVW+0bWTRss2SZnlFEOez9nWfwPApFPJfc0sL8CR+13B7XRrMkkuIJQ4G18mOKd8EkIcL8CR+13B7XLlk89pyoh1QKcIdUpPLmJa56w8vceuNo4F4nVa8gglKC4M2ldNdvvV5KwHOLh+21qcDEz+c0ePOLK/sUI46V8YdjS8RXNV4pGindyFNVcwHLUIS46No9mzCUn/khgvDJq+9yLK/bVb8pvPZIbEufcGnflm2GWPztaDHA85r5sJm5fcLCHADv2jAgLGi5HPbDIIvT+UNORMQ73kiJl9dwNPl0uiV+r/FjwR+mm+pxTPoBq8OYNNE4kYg0Q48qDxHc4iaT6/CfvQYwICxouRz2wyCL0/lDTkTEK6IzqKwTYCIC9JBI3SCKF4DNUCqI9DySWQ6MbX8gbuQVBFNCDVDPUKM1l0e/dWYvXgkDBylGzbClaqHQ6HYhZQH9bAy+mJtKRvgfyGsBOHiLfZg5JfrVqDGTzC+tFdi17GNtU97kTE2foAOLnMoIHz8BqKRjeRUOc4SNAPWFs2eLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhSZQ8ZfcClobgL0kEjdIIoXMucqJyHgRfI6Sgfx+Tritgwdk2R1rKY96mycOFNXsoMgZH/Prfb6w6VqodDodiFlYX0HiBSNyGJCwH/1ob0ps6YNRCoV/0fFnrgr/BC+fs5OQZIm7+zr2MLg4TLFSlMPYX0HiBSNyGKf2Heakqlos6YNRCoV/0fFi0kWLnusckK6maR0RWksW+zfWsfwbxlzfkxUkNGCvYC18hkiP87ekmOO37jkgFi5zRzg0OEb2CI9KaVxMDNcjFrgSNBvfq0OZf11sV/DEVQDa4kJbwkYlvbzb1lLp7PunKHfwMRrctgB2E5tBALqlk3Ptiefzb1PoSK0HM6L9mKCKTvWZGskVet9eWbiHM1yewPNu32f/eGo9dkPDMlP0jAngQRNwEssM834MV6TY9v1JtlJcy5d8des3WPu4Krnv3T+/Q7PTTnsK8azPaeTkABfKVnhNsPIhFirMnppqO//d08rqXGXmEW2fhbObAR4bzSnnY2x+Yp4BhY7c6QzjPk8PMF1R2mfOyYrnOJScS4Ya77f8vmAHcBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwaPuY0ytJXcySg1SyullYXXGYp0zPErq9eAYWO3OkM4z5PDzBdUdpn+7jKr74ViyVhfo74iCpZsk6MWLd6UpJ7OEZWXg5HIFIRBEBAAoExafML8H3LkfDQYzD3wu+7NmPzF2hxrsUvM6hX4d2A5E09s8cNhpUJS1Zxj2xuG2LhpYfAajdaw5w8QBfKVnhNsPI+gshURdqOAnXSXFVIez/dFLq7MkKvgJaRNPy8skmeof/d08rqXGXmEW2fhbObAR4FDV6GVp4/5FyukvJ0+dhsEjC3ppNPqoTs2S83Bnryq19KBwt6lJD4MkdbbcYtd+SRV+i6eojCUJk64UZfDY39vqQ+hWjUfbwJwKbmEPoM8SSN/EuPlxUHgPVsgh3Usnguksy08lWUwVGLlxj2xmhcW3gjXOEok0S/OhIj0EhripiYAEqiFN1AvFoG5ZSuGPqCErNTdvdysljjt+45IBYuRVzQSmWmZlSQuplHocf5yYg8uqjQXuUidqaSN1t9yqBmYE/UXFCwAqjCWgfZ262/Ztd1mZMstlcC9oKjZhmr9QOzKo0Xu8noCjj+QYG2XPPnuj2nkTy9e2LcIkEMQKv+fpVTXQbzA90jMPfC77s2Y+cn3x0dVFB3kGm6u4OelGMNrBKvbSWGzj6iRtWQCv+LQUlqpEcmZ8nt2gndgCcCtgwJ4EETcBLLNTApZCDPiz2gvDzF9jLR6zpHCFgEF9jCJqOfUlpK0V+FQRTQg1Qz1CuXpj++ES6Sy0ZgNEGYsaRLbgcJk9oxelF3UsQto3MJFK+mLs1oChWDrRzo/JitRdB/UCBUWZncGREETk0GkowQ8IRKH16JozFhL8CoTHuerPhmr+Q3Q/WvfleZEDxrLHUS1KTpfKmbIzD3wu+7NmPcKiq3FWcSYmVONf5mDWVfAS1GUT/Suh2kd3rXe3ilhk/AaikY3kVDgTcJnJ/jBGkkg4zGKjvv/obqH3qqgQ2LeRo1Ob49F/c6RwhYBBfYwiajn1JaStFfv4ndrcguBFs44hnMX4wIfxJGyiU+VvebsRP+C/1wxb15ZYdkWGV8rjhMf1Ln8wqS790/v0Oz005oTxY4dMToqfJ8kit+cIxLPvExV7KRT08tJK+QoSfhG+FdixWTs9WPoEGC/GguvaFzmP0X2jn7KB+RwOjSEzxFcrWEA3SqQuEzFtgQS+9kzZtdCwTRMZsej8+JvQ8lPkY9bMpVXuOVT9YggAh2zYxKvJMoiRRwIwd5CMOzvxG0FGjw8gZK0E0BpbwvYc4DSbFqOj0f8ciNYT/fCB9ZwjXIzSgfDBP+my+ICPNTACKZZ/sY21T3uRMTZxqJIHSnBRTkAF/GUCkG+aJrvqYPJMS5Zu0avgPbwcJgQYL8aC69oUo7JHWSEB+p/Um2UlzLl3xQEECCmIQDytr0IpCVjxOwrSSvkKEn4RvhXYsVk7PVj40pQm4AXDhtV9zC0RPBePatp4a0882wVTd8Hgz4f75dmrP1mFYe+i8NWYnM+lVTIRm6G/a65dI8jcjzxRVwwq1a9CKQlY8TsIr5MLZhS3k9iThiTasbWyXszV+Z4wJGpGbtGr4D28HCTSlCbgBcOG1u5w9Qbsfw3tS6uzJCr4CWkCS5vMSSEZ04cMmgMS30D35mIpPSMlFC5ABfxlApBvmMHiwATbD+KiXv44E5MyRAM3NonL3dWzR2rxXc96Zmxf6KLPnMlXaoacvZLBp3aKYHEcuJ+RvSwbI81TG9lnq4EFugNZPx3MjCsjKg6IEBFjCCD8Qa/jQUD8+JvQ8lPkY9bMpVXuOVT9YggAh2zYxKvJMoiRRwIwd5CMOzvxG0FHXK4QqZNaQc5rAIJABuX9nLa+WDqSMtRq4TtEeILw6IuHDJoDEt9A9FIjp1DOt+yfCJY3JM3IuJLibRfxGCr/OZH9vVS/7bAGtQfOO4jKx5jjgq5bS0R06bUXfYiX6zhTbA8chY5Tt3EhjM9vrnmdlm1zwakYfGRWlaqHQ6HYhZWnwF2qWDbObnQgpUI7ZC5rnMUy2k7tYkVMbIkusOU862QzUkp+X7SH4Wi2hEgoSyP0QyDeUmpFxveE2zz16lwirSgwwyJbaSdBGcNUDt/muS1VycFim3gpUZYUlQ5iaO5wJ6kWNLc6Zl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGaErZAzMptxgnEnTUb1FH+KDsgvF3nGagSG+j61Ycz6yVvOJnWltAuqG0k6pUgkH6tOL1NY5DSjnNgfS9N4r2RG6JGTmRR9C+axQ64GUsiZufL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyBhIwYo4qRNaCZjDQNugQQmXmk/7/DktWDwz9c8cX2oM3yHCRp5cv16eTMFa3S0m1hjmtOXbiPubZyvv2c1cYHFw6aU7RrgfF+63ZBBxfwvJJ9oJZfkDoldUAFim1hatMyXMOhhyiJPO8RlGCmkrijmCvd46Ibw8xuQ0mWUflRQkls+xA17uAZZ2tvUCPKMVBhr7OOWvkYN0AsFHOGGwbhDtJ7+F4mpB1Bid/nW4qcwJteNV0/W4f+mYftLJ89blVXbJEU00B7VPSDbOaea6xql5RegVUkdwR/8Z0yzxMB+OMKA1BJV2ZMjVjUK4txKY73CdZDM6AY8u5WmZ88UzVNwD3wNVtyCHZJbPsQNe7gGWdrb1AjyjFRZ/ErBoEnXnA89BbCQ0q9iyJ+jLd9gKjscM6uf5mBuNu5uHUzdNVg9yriECxML5w4OIP14ws2c9Ursi40Umn/4P8u3sezvxz9lHM0qos8cp7gUWOm1eVjvlXhHrqX7elJ4XU5FlvXWO8jen0O2p/Qg03FDXJR2t0WEnLoLATm9WPXs2xkcBdL4aSMqIrfVMHatZBcswRyPRmYp9OqMX+qWyQZBY3GfwFW5H+ZH7cBlayULZm+6+01MIwD8/MKoQRsJCRCunbjDzsBYLB37rmkwrJ/D92II+WcHTEiC3jvlSu9rQ1hbg0cdsiV322FEdL8uJTprYXRIo5255HY1yEwj5vyo4OV1XgcHswTrC6E/5JHOYmQajUx1+lhaxBHFM5Bg1MtGwBlMyFEJZt5I6hoNu3BxnJnHGi2Bd9N+G538qprs6rcE5ddzG6h96qoENi0OM5w1TIwwXrbHAWzGVQpXYmABKohTdQLxaBuWUrhj6qEitBzOi/Zigik71mRrJFV8xdfIHXy2z96NrpMPieZ8Tq5A4r2MI17e27KfWpZ8p/oos+cyVdqhpy9ksGndophAvDiKK56g4iHtmpgoIVG9yjTj3Os72sZAUjqf8aFBxTVmJzPpVUyEVH+pzO2S/SEBP4Lg3ltyKuxjbVPe5ExNMHRKiVWorhuZW8Gn8vZC/fW6vkyqMkRTPS2honXOFi8dJ1GNx+38IpU41/mYNZV8Np+ipJFgnO/C4OEyxUpTD/7rFS/YCcMmaIDJFYGPRH+z4syGXyZvxXsiK+IpNkfCC7NMwSseYju/1e7Op3Ii6MtQhLjo2j2bMJSf+SGC8MlYggAh2zYxKrOm4GNjZXJtIKLVRP+gR5CiNqZbc5+5EoT6EBJDziQgVYL83Ne2Kt/X0r37z3x1nwePxLG2o3WY6dZEDtKimZzAIuzossqYtsLg4TLFSlMP/usVL9gJwyZogMkVgY9Ef+of69PyB4yi/wEAvHr4WFPFw6aU7RrgfL/V7s6nciLoy1CEuOjaPZswlJ/5IYLwyViCACHbNjEqs6bgY2Nlcm0gotVE/6BHkE7868HnqpxxNrBKvbSWGzj85jILoHNoPoa31l+4dBcLB4/EsbajdZjp1kQO0qKZnPECRoXGgzTE9SbZSXMuXfHQpQ+QOt3fsANccOO/XLE6ACDwf94yKK4fESbyBRa/NKaQYPfgt28Z3fB4M+H++XZ9qdnVXZZL80XLU2IJXChka+7Cg3u9XBOrSatxI69erOb98+AaJaEDsG+QROCz5dYaeSEc5Yud15hSJ4nVh6Bl2K6hMdSPTRyyImF4gLRZATzPzcml80oZGRW7GsgL5aHMimULbhc2vRyNyZstNr4d5xdqc9Y/tkcATCfFXsIUI6rSZnPjhQ42RpPP13lyeVCnQKsaPZyf3LKsUXOyLGy7jI8rTYbbMrLVlP1PCMWiXMXDppTtGuB8VJ+ODj1Mf0QDDmo0qbnltslkgnfFIyU3AlmaCC1zlCkXNXmvhcYZKTkO9kUm1bA9x/xJJGMtS1ySWz7EDXu4Bq/7/KyzDUpMLor9W2CqgTboj7CG+iia2YMqS9j75lvBcfToHZ5ByWcbfKdF9AnQ9s15nwEletwQldmD65voKkpAhoDL61JMceRAr9Y3JhT7GmM340wuvpHo0u8+V8CORoASBrsEHIC+EGrHYIrLZhM0nN0fx0OZ3Tkh1dWah2CZUQlm3kjqGg20C28BNr6eaRt8p0X0CdD2SGMz2+ueZ2XSMuyhLR7IujQ68/3TNPUeGmM340wuvpGzpuBjY2VybfOoYXf/L/aGpxk0KAaU9eZuCUJl+r1Ko6+dhSVvWRZXV5gHmKglRiDMQT5ndyMiZzssUGdd2NvHgfEidBKHLafLk+ksSBii9Bhrvt/y+YAdZAVMQmFAh8emOUcbe62Sr8woYQPPigMRpexnL9SFCK3AWCwd+65pMPW6vkyqMkRT3ic5f2hOStc4cgLTyWb6yxMY7OSSvyJ2mQ9nw64RHES/StlC46lljpDRDzKAm9d6Yfo34/iLJxnvfAdTI+c+lH9UT7T+OlhGTtQr8I3+EpweEzJ1Rft7PC2vlg6kjLUag7kH7mhM4ejAWCwd+65pMB/NbgfH5clPHCY9gQ3NYJ2gnDVviL0CU0Te3KALTTmkSPSFldJ3ZOi8J65rEhuGBAyrarwHiLkNKAHh+NiMl4WSqL0g4bTQTBaRCtxdtd7SCus+RAcYvWhwjdJSWIVmBhp+hfQ+PJsIqDXxlkXGyt8pYDUFqKqyA/0UdzWIoAMcwZKHy/0/qrjmIqollrQmags+P2oLxFqD/RR3NYigAxxK+Z0XG6AnAP0UdzWIoAMckNEPMoCb13oLPj9qC8Rag0JD9RYEgn3vSvmdFxugJwBCQ/UWBIJ97wKB52gK4D7dRIoLn9egg/ArEd7yxJsnBqEf2l0Bu8dR72dsWBzBmp3Si3gnwT5xusJX7uUHYWcKoO2wwvuyY0Pmztp2apEI7nPQZQnBDMuFLzZqVUL5auoTnsUja9eUNqeiLfW6pi7ZwFgsHfuuaTCwIunSMMCd10Gm6u4OelGMPmrlMZOYS83w1hsUko1HBOvRIGFWSMHaNKUJuAFw4bUOBC1gLbvd1CnubR2ge3LotRWHyiFd5srPHH4OqAA6G8lkgnfFIyU3AlmaCC1zlCnAbqTKb9B6kjkO9kUm1bA9sA5DAM10CJtBpuruDnpRjDPMU9AxELw6np4Co0zf3UEYa77f8vmAHb23f9HiueSywFgsHfuuaTCIR4RxGWJ3azTXYXW48vaygTJ1LC156Wv+EyL7+ZhGMDPMU9AxELw6np4Co0zf3UEYa77f8vmAHWFmjN23bm9wqDXxlkXGyt+zamv/jJz667vlGl4H81DaxFePoirR2O0TGOzkkr8idlEAxF+JRliseCF965vPs0iJrvqYPJMS5XrjUnefVCQ49bq+TKoyRFOq953i5K6w+sBYLB37rmkwJgIAUn3Gw1Pdoa3lrlIzwALDpkyH5wfQ6oXWQANZxjEUOOFHUaMkut37uleBhS0UHHLMwdqMmmHAue5f9HiTip8p6JMQ3XndwFgsHfuuaTBCfMFMEwschXi/yLeLHPT7tccbtgzf6+pw3FUTCW8A9lKFmMSKGaCwJyOB5VW4Jdu1jYKECFFWP+ihfLxs7VlNe/nBiB5na9xaskvy1xDrxKcuF1TNa80s3OQdDSq7j/SoNfGWRcbK37kMM64Mxs2Vw2LdJVzzW0CuxJyd9LM6xDSlCbgBcOG1j+3qyr92AyQYrjiRX62t5KZhREc2ssOT67Cu6nIIXDYRDR43DzY5nk7Jwm3dUKv/RzlYZGU0qPqnbmeHkoMiQJVjm21wmymOGGu+3/L5gB2RjGUlDW9J9JRJ3ikEEnNVJL423q32qTBJFKY4b6NEVpK59SuWVNe9wFgsHfuuaTDeBViJgfCbUV0wzV75UBq9UoWYxIoZoLB2fQ0iqcKd+ETS6iLNamGGFh9/NNU+J0NXtqiBWW1lAScjgeVVuCXbwFgsHfuuaTDUijC1zL5WzvqIgTbdtdqmhvShEzA15OCVONf5mDWVfOsnWQqqc1EEy5PpLEgYovQYa77f8vmAHbWNgoQIUVY/xP4Nmi2XI7B5O0BAuyBLQqI2pltzn7kSyna7wE1bGzUc+jjnQlct5ILUi61PmdomCTD3uyIZyiwnmYYVTfNizFtTz97zD0D34vTbZ33JAvjAWCwd+65pMBSozNhxHwPCpoq1vkhTVUBSiM6w2HhbU94Kn5TsgwG/fXPtOZpTyA1mDmarMzI9a2yvZaajuJ026t0O1kn+EIo3CYt1TbICinbi6/K4P281GGu+3/L5gB21jYKECFFWPw4znDVMjDBeKHRZd9woXk89Pq7ZrlHYsrDJDPOfVY5omTQgmaQbsiI47qdjr1XbgHbi6/K4P281GGu+3/L5gB0xfQfSHVsrqLEddF643SlEwFgsHfuuaTCiNqZbc5+5ElXEAhZyE9IZyPSIS8uAc1LIwuqCJ5NKbetYAVL3aqqGoyBnbjeew191q4Riu/t1O5kASTy+i66UrxcNN8+D8sdGXKBF50gPHcBYLB37rmkwfC6ZEX19VS7eCp+U7IMBv9D+MdSntkCq6KF8vGztWU3XPZKLVGOY7BdT29xthLS5th44Q9DV70tBZE4CG6RYfJFARHmKW6eCNEfS46dJiQ6Q0Q8ygJvXesBYLB37rmkwojamW3OfuRI6V4PjRFHYJsMoYHudomr5uY06uMvU8st9c+05mlPIDUYENejXyaZ0NEfS46dJiQ6Q0Q8ygJvXeuxn4cPZRGabNv1C5IcM117AWCwd+65pMMdVtoj3JR+qG6CItCHO0RTAWCwd+65pMLTno2L+/ylGO8RlGCmkrigMw1M5J4o8Qmz1ByTIRx4x1a0eNY3QydQo7stvTR0s7eS5DQPA8zSVzvHgUE2mLXebLY7hnTYam6g18ZZFxsrf/RUmdUyx32wUOOFHUaMkuoS3DebhqcD/b4a64CejUfFg3JsG8RrWj6g18ZZFxsrfSvXkPabCstbFq37GJecbAoM3yinTYVCSK6AenPDDrkN2TgjiseEewcBYLB37rmkw1i5t3ireDk/AWCwd+65pMLkMM64Mxs2VStY8o/yfKK4++7088262j8tQhLjo2j2blopKY2Hp5D+oNfGWRcbK372rBUoGQrMwXWjfuQUjOLfAWCwd+65pMFDZj0W8HCXeD/+zzn0zT0E6O8ok+edEzFgOp7WWQNPu5SGockr4K6v7J4q03ufsn5DRDzKAm9d634OWJ6JCNDDr+fwwUr9VdAj8TPytperYnHNxHpyGcn/ooXy8bO1ZTRlTHfb2JHdTgdI7sbSXZa/AWCwd+65pMIhHhHEZYndre7yimUIEs2nZ2v6UzIAJW+tPYZrebgGzrB0lvwJpNQcfESbyBRa/NGAk6ZHNFtR8AEpUG6CU5b4S7mzIwwp3t6g18ZZFxsrfnmWzE0u/IKAFF51IrDAs9F2v4peCyWbJ/Wwq7SmsOmoDEBaMCddpERhrvt/y+YAduTXTDWFt4jK9P28sza+jCo0HNlT3nUEOMHiwATbD+Kj7uk6ahXm2yjB4sAE2w/ioQ1LmQfYlGuEw0mP3skyStMo/BfxkaL9tPwGopGN5FQ5Lybzp4Lcz84MqS9j75lvBvoiGCRllu1QQ9BMUbPYIWyzSrZCTRoPluBJBuMQkbczzl7xfWbVB0hl4xHnoc5F38v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLeZQ8ZfcClobg5jHkNozGqj8G0q9x0qsieJmO+09QPdxLNqa/+MnPrrH/HxnvP/lOmjw8gZK0E0BoBVgVE4wPK4b4a64CejUfFAgn4KDUCApRo7msUUe5bKjQc2VPedQQ6JrvqYPJMS5dXyZBsWXoSR9pW8s4hEntwf/GdMs8TAfhRHjNQxttQBjQc2VPedQQ7Fw6aU7RrgfIBVgVE4wPK4b4a64CejUfFAgn4KDUCApbk10w1hbeIyEhLNw8lwO8JIYzPb655nZaKdQxa98qI6+iiz5zJV2qGnL2Swad2imEC8OIornqDi8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEfUWerP1bc53CJ01QkFd/5eWgKyvsf7EpaXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZs/9kpa7wtawR07EIzlhgQPrMDTBmluIkfxScREvltrsHDZMRgFfe1OrGISi5pGmyy8V8b58GG7aywKTkKJerd+XIk1JlZdjcvlb6sRvxeiu4SSlnUTC2QhhfQeIFI3IYkLAf/WhvSmzOuf5rG3jMzNs/P9zr8kn/aI9EAkCE4YeNV9NkJ3IgcyJxj1tFS/ZF7QhuTs8tQu478bAujZ95coAYoTweg/wSORo1Ob49F/cx0TZ3feVhsRhfQeIFI3IYjxStOXLI6x8FuLOxxnorAUvB2RBqE8Qg/GED6cYfjdoNrlzvRZ41imTysGfIDZrZ5jY2T67Es+9y5PpLEgYovSzxO7EBtu+KLFItsraew8YikQAyWKXI4K/EUKWXiWm56g18ZZFxsrftG9I2nhppXmlVI5U9r6HGjpHZex+pcjKf2rv/Gw2j9nmAJNwG0YmvbVZ5juEEmmIyXyCHvmHys4YQWCKOqYQjTh5YBq8SNcBiH6yES2OC0Yvdm4Kr7872HKbnuut5hseg1lMb6Hbfejaw8arIkSo29TtvjGD9yErORlBy7+DbHPwJRVuVusUmDbwBM3rVecmDQf04/DAp2aCGooMjoDh8mDd+iWbwezwIuM7HDgBzj20OhnMHWApzBhrvt/y+YAdjfuoxOiR3gu3FdIBL16rtR7Tp5aGSSXNVMz8s7lE/N3Y6989s6rHy/eN6Mx3/cp0np4Co0zf3UGmYURHNrLDk/e1y6LjoC5l45v5ZAv/X3pzrAuY07l19raO9KF4fSqQFRVF2VN/TwK+Rctm6CpnDWY8kpni2j7KDB2TZHWspj3vEqVN/T2s0jSiIOJ19PYD4+UXIMII0IWwpGBD4G1YcxYAy57wk7ci51GHfWfElCG2Wc5osDyA88/zh0bfFD3m0yuXRCCceOY6/ObjqhPDcbZZzmiwPIDzwyrO01hlSvXAHFbRcisv+xU9K49uQlVwvasFSgZCszDjdhVjvvgpIWFmjN23bm9wM1ILnQKCFfPmjKghd4lsWyhQdezf/DTwSUvhi48fIltZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyqDJmsR/9kWohz+Pg21Gw+w0zB9aWHlcmao00x1enIKFJVOS/zOfjAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctBWUqh8ccsm2utZi+wc2cjOx7LgKysZ1ioEByRFu5q/m9ftHBTauKeUesELTuRK270nmAeVpWqKqvgwI9x/utdQxQ/1o3LCLDdI9OVRdvOOQbCAZ+BPqWvnBu5IeiZ8zAIkzSE3MYmJrprAqF0GgyQoZUSBv4ND0i492tamatT7f+RcPO0h2oArzA5qdqOTH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LxrFahAkPT9XzCterMAWpOmg61dEmrqcrGh5U5irJnyoBYNAncoGkg3cEuzEuWPSs0oCK5Nw7o/GPmErSoWFZK71siqWXvrBM16nabgm2gyiwjo6nhJm63zYNGTiJQjXZL/eE5UpRoQl42s7fuq63wfiqPFZR5iDogngZTYpYIfZh/AK6jyUPseuPkEySJxGdygDEbahTo5nXqdpuCbaDKBQOrzNqj4aqZ+Zcvc8YqF7jOMYv62/kSFtcKUm8bHtczoKtO3DvU++IQUJKyK6p0MBYLB37rmkwwFgsHfuuaTAM9uQHNB2YXgLcbJ4q7WwDK6IzqKwTYCISV5hreh9iBVSvlQqotonlmAjSQz3kM0hiBli3GwHjRi8C9IJ9QG7LcZinTM8Sur0964hux0Ylenlwjxm5HlVHvRmqVUEb0horFUcWgliT4Fh5E0gkpomTYDx0oL8iJkpmAmFR3LKaecIKQH9xapKWm5wIy7VEbo3tIPi8/JGwoF4JAwcpRs2wpWqh0Oh2IWULQ66nxKXucZs1xOkrv9moZgJhUdyymnnCCkB/cWqSlmpGPxRfAM1oi0ObZKSgLuZWYuTZOUuk8Bn/DST+uUdZEtRfj9IyqtXDHdoXX4sTnXFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/xMY7OSSvyJ2J1AqBPke3MF1YKbw3tpRShxHLifkb0sGc8rFJQKPIgNsR6DJqCUVytkjreHqRxKOnvPZszYH98tOQZIm7+zr2MLg4TLFSlMPXOLFD8ojL7/gLG/13Fj1hQq3p2gYMGjNvayS1Gpqmxf+J3a3ILgRbPmQvJ/Gtg5qj2idcEsQWxpTMzE3dlWywDpKB/H5OuK2DB2TZHWspj0NR6n22uP2ckngnZslNY0/aczFCQcL25Jr0IpCVjxOwjpKB/H5OuK2DB2TZHWspj2TbvQI0FmplzGFM4H4efwuTkGSJu/s69hx2YiI2TiMCPrcjZNT906bnE1AManRRv+PLBAAhEo5A8fgTzjkOKH6vt0W25erGIQD9tcnMj9RLqKxb1vVW8iGaCZjDQNugQQF7pVL7p7RG2lAqlLKErBpe66BPmKRG8XRDKF8K3NC1sIKQH9xapKWFIjp1DOt+yddA2JupV+0lE1Wmj6SnQZ1MDvPQvnae4ogi9P5Q05ExEFugNZPx3MjzRzg0OEb2CIcAhLKadUm31TM/LO5RPzdKL4bTgl9GUBUVhyWEPx3h0FugNZPx3MjDB2TZHWspj3fXDudT0tJURFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHXi2iAYDnChVzSsNPYwSujabXPBqRh8ZFaVqodDodiFl50r/6zZg8Qk+YCwwdvsA6leJkUNT+OJOKX6FkM9GFm5kddk+/b2Dhm1F32Il+s4Ub7CKGgQd+ImJxj1tFS/ZF5suLqNLo4djdWCm8N7aUUocRy4n5G9LBg8LfDEP9VEQZFdkSnhQ3bfy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR3+OoqL6yzGhJJGOGqiptanNHODQ4RvYIjpHZex+pcjKOZfAmSNmqnk6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcuQ2U1QDlmx79vNvWUuns+6cod/AxGty2OnTdwMBTJy+3LJBrkcxdC4ILsV8cKYvdWOO37jkgFi5zRzg0OEb2CJZGp/c0A8lBm2IZAJuaxDkRtVIfZAaxOLItndgTluCaUTS6iLNamGGFh9/NNU+J0MnrWRTas8+L3GYp0zPErq9PeuIbsdGJXoFsPDWrVvcYK/78KYYJzZNaDHA85r5sJlgPHSgvyImSlqk89/pi6AIv9281ooBjDYfILcYi00x4h991K5Rjd5QAgRr7UzjYUyoNfGWRcbK35TK09xkZJv1pfANeIcqZovDHzwZbJ7YC6FGpyom4OYrK6IzqKwTYCIC9JBI3SCKF4DNUCqI9DySWQ6MbX8gbuQS1F+P0jKq1cMd2hdfixOdJj0S8EAQi+b67pZhSX17SGJPnIh31XTulXeHI7I2QVsQ0gqCcU6w2oZD0YxFx+dr2OyoS+nYr+kvufeYUOXH4tAYj6W7Itm6WdDQ+ROdZrRCQ/UWBIJ977/dvNaKAYw2SQAYMCrv5UAotEvnc1rbYrV+ecwszI8EYNTLRsAZTMi2Wc5osDyA88VCgDEWvRH5UdHwA4jDjhhNVpo+kp0Gdb/dvNaKAYw2jfuoxOiR3gvPDmkjHL391FHR8AOIw44Ypsi835K/y9pg1MtGwBlMyLZZzmiwPIDz6Azmw+1XRmUMHZNkdaymPcTd5fHu6/15l2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkzn2Cf6wkDYmKavPtvrnwfrfqT+rxMHfMKhyurFjgufo8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/Hv0qNXg0VreFvQbK+WNpjgFObksMIQgJYmf0g7T8uikTmdjCz+epvdf0N2LXKhc5+a7Oq3BOXXcxuofeqqBDYtqGOBmnrDSvI4QVPq91Hl1YtJFi57rHJCAYCZgsLQ7uYUUFR/hCG6sq+Y2yg9NPB0nOqsxBXdWjavKRGwGO3hRS8V8b58GG7aywKTkKJerd+XIk1JlZdjcvlb6sRvxeiu4SSlnUTC2Qh2nX0sT4sDZ01Wmj6SnQZ1jRBmQQXz8GWoNfGWRcbK3zugtMZkamNKVbLK0jOxrG9RCWbeSOoaDeYkZzDDBaT7oSpQgBt0sRKf2Heakqlos6KPQswpnKzVQIaAy+tSTHE37Nk97b+6rmi6syZn5bD0l7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHHgsHxKdieRYWfoJvbUlc1kRdAmZwNaOLOEkpZ1EwtkIDwER1hjfhgb9VENR8xGz+RtqV9Udff3tL5Yp8WHpb8cVPSuPbkJVcJG7d8H0C1oz++yN/aFB7gkihr1LzG9HRfvsjf2hQe4JcRKQcX8ymmvjwuHDWjtEoZDRDzKAm9d6IhBYHCkvNIxaPyaFsoTw9LPyE9mT0B4Zu4I3OO3WRT6oNfGWRcbK360yD9MfwDAwgz5oQLaYuGZrHszq1lh4rvaK6mWAIB6b7sy1vrLm5Nvvbnyv/ffBBsF42tLIfze/WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm/AB1JrK16ldGxnewAZp2u53Tw/0vx8AH8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTIGEjBijipE3rdOz8XSMszo2y6sStNCDlhX9ZTeqm6mvtnfogXPL9BR8gtxiLTTHiIv7VDZlL2+XET/gv9cMW9eWWHZFhlfK4gPPvH8rhYwxTNm7vlhR09S/pdx3ngm+DIbFyY6T+wx8L73wTv+yxejc99kX+ZhHEpAYxBvVfzDgxTV3dvNtBTh9TFW4JdLljfY+SK17iu0YpD1cpko4vTY1VxarjbYSyYNTLRsAZTMi2Wc5osDyA88MqztNYZUr1dqhif0+tzjhmPJKZ4to+ygwdk2R1rKY9y4lJBcjT3OBAhoDL61JMcTfs2T3tv7quYNTLRsAZTMi2Wc5osDyA884Z96hw/mQcJV9ui98xHoMwwgxUJiDsGYBsBZkJMrW4D9c4l/IXVcNjewISjbwVy3wn9WtT2F5ray7Eodh8NsXhJKWdRMLZCLBvkETgs+XWwx88GWye2AtCYFiyHqgz6XEK95r9tEWsOvzm46oTw3G2Wc5osDyA88MqztNYZUr1Gm4I/d+gjR74Fbsq/pafJxhrvt/y+YAdjfuoxOiR3gu3FdIBL16rtZyW3lcNsW+VH3LGZz3tJ1Ek2F/s4q9aYBVKofLfQBmcs6bgY2Nlcm1hfQeIFI3IYp/Yd5qSqWizmJ67Ysv3txgdu62tcw24o7Z6L43c2d3hEPQTFGz2CFt3DCpm/rPLLq0yD9MfwDAwm7Cl/JGm4dRMzOo1oB5ATet07PxdIyzOPzURCNT9pGtwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3K6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiZEfwOqUUUJloUkXSGwKudVVE8Ebn6RXJynRi6WSalTmzMlfuRRpczm8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEdU8aqrXQC9Q2+x7ws0qUSn6mvGigMRpsklIg5uEtIbIYoTLfhodikQO6C0xmRqY0rgxDVdCuODJi0kqj/EritXUlO5TcmQkUge44zjqqXVT1WkSxWC1g6vivPvFHm9msvQrJURgKNO+4TkHZ7hGiLD8tbuCI8byk7y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPJto0/qBvL6+rdgUVHazgAVASjzdxlBBaX+7Hktoq/ItK7k1fdUmQuH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LiSreys3v6nxINhgRlnaevm2uLWEhhru+oOllZc3NZdKTk6TnAYGgqFxwAqIx4LVlsXe5TYf8MLJA7xnFayTiUrVt+Te0tbWDf17ZWwanxfT7j0y4SADvom01ow5XS2t4DZ82SMssH6LKoosXlmGqZ9m0sv7LJtanH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LvOELWtFYaJAxkL91+oXh1AAHKLhj4L3RjWp4X/fEthWNsdqxvyc0pvvhO+I7b9wotfJjinfBJCFC6f59p0irJG04IHWlU/9ghV7vicnp53OJ3RH1LBpOW8EFAOSDxDes5D3OwqTwAiJ1dCgW/W9lYAOWEQORr+Oi6pOtkR5QI7rnkyOhxNuHYrGs3fCXspGa6pOtkR5QI7oqjDr0IxGcVH9HBliQU+fp4zjGL+tv5EhbXClJvGx7XM6CrTtw71PvyLZ3YE5bgmlE0uoizWphhhYffzTVPidDNrBKvbSWGzjI0bp60Zfoq9nduMQ1dMye9xQVVy563YWC5AMwbRJL6V4JAwcpRs2wpWqh0Oh2IWUqosG7fI4x2ji1OZ51LoAHMCAsaLkc9sMgi9P5Q05ExKXZ7WLKC+D7uwWlpXTkn4NeCQMHKUbNsKVqodDodiFlHMiOaRE+CGpcxnIcGr//zB6lCDqYs98QPqMP6+KpyBpsR6DJqCUVytL4OQ7x9ikxZgJhUdyymnnCCkB/cWqSlqdxdvymQ2Ut/RR3NYigAxz/N2MTaHVG9xFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybRUEU0INUM9QztrSBB49v8Q1Zicz6VVMhCi+G04JfRlAVFYclhD8d4cH35e84+ZjqFAwKmLaU3muxLDbbahrs+QG1veh2UF/KpucCMu1RG6N1Q7YygwOAJeLfZg5JfrVqDGTzC+tFdi17GNtU97kTE0INkwj4mslX0R/A6pRRQmWdkmKu7UoUjSK4FmsDQU7Vvj10qKusZM2iMSlA/mF8JWO1CIYsmAvm3HO1gemEq84IIvT+UNORMSnC3EK7+Fb/MbXe09SFZZkTCIv7ttHc24RaygtE5naOViCACHbNjEqs6bgY2Nlcm3+J3a3ILgRbO6hN6M8acG5uQ6xY9qr2zkomfIY+Y3JZqAzJs48yu0oxF5kW0MLn8n6SMPtcQvVilfVkVgRs/0NPSmlcTAzXIxa4EjQb36tDmX9dbFfwxFUy8qBmrgwNGmInzg5kowD7X6O8+JEslxo8nr+ei788bHHVAfh+xg7tidJMmXJlwDjrjkwZ5Cn8miG71p5NFW87CJBkOvS8wY6Tc+2J5/NvU8X9jYeMTbpPvaVvLOIRJ7cIjKBsWRuLqiajn1JaStFfvGmdSC3aPlHgik71mRrJFXFpzMnvL9da0c5WGRlNKj6p25nh5KDIkDWNupr41iVFwePxLG2o3WY6dZEDtKimZzDPI4Y22ZnycBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwwFgsHfuuaTDsTHK/kmT+qR8J4GPXWCi2zDKA1INdVVkHj8SxtqN1mOnWRA7SopmcPH653q9/13op6lBmB0/fidwCF2aYxLYwCaVW8zsyS4fmT5kXDwJhhCpKXpL+hAWKxE/4L/XDFvWlC4hKO54XarYi1YtYrn9Gq3c5KWsu12iJWbp1N0EuiqEitBzOi/Zigik71mRrJFXdyrFR6viX/RxyzMHajJphwLnuX/R4k4qgN/I0+LGm1Uc5WGRlNKj6p25nh5KDIkBdS2xcwXwl6Kk5bc6diVZrkMujtqL7OAF7yysvY6nIChMDweU+f6Bsyp9uEq4Omqkk07wBT3oQ7VU1ZKlbjpVkHA4GATC61rStRKzJeyFCyOn7cWDofmj/yBAEFHCNZcZ3MXLiGV0fsIzD3wu+7NmP8ptsKVXQFSWRcaK7fovuTQAB4LgJfBifAZNoyurJazlDtJ7+F4mpB1Bid/nW4qcwkw9B2QNLfK3kWivo1U1Yp7AEOBFS+2GB4Tdq4N/b06eWLjqhdv2I2U6eP+E3qtBB5xpDfn//+Uft9Bl8kMMdX/o+fz8W1uhtYQ7X/ACpg7r4TadN8gbjjmz8/3OvySf9yPNUxvZZ6uDET/gv9cMW9WN7KwF4fRmivNhTaq7tQKS/dP79Ds9NObhwThsQ6qwMJyfLx6uu7u5AvDiKK56g4k3Ptiefzb1PxYJ6pTyEyFfrlznYlwOP6Kvvciyv21W/7gHEPwh5ar79FHc1iKADHPvExV7KRT08jMPfC77s2Y9wqKrcVZxJiZRt8y+CF6ptWaFvxr0W9Ot7A827fZ/94cqhlJEpWxCkl1Mr+8umKcdDdV7LVAvMyBTqe3BHol+9kk8EuEu/ErW+tfJPuegbDM/0HdKJTlSWkbvIgdlVIt18NHwseggR9MAyNKe6dMx+IjmEWfL9binOGbTydu4IPhxVLQR2X9QsbPRnFTdgewvzOIRj6etOhG3gjXOEok0SVH+pzO2S/SFZoW/GvRb063sDzbt9n/3h/WlzCa9iPRej6/LztCGn+2a0hyY5UrrqxE/4L/XDFvVhsmma/KpopeEx/UufzCpLv3T+/Q7PTTmdM4yGuwpymLl8DHo5Q8yKMMiP6IBLoQIcEwbZv3JZJMhZxK5Vy4qPevDVQLF2eNGboeu1t9+TNvlU3LhetGt5UlBsfAG9u8PzKkzrlEAfI5rAIJABuX9nLa+WDqSMtRq4TtEeILw6IuHDJoDEt9A9FIjp1DOt+ycvJ3O7SnS9UnwVJOu/RyyReyIr4ik2R8ILs0zBKx5iO4BVgVE4wPK4b4a64CejUfFeSk+xn52dIcLg4TLFSlMP50r/6zZg8QkaO5rFFHuWyrKbpNn7hkAvyFnErlXLio968NVAsXZ40dXyZBsWXoSR9pW8s4hEntx94Nz/Qo5rqysE6EgXdjLiHBMG2b9yWSQY1vbGF1Xl+Zb7Aw3YhO7OBZWaL8uN0xipc+ZvG0MyEd3DQ+tmxbH7pbqMC1Ds1LNeFCdKeXw5VtQpwH9+dJ6NMNJj97JMkrRUVhyWEPx3h0FugNZPx3MjFEeM1DG21AGym6TZ+4ZALxjW9sYXVeX5Z8qbqWlICMYccszB2oyaYcC57l/0eJOK2gvpG5cakkDRihv8bQ+HvedK/+s2YPEJuTXTDWFt4jK9P28sza+jCjA7z0L52nuKAi5nyDP1E0DB2Ap76lYpcPUm2UlzLl3xQEECCmIQDytr0IpCVjxOwl4ruVEFfBRD5CMOzvxG0FH555utOKn6I5rAIJABuX9nLa+WDqSMtRq4TtEeILw6IuHDJoDEt9A9FIjp1DOt+ydmk281ISqwQmO6ppjjBwmOSHmEoHtvgyx5xmXMo05cKjjgq5bS0R06bUXfYiX6zhTbA8chY5Tt3Oof69PyB4yiwgg/EGv40FAVUiE4dn+J1wE/guDeW3Iq7GNtU97kTE2caiSB0pwUU5ABfxlApBvmozWXR791Zi+sPWg6FSenyPx9q8/kPpTr+VqsHKyV31SVgGI+c9Ws26g+6chaHiS0EOfZEhOIKBMKvCL+HSA6aIE+jOBsGK0KE/34Z3y6pIThMJn9uVyfBiAtZkpLXQwg5DHa5eRNiiSFoHLQX6IZgvrzcrVPrhZXcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JiL6U6Zk7fLnIWejdBnAPYSxPDXWZ5bBHqbkncCzfQVa9bpiag0QICsGTtZFa3mIkP1y0YwqhtmTFJfCH5ij0a07s3gEvQ0hfnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTuvFlDLeVAgxaPbESEh6WniDxBDjrObGCRYbPk+prwtwaeSEc5Yud10znYrpwLeLrmVvBp/L2Qv31ur5MqjJEUw5XrNsX18DpHSdRjcft/CKVONf5mDWVfDafoqSRYJzvwuDhMsVKUw/+6xUv2AnDJsyVYUpSVWm2QkP1FgSCfe+Sh6M44dDko41by5HOo3XR1MRa2IZWQ1EcRy4n5G9LBnPKxSUCjyIDk7EXRx5S7nqVE7mAPLgIqlIjgPmtbR7lp7nrzt2/8AbgKQSDyK4n20XLU2IJXChka+7Cg3u9XBO16FJIz9mmD+HDJoDEt9A9G5ijMvAwQDKo1fNd3oasbXxi8NXJzKtA/wEAvHr4WFNLihmy6c4c8jR5O0NE/WMyRNLqIs1qYYYWH3801T4nQxxHLifkb0sGc8rFJQKPIgOTsRdHHlLuepUTuYA8uAiqE/zFwvjNPJsOM5w1TIwwXpnbKXJWyZ75RctTYglcKGRr7sKDe71cE7XoUkjP2aYP4cMmgMS30D0bmKMy8DBAMqjV813ehqxt5MkfMQRqqbq/dP79Ds9NOXCuVTJSltfSuEB5IxjYcuZE0uoizWphhhYffzTVPidDwU56OYAe6ZX2lbyziESe3LlG6tYuc7o0J3ow1ybKT4yRDf3vuHb674uvUqjSo744NWYnM+lVTIQovhtOCX0ZQFRWHJYQ/HeHJ3ow1ybKT4xDo3k2/UqVZkrWPKP8nyiuxj2xuG2LhpZF5/BHLWM01IEwRvSjn+e1cZinTM8Sur0964hux0YleruMncCERbo8H1MVbgl0uWN9j5IrXuK7RikPVymSji9NjVXFquNthLIbfKdF9AnQ9s15nwEletwQldmD65voKkpAhoDL61JMceRAr9Y3JhT7GmM340wuvpHo0u8+V8CORoASBrsEHIC+EGrHYIrLZhM0nN0fx0OZ3Tkh1dWah2CZUQlm3kjqGg20C28BNr6eaRt8p0X0CdD2EUvLlnOefzXIune8Z0CxayVfbovfMR6DiHgF0XwIjSVkv7zXjDWslqyQ/Esv7yB9eCF965vPs0gweLABNsP4qJXZg+ub6CpKQIaAy+tSTHE37Nk97b+6rmi6syZn5bD0l7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHHgsHxKdieRYWfoJvbUlc1kRdAmZwNaOLOEkpZ1EwtkIRN7coAtNOaT75A5d2KZgpymd1GvVwYIvVqGf7On3equX/Jd7sV/2dQs+P2oLxFqD/RR3NYigAxz/aPKDhBFzBg+gAXJbUtEK1g656/vN9ExUf6nM7ZL9IeiPsIb6KJrZwFgsHfuuaTD1ur5MqjJEUz1EgwgHGusWOHIC08lm+svQGI+luyLZujdFUnsP+5v3v0rZQuOpZY4CgedoCuA+3ZGMZSUNb0n0bFRpQnGlMxFYFOviZOqSnQLDpkyH5wfQZXQwZfR4Kjv0si9j1ltMxMHXYz+qP8poFZBGX3JVajOI+ghwMAM5XMxBPmd3IyJnday3vixe3DDNwuxPM/nWGyavtMRTLpLjwFgsHfuuaTBrdsX1B/aD/c9OQFuQqdpjehXa9V+jopf1uGjNuwcQNw2TTmFZXfuKtuUiN79YLGTAWCwd+65pMPW6vkyqMkRTw2V3UuBe0+b1ur5MqjJEUxeAIzzXgm7ZwFgsHfuuaTD1ur5MqjJEU6jXxEDppD639bq+TKoyRFO4o+rELtG0r8BYLB37rmkwkzlWvFuAZI3LOFgrq2wV8PXRHYV2QqsBy2C3pgvuo/OjjpqyTTRU77l8DHo5Q8yKsSw4+KysBeFYdGOsdmkCHIGKpp/33etHy2C3pgvuo/OMJOVZbqIUirOm4GNjZXJtb5lhdorn5WioNfGWRcbK36MhehYK1fxki69SqNKjvjiUr/b5CKimEdyoqaWzVIAC7Gfhw9lEZps2/ULkhwzXXqg18ZZFxsrfbpRsWACL1BN+uToH3eEJp4N8NW6mtnnw3FQqPpfDZI2jVwAI6174Oww/Gicvg9ZzQvZOoeWO9V+TOVa8W4Bkjd/P34Mge7YUQabq7g56UYyzW4QGgJqqnxhrvt/y+YAdgBIGuwQcgL5a4fNC4Bg8vFFHe/pf8N1kPwGopGN5FQ6yNcfwmy5SoQo87QNhWHJ8WrJL8tcQ68TAbqTKb9B6kiAlcEigg2iTLcJ6k6ujQLsYa77f8vmAHYASBrsEHIC+szV+Z4wJGpF/8ieeW5JAectgt6YL7qPz8n6d5dFRJkoiEL4cDCPslG/qpTA4Xawkb5lhdorn5WioNfGWRcbK33ghfeubz7NITDZKaorzh8J641J3n1QkOPW6vkyqMkRTF4AjPNeCbtnAWCwd+65pMCkURaCveb8IKjhT5iFHbnotIpsMLz7X0GWxPwOOlMm6qDXxlkXGyt94IX3rm8+zSMXDppTtGuB8aflC5wiB8yWTOVa8W4Bkjcf9eelcGFYNAEpUG6CU5b7JoXTMz08Azqg18ZZFxsrfTlP+WC4ayuxYDYjolo9NWCe8p23olab867Cu6nIIXDb8AFsmM+nuQu+ylNhH2VvCyqqQM41WEGRvhrrgJ6NR8f3NwfT5Ma0xqDXxlkXGyt+5DDOuDMbNlXO8DftZah7w5jFX3I/rG+5MNkpqivOHwovaLJTCYZnvUayQE/Mkam3AWCwd+65pMKI2pltzn7kSbuSKFBqhomoaO5rFFHuWyg//s859M09BwCoSVQoN0XSzpuBjY2VybUr15D2mwrLWFEeM1DG21AF7+cGIHmdr3BFLy5Zznn81TjV0yQLpoLP7k3E6Mz6SDgKB52gK4D7dzlQhkJuH3CkW+LSVy/V3Aa1XhbOjYyqMRctTYglcKGRr7sKDe71cE5C4sM5EnVlKzzlVju9HVR1Eiguf16CD8Dn9bRoAI4fNDy+psI5VfGSq2ejs9QVP/dkFuPehYP7oGGu+3/L5gB1QBtKNVwBE6TNDkC7ElrZUi9oslMJhme88JLP2Ojg4u0c5WGRlNKj6p25nh5KDIkCtvyqOrrmVi1GskBPzJGptwFgsHfuuaTCDomWkfWEtaxRHjNQxttQB1z2Si1RjmOweXE2LgPCRi+YiqiWWtCZqwFgsHfuuaTCiNqZbc5+5ElXEAhZyE9IZyPSIS8uAc1LIwuqCJ5NKbeAEFvbRl6/goyBnbjeew191q4Riu/t1O5kASTy+i66UrxcNN8+D8sdGXKBF50gPHcBYLB37rmkwfC6ZEX19VS7eCp+U7IMBv9D+MdSntkCq6KF8vGztWU3XPZKLVGOY7AbQg51J7QBcth44Q9DV70tBZE4CG6RYfJFARHmKW6eCNEfS46dJiQ6Q0Q8ygJvXesBYLB37rmkwojamW3OfuRI6V4PjRFHYJsMoYHudomr5uY06uMvU8ssppp+CeqsvfEYENejXyaZ0NEfS46dJiQ6Q0Q8ygJvXeuxn4cPZRGab/gWHRCvm82rAWCwd+65pMBSozNhxHwPCyMLqgieTSm1SiM6w2HhbU7GGVJChd5jgfXPtOZpTyA1mDmarMzI9a2yvZaajuJ02+oiBNt212qY3CYt1TbICinbi6/K4P281GGu+3/L5gB21jYKECFFWP+ihfLxs7VlNeTtAQLsgS0KiNqZbc5+5EoiOLu47xHfsHPo450JXLeSC1IutT5naJndgPjag9ge7bzu1PrvH+lxbU8/e8w9A9+L022d9yQL4wFgsHfuuaTAUqMzYcR8DwgfqmHqo8OWMFredfviJ3yoUR4zUMbbUAdc9kotUY5jsMK3N7Vf5hfYyS/1ZWcMwg+L022d9yQL4wFgsHfuuaTBhZozdt25vcKg18ZZFxsrfvasFSgZCszD5DAIG3fAXXBhrvt/y+YAdVbGraVyvYPQaxvwn/FNYsPNryEScwKMMjQcyNxXba5TIlWv+CmAf+MVW93s9vRKe4Yqd+lhQJBUFw1dSiTHJcJrHPf+Kbf3stwBulidXhNXMQT5ndyMiZ/wAWyYz6e5CBnNzNC/yWdT1JtlJcy5d8bbrCdK9iLZxuWDl+4FOsmjAWCwd+65pMAkw97siGcosTBMvOg2KbBo1Unf0L4On4mPe7K4RrctTqDXxlkXGyt9vmWF2iuflaKg18ZZFxsrfSvXkPabCstbFq37GJecbAtiAcRzVt4ZOcZinTM8Sur0964hux0YlelEAxF+JRlisgypL2PvmW8HT9cMkv92kqxhrvt/y+YAdgBIGuwQcgL5a4fNC4Bg8vAbQlShPjyqnZ/Xo0lhR9YXWjCbgGj7hFx8RJvIFFr80YCTpkc0W1HwKPO0DYVhyfFqyS/LXEOvEpy4XVM1rzSx17TDl/mvDrKI2pltzn7kScCWhfBWHo6ALnISQUnHalhhrvt/y+YAdgBIGuwQcgL6zNX5njAkakYvaLJTCYZnvf1XS8CNl+8IUR4zUMbbUARlTHfb2JHdTgdI7sbSXZa/sZ+HD2URmm5Yh+oizR4En4+UXIMII0IWRjGUlDW9J9MwvwfcuR8NBa3d20xoMxisX9jYeMTbpPvaVvLOIRJ7cFl+B2vyhbsx4IX3rm8+zSDB4sAE2w/iosBKvXvYz5JlIYzPb655nZaKdQxa98qI6SGMz2+ueZ2V2zXhKidh7YQf9De6l7YFLghX4L1x80hEXIxaAwuMe/MMd2hdfixOdkNEPMoCb13phZozdt25vcB+pBQUd/IzhvoiGCRllu1SRftjjGWJHTVyT4dfEL/inzN5EASkXmzE6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcsGOdbJ9JQtTVl2Xft10DA5koR7mAtx2FjvEZRgppK4oPo/jL+D3l26c14GdqdGddc62LhWsI6cm/3wgfWcI1yM0oHwwT/psvoY3RYaS4wOcPgCgf1i1kniaHQOi5kePv1qyS/LXEOvEKOyR1khAfqf1JtlJcy5d8UBgGExWwI04747LcN29Z/DvEqVN/T2s0hFLy5Zznn81/3wgfWcI1yM0oHwwT/psvoY3RYaS4wOcPgCgf1i1knjDKs7TWGVK9cAcVtFyKy/7CnfuWxyzru+AVYFROMDyuG+GuuAno1HxkLaF0j1X2V5wIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk6ufWkn8g78DyNnU0wlPo3tjbthrmLPRRVnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTEsgv1MXXJoi181pf0kIuOCW2/Bop+dbdIPEEOOs5sYJFhs+T6mvC3Bp5IRzli53X5CRqz7/gFKofUxVuCXS5Y32Pkite4rtGKQ9XKZKOL02NVcWq422EsmDUy0bAGUzItlnOaLA8gPOp8akuHxFzA0CGgMvrUkxxN+zZPe2/uq5g1MtGwBlMyLZZzmiwPIDzH64dY+z+8hJAhoDL61JMcTfs2T3tv7quYNTLRsAZTMi2Wc5osDyA88MqztNYZUr1dqhif0+tzjj3GKSbJQo2s/eBG8KWa740kKxaDasfPpti/QZxTA2ygikJuMch/Os1uWDl+4FOsmij7dfjcyhJHpkLg62wnfIElpwAZIX2MBvYrqEx1I9NHJGMZSUNb0n0LFWd+K4OI5wFbSMl/7gRZL2d4PrZZro1ZjySmeLaPsoMHZNkdaymPRUq/8MmgNJgUhP6NUz+uHQZ+O7mgQFcx0fzCHzVovFB8j2157ZHbB+Q0Q8ygJvXeqcLcQrv4Vv8TFc+ZFbYaF9scGRP3anPN6ZxFZnjBa/UYGaqsJzbjYaUbfMvgheqbeiPsIb6KJrZqDXxlkXGyt8L2l7RXsFjRvJ9qlCgm7F6K5CC5OYwi2mIxKUD+YXwlVjYvCkiKJEQFhCPWhSUC5k1X02QnciBzIjEpQP5hfCVEXU8sh86oYzhMJn9uVyfBtMX9XZt2jt8EPQTFGz2CFt3DCpm/rPLLq0yD9MfwDAwm7Cl/JGm4dRMzOo1oB5ATet07PxdIyzOPzURCNT9pGtwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk9q++V6uymFYWuBI0G9+rQ7yJShURQtb/ADKuVfSCivqH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LmmFES8+Cm8cGkhh4DauPmQGCFICShv5G1xg+mXKd5vkWAwRWLohduWwWyFLGq9l95dHXktQENbxD23+ziOLLX21Ukx/l+oXSo4f+2AKQ/RJI9cV2ZZxh2/0WQQjDWNreKweuWjCXiFaUuAH1jBo4g+inpX6f9thy2jmz4lCH4bEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsvZXzvFjDk/E8jCmrTA34ECueWGoonK3GY9BCSCKyXy1idipxlUuI0S33hUU5oIdEEWH4+LwrdSY1qeF/3xLYVZd6RBKNM6Eip9JBxvAjUF5wM/7WNDT+Ht3Ho6t/zr3ksoGaY57rssjtPolD6Gk0RojRR9jbQ+n40bOxDv8HmnztPolD6Gk0RFfsFXngExvN532mKjRs8Ag1fLXh+Rnpy0CNhofJt4MQSNujLFNzqC444+Osj2RCb0kJlNbXTHL7SSkFLmvgtji8C9IJ9QG7LKVP553NK9K5gx0wYE6lyMwz25Ac0HZhehgs3h8vaW5sqn4zMQnkt1w8G5+oIPR9Y6qh1DAeJ70oBYNAncoGkg5+gA4ucyggfGnkhHOWLnddxX2xf0wa4olMzMTd2VbLAHYNbLmfROv/kt3c7HJH3bJTOxVf6qMnZwWFEse2vnPZYXgyXk/raPQYIH6B0tKsptzdiLT7PbX7sY21T3uRMTZ+gA4ucyggfpaphVYGdTD5mAmFR3LKaeZ0aURK7nY7e099qJPs6ezkcRy4n5G9LBnPKxSUCjyID2DJ/p/4Tr3tmlFr7uAIXDJTOxVf6qMnZI4vTKyHBGc/8kzRDBuhudXHZiIjZOIwI+tyNk1P3TpvQI2Gh8m3gxBI26MsU3OoLPwbE5encBDLzuS3Svt2/jkt3HUvKPCdEFhfroqXXX8/55DKxfQFkEF73gOFfQuTIgtNdqGRakgznSv/rNmDxCet3yHn2palFrD1oOhUnp8h3gCAXaX5vsZKWQvmIGPZ8yxo5cZjlOmIBYNAncoGkg5LFaicXcUrcYcOMnvWkCBVUVhyWEPx3h0FugNZPx3MjS3rGKaw8lmcUbc/kH1brCpTOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMP50r/6zZg8Qk6woJNwQZhHt6SCsQy0uJ9lM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw8yxlfjqWOYzCnN+csYvfzxSYsnW3mFb6Y0nN0fx0OZ3WS/vNeMNayWFF+xR9syirfTgI+gsDxqVRF6KSzOPHtSJV9ui98xHoPTa9jgkAF3BCFPzo8BU4q9+jTmS3i9u2gfILcYi00x4kLLskYAyzFiahRfk6bD6m3oi9Fx59gBq54dOTwQP7uSmYgTZeB7vbBdaJa0dikXy/x410QcAsZTqN6SPs8vLOUl+o9tVuEAMtwq0tqJqU4saoTYGcjqaQqT6B1O4TU1gpJbEqlIN8KV1QerqOHafmx9m4/ShG5EHZTzd5+6i/sThzNo5wJfXC23kQ9N5RX7TefUh0ruRNVkrHEBNYVWkOfy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8dzcra8DF86tesx3hjZLBFUtqyQSO80OH+GczrbjADL/uE0MMnb24ImruyKeBbqLSPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4qWZ65dJunQWmgBv7vT+q0r9QUtczyfvs/35yBET7Vl3LJBrkcxdC4nHdTzrUUV4meMi5QVhkeDKRn1IoBQOn15PrdPzcq1a8tGE+AYWW3n0Kur71o/fuioNfGWRcbK3/u1sGvyizUfZ/nY7DOAj23nqLrMhomH+6i0zr5RNq4L56C69irDlslcv5nF8y9r8Rew4YYQevj+Sbhhe2Z6yRRowroLdcVxl7Ai8d3XbgyIFP4Po2mVehQTu8InJFdn3bFEhaeFPiNRdHZOMwzPULOUzsVX+qjJ2SOL0yshwRnPmcMADL8wR1G/3bzWigGMNtBCLtfkL/wdxPY/UBscfai+i47LNHaWlxaWeXv5OvXPMVoCMusb8S3/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk7TizYXxkptynHPfy+yGTjEo36jxjcHPC0RVGXD4Jha91wH27+pZglAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu4HJ38+96tAVqpLnfMG0vyGctd0h9c7W82lBBZ/ke9hT56hrqsU0m79BIfZhkVbfEV4TpnKmhoV9tabHMeVL1c+Fj7EA8Hh3eSCBV9piJ57cbjNWw+J3PGRDI8TqCS5LTwibdg+dXfa7cJYGK8HkqvEe/b7W25f1cC+Y9M7rTNLcd6fD2g1eHbJ5Kx5WsjPmjwzW77YErt8wa3YSKMusR/KO7Lb00dLO1E9oJN6JqfTZt9xwZbyvg6+wid7RW4sFiPWmwhxVmcAAiymnrTvhIPs9+PuhfGXttSm4BJAkwFRr4g894j7oqZwx3aF1+LE51n0bETR3OxmwDKuVfSCivq03NQQFCgtDwfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctPT/IbYgO2uVnwg/IMu6/6X3GFc3FY3ZPv+ggUqaEPvXOGXMNJvXM3NonL3dWzRS56qn3s1umWY9BCSCKyXy1gWv4xlzFUdpfSZQ1rylVvtG1k0bLNkmcbsJ75bYd9xRh2ETxdgzu21CG6JrnhRgdyZ5m3LYOxnpIxKOsNBr3GB6DBkVbuExDCfeTM9uG9xWWIE7b+X8v5SuZQYSsVEPZ+EUGJMpfqGhRrtvJVIUMOqR6tv3/Q8l8xL3s+sauxfHE6bSg8iThwM9uQHNB2YXuPUXcOGGOvVi+1qtVxWkYo8C5TsJcQtQdhFiScL0SeMURK2DxrwY3tYeRNIJKaJk2A8dKC/IiZKZgJhUdyymnnCCkB/cWqSlpucCMu1RG6N7SD4vPyRsKBeCQMHKUbNsKVqodDodiFlAf1sDL6Ym0r67pZhSX17SGJu0vDWy4qIlM7FV/qoydnBYUSx7a+c9hUEU0INUM9Q3EyAkAB+q8snp0XjP9MNUfWzKVV7jlU/WIIAIds2MSqzpuBjY2Vybf4ndrcguBFsrrYg5rBMpD0I/COA3pkEMNTEWtiGVkNRHEcuJ+RvSwaFY6DqIinVRu4OaKttStUSXod8D+TP6M3w5c7QuZaHtuSOCFwaOINhKN+o8Y3Bzwt1Q22CFKYv6xxxThBinnoiqxZl4MVZrJHET/gv9cMW9YSrYjXT0gkMW/bAhgJ5/Mk2sEq9tJYbOJc+dHZT/9fZ82yugDb7RNfKScVTKdMiUCXWKDmY9kDviU8ROYelXI/RZ++3QEqeiahB+B1OU9B4Tc+2J5/NvU+1bBl0nxBb95+yuUrJiANvewPNu32f/eFbNVwl9PhkPOonEreOqp1/PQmUO3tK2+jryURPHxh3SBYAuu0FrzaXrYuJOWYBPJWeuCv8EL5+zoiF1OttsAwHVFYclhD8d4dBboDWT8dzI64UwxpT64E0Qcj1oMvj/BODcSDGIc5qe+HDJoDEt9A9FIjp1DOt+yfdv7czRvnKL/3+YEl8JkNJ1ZmiKIU3ioflGPuPLedAvAE/guDeW3Iq7GNtU97kTE2caiSB0pwUU/VvfHslr74/zdDC8HvBEJWsPWg6FSenyOpt2ZyhBio8Cg6Y0RWO1So2n6KkkWCc78Lg4TLFSlMP50r/6zZg8Qnrd8h59qWpRaw9aDoVJ6fId4AgF2l+b7GISx6ocjkhJy6YNHca2zaUr4ePFoHgHvitHnTxlMad0dqlJ2PnUq85a9CKQlY8TsIr5MLZhS3k9sav0b7CzNyrFSnZpTP6WO7NzaJy93Vs0b5cQk7uFTrLOB129t1fowXRihv8bQ+HvQq8Iv4dIDpogT6M4GwYrQrxqVvfncEIrr+wWkWw+s+WTThqgOn59/4Cwvh5baNINkqelBsHOmpc+YvP2ifTwKmGemSMar/2gv7bR5f4GPKte3e9qzTxDx7NqyLGdo9RMhhDbO2fqMew0GaT9Geh3N1y6SUn/IOb9WPC5sDZ9s7TjfuoxOiR3gv+20eX+BjyrXt3vas08Q8ezasixnaPUTJlj6QQZq8aMgUUd1BPN1gSS3rGKaw8lmf+iguvnHiNm2z8/3OvySf9kkLIFFgqbo06woJNwQZhHt98dMw8FrEEbPz/c6/JJ/1NtKJ/2XzCN7SSscdUz+ZfgveUQAQXBCGXIk1JlZdjcm8c6tWxl7r08v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEdu+Qhalpct8FefWnp2D8i5yZ4JHOwzPVry/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTdE3sIX0nm1Wqc+lDkYz2Pn8UnERL5ba7Bw2TEYBX3tTqxiEouaRpssvFfG+fBhu2ssCk5CiXq3flyJNSZWXY3L5W+rEb8XoruEkpZ1EwtkIr3rQq99JZGJbEXdj+KLarkCGgMvrUkxxN+zZPe2/uq5VW3DiKRkzwq8tDEIZIuYMC+98E7/ssXoBJdeeMgT0Rx6dbQt3lImQtJelJ2P/PoEETOWt0KBunJJ3ezUKUQNvZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYcQr3mv20RaxC9k6h5Y71XxUEU0INUM9QxUKAMRa9EfkRO5zafLLM3OYiqiWWtCZquZZz/4Z84tit+0BpznpsqZ9OcakrJ0vrNiuqlYYkE61o+wnX0rc+pyNfAgFX27DVr6fZWZARLBrSWgC+kGOwIol+AN5C2/Sh03Sz3ydk7jMYa77f8vmAHaj8oM52ZaSHnaGT9cmZifG+Mcaf1n580nhkJL9CnTcCKnMAnFLD5Y0sOfrV7MRNjfPL3+hxaK4Of1tRnnB54EnF7hPlgASfqbVsGXSfEFv3GN3M34HftB7mIqollrQmak/bigXIRUzqNy3i5SNAjHMlX26L3zEegzDCDFQmIOwZqDXxlkXGyt/WLm3eKt4OT8BYLB37rmkwMGtidvOZwgvgpVaY4aXfF8ogeBHo18wvkNEPMoCb13oQ9BMUbPYIW3cMKmb+s8sur3rQq99JZGKDdcb3nkuRxKlZBRlHPBlhl+VJtD/uv6A2/ULkhwzXXr2rBUoGQrMwvnE5wKNaMBRiCjv/vpJYcMlrwpfsw6JL01+Hv04jZPQ6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcjI9RKJpATlw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/E6tOWoUnQI7Yu7X0QlN5LocCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNwY1qZHZMRiPsDCQkGF5TbBYQtlT4HBvMSBx+ApnC1dtyyQa5HMXQujpVvpgKf7cqetr0qG8sR2mdwJ68rjScMCtziW64KHAIj8G3eo7Q9Cu89XmVsQ5oR8LSRLM6i0pLhAiuoYSpfrNWZoiiFN4qHbQjASL1/A75mpqVKariN8txDu4MBCLEPXvpQWOSvxX24ZTogSJ81bgIuZ8gz9RNAnCa0GVLU3TzCFJNutzl2trfLjI/IcF+8qxHeJ7Xm56mdGlESu52O3gY+nSSN/ImOYZuXUTtMp2CoNfGWRcbK36jj6n5cKKkIj5IASVMIQbJ3JjemjG0NjEcuyxcVE9VcpWgH+DiJO1DS5B+HQuLItdxDu4MBCLEPLrzc7vG4bof0WRP9/7dMbG8VngA/qpziqDXxlkXGyt99QFCbsEdS9Dl4MXeNpD747z1eZWxDmhEtVDuLVhKgTT1N9d+fX7PwqDXxlkXGyt+WfTcDF5dBVCrYVflocTdqwYVIDFJRxvEr6UhuhHB4P2LX+CPbZuWdj0/592s/krZZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk0MSw/dqK9HHl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZMEaEGcGD5BKOCQ/Wta/Mur5ehiWYEzfDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8SB5AWeCzcNbVd4zBPYCpUI2jFsjiZ72mKZkUi6qw8jhgOtc6uS8kSgAzRUxw12Mz+b98+AaJaEDsG+QROCz5dYaeSEc5Yud15hSJ4nVh6Bl2K6hMdSPTRynC3EK7+Fb/DMKcO2ojSZ8JV9ui98xHoMwwgxUJiDsGag18ZZFxsrfhnpkjGq/9oIVAfLsSgeMGVEJZt5I6hoN5iRnMMMFpPv3GKSbJQo2s/eBG8KWa740kKxaDasfPpti/QZxTA2ygikJuMch/Os1uWDl+4FOsmixRWrYwzwlswVKXuPBvFInCso1jRkOTuBXmAeYqCVGIMBYLB37rmkwhnpkjGq/9oLbFNRAIs3wWx3A0fnE+ogdwFgsHfuuaTD+J3a3ILgRbHJVWGQFj9RmnSyC4YlbfY+PT/n3az+Stqg18ZZFxsrfrTIP0x/AMDCDPmhAtpi4ZmsezOrWWHiu9orqZYAgHpv1CkmbGnx0QtSMm8EQGs7zxM8HcI9XT4yXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZhmbc54Qbzm7vt0W25erGITJibuQ934z3OZsPEA18kKxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Lw77OF9d4rOWvl9lNkq+IdrX6T0NpFxbWIc83RD0iU+Wvu4K8NlLooedDa8/RTQEBD69i27DxUHP/OYV0R4td6r36mE7lWClZdLuAG7fM0+01lFoJxGMUvk5HPTRxwHNcLPe5OJbhzw21+ji0q/01SqEJHBnRAPIOVXok0c7Slo4aONrE5vpAqyiIEDQJCrR4R0vkTx8jAuHyB7SGLKppN4di/BW5rpijdr9OhV3OvWu4YnNpOZCyWtjMikXbcoiX2bSy/ssm1qcfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu84Qta0VhokDGQv3X6heHUAAcouGPgvdGNanhf98S2FY2x2rG/JzSm++E74jtv3Ci18mOKd8EkIULp/n2nSKskbTggdaVT/2CFXu+Jyennc6YKtC1om99Omcg3KvWmp5fHyHG/4bYl62fgrpUCcPDtPSYisw/CJsfbd+ErbQ3haY5ylQhF7i9w1ph9EJwygYpWj0KFx+ag3+SR0MqJ2L1KLoDy6LMmGU1U2otzxEUoZFuLLdvgaFIRdjU2j4ISnB7w6UokcnK8ntO2bz/z2G7xuKubYBgw9zC+MQYhrirnU7B4b9+WeicmLNVi6kzY6FitEZK7kisEEh2DWy5n0Tr/BMlZKI/I2EqsPWg6FSenyE7slFv/HsQ4HyC3GItNMeIa+4JkKGk8XJTOxVf6qMnZwWFEse2vnPYVBFNCDVDPUNxMgJAAfqvLJ6dF4z/TDVH1sylVe45VP1iCACHbNjEqs6bgY2Nlcm3+J3a3ILgRbK62IOawTKQ9CPwjgN6ZBDDUxFrYhlZDURxHLifkb0sGhWOg6iIp1UbuDmirbUrVEl6HfA/kz+jNqHAA82TVfxbkjghcGjiDYSjfqPGNwc8LdUNtghSmL+sccU4QYp56IncB9p8tbHpLxE/4L/XDFvWEq2I109IJDFv2wIYCefzJNrBKvbSWGzgmtgEXIx//ifNsroA2+0TXyknFUynTIlAl1ig5mPZA74lPETmHpVyP0Wfvt0BKnonALizluSC12j/OY6jMdBxTb/4eFkoXysEbqH3qqgQ2LUuOPRgIUequX32Qm+hTO+aajn1JaStFftQ1gA6qolsK94u8CSrPQ/1b9sCGAnn8yZxqJIHSnBRTWJbN2Q86ef1uVZtPPGIBbpi3nmW7jCeRHEcuJ+RvSwaFVSD1FKcXtP9CJj5CZlsarYuJOWYBPJWeuCv8EL5+zoiF1OttsAwHVFYclhD8d4dBboDWT8dzI+4ZC1Q/KF70r4ePFoHgHvitHnTxlMad0WcDgnFz75b9uE7RHiC8OiLhwyaAxLfQPRSI6dQzrfsnp68vGoAbglJEIb26/dclaQFg0CdygaSDksVqJxdxStytQfOO4jKx5jjgq5bS0R06bUXfYiX6zhSnJ6defzt03atESo6vr1MqAWDQJ3KBpIOcaiSB0pwUU5AEldLyOmMlEzQiZFoHye2UzsVX+qjJ2SOL0yshwRnP2W3a3wXw4fbC4OEyxUpTD+dK/+s2YPEJOsKCTcEGYR6lNWOPJiOWytWZoiiFN4qH2kkRKKA5QvZYggAh2zYxKkC8OIornqDiZdsjXDviZ5zzIKTcp0Jivoy6NTgOShUloNbk+aiHxqVp8Bdqlg2zm50IKVCO2QuaA6ZAmpajGJ8gLDtzz5ZwRbZZzmiwPIDzWXk+RRG5wTDfAAkN/fGIzPiPl5MiZhQu2QzUkp+X7SH4Wi2hEgoSyO2wQcP6lym6LBEHGUH8dAy2Wc5osDyA81l5PkURucEw3wAJDf3xiMz4j5eTImYULvrzcrVPrhZXSW7KL2E8xzEumDR3Gts2lDSc3R/HQ5ndSJzf7aYh7pwUX7FH2zKKtxJXgTipY6moNJzdH8dDmd1kv7zXjDWslmHY1KyzivUy0Jfc4AgPp/TiXFvp7Ix3TgFkCn818U6ycrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Jq25MXY5NEIz6g6QfGiE/1dZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/MPu5duQKtzKx5ZD81sWasmXmk/7/DktWDwz9c8cX2oM3yHCRp5cv16eTMFa3S0m9JH4RiFSfrKeCwfEp2J5FiboR8KKvMtE2OfTLT3e9rBuWDl+4FOsmj/09byjs1c/z4+0sgCXTvPbPz/c6/JJ/2iPRAJAhOGHk/bigXIRUzqNy3i5SNAjHOE99qa8Zlz1w0KDdauuoRlGHu9cSXeg1vLcOzAH61pHGi6syZn5bD0l7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHLmWc/+GfOLYrftAac56bKmfTnGpKydL6zYrqpWGJBOtaPsJ19K3PqcjXwIBV9uw1a+n2VmQESwa0loAvpBjsCKJfgDeQtv0odN0s98nZO4znwDziWeYZMyLzKGYDX+EQcKCoYvRrkw+PcbXn57c+przoFW6yuS1OvDFKejzwt7G4gNyZ6YCVLIrJgj0vjeWlNWlReDBnF9nPlI7GciR+cNaMQZnlv49VQVljdKlLijEwFgsHfuuaTCuFMMaU+uBNDSc3R/HQ5ndZL+814w1rJYvxMuc4I56TpvhQT+f1furGGu+3/L5gB0enW0Ld5SJkFz/aSx3XfJ6Or9v5F34ZyKoNfGWRcbK360yD9MfwDAwnTBiBzuxSrQOEEoSOPCNxvT0tuiNCFmwLnux/W6aseatMg/TH8AwMJuwpfyRpuHUTMzqNaAeQE3RN7CF9J5tVlBtg3yQrquH8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTbAH7uH46mzpwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk65y/SiHqTyWq3eWrDuRRrChFf4W6s7mRvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxO3sUjWBOwNwKhS42MiSYR4X0i1k4boFv4kBOEElYdWzyP5RBVXdjdRxxThBinnoi69sQejztKcsUl4pP7SE7y5rgHTNiKjwkRtVIfZAaxOL07LtW3s2cqHR2TjMMz1CzlM7FV/qoydkji9MrIcEZz+HOpWpJxAF0K+lIboRweD8nl6Af+wRDzXuZeP9gUJIJAWDQJ3KBpIOSxWonF3FK3JVTmqiZ/tUYv9281ooBjDbQQi7X5C/8Haw9aDoVJ6fI6m3ZnKEGKjx8aWSUg45QJ9Wa+2SQ2WBb5irLF9XJUAPnoLr2KsOWyb7AJY8LvE71C1/hnQogtm9/piXYAzy7Kz1N9d+fX7PwqDXxlkXGyt8dFcJkhgsUvirYVflocTdqwYVIDFJRxvEr6UhuhHB4P+T2sOlR026GXFYIojpz9Ve/3bzWigGMNkrlJ4aWn+UVulhRBnYeT+x4Y8XqlYotK3HdFrEAEIc0syuQPp/8Ye3TgI+gsDxqVSzqycMxuT6Eqk2qWKPfuUUuxPUN2+8SQq4ff7MeCeGX8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTbAH7uH46mzpwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk65y/SiHqTyW+68sS9oZr4aycgQVUd02w5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmDX/aUb2X9hazgeWK5JirGg+/b07x5zgSoWFgEdetSo1nauqvuIr+zGpQqLKO6hlOJ6b+11OiNzEAGkuTHgN5IB8gtxiLTTHixi1yExziaZRxCvea/bRFrDVfTZCdyIHMN5EYmtNJnq80OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm0avIGz3q2D5jMKcO2ojSZ8JV9ui98xHoMwwgxUJiDsGYBsBZkJMrW4D9c4l/IXVcNjewISjbwVy3wn9WtT2F5ray7Eodh8NsXhJKWdRMLZCNZbUSIgt1qhN5EYmtNJnq8mxq/GMTx/a/CDAdI6K1zo3PQklR7DhT7Nov0IX6w357j3SPMcAYeAtlnOaLA8gPOzpuBjY2Vyba0yD9MfwDAwm7Cl/JGm4dRMzOo1oB5ATbZZzmiwPIDzlBlwTxqYgv5ZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8dI9QfLeS3idmx6myoLZxRzI/wsCS0pMUKH1RpANeJ/UMc8eAUmMqAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsAyrlX0gor6tVKtg7aPDoVB3ByGK/VBOniK3a0yLM5mRQQDm0+FyW5cCrRrGz4N4rFPwThf4xO935KcFXXGVwNLFN64LgH5CMAyrlX0gor6r9bgnYkdWlIlLgB9YwaOIPOoR5mYSh/MdznjNahCgxJJtrrWYvsHNkfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwuww3/rjHvIFDePOF6xG0Bh8pwSfM8eXNQ9RXqivQAlT+abRD+5p50oQYXB1BpvjBwak08m49SkB+iUB+Pgbq2QzfePEWZj9IYLc27ZGf6M1HVODk2HTHtwJwwMAKj03N7amJweZoQIdS44skmZi9WoTXyMX37/h6NNz7Ynn829T2x1FGV4L1RoRp3Z+BImbXi/dP79Ds9NOfFXIUJXT+yExE/4L/XDFvWcdeoVq6McDzw6A7szFSFvxj2xuG2LhpbxIXdoVlZMAozD3wu+7NmPFy9RLzcVy2H9nzC7v1nHd0c5WGRlNKj6rjkwZ5Cn8mgAvyhrEnYLsXtGVKQ7oCj/beCNc4SiTRIji9MrIcEZz2OO37jkgFi5WQ/Sa6Ht3HC/dP79Ds9NOT91/aHKeIcRxE/4L/XDFvVMrpf4fjuRQ2OO37jkgFi5WQ/Sa6Ht3HC/dP79Ds9NOZF0Py+LSCPmRvIdFJb4qjDube7gCSjRHRI26MsU3OoLPSX+5s87cFdwukwNlc6T+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3eCMgS2aQYlSf8lVN2ZZgfoxCFMy3ABQrty9SLWj9MahDVHhRSEtqXSdRsYz5JZBMnmvXHN8NcKUL5H3JR+gnQZvxh72Y6FA+VPnyoAOCdrJtrrWYvsHNlUFh09Ch4hbnzLmZaGtklfhrmggKLGSVOfHOCv+mtTwMLT3JSAFfVg2jmz4lCH4bEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsvZXzvFjDk/E8jCmrTA34ECueWGoonK3GY9BCSCKyXy1idipxlUuI0S33hUU5oIdEEWH4+LwrdSYan4nrK5j1oJfQStDLFQ01WNbV8zjtZu9Fp9CoamTipsFAU5C9nfKJWNbV8zjtZu66BdPt4ta9+W5wwOVSASsU0Pn/VgPsBD18+HpiKWFvZCqlntSoAU7cJuaglfeAYm563PkQGIyQNEAGbFVIr1LCkyA2VBukLUFfZITtU129QrPZi+i+QC1gUiOnUM637JwO1EyZzJsbRI76HSrUmNBv9FHc1iKADHK9pzNU3Tj8aSD2I43Q5NToMLtD4gPUc+kFugNZPx3Mj5up/OZQTrX8hW5crXar1Le98B1Mj5z6UGmzRe6RhG4gtMZHWzYyLJ++4Gv3Cdn6ZIULKBjHbC9aDnHxxKtmNhOic5viU2SKBpmH7SyfPW5VZspqzcfZdUfJMoiRRwIwdXIigbRpCe1exCSNu0O+EHb/ux4kGVmNUGmzRe6RhG4gtMZHWzYyLJ++4Gv3Cdn6ZIULKBjHbC9aiIcDNDHyPQGoU4qDWArjTkMABQU0zL8vM+OWm9Bv/ZhSI6dQzrfsnzipsXfjRAZ/4A8kpkiKbhK9pzNU3Tj8aSD2I43Q5NToMLtD4gPUc+kFugNZPx3Mj4zAgiQwcdlsl5L/8f93KWQaTyGEi2sMJo42UxL+43zq1wem1vSaaXCvkwtmFLeT2ENIv1RfnlJRdUSTZQAKh8FtprfyFIurTjv5IIDcgmHJ92cTxFwWkp+dK/+s2YPEJa+BsP8xrvrS0AeUQkzvyl2JgASqIU3UC8WgbllK4Y+pjvMEvk2JyMG+wihoEHfiJYiXjVB/XWYVm6N03kOe76VtprfyFIurT2Nw4dCbyxOa1wem1vSaaXCvkwtmFLeT2mYjM42BnfnVaaAG/u9P6rd5h3/0++q6msoKKioP2TabxaBuWUrhj6mO8wS+TYnIwb7CKGgQd+IliJeNUH9dZhWrmsl3HZ+TuwnVa7oVxliv8ShOLWwn4xkg9iON0OTU6DC7Q+ID1HPpBboDWT8dzI10QQrtbgdatCONgulB3uAaQwAFBTTMvy8z45ab0G/9mFIjp1DOt+yelN0crhBSppkjWtpFKgZnKAAHguAl8GJ9hJUIiNX81b5xqJIHSnBRTtZs5Ri1VsAqFPJUxZTNeEzmLk6Ur368FUiOA+a1tHuWjjZTEv7jfOrXB6bW9JppcK+TC2YUt5PYpZGx5Ak1/OJQbQlB/29fgPwGopGN5FQ49Qrf25DvhdpDAAUFNMy/LzPjlpvQb/2biV2Iip173FdeCiZpZemRCmxzv3OMGq/pICbUolqPW/t/tTbF4kMUBy1MeSZtsoFZywW88GIzBey0xkdbNjIsndayI23t8j5ZBboDWT8dzI+bqfzmUE61/nMLmC8e/7qJOoLBj7nZ4mIxXewkyAg4w50r/6zZg8QkWNBDZldmkxocqqiDGcCkS99GvZaLhYDteGO/gp+2qSQo+otmfV1RcK+TC2YUt5PYsIxenHftXO/FDNmTI2QuXJEFN2uPF39oH4hDXtDroPZtBYU8vr0+0K+TC2YUt5PYsIxenHftXO3zG6KXCFf9gKklPVvhIMMBWkusaBbGR6NI1YI3AIDQKnGokgdKcFFO1mzlGLVWwCkDeFbQdyaYIODzP2boa6B5ywW88GIzBey0xkdbNjIsn+FLSMoeflC4hQsoGMdsL1gBCcn4GIYDutbsoW7d6GISX+GA/l3fSWMVy62lIczC8YSVCIjV/NW+caiSB0pwUU7WbOUYtVbAKJw9YlomiUp8tRTqHjCyh8oTfLYjdTFy/tCwUm+iC4cktMZHWzYyLJ++4Gv3Cdn6ZIULKBjHbC9YAQnJ+BiGA7l73gOFfQuTIgHZAyG88J4n8ShOLWwn4xkg9iON0OTU6cV4ughi1LB0UiOnUM637J9GZYB0BSKJQFEB+jvEgReFAUjqf8aFBxdaYfRCcMoGKnGokgdKcFFO1mzlGLVWwCuTjfgXGuW/LQkP1FgSCfe8M9uQHNB2YXkF1/DjXpATYIULKBjHbC9bEM6dtEg2/A968EOBIB9h6Vw2+x0N47+cMq/0Q2lYh/0FugNZPx3Mj5up/OZQTrX8MHZNkdaymPRCI7jomL2c5DhLedypjXa0UiOnUM637JwO1EyZzJsbRqORYhzctgv4uktl9KR8Xm9aYfRCcMoGKnGokgdKcFFO1mzlGLVWwCsgAjJdbGzIuRTbr/KAiek0M9uQHNB2YXkF1/DjXpATYIULKBjHbC9bEM6dtEg2/A3kNXIfeKigvVw2+x0N47+cMq/0Q2lYh/0FugNZPx3Mj5up/OZQTrX8MHZNkdaymPRcxHTrFz83oDhLedypjXa0UiOnUM637J9GZYB0BSKJQFEB+jvEgReHG13tPUhWWZEYNHhdfKXcB+XkZao+zO25ciKBtGkJ7VxM3fs/sBgyjDB2TZHWspj0HnJvSxYDypQyr/RDaViH/VPGqq10AvUNvse8LNKlEp+prxooDEabJk0Zf5TxnF5p1OluoqQqTLc7W+/RZJSOcly6IveSStcCJjSURAVkO2uZsPEA18kKxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Lw77OF9d4rOWvl9lNkq+IdrX6T0NpFxbWIc83RD0iU+Wvu4K8NlLooedDa8/RTQEBD69i27DxUHP/OYV0R4td6r36mE7lWClZdLuAG7fM0+01lFoJxGMUvj5qAU4OLm+bNy+Is2NkTwvR4NJ8ws89SlLV0lODWjt8YHVji4eQbrcNfP/1CBud8czmkN4NvJP4ziPleY1lNnw5M4JeSPOmhkTMjO1CNQCPWfW+PJc4cI/xsDZNQf5yfinQCRuSRe17kgPndk02HPfBKAUQhYItKliSMtNc9SEvekvLbDDl+SqEICzdOI5KsZwNIS8zqKxsbJ2mK+eJVY1EVijxvDsK31nhIRslsGhtrDl147+Zt66+ifnZ4SKPdvsqArPxcDnjP7GjsmFwY0RkRcQw8S3MqScEHHnxd1EGcSbaa481Dxg52Ev6fZfk5bTOZoYotpWm9VrgRT0bneYRFGZ8kD+YFRB2GOqBjCWR0xkwnC4cf8+AK8wOanajkx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC8axWoQJD0/V8wrXqzAFqTpoOtXRJq6nKxoeVOYqyZ8qAWDQJ3KBpIN3BLsxLlj0rNKAiuTcO6Pxj5hK0qFhWSu9bIqll76wTNep2m4JtoMosI6Op4SZut82DRk4iUI12S/3hOVKUaEJRnoIJ9g2lpY0Pn/VgPsBDy/3hOVKUaEJeNrO37qut8H4qjxWUeYg6IJ4GU2KWCH2YfwCuo8lD7HO1vv0WSUjnJcuiL3kkrXAed9pio0bPAINXy14fkZ6ciKkk5GRrj0R8Zi2qBAyTsfSQmU1tdMcvtJKQUua+C2OOFTpMzY6wska/bmiiF27WU+R6vAG7XITCOor9i3pSbRihvvBdVc3zeD/R358veDxiFiQ0ht2FeFYN5Gu44AJkf3xP/3CDHj6BLUZRP9K6HYcT4NCWvNKVqwcV0A9sL6eH4XBOP/gst8ISggg8rXMzpTOxVf6qMnZwWFEse2vnPaXIk1JlZdjcrInvCB4XJTTAWDQJ3KBpIMINkwj4mslX2dAD0Fzenj9s/fOdT+1++tQgnJmgVSSnmxHoMmoJRXK0vg5DvH2KTFmAmFR3LKaecIKQH9xapKWp3F2/KZDZS09R5QN+j+vQlKUnG7T12N5f5Lu66NXfxGncXb8pkNlLT1HlA36P69Cc4SNAPWFs2d/ku7ro1d/EadxdvymQ2Ut0xfoFCmg5eNSlJxu09djeX+S7uujV38Rp3F2/KZDZS3TF+gUKaDl43OEjQD1hbNnf5Lu66NXfxFqRj8UXwDNaMOcPsm7HRZy4Cxv9dxY9YX5+7dLcygsMP4ndrcguBFs+ZC8n8a2DmqPaJ1wSxBbGlMzMTd2VbLAOkoH8fk64rYMHZNkdaymPYCZ5+GacpKgNWYnM+lVTIQovhtOCX0ZQFRWHJYQ/HeHpwtxCu/hW/xMVz5kVthoX0wiL+7bR3NuEWsoLROZ2jlYggAh2zYxKhG4sbj7Agur8HCdlyZMBoCZzEU9ofVWWvViczpsTdN7rgZrXgA/9JBzI/wsCS0pMXRTrjGD3MY2bV3Sg4yPP5eaMs1s/8Z3eBuofeqqBDYttuPIRceaHpVniK0mrBLjvIlZunU3QS6KbEegyaglFcrJHIii8Cp914pdE0Xytk/cFQRTQg1Qz1CrZxDcwVVlEjDIj+iAS6ECFIjp1DOt+ydgTG31GYr4clBamQfZC6JdnlHUuVejHZmuXpj++ES6S7hO0R4gvDoi4cMmgMS30D0UiOnUM637JyphNYfoJ1rNUFqZB9kLol2eUdS5V6Mdma5emP74RLpLuE7RHiC8OiLhwyaAxLfQPRSI6dQzrfsnyaBgzyaeI9rYZLLjYfnGANMX6BQpoOXj1OAwv+4oT5w2n6KkkWCc78Lg4TLFSlMP50r/6zZg8QnxDoMZIVQ0xsD7L6jdjs6tT5zqLN228HOojmkspMCESTDSY/eyTJK0VFYclhD8d4dBboDWT8dzI4+SAElTCEGyCnfuWxyzru89zQjfrwajONWZoiiFN4qH+bPzAzu/mfq3BrWU01tJZinBQ55mE3EBtW5qi9YbEZtcrVE31n15MZKHozjh0OSjpcKnjDbnXtGZkLwGqEuUb1CRrP4WjxKEHEcuJ+RvSwaFVSD1FKcXtLVuaovWGxGb70Qkv4MmFaGSh6M44dDko6XCp4w2517R9O+4qWJ17/9Qkaz+Fo8ShBxHLifkb0sGhVUg9RSnF7S1bmqL1hsRmym9qAc5ZTKvmsAgkAG5f2eWpgbSIG28zbhO0R4gvDoi4cMmgMS30D0UiOnUM637J2X3odZT/uq0r7seiTCIRK3ZqJ9e6J+oSWxQpMAqVKTVNp+ipJFgnO/C4OEyxUpTD+dK/+s2YPEJBmrZPIZVucie6bg/l3CVrthksuNh+cYAPUeUDfo/r0LU4DC/7ihPnDafoqSRYJzvwuDhMsVKUw/nSv/rNmDxCQZq2TyGVbnI9gUipQkD7bTYZLLjYfnGANMX6BQpoOXjoLAobAf76/82n6KkkWCc78Lg4TLFSlMP50r/6zZg8Qmlt+S5qb0aNcIIPxBr+NBQ1yMqcIwIh8X1sylVe45VP1iCACHbNjEq8kyiJFHAjB3FTczZP+QykPBpgJ3l7HJANWYnM+lVTIQaOPj4PTgm7wE/guDeW3Iq7GNtU97kTE0pwUOeZhNxAbVuaovWGxGbDCRDcuBbj30m/iT4JatGqtmon17on6hJbFCkwCpUpNVtIpEPypiDT21F32Il+s4UpyenXn87dN26NMakaRBDLN7Wo1mKhDIgmsAgkAG5f2eWpgbSIG28zYGpI4qOFrpUDWHYV3mAVRdYggAh2zYxKvJMoiRRwIwdk4ifbidJd0QxlWNEPFtMgf3QKvhcCLHPgQu9lTzYU/Rtymqjqiczx4AWpEcZWSK6gCrGIzHFYIhr0IpCVjxOwivkwtmFLeT2zjCnzIV+ujYKMgEhYlMOs2MF9WizK2bj7NlM8jYW2XP98T/9wgx4+jafoqSRYJzvwuDhMsVKUw/nSv/rNmDxCZRrBTzSNecVs6G/BDHDNQDCCD8Qa/jQULj5fWs7R8UIBoOOv9pjoLY44KuW0tEdOtGKG/xtD4e9MsZX46ljmMy/Wj3bDqhdafseG3UkeS314CHzjZkiXGuMwrZJ/yLzJSdcGS34ROwfURkdQH8hEA5/pyLGzhNc8rDtGY9Am3FmfiNFTT+VaudqFF+TpsPqbRUEU0INUM9QnNCBgNUyzNd5WG+GsrYMT0qiFeKDhAZklBTHdywkrueBUrBZWb2wUHdiE9pG6vdXl4CAbPrlNdxO3yxKl4AKizQxVo8xf7fMhzHrICdZBilwdldpV5luxThVOIfya3Y9WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFl18o4pr30NylAjpnoJBn29A0AJGzHDO6CO2xsS3BLGbccCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPoqIeA1IHCv6E4eVTGUE/G5oyoIXeJbFuwNu9pJr5KepciTUmVl2NyLaph3YSB0q0NBQUlLIPgxU2EM6jlg+dX8wvcQ79a/M2OHAgZShzLsag18ZZFxsrfzEuVWm/9dEFRCWbeSOoaDeYkZzDDBaT7wAFqnNEY7AP2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTLMCHQ82jTpQLtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXet4ukHksUsx5UQlm3kjqGg3mJGcwwwWk+/cYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaLFFatjDPCWzBUpe48G8UicKyjWNGQ5O4FeYB5ioJUYgwFgsHfuuaTDABloB0liRbp5R1LlXox2ZF4AjPNeCbtnAAWqc0RjsA2sf3ioWwd1cCOUu/aT4tHRMpVL58MJBQswIdDzaNOlAbEegyaglFcrk/Zu1ZGtBjxhrvt/y+YAd+z2vst+xJ0U/AaikY3kVDn29qKkoTGZVMX0H0h1bK6jmop/JDB5dF7xiooMp8WxaCydMKLoRPvEpCbjHIfzrNblg5fuBTrJoMhyPmT7y/3vND+i0phFmJue7kTKg4X1c7H665ic4bwuoNfGWRcbK3+gr7T+/E27juHkcmlnxQWBqORwzQdMkxZDRDzKAm9d6wJQiQW/mp7erSgwwyJbaSegcFQfpx6So+u6WYUl9e0gY8N6x7csw+o+SAElTCEGyCnfuWxyzru+sNWZ4XQCGlRxHLifkb0sG791WEgQYy70FSl7jwbxSJ8iMzdoDpUuKajkcM0HTJMWiAiNHs4agN4V/WU3qpuprnR2HTmeWNsrkSCKtN6j5A/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8WlsSdjcKS3WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFl65h9eL/S1rLOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHKGpZjCaHs19eswNMGaW4iR/FJxES+W2uyJSqCvee3WvmRXZEp4UN23eQ8qM0FyDJNmzfnCvpTk9bhdDjKl/Ez7cEVQvmZs4ZhxCvea/bRFrDde8ENKgQJ/Q8z2P5ELsBXzIJTRiSvqzN+4z/c88WUg70Qkv4MmFaG0JRNmyAH3Tt+4z/c88WUgdJicLigQEwimhxB5IgR7KLSNxaIJSBYOjtAXWQkz4pWoNfGWRcbK39Ctw/+nHcWLJloUTGTMtyXn/wrFhQhdymo5HDNB0yTFogIjR7OGoDeFf1lN6qbqaytVLw03npJYWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmxENE1poj4uOAJ5tY+/uqVvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx/UgfHzaSbJTFjldOYbCwsMORnsnb0fiwFEGJTkliJ3M98F6mH17CrexznlZe+itMGhSVUHuwHBahYWAR161KjU6AUrJpye4vLxXxvnwYbtqzxO7EBtu+KPeBG8KWa740kKxaDasfPpti/QZxTA2ygikJuMch/Os1uWDl+4FOsmhvb3i9iLwPrAhvx0ijQI5jzQ/otKYRZia+rgCQwqT6QU3MX6j7b5BtINPA6NourjgYa77f8vmAHaW35LmpvRo1dlwxxC0lfUYsH6sQ773h0N+pvYkKN7aIfDoUb8+Ic19fgIcbEXWDEwnHFDSwH0LLjaf8vjpHQYGQ0Q8ygJvXemFmjN23bm9wH6kFBR38jOG4EkG4xCRtzI6ubadH2ZK3ogIjR7OGoDePoZw8slvU/kc0YbXtPhqQcEXaU1pdjBZgZaFwY9tdizTPbYcyauupi1zrjXFtghQTgIHSttikSyn1TzjdVQn7GrSgLn7jD9CK68E6rjNXlLcrUtDe9UIQJV9ui98xHoMwwgxUJiDsGTNSC50CghXzZQ2ksFQBW/t20QnqtGlOZAm19uk/+xnMcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxH0nTDT+te3dYHeAmQafCVbWtHAtZ4q5p2bDWNQylDsBho1fMGbEvhHX51YzsqrFPgOVWtiUR6FRvDQ/OYk+OUWFyl6R4uu9tIgpIb7wqtWT8H0IhXtfXRQ7sCtl6ZHmMA0zE+qSrLhG90u06ezkn1Wp5L/I/qh8qw6H5bbxwJVMDyGzSYE4mShCAwT+5oJzE9kbV1of0WE6by/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOys1ZhDP6lMOpbTdG2Xipm5oyoIXeJbFuwNu9pJr5KepciTUmVl2NyLaph3YSB0q0NBQUlLIPgxU2EM6jlg+dX8wvcQ79a/M2OHAgZShzLsag18ZZFxsrf8bMZjqtUqowuL5sqWKTA6btwcZyZxxott1OLXHeZwhgETOWt0KBunJJ3ezUKUQNvZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYcQr3mv20RayRjGUlDW9J9G7WfqVfTgE2papsv/i+Wjg9f3OXpzhVf6g18ZZFxsrf8bMZjqtUqowuL5sqWKTA6XHz9ibeNGNAiDDGWXs9z8gaOPj4PTgm7+u/XPT3GtuzoSSPfVvb5wjSz5J0sMuXzmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa3AF1QC2M35c/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNbwb5RoGmEZTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyUf7ZcmeleQMxixVXOneoKVubSshGQ7ITl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGbJW+t9q00ZtJ+VC+Kd0F0sjGH6zOWYYzwg8QQ46zmxgkWGz5Pqa8LcGnkhHOWLndfeHv5fPyuFQSCi1UT/oEeQjtyOtybz4Xcl5fQLzHD7DzVmJzPpVUyEGjj4+D04Ju9f9txzzDmrqQpjuIPb3Eq52gvpG5cakkBtRd9iJfrOFNJH4RiFSfrKeCwfEp2J5FiboR8KKvMtE2OfTLT3e9rBuWDl+4FOsmjH9CKzhSnTcdPi6uk0GLKYNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOyNdPK8gvM7bZiaoqzMNXVvaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMuOdoOv5H15gMZVjRDxbTIFfzlp9Qg9NWVEJZt5I6hoN5iRnMMMFpPvxrgyE9IJwdgnYdX6mqL8wneP0N/uBkPMlX26L3zEegzDCDFQmIOwZgGwFmQkytbgP1ziX8hdVw2N7AhKNvBXLfCf1a1PYXmtrLsSh2Hw2xeEkpZ1EwtkIlhjpoPRdHjNN3C+LzYQDrJrJYspl083thztHQJ/KRlQ03iPskC6pCt69z7ciin8I3L7iy/OqQ2MEvkU6E87rjtI92U2r37AzoIEZQg7ASVOzxO7EBtu+KGqObKHokHBEMHiwATbD+Ki8Z0nXPMNMRhE7nNp8sszc5iKqJZa0JmrI108ryC8ztoG+aJnn+DCyAhiVuCSSNr803iPskC6pCpDRDzKAm9d6YWaM3bdub3CoNfGWRcbK3+ain8kMHl0XvGKigynxbFot16fYShoRjikJuMch/Os1uWDl+4FOsmhWOlUA/aj4U+EhI44TOkECrWusx+GLzYK6NMakaRBDLPCDAdI6K1zoajkcM0HTJMWQ0Q8ygJvXesffPy3ykWGRwx3aF1+LE53DTSEmGMKZ45acAGSF9jAb2K6hMdSPTRyVGm2Yy1/pRSUBzTIx478jlLE36kooLTC0pJAd2bC8Mk+hLtsQRDTUk0o6WrXnH7r9wJtSRXW75NWiqZnaehAmqDXxlkXGyt/BsVTG/zAj6tmJqirMw1dWdg+mmYluNhwCoaK7N09e5DTeI+yQLqkKHW3/B2Qb5M/tDesA38ry3ejxlboWU3JOAEpUG6CU5b5rHszq1lh4rmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa+NZzxld2Ok1LNQhPTsugXpMpw1WPUpsr/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8WlsSdjcKS3NrckhA6IJLEpJJ5d/icRvuzFx2oeyBToH2FmcHgzfk3Q57pjagUkkTxStOXLI6x8Z+40czJexoYFSl7jwbxSJ70/byzNr6MKaLZ21VYfjxH+J3a3ILgRbAib78JuTJdWj6wPS/y3dBqVkhSa32cs4NOZgk+wyD5DTFc+ZFbYaF+91ZxjHmU+SOEhI44TOkECl0FgRYVgViGcc9/L7IZOMSjfqPGNwc8LRFUZcPgmFr3XAfbv6lmCUB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC7gcnfz73q0BWqkud8wbS/IZy13SH1ztbzaUEFn+R72FPnqGuqxTSbv0Eh9mGRVt8RXhOmcqaGhX21pscx5UvVz4WPsQDweHd5IIFX2mInnt1qH4OPNW7bySbCzhGks5OI7l2KdYD87KAMq5V9IKK+pri17tNC1sPqIc/j4NtRsPE/NKE87MWDeH+mGfOlMxOW1llzl18M+pXv8Xy1b5U02+zpQFo/6qwFn1vjyXOHCP8bA2TUH+cn4p0AkbkkXte3egLM4xhJHAwSgFEIWCLSpYkjLTXPUhL3pLy2ww5fkqhCAs3TiOSrGcDSEvM6isbGydpivniVWNRFYo8bw7Ct9Z4SEbJbBobcCmF5t7JD4S/yu4BfH8hPz/Pp+HPOKCEry+SbxqXfl/B8Q3rfPNbTVyac9JRRGayDObwTl5Baxp8ycPavsZ2M93ksUDmdYbCs1QTucivDx91rp65cg9fUqCJyiKIRzD0/8ruAXx/IT8y5Zfu2CAIiqcFmUMNY9FzR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/X0mFXQGDwUBfxxgLW/DpkietI52dApanS0ZwazF+DSia1Dv3sAhvWmfnNRqgv4UiYRGFaybmRCQWc02j3u+2kOy44C5ZqFQCn5vz96kpWbarmDIzkr822b6s8qwQE970EPDmeXSehv1knBXlhDPOgjbPf3JibGS9KAiuTcO6Px1knBXlhDPOidKCAKe7ioPLBQFOQvZ3yiVjW1fM47WbunY+wI9aowrgC6kcQC+v+PygDEbahTo5nXqdpuCbaDKBQOrzNqj4aqmcxFPaH1VlpawYxusTCt1k/fZCzPjHVmaDHA85r5sJm9Zexg2eOYx2FtdDrFhFIv9215oa1VU9xmida45vX90O0N6wDfyvLdZ4itJqwS47xMSjw2G8mDE58DpgLoxhi6Ik2IJ2hGPYqcLahDynC0qMEfppvqcUz6AavDmDTROJHSgxLdGV0Lwmm2mMkhPMtOrD1oOhUnp8hO7JRb/x7EOEiy5SHYswRMpVSOVPa+hxq0//yLJZNFE5V3hyOyNkFbNXqcWlKuB7g28Aqfjb0yfgFg0CdygaSDn6ADi5zKCB8/AaikY3kVDl2ntTTj/8rdnvPZszYH98ufoAOLnMoIHz8BqKRjeRUOEIjuOiYvZzme89mzNgf3y5+gA4ucyggfPwGopGN5FQ7kR5TJwQr3X57z2bM2B/fLn6ADi5zKCB8/AaikY3kVDowOtu8HfkzsnvPZszYH98sINkwj4mslX2dAD0Fzenj9JxySuyuWh3sjy/wmmqpxBtz0JJUew4U+IpwhbRLiR7iPsZ4QF178O5TOxVf6qMnZwWFEse2vnPb+J3a3ILgRbHS3mX8pJVcMuQ6xY9qr2zkomfIY+Y3JZuHDJoDEt9A9+PXSoq6xkzaVhqsillAnUpOIIHKIWQiri0kWLnusckK6maR0RWksW+zfWsfwbxlzfkxUkNGCvYBgRgpuDZ29GNIKA7Ic4jbmrZk23b3pB/JUBKPN3GUEFtb9ASa5UQIg8UYeBz++Lb4SGMJtKTdcZ03Ptiefzb1PGHGCofMyG21ZoW/GvRb063sDzbt9n/3hhk+GvQexBgo/AaikY3kVDoVDCvRAw4KkJh/574MxbuHTF+gUKaDl49TgML/uKE+co3ZuRfEeRrlt4I1zhKJNEuQWQJ3cl6QlZ4itJqwS47yJWbp1N0EuihhxgqHzMhtt9Ibr4nY2v1Rxrby8Y+blW3GhHSdfPuNhcQJL0/6MrJKeBXXxYHpQ+/WCKtFaAB0psG8Yb2H0+TaawCCQAbl/Zw13upk5y+2NNp+ipJFgnO/C4OEyxUpTDzGkUbScpd8XjnbZ3QkVxUmY+J4/Sp0GR/vcFuOei2kg1q2+TcODnANtdCwTRMZseqZ0ioxXultPAT+C4N5bcirsY21T3uRMTZxqJIHSnBRTBKgVltCS8e4D64a1JkBbq4522d0JFcVJ71BnVEfb04JpQKpSyhKwaf6OBdxXWr6KkGPFOpO5PQmmwDx43dJ3DQS0SN/g8i75+u6WYUl9e0ggLWZKS10MIK+HjxaB4B74rR508ZTGndFXX4rD7vXyZrtvm0WReuEKFIjp1DOt+ycQi9NfGZPExrTEI9OwCNNcyD7Se0O1dg55xmXMo05cKjjgq5bS0R06bUXfYiX6zhQLyDUTgzT9Ni5sD1/aEdimwgg/EGv40FCmdIqMV7pbTwE/guDeW3Iq7GNtU97kTE2caiSB0pwUU3Ntylp2zkP0koejOOHQ5KPzEs97qfveGssrSF7kR00hyE4aJiUCGxU2n6KkkWCc78Lg4TLFSlMP50r/6zZg8QlTxP7IE+yf6ZKHozjh0OSj8xLPe6n73hrLK0he5EdNIchOGiYlAhsVNp+ipJFgnO/C4OEyxUpTD+dK/+s2YPEJpsQtPC8UiDcQrexD2QBexprAIJABuX9nDXe6mTnL7Y2V/wgWEVM4l0NxG3YQWDVJa9CKQlY8TsIr5MLZhS3k9gfe7Ma3sYMPuRPLKQUmcjw1Zicz6VVMhC9Lz6GPyonWGfnUZFm/vqZ+cDlC3s8/tViCACHbNjEq8kyiJFHAjB2TiJ9uJ0l3RDGVY0Q8W0yBf65pTgrPqZHIPtJ7Q7V2DhIaA38op9sp5BZAndyXpCWz/6I00m5OwNx4dRtVkKtQHEcuJ+RvSwaFVSD1FKcXtHIM07ImKul/NN4j7JAuqQo9LaGidc4WL4FEj6WZn/ACCy2C9Wo5yIDTC9EFpUA1GF/23HPMOaupCmO4g9vcSrnaC+kblxqSQG1F32Il+s4U2wPHIWOU7dylkMm60A9Ng/7+DyNDUNSsCPwjgN6ZBDDrdOz8XSMszvWzKVV7jlU/WIIAIds2MSryTKIkUcCMHTj19FbV2LuYJQHNMjHjvyM9LaGidc4WL7HNsaUk+PHs7Q3rAN/K8t03I88UVcMKtWvQikJWPE7CIr3eDC7WCQEgFxsc7HdT9fL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZdx45Dw2/ZuhgoGYRI7CS9JdDD6unk4J+eUZT5ooO5sxZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk7T7055ep4FkQ78dBCdzO2PrMDTBmluIkfxScREvltrsHDZMRgFfe1OrGISi5pGmy8GeX39/rGN/heG7408NWDUq3tQQowV1uJKHozjh0OSj8xLPe6n73hr1sylVe45VP1iCACHbNjEq1qk6FYBnBqZs/P9zr8kn/aI9EAkCE4YeUaXl6z3PdmRq5SZSFuyRgxb9ZF9SEVwiwgg/EGv40FCmdIqMV7pbTwE/guDeW3Iq7GNtU97kTE1Q0Eb6lzyhsxPXNYKURi0fhcuOI5OOxTLSR+EYhUn6yngsHxKdieRYm6EfCirzLRNjn0y093vawblg5fuBTrJobUiOaRHZTlOnQedCAf46ilEJZt5I6hoNu3BxnJnHGi23U4tcd5nCGLOm4GNjZXJtbUiOaRHZTlNBUGHLZoXd0FEJZt5I6hoNu3BxnJnHGi23U4tcd5nCGLOm4GNjZXJt1uhkf50lBKQweLABNsP4qJXZg+ub6CpKQIaAy+tSTHE37Nk97b+6rmi6syZn5bD0l7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHHgsHxKdieRYj5IASVMIQbLUFI/NHsjw8MuT6SxIGKL0GGu+3/L5gB2O7A52IMODWZ4Usu9uqZ+vRyJFwQgHYwnZdrxFpecIx14A0YV60dR61aKpmdp6ECYU19kUAs1f2hhrvt/y+YAdjuwOdiDDg1k+kHD7dnMnelLeZU8aZXW00xfoFCmg5eMHLaZSE65mbr9K2ULjqWWOYD1RXhKmNewYa77f8vmAHY7sDnYgw4NZPDyN/gyVX9VHIkXBCAdjCY0yqzUs37pLXgDRhXrR1HrVoqmZ2noQJnZwyyiJJqK/GGu+3/L5gB2O7A52IMODWYn8BfXoPIeyRyJFwQgHYwmNMqs1LN+6S+0uCSM3zXXZEYmgfEdYGnqyqDSVLaF7LLXFtL96Z4yoHra5KgNSpAG8xWw9WDkBHDGc3nODWG+mq3MVcwACw5XGDUrUHXao0T8BqKRjeRUOeuDIlcBEJ0vIThomJQIbFcCWchPbR47aPUeUDfo/r0K6TPTLoyrwdj3jkIDRspA8/1U4QQ+VIc9NSMqRA+KwwA5GE/InM25D6vikZ+3eQoiJVWE6BiRSTtpyo8QcEA4bZa5ncP6fE1YVBFNCDVDPUKZ8yJQvahrPVNHrwZG0oFCoNfGWRcbK36l8+09yWfa4oSpQgBt0sRJo5LJa3BdcWK1ZZsWEi9vE4VU00TfRW40T7biyuzy8kw91bZfIhUf8gnh+HfoOrPn/VThBD5Uhz8EgPNE3qY0XOL9wd2D6GbUGwJdCtvbRNo7sDnYgw4NZMZwzc9sXDe8Nu9GXfU3btYMqS9j75lvBvoiGCRllu1SSoGtWHrMQoDV6nFpSrge40jLsoS0eyLpgbHE/GW0UATB4sAE2w/iocXD5fgOfVn7DHdoXX4sTnRa7zoMzwU8uQYrSQJBv7P4m4Cs6NtgPEWxHoMmoJRXKJ0AGsvHSsBgfqQUFHfyM4b6IhgkZZbtUkX7Y4xliR01ck+HXxC/4p0O/HQQncztjRK3rZqU420jy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNsAfu4fjqbOnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTDSn00tWjyqnbBQ2HJfFxAo7l2KdYD87KWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPzD7uXbkCrc77a9ocBJ9+mJn9IO0/LopHDt6XhPrImaub98+AaJaEDsG+QROCz5dY2uXO9FnjWKZPKwZ8gNmtnmNjZPrsSz73Lk+ksSBii9J7WNoaMRI3YQw996IZF2ACn4qgYoYLr4bMdxlXKnJPqntY2hoxEjdgubA9f2hHYpqfiqBihguvhBXHsXM6KekKe1jaGjESN2K3H4DQRhne8Qw996IZF2ADrslX0in546XhYonbMS0/WiuvBOq4zV5SVlU453hhBKUf3rTN19VgbYWaM3bdub3AzUgudAoIV8+aMqCF3iWxbs2P2dk0hyehwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk5ObRzSM0cQs8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEfSdMNP617d1gd4CZBp8JVta0cC1nirmnZsNY1DKUOwGGjV8wZsS+EdfnVjOyqsU+A5Va2JRHoVG8ND85iT45RYXKXpHi6720glzZ3aJTg6SSUBmcxnxZa/2m32fISQbGlixpxRaEIXoDObwTl5BaxpH2KmNs7ClyHdGk0cRHYrFTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyDrBrJ/SkkFFsH+k+A/rBfaFhYBHXrUqNZ2rqr7iK/sxqUKiyjuoZTiem/tdTojcxABpLkx4DeSAfILcYi00x4sYtchMc4mmUcQr3mv20Raw3XvBDSoECf/JLt+zJ70279qoHINnqNTQT1zWClEYtH4XLjiOTjsUyb294vYi8D6zb1sn3BQ3qCDSc3R/HQ5ndZL+814w1rJYvxMuc4I56TvGED6cYfjdoNrlzvRZ41imTysGfIDZrZ5jY2T67Es+9y5PpLEgYovSzxO7EBtu+KGqObKHokHBEMHiwATbD+KiBCNICj+LaXxE7nNp8sszc5iKqJZa0JmoRoNO9lCVJF6Jl2iG0D5ONImHH5zsj2+ln9X/6UGEpdr3j9ojp5x60eAn/Qv5qHLuQ0Q8ygJvXeuyRsxnBe755BUpe48G8Uie9P28sza+jCjmpvvq5gyAjV5gHmKglRiDAWCwd+65pMPGzGY6rVKqMo9RQUZ2e7ZnQ5YzjkTX+phFPpUd10VriKJ6LZqHVfyMASlQboJTlvsmhdMzPTwDOzEE+Z3cjImfAlCJBb+ant6tKDDDIltpJXRVbE9BqVFm/EUKWXiWm56g18ZZFxsrfVHAAl8ubAFhjLo2ZatRFW3Hz9ibeNGNAgH6LEA/RlEy7zba5wbSWgGqzsYFhmHXtqDXxlkXGyt8EGIkuMMZSUPrulmFJfXtIGPDese3LMPrGkgfxe4lqk3EK95r9tEWsvq4AkMKk+kHQ5YzjkTX+piZeRju76fKYHw+rdA37MM01nKCnelJtRjwu599uOMKZvasFSgZCszDjdhVjvvgpIWFmjN23bm9wM1ILnQKCFfPmjKghd4lsW5bTnVvoBnDXWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmmUPGX3ApaG7q7nKCHnP/5b5Fy2boKmcN8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEfP/ZKWu8LWsLQI8txV7R8uhnFgLqlqUlUmf0g7T8uikTmdjCz+epvdf0N2LXKhc5/X88nixuUVIMk0flCMwg9o1dZ0prWwPdDsynjmpITlE1eYB5ioJUYgZjySmeLaPsoMHZNkdaymPV/OWn1CD01ZUQlm3kjqGg3mJGcwwwWk+2Y8kpni2j7KDB2TZHWspj2+c8SO015jYlEJZt5I6hoN5iRnMMMFpPv3GKSbJQo2s/eBG8KWa740kKxaDasfPpti/QZxTA2ygikJuMch/Os1uWDl+4FOsmhUDq0fdcnxCjPWMftH2FdgCcat9FVlXW6SHPgP+RzESzV6nFpSrge4SylxqcmnpefvO9a9FEIgEOEkpZ1EwtkIZjySmeLaPsoMHZNkdaymPXQH2NPgWfg4Awl+HhDg0WgH5xJEZfU2wQwkQ3LgW499JNHBwqklmOSCEpjJXQAJNHNJniceC2vC22RPOjd1WnezpuBjY2VybWF9B4gUjchiHNYQoPY+k1d2D6aZiW42HMl6oOggoczfE7EHPXDb1nxYAntEFGTxwNI92U2r37AzwyhKE9kaKyX9wJtSRXW75NWiqZnaehAmqDXxlkXGyt+tMg/TH8AwMIM+aEC2mLhmax7M6tZYeK72iuplgCAem8xp7Q1cj/59xu8wRnKuEEyLVA/mweBCLjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRywY51sn0lC1P5t6Y7pHXqS5mo1m768rOuk0T5NylBw4o2za4ndYsaWbZZzmiwPIDzwyrO01hlSvVgbHE/GW0UATB4sAE2w/iouQsuVmomRn9FAomrFMgR/1rgSNBvfq0O8iUoVEULW/wAyrlX0gor6h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC5phREvPgpvHBpIYeA2rj5kBghSAkob+RtcYPplyneb5FgMEVi6IXblsFshSxqvZfeXR15LUBDW8Q9t/s4jiy19tVJMf5fqF0qOH/tgCkP0SSPXFdmWcYds1ELDnURHRIbyIU39K9JJ7/O8bOCILc/n7f+RcPO0h2oArzA5qdqOTH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LxrFahAkPT9XzCterMAWpOmg61dEmrqcrGh5U5irJnyoBYNAncoGkg3cEuzEuWPSs0oCK5Nw7o/GPmErSoWFZK71siqWXvrBM16nabgm2gyiwjo6nhJm63zYNGTiJQjXZL/eE5UpRoQlGeggn2DaWljQ+f9WA+wEPL/eE5UpRoQl42s7fuq63wfiqPFZR5iDogngZTYpYIfZh/AK6jyUPsc7W+/RZJSOcly6IveSStcB532mKjRs8Ag1fLXh+Rnpy0CNhofJt4MSHKqogxnApEmfgrpUCcPDtPSYisw/CJsf13HsjB0ZnrYpceYJJa7kCwFgsHfuuaTBcKPIkz14E8/yckXe+72PbXrgAWuYSn8biY+JWwK8YF2G6OTbX40yT1ph9EJwygYobyVvPnftlh76J+dnhIo92wFgsHfuuaTDvLBREZBsyKSznCTT1KMwT+BzPnHQ3hXBu0UHDi+og7FMoHBO7CYg09dx7IwdGZ62ZJKYLkt5Nkm3kfBhmCLGRXCjyJM9eBPPUqcS18oLPlSH/Az7EINaUyCsc6J41TV1CVpf0fc8K4MPxbAaJM4pXVASjzdxlBBZG93gikoryXwjqK/Yt6Um04m/RGRXCtaaKH4/yj+If+fawMr5DqsStZYPMjwdNq+CtEZK7kisEEh2DWy5n0Tr/BMlZKI/I2EqsPWg6FSenyE7slFv/HsQ4HyC3GItNMeIa+4JkKGk8XJTOxVf6qMnZwWFEse2vnPbpG4jXwUtOiPEZM0BP048II8v8JpqqcQYS1F+P0jKq1cMd2hdfixOdcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/GiMFB2SyS1+ILfK3xQ3PksEfppvqcUz6AavDmDTROJES1F+P0jKq1d4SNc73+P83Hdtxg6oOGCMomfIY+Y3JZuHDJoDEt9A9p3F2/KZDZS1CQ/UWBIJ97/83YxNodUb3EWsoLROZ2jlYggAh2zYxKrOm4GNjZXJt6RuI18FLToiYAIPUc68MBrT//Islk0UTpwtxCu/hW/x7roE+YpEbxffIsUQ0jlrJrD1oOhUnp8hO7JRb/x7EOI37qMTokd4LNDt7WTzRCmcfSSbQfgTQYg+w5CPuIzPya9CKQlY8TsI6Sgfx+Tritgwdk2R1rKY9KyiyGAu62Zo1Zicz6VVMhCi+G04JfRlAVFYclhD8d4cgejfQK7nsB94cP9e35gy3vtXhiXMQYGMSNujLFNzqC+00Q4dWDA3cYqUN4zQ2F0vCCkB/cWqSlmpGPxRfAM1oq0FBeFAOCWIe9p3K6OuLN2xYNjq+U59gvlkP4vG3jtSioOnn/o5+eWUx5hnADsYsrD1oOhUnp8hO7JRb/x7EOLY8xLkcGBQ5WmgBv7vT+q08FF6EgV4/kC/ErR5R46vaNWYnM+lVTIQovhtOCX0ZQFRWHJYQ/HeH5qBEytoYnUao3pI+zy8s5SHVh5/7SJqNZvp0Q3jUzh1xX2xf0wa4olMzMTd2VbLAHYNbLmfROv/wNH0AApHhwBI26MsU3OoLq7g57ipYIsn/N2MTaHVG9xFrKC0Tmdo5WIIAIds2MSqzpuBjY2Vybe7lwxehGWA3KVP553NK9K6jwTGB+vCg0JRSCAJFZ3PKMCAsaLkc9sMgi9P5Q05ExOagRMraGJ1GqN6SPs8vLOWKRO9tjjAS+LKJd520tkKhVMz8s7lE/N2Bxl0y+KwUu+zfWsfwbxlzfkxUkNGCvYCVoorist+nqiHYJrK0pbyhkTk+9SxN4FUNfP/1CBud8VW7inPYRzEO4m/RGRXCtaaWZgZUdK9YnOdK/+s2YPEJZjpuluFYR5HtNEOHVgwN3Kw9aDoVJ6fId4AgF2l+b7GSrEnbZljYtsNTk/uijlr+yq+cHCEUHmxTMzE3dlWywCvkwtmFLeT27aAMEjQ9WoLjfxYuAdBcF7KbpNn7hkAvlM7FV/qoydkji9MrIcEZz2IKntpxNMntDbvRl31N27XnSv/rNmDxCWY6bpbhWEeRy1xXY9xNG3iXv44E5MyRAM3NonL3dWzRF/O8s64DUvI44KuW0tEdOnt4ahAdjknfyNuIjjJNURikoWTY0fIsOZlzPYM1YiDBmLeeZbuMJ5EcRy4n5G9LBoVVIPUUpxe0kqxJ22ZY2La1uyhbt3oYhKcfSSRK3+yPPc0I368GozilaqHQ6HYhZedK/+s2YPEJkshNSmg35UieuCv8EL5+zoiF1OttsAwHVFYclhD8d4dBboDWT8dzI+Jv0RkVwrWmWnw//gC8XDqZ7giR2adr1gFg0CdygaSDnGokgdKcFFO+TTt0tEZq+/jYJ44oWZlsMDvPQvnae4oCLmfIM/UTQFNZ+VBB5qxL7GNtU97kTE2caiSB0pwUU75NO3S0Rmr7LUU6h4wsofL9/mBJfCZDSdWZoiiFN4qHeSpTVUvYTNRYggAh2zYxKvJMoiRRwIwdaUCqUsoSsGlRUvaLaCwGKv3+YEl8JkNJpWqh0Oh2IWXnSv/rNmDxCcCUIkFv5qe3f65pTgrPqZExk8wvrRXYtexjbVPe5ExNnGokgdKcFFMEqBWW0JLx7s+Bd63Gxh9Fi0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+In9FHc1iKADHLKbpNn7hkAv9KM91k9syYt2IyXcILkWAA270Zd9Tdu150r/6zZg8QnAlCJBb+antxBqx2CKy2YTSX1eYZ5oBk2JbNXR2Y2XTvEae5HQ/VvXK+TC2YUt5Pa0kX65q+MC7v0UdzWIoAMckoejOOHQ5KMomfIY+Y3JZuHDJoDEt9A9FIjp1DOt+yevlaxpygmp0mVsn5R87rmOwgg/EGv40FBOQZIm7+zr2MLg4TLFSlMP50r/6zZg8QlrMd5VsR3PnWMF9WizK2bjD7DkI+4jM/Jr0IpCVjxOwivkwtmFLeT2kMFwoSn84t09LaGidc4WLxFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHWlAqlLKErBpe66BPmKRG8XRDKF8K3NC1sIKQH9xapKWFIjp1DOt+yfdv7czRvnKL97Wo1mKhDIgdWCm8N7aUUocRy4n5G9LBoVVIPUUpxe0BLRI3+DyLvkc1hCg9j6TV5KHozjh0OSjKJnyGPmNyWbhwyaAxLfQPb6hnFtLa1bd+FotoRIKEsj9EMg3lJqRcQoI1NNC5RgMawxBUxCOB3ICwvh5baNINk3fSaLMZtg8GVad2lsJriRFA+yTu5xiG9BGcNUDt/muS1VycFim3gqgczzEVznGKWXbI1w74mecNIPm9GswZnNcQ1fuzhGSqtzUcTNyiZjlOU8GPMsjGFGJPQOlYZmoO5dHmN06ubPPCrwi/h0gOmiBPozgbBitChP9+Gd8uqSETaNQq82vaebm0LJaASIpe9BGcNUDt/muS1VycFim3gpUZYUlQ5iaO5wJ6kWNLc6Zl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGYC3xAKIihfAiXJ89E6gY6/MTI7bmQ0eUTy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8cUnyYHq+c4njb9uZP+Vgro2jFsjiZ72mKZkUi6qw8jhgOtc6uS8kSgAzRUxw12Mz+b98+AaJaEDsG+QROCz5dYaeSEc5Yud15hSJ4nVh6Bl2K6hMdSPTRwa6vwQqgvpQldtJhXraTA6jRBmQQXz8GWoNfGWRcbK302jUKvNr2nmzYpwOScyB0cvZwDlzKIgxFKtq1msf1HBa9gNWpgrzmv1MOfjYH6b/Gz8/3OvySf9oj0QCQIThh5SratZrH9RwWvYDVqYK85rRr8y7cGcsx6NEGZBBfPwZag18ZZFxsrf6tTBORoJzQk994SG3n+PW2g3zfMriZWNUQlm3kjqGg3mJGcwwwWk+04QzMm07qCpw1OT+6KOWv5H4j/NjnSpD/aqByDZ6jU0E9c1gpRGLR+Fy44jk47FMvcaLydpsQM0S7519g7oX491FiiUOkfRs6a35DOqZ0CrvxFCll4lpueoNfGWRcbK3ygeu7196rwDDzjExFhGseGwtb5ZwCsOj0L2TqHljvVf8/TVDKwR8YQk4Feq0u3fyzLFtLit8MJf2K6hMdSPTRxSratZrH9RwQ2H1U3V6ysbYhuij7af+rR6c9O0Bg63VvcaLydpsQM0FQRTQg1Qz1DFQoAxFr0R+RE7nNp8sszc5iKqJZa0Jmp4LB8SnYnkWBojBQdksktfWcJ2ZgASfSjLk+ksSBii9Bhrvt/y+YAdGur8EKoL6UJXbSYV62kwOjWkPv8rdyGLqDXxlkXGyt/3Gi8nabEDNGrmsl3HZ+Tug13y4U0eCPGo3pI+zy8s5SX6j21W4QAy2oSI+CyoNq+5YOX7gU6yaE4QzMm07qCpJgudxL64SCh2E10HJA9hjS8HZEGoTxCDAEpUG6CU5b5rHszq1lh4rr2rBUoGQrMwXWjfuQUjOLeRjGUlDW9J9BlUettiSmAiC4WuZKNK8yMoh5adtxvxRSgqkwkNb6LvKVP553NK9K5gx0wYE6lyM+ejRt2PlbZPcK8cDIAbFwJUI5T45kDfWmlSVly39FTMXGq8J3GheZQsJuhlHhzK0QVKXuPBvFInuFiUdEgxo0WQsMYuPSU9lSC8SwZAElO9DsnVn2RtsT6d01DZW2UQ9EC8OIornqDi1LuuQDvoQhaYb4ED1lzpQg9G//g/VOp+wZqTHdpFJLBC9k6h5Y71X/P01QysEfGEJOBXqtLt38syxbS4rfDCX9iuoTHUj00cUq2rWax/UcFr2A1amCvOa/Uw5+Ngfpv8bPz/c6/JJ/2iPRAJAhOGHs5UIZCbh9wppKFk2NHyLDnoT0ubfAasdgKGUQfpLO4WenPTtAYOt1b3Gi8nabEDNE2jUKvNr2nmikQAyWKXI4K/EUKWXiWm56g18ZZFxsrfOCFIyjl+ejg8CJDEOXPWVOcQNKBewy0XFpYxxog+HqZi7mYxX0WepLTW8EUofh6+PAiQxDlz1lSYN4jpzhzDkb8RQpZeJabnqDXxlkXGyt/XyBR0RCvVpqShZNjR8iw5ekUSMJC6vfrib9EZFcK1poofj/KP4h/5Ipffuy3PPvHmIqollrQmas5UIZCbh9wppKFk2NHyLDnkXc2CYPoNbUCGgMvrUkxxN+zZPe2/uq4Ya77f8vmAHVKtq1msf1HBa9gNWpgrzmtGvzLtwZyzHo0QZkEF8/BlqDXxlkXGyt9vmWF2iuflaKg18ZZFxsrfThDMybTuoKm1uyhbt3oYhMrp7Sbh0xddtbsoW7d6GISPIc/w7vkqDRhrvt/y+YAdEPQTFGz2CFt3DCpm/rPLLr2rBUoGQrMw43YVY774KSEQ9BMUbPYIW9LsE7Qbac9EaPuY0ytJXczRZoACPjE2sUkv8pu6uoVyzasixnaPUTJ8gPwsN5c8KmY6bpbhWEeRy1xXY9xNG3iqIgN1+xvhieiqBtroy0ISzlA6TTOMdUHpORwM1115KjmXVBfK4hJZ3KjZPqsRiGA2n6KkkWCc76kKusz0wYsi6tTBORoJzQkisaKtRaw2LE4QzMm07qCpw1OT+6KOWv5H4j/NjnSpDysJ27ZaK3LWXGq8J3GheZRkVmFlVn+Xw+ecPZrntmq39++9kYXAo/KsNWZ4XQCGlRxHLifkb0sGlDo5Px/c7r1+nGsLM3sBVEyLPyOhi5paEPQTFGz2CFss0q2Qk0aD5bgSQbjEJG3McCP3rumN0oVNOMIRwaIAjk5RPjL/18fI8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLe+1eGJcxBgYxI26MsU3OoL1olBKSbFPD4Kn9CGb+fOCAqBlTDmmLUwcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JnpsG2pPCo720hUZRbtecSWFCRKV1Rxd4yEJF6wmy8A6Ap8bN8Q6wMSLM2iYdad9RuENbGpoR1eDl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGaru9Aw69EZmsm74WPAGRdyJl5pP+/w5LVg8M/XPHF9qDN8hwkaeXL9enkzBWt0tJvSR+EYhUn6yngsHxKdieRYm6EfCirzLRNjn0y093vawblg5fuBTrJoACNE63M4AbY0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm34sB73nkzKpqShZNjR8iw5dBgKUas318N2qGJ/T63OOE4QzMm07qCpXveA4V9C5MjWWMjqyhMq4FEJZt5I6hoN5iRnMMMFpPv3GKSbJQo2s/eBG8KWa740kKxaDasfPpti/QZxTA2ygikJuMch/Os1uWDl+4FOsmhyErauFowuZs0hhN5Hi/ZjauayXcdn5O5Zb/h0F1jGIpFfYFLIqsKzcQr3mv20RaziRElPR3NRSlA0dNlUkkQR6aD6fpe+v7CEHKK/IN9j4dNfh79OI2T0FpziG0dVJueDKDWQOh0cR8zJKgc8CRuDKwnbtlorctZ9tMtbL2SDlJDRDzKAm9d6YWaM3bdub3CoNfGWRcbK33alVH2frhx/O7+61WV8WGLgKtLGyexHBMklwdAJMwiZFZtQw4g9x3914vBOSJmnnLEddF643SlE+eQysX0BZBAh1Yef+0iajUXC6VRVMyaDtjzEuRwYFDlaaAG/u9P6rTwUXoSBXj+QksjuLPTqop6zxO7EBtu+KNZn81AuN/xX4m/RGRXCtaZafD/+ALxcOv2UEWSsyzn/KQm4xyH86zW5YOX7gU6yaGlSVly39FTM+NgnjihZmWxOQZIm7+zr2FcxK65ky8q3rD1oOhUnp8jqbdmcoQYqPN9yIvxc5OLJ4m/RGRXCtaZafD/+ALxcOlbCos4995JpgypL2PvmW8G+iIYJGWW7VEL2TqHljvVf7uXDF6EZYDcpU/nnc0r0rqPBMYH68KDQsExWvmX7W5O/EUKWXiWm56g18ZZFxsrfOCFIyjl+eji2Nm48XZHuKjjgq5bS0R06g/pCOhWYIWqUzsVX+qjJ2SOL0yshwRnPCf5gKa5jLihaaAG/u9P6rTwUXoSBXj+QfBhpIwv57iIASlQboJTlvmsezOrWWHiuajkcM0HTJMWiAiNHs4agN4V/WU3qpupr0k5NefRgwv7zhob8+jNnK3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR0llztVWLnrj5DYxCpQTR4IEyrp6E80Nb/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk82Mu6gurrCcKVP553NK9K4DGeepNR2vsgsie52kK+VirCWUbDj7YfvR+4b6V0VfM173gOFfQuTIIHtFAGNy5RJP32Qsz4x1Zg6OyG6bnoLJ5S7VhRRSwLjib9EZFcK1poofj/KP4h/5+s5+HqB7x4fib9EZFcK1poofj/KP4h/5T/rcVjJhcFaa4B0zYio8JEbVSH2QGsTiJqWbEMG9PrK6WFEGdh5P7HhjxeqVii0r0oMS3RldC8LQNO+VCg0OpRp5IRzli53Xv9281ooBjDbucdi+/J2AzvnkMrF9AWQQIdWHn/tImo1zGNq00RZwIi+595hQ5cfie+rN2J8ozW0uR2p43GIz8LyqTLJtk8MmMfPn0gsZUSBmOm6W4VhHkaZWQltNOn7SZjySmeLaPsqdTLLphyYjxC2ZCH5A5EhFpIA1GoM5+83/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk1vBvlGgaYRlOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHInM2jdy/gRAgL0kEjdIIoXBt0iTwmsIN7Vguiwp5cHh/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk7KzVmEM/qUwRTtjj2C2kY19M3ZqZelGvoV/WU3qpupr7Z36IFzy/QUfILcYi00x4udtI/0UeRgdZFdkSnhQ3bdyErauFowuZk/kMqEp6+Cp4YUHeRv16uTmIqollrQmasCUIkFv5qe3gXcylQpMNl0vZwDlzKIgxJKga1YesxCgQjEwLog94FU0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm3W6GR/nSUEpB+uHWPs/vISQIaAy+tSTHE37Nk97b+6rmFcV6pKQIgY/RR3NYigAxxSQiTI9fxSyrtwcZyZxxotq7z0WNseUXcT1zWClEYtH44v3PQhoFfMkqBrVh6zEKAjuQen7Od6z5XZg+ub6CpKQIaAy+tSTHHkQK/WNyYU+xpjN+NMLr6R6NLvPlfAjkbxhA+nGH43aDa5c70WeNYpk8rBnyA2a2eY2Nk+uxLPvcuT6SxIGKL0nwDziWeYZMxCe3/bKBZ8AzQAkbMcM7oIa/Q6B+bm9wxRia9YFK/dPm6E1sTrkWhZ4z2RP31HeuNC9k6h5Y71XxUEU0INUM9QxUKAMRa9EfnUk8RIO/7+OmxHoMmoJRXKLwPt1CE7JrEHEpJl7xtSvrqxCJ9pMY+inQkzyS0WZ/xjn0y093vawblg5fuBTrJoMZzec4NYb6ZigEUXHcYdrmxHoMmoJRXKC15MEywTNkD/VThBD5Uhz0JD9RYEgn3vax/eKhbB3VxlsT8DjpTJuqg18ZZFxsrf1uhkf50lBKS+YtTgXdvGiziTj5XxuRg5FpziG0dVJueDKDWQOh0cRzGc3nODWG+mndNQ2VtlEPSNEGZBBfPwZag18ZZFxsrfrTIP0x/AMDCmYURHNrLDk3pmPJjHlS3Ifc1LVKQQE0E0PjlidWHKn4szaJh1p31GKw/ZqTnLgIw9SfT1XUhXsp8tqvscB90rwJQiQW/mp7ebmzzPUPBXvZJIJff7NywdUIH2xnbSDJLThEiZfzyVFkw2SmqK84fCWhfB7jTkExej9a4NkQvW6W/yrwRR6EI6WbfkqibTtoChKlCAG3SxEtzUcTNyiZjlyLp3vGdAsWvQGI+luyLZunkJ/VWHM2iFQkP1FgSCfe8Wu86DM8FPLkGK0kCQb+z+JuArOjbYDxHAlCJBb+ant7I1x/CbLlKhYWaM3bdub3AzUgudAoIV8+aMqCF3iWxbbm15BjSpSR7NqyLGdo9RMv+o6hWtmGM88v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTI9fIwYzQA4GVNSsNNAgsEmKARRcdxh2uwJQiQW/mp7da4fNC4Bg8vFLlH1vJXaFHZQqq59hX/k2CSKAiy43mJtAYj6W7Itm6N7q27ssNaShAvDiKK56g4pYlHfB/zqZzxAHZv+4XFSx1U6N+5sUz+mB3XgZZNAPjTkGSJu/s69hx2YiI2TiMCMMb/Nwqih1HIdvHuI01VL7bRUNtURyxAV73gOFfQuTIaaL5U4lIBgMIozZ/XwlqSN+3BFUyRUa0rihNi4/CQUi8keP8cRkN9HZsepsqC2cU85vZefzHUMKRAexMN6ip3gfwF0/Kq6EVi1zrjXFtghRcq+c37hWj0j6TwSXYrcQN5SYuCB4yNtl5Dw8YqLlE11jRn8kLVU1sNHvHthUY5liOcLDd+unG1ZnMRT2h9VZaT74LuhviUVPcmeZty2DsZ0lu4sES4sFVGGu+3/L5gB10T/hMTF3EP2WFBpwGO1URuV9MKuzNnxuoNfGWRcbK32Z7m4twi7zVraPLyK57K85UgqPyJhcdmA/qKq6oXwI963Ts/F0jLM7ciwrbHiNyxwaiOcL9xq9I2tWZ4ublbysOjshum56CycBYLB37rmkwWLfuNP5FCVhn+djsM4CPbRhrvt/y+YAdHyC3GItNMeIffdSuUY3eUAIEa+1M42FMqDXxlkXGyt/q/B1JkFXPe8EPr1I7wXY8zUXhaLMpmYTAWCwd+65pMBUEU0INUM9QxUKAMRa9EfktmQh+QORIRTrs7IZ1ypQho/pRr7mP7MCoNfGWRcbK3xLUX4/SMqrV/oZqqYq6rbMaNf+4+Qw0BP0UdzWIoAMcv9281ooBjDaVd4cjsjZBW8N9WS0N3Ar0TKtILK4VGM/QGI+luyLZukLQhhfkIQJ6Af1sDL6Ym0qNMqs1LN+6S01KMv0xgpOsqrSHE67+NZ7AWCwd+65pMBUEU0INUM9QEW9fEec7vvM6k+0KUa+B4kLQhhfkIQJ6lhjpoPRdHjPDhxg6ak1chom1hyBT2RJQij1RmOdVVdanC3EK7+Fb/HuugT5ikRvFiS3oK3vtfvM8UrTlyyOsfL/5cgVXFR2tZjySmeLaPsoMHZNkdaymPaxKI6Es12nE1IybwRAazvO/3bzWigGMNqcLcQrv4Vv8TFc+ZFbYaF9ieCBrHGhoxvypk2T6X22ojl5YD7ZmhyYIMEmt5aG1PYYg9jBaTAs0l/rJHfRkNDh2IdBu8jtk4sRorHQ1ijfAj4RU5H9cQomF04Og1lJRyaKZnONASFztUzThJ1N5BVUatKAufuMP0BJXiytiAP06gOPwyC6p4zLiQE4QSVh1bPI/lEFVd2N1n7/xfjsn7fyoNfGWRcbK36Prf0CC1QVuj+K97Q/MpF8P6iquqF8CPY8RtM3IA8uKXZErJTMi5gSLGTIcb5Bh23etRIiY0bSldzdvGzueikSqkcf1AhnVK94e/l8/K4VBmuAdM2IqPCRG1Uh9kBrE4kWyOTE2UwNchBdE73GNEXhycn0fczLPWC+595hQ5cfim6EfCirzLROsZa5+kF7nponHHVYrktigRIoLn9egg/BnQA9Bc3p4/bP3znU/tfvrUIJyZoFUkp5PWdlcJT28jQVKXuPBvFInuCMKRpSZEwXnnD2a57Zqt/fvvZGFwKPysnbOiShnZxti7mYxX0WepD8BqKRjeRUO6MkBiFfvRKmVNSsNNAgsEtjsqEvp2K/pwFgsHfuuaTAVBFNCDVDPUCu96RyF+yv5azCcevyCvg+kmn8ia1Gt/Bhrvt/y+YAdbEegyaglFcrLyuPmr9FUIB4C6/8yiKr1UzwCUlzmNrNPWdlcJT28jdMX6BQpoOXjOaTkjrgDvn5583upOJS+Ixhrvt/y+YAdSLLlIdizBExC2906JuabGs1F4WizKZmEwFgsHfuuaTD+J3a3ILgRbPmQvJ/Gtg5qYnggaxxoaMYP/9hTuIR62b/dvNaKAYw2pwtxCu/hW/zG13tPUhWWZGJ4IGscaGjGatZfxrEvPYbAWCwd+65pMP4ndrcguBFscHvbVgXuI+EMHZNkdaymPZgbWnLWx/bOQmYYXfngN8oBF5x/e4AMjYZw6vEYBeTFcOqfqeMO22XTmYJPsMg+Q3uugT5ikRvF/kwxXrSm9rQ8UrTlyyOsfMiMzdoDpUuK/id2tyC4EWwIm+/CbkyXVgwdk2R1rKY9LOfCKS/iSj+2Wc5osDyA85qxY4lWWZMXlYarIpZQJ1LIGhYz4H/XH/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHSQAYMCrv5UCV5knami9wwVVRwMjhBTMPcMdlhAEq5i2rC+8KvwcIAjokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyivPvFHm9msvQrJURgKNO+4TkHZ7hGiLDNnr+NhM2pvDm6n85lBOtf2rmsl3HZ+TuOCXu1KdUlzFI86syL14DAbdfVTkQBuvYepnjTW5Ing27ZNdaujmE8lyZgTqkRGwLvkrkzINfvkq0/SkN6W5/RiSJw00xaEzAYicsrb8/v1TXj8uhnbttMrkgDO/3EBpmJ+I52+u3kOh17TDl/mvDrBV1/Sw/wYuve1rR3etR7Ep1U6N+5sUz+mB3XgZZNAPjTkGSJu/s69iGgXcP+zjV0ri6ANeDp84/Jw9YlomiUp8tRTqHjCyh8nMpfrDdyM6iSPOrMi9eAwG3X1U5EAbr2HqZ401uSJ4Nu2TXWro5hPJqmCwhxzfuO5JYomVfwQ4v3u+M/mYh2Qlhw4ye9aQIFWnFbCNmqEXLuLoA14Onzj/ib9EZFcK1pk3A2W623f1m7qCe6H9mcHnKq+3P0DMDjPeEwREjpXKcmv7G03ZpvcXsi8kDgweUqSOGVo5Wlik9tP0pDeluf0ao3pI+zy8s5bLRL1Fn6wTBwCgKozFLP5kzrrAH+4kYehAkUmrpBnV2wm2ChLjB6jSLhea0A4YkNRzWEKD2PpNXrh9/sx4J4ZekyA2VBukLUFfZITtU129QRXYk5FthMQU6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUckUCiasUyBH/WuBI0G9+rQ7yJShURQtb/ADKuVfSCivqH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LmmFES8+Cm8cGkhh4DauPmQGCFICShv5G1xg+mXKd5vkWAwRWLohduWwWyFLGq9l95dHXktQENbxD23+ziOLLX21Ukx/l+oXSo4f+2AKQ/RJI9cV2ZZxh2yxTliixcR7s6zi23tAF6jPKoosXlmGqZ9m0sv7LJtanH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LvOELWtFYaJAxkL91+oXh1AAHKLhj4L3RjWp4X/fEthWNsdqxvyc0pvvhO+I7b9wotfJjinfBJCFC6f59p0irJG04IHWlU/9ghV7vicnp53OJ3RH1LBpOW8EFAOSDxDes5D3OwqTwAiJ1dCgW/W9lYHnfaYqNGzwC5D3OwqTwAiJ1dCgW/W9lYAOWEQORr+Oi6pOtkR5QI7rnkyOhxNuHYlElQzqmYXRQIIlNnRYNwXE0Pn/VgPsBDy/3hOVKUaEJYvRgjO8tDxUiqunfEojG0IJ4GU2KWCH2YfwCuo8lD7HO1vv0WSUjnJcuiL3kkrXAed9pio0bPALkPc7CpPACIoG2zufW9P1rC3Nu2Rn+jNSwUBTkL2d8oqYKtC1om99OahAKxjmqWbfq1ME5GgnNCU/JXYZX9iYtT99kLM+MdWZoMcDzmvmwmQQBhARakHBawFgsHfuuaTCdtGpEtXPBKyDzcsAxjJBkAt8QCiIoXwK4I23rzbbn29A+NHFVdvIm9dx7IwdGZ61FLLB3V1f6P8BYLB37rmkwXCjyJM9eBPPUqcS18oLPlT5qAU4OLm+b6BBpsssZ2S2SA7eP8fIZ3WpRpCfou/ahopmc40BIXO3AWCwd+65pMEYNHhdfKXcBptzUYUBdAwCDEjmNBHtvdiAqB4HZKmo+tGH0s96rTnJ2bHqbKgtnFIU168w1ZvWJzBqYhmgMdqovAvSCfUBuyylT+edzSvSuYMdMGBOpcjMM9uQHNB2YXirPy6PIIrxXs/44G2kt1zGjDDW0uDLVV8OTG+IIjGLQmxGMR0e8xl/ItndgTluCaajekj7PLyzlcr/b80ORl+lGDR4XXyl3Aa/LIV9FZHR8gxI5jQR7b3bheYWBHXXXQQLpWSLblckQ+zOgBxJIwHmfA6YC6MYYuiJNiCdoRj2KnC2oQ8pwtKjBH6ab6nFM+gGrw5g00TiR0oMS3RldC8JptpjJITzLTqw9aDoVJ6fITuyUW/8exDhIsuUh2LMETKVUjlT2vocatP/8iyWTRROVd4cjsjZBWzV6nFpSrge4NvAKn429Mn4BYNAncoGkg5+gA4ucyggfPwGopGN5FQ4iX4kqsYiFwjAgLGi5HPbDIIvT+UNORMSVd4cjsjZBW0BSOp/xoUHFyVCHDB3/kewPsOQj7iMz8mvQikJWPE7CHYNbLmfROv/QGI+luyLZunJ8W3W2YQJWdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDSLLlIdizBExC2906JuabGs1F4WizKZmEYX0HiBSNyGLUjJvBEBrO80IUGh1sl2hPqpAPer6kaNEcRy4n5G9LBnPKxSUCjyIDjfuoxOiR3gsx3A7vFzCo2x9JJtB+BNBiKYpuXYGa4XRr0IpCVjxOwjbhfUs2/G3P1eHKnnBEGecZ/QxobMKWYN4hiMQSDHqks5Fu2nrxOvfEhgseMfYZ4x1ULW2AWLCOOWawsYKTQp1YggAh2zYxKrOm4GNjZXJtnhuXdOrQk/5ohxrB88qpuSlT+edzSvSuXW79BE0ttx5TNm7vlhR09bmYpk9pEF9gwuDhMsVKUw8D4M42fjKU8ZuPg6MlUyAVL/w0K43rQfgIPi1IK5tHqKw9aDoVJ6fITuyUW/8exDhxR2dWpC/g2OzYGEHdtxiF0GKme4j8TC7dPeo4uc8BXXFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/yWoe/lNCs/AydBnPve1Fd9/y1pHgzmXG6w9aDoVJ6fITuyUW/8exDh00pwpiy/KVzFtSD/oT5P8WeKdmTkEiU2cttEH0AG40+7lwxehGWA3KVP553NK9K6jwTGB+vCg0FKUnG7T12N5i0kWLnusckK6maR0RWksW21F32Il+s4UwU6UqoOkzCjib9EZFcK1plp8P/4AvFw6/ZQRZKzLOf9mAmFR3LKaecIKQH9xapKWm5wIy7VEbo3NIYTeR4v2Y2rmsl3HZ+TuIrFPH/HX6kGLfZg5JfrVqDGTzC+tFdi17GNtU97kTE2foAOLnMoIH+mg+n6Xvr+whByivyDfY+EqEHNKcJDhm8WJtc9KKXbvwR+mm+pxTPoBq8OYNNE4kcFOlKqDpMwo4m/RGRXCtaauhT3ZL8d6DhBcYyRrjy2PmLeeZbuMJ5EcRy4n5G9LBoVjoOoiKdVG7g5oq21K1RL55DKxfQFkEHsyA0WfWJdQnTLGBsENvg1Ldx1LyjwnRBYX66Kl11/P+eQysX0BZBB7MgNFn1iXUA2z5EyYI0PSkqxJ22ZY2LaioOnn/o5+eWz+KYrx7nU/MDvPQvnae4oCLmfIM/UTQI52DSEcWN0i+dEk1VgbrDmuVwjWsxhQeRxHLifkb0sGRVxgon0onxzHSRu3sbgOzSlT+edzSvSuE/FFlgC8lHyjNZdHv3VmL6w9aDoVJ6fId4AgF2l+b7HHSRu3sbgOzSlT+edzSvSuE/FFlgC8lHzsoHWYm7luenVgpvDe2lFKHEcuJ+RvSwaFVSD1FKcXtMdJG7exuA7NKVP553NK9K4T8UWWALyUfOwExx7u8RmsdWCm8N7aUUocRy4n5G9LBoVVIPUUpxe0x0kbt7G4Ds0pU/nnc0r0rr/K1Pyd0vS+D6f8dhzI3MUBYNAncoGkg5LFaicXcUrcWw046j9A4ZopU/nnc0r0ruzApkkoaMDp4cMmgMS30D0UiOnUM637J0kkFFBrL6/VzQS+GzP8/IY4w8xMhWprnhQshgLH884krD1oOhUnp8jqbdmcoQYqPJw6Y1Q2JCn54m/RGRXCtabgoEHWaoQv5OxjbVPe5ExNnGokgdKcFFOK3PbAXe25NBI26MsU3OoL50K2YSXp6+1d4o5hpphkjZ0aURK7nY7ejcwIAu0rX9LRoNlryl3GkKD6vHWL1wQ4MNJj97JMkrRUVhyWEPx3h0FugNZPx3Mj4m/RGRXCtabO+NPuy/V75v3+YEl8JkNJpWqh0Oh2IWXnSv/rNmDxCfnkMrF9AWQQLOMrJ8XLATF7roE+YpEbxdEMoXwrc0LWnRpRErudjt6NzAgC7Stf0tGg2WvKXcaQoPq8dYvXBDgw0mP3skyStFRWHJYQ/HeHQW6A1k/HcyPib9EZFcK1poZjdua1PKtMXIRzBshYOV4qCfVaE7GUfe9+J4k0co/Kcij4eRVyAumEHKK/IN9j4UHjZbYbHfxHwuDhMsVKUw/nSv/rNmDxCfnkMrF9AWQQLOMrJ8XLATGry/VQ3f7pbTWDp3sTkzViY6+9Vgqh0mtbDTjqP0DhmilT+edzSvSu7MCmSShowOnhwyaAxLfQPRSI6dQzrfsn1bOEkfe2txu2QIDgYQjo+IQcor8g32Php8rEBx2amh2vkRBUqqUmZ+xjbVPe5ExNnGokgdKcFFMOYYRW4Am7qjmXVBfK4hJZ4m/RGRXCtaZl+9ywoPPKHFTM/LO5RPzdCa1xN53e85ZtRd9iJfrOFNVVQjB0a0gQ/jJqw1iTxNXhYV8uIm1ggnarQEoD4YkIUzMxN3ZVssAr5MLZhS3k9vUPoFgvuk6oiM2xviRG/p7T3UDwJBQZLAFg0CdygaSDrHEBNYVWkOfwzVGbaYcUaW4zE280kuSmBDEKRORjQV0C1/glDwNc/q87vMSgEn5jhIyIakpn0vqnErAoUKDlkU2JVifYsCFFv1o92w6oXWnYjk+07m1SDj77vTzzbraP4m/RGRXCtabiN7L9OTBPDU3Ptiefzb1PmewN5sq8lH745izPgrZskPZBDo7ojZhfZ4itJqwS47yJWbp1N0EuirxRLu0XWMpKfUPEHPklzSj50STVWBusOUQbXBuFTLzoN4fexfEEdr8bqH3qqgQ2LVqzlgMXMBfClqKrgZ5J5W+j/1mV2MnOXRGMjse9BLD0xj2xuG2LhpbZskpmnJ1QIoMndA828MhL0aDZa8pdxpCg+rx1i9cEOCMkpe6qB+YHftEYEflCOY+WoquBnknlbx3x5pE/dG2tBZWaL8uN0xhPSLdtgZP+k/Cuqig44hMJoPq8dYvXBDg89r+1I0uw09hBgqonNW5qghX4L1x80hFyTS01Zgw1yc8vlkdfr92o8K6qKDjiEwmg+rx1i9cEONTEWtiGVkNRHEcuJ+RvSwaWOe4Bcfllvvx+I2ceTHUviGd8RVhhBBpWc2yTwbGGAuyq74nZmlH18mXlzgE5ISMIfqW0OanmjfUXWl3DoGvHnkwVsyySTqKIZ3xFWGEEGlZzbJPBsYYCnGokgdKcFFOUqPaLiv7Tb8UCSf/U9xrs5UHA9E/nuzM+UmFgsZzYyvjmLM+CtmyQ8nCmN7WTh3DijYfou0DdSrIsYSM3OD0sxQJJ/9T3Guy5+YnxQteqre4hj4WKLxruWIIAIds2MSpAvDiKK56g4vOqxRniGbE2AAM3ZH/iRBGAkpUjEUlv/7gzMGFy6BD4TkGSJu/s69jC4OEyxUpTD+dK/+s2YPEJZwI+BXKoCwDU5dGKHUkizHu13ZHOc98ksJ1MMFbREzxr0IpCVjxOwivkwtmFLeT2dWkHK0r7GzRixQY/UNc9Wzttpl4jd3JtbcuKYkbpcAjsY21T3uRMTZxqJIHSnBRTr6eZSHK2PKpTwocHwt0Z0YQJ++a4CdtoAvPpyRBLFg9YggAh2zYxKvJMoiRRwIwd5syRnZ8RWQNX6BfnfckxRyoJ9VoTsZR9VS5u/JGrKcQcRy4n5G9LBoVVIPUUpxe0pWGb78OwoqIcbjQx7Ks7jzWDp3sTkzVi97HLe2eeQZ84HXb23V+jBW1F32Il+s4U86rFGeIZsTYAAzdkf+JEEdASKNxWIRJorMa75Ri0Knjm1fRD6ARM91RWHJYQ/HeHQW6A1k/HcyMsn5O2x1G1nl2g4MYwsO3XQ6k9Q0JCWmP8BVvBnRzJscLg4TLFSlMP50r/6zZg8QlnAj4FcqgLAE5+xJfPT11PmFTPSoac78AcRy4n5G9LBoVVIPUUpxe0pWGb78OwoqLF2HimQUuPLGO6ppjjBwmOa29RXdEmURdr0IpCVjxOwqExlKxSUW3tOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2W3BEcGDMyMTUMVJnXwC3aim57Lg57LxYpdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxmk1WLWR4tywks6aP75sdn0d096ji5zwFdNoxbI4me9pimZFIuqsPI4YDrXOrkvJEoAM0VMcNdjM/m/fPgGiWhA7BvkETgs+XWGnkhHOWLndeYUieJ1YegZdiuoTHUj00cGur8EKoL6ULdPeo4uc8BXVJCJMj1/FLKu3BxnJnHGi23U4tcd5nCGARM5a3QoG6cknd7NQpRA29mzfnCvpTk9bhdDjKl/Ez7cEVQvmZs4ZhxCvea/bRFrFKtq1msf1HBZd/yTly2zIJx6rBvn1PN5i3UKe2EAR7G3T3qOLnPAV0/nmWvzkud8KKg6ef+jn55bP4pivHudT9aF8HuNOQTF6P1rg2RC9bp1UH3Z/V+LjCioOnn/o5+eRggGvnT1dc6ajkcM0HTJMWiAiNHs4agN4V/WU3qpuprXhkWLTJ2+6xmHE1i6sjYuXXT8LRrcCLGWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxmu+GOtlB7MKjR03DvDUKeAXT/O9OWBsaTrnL9KIepPJbrbSGOSTpH3cpqRuI3PA+1afhOdFPQTsdwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkxFfTelaJJvDKVP553NK9K5X9XD8eD9cip/ASs3EKJtG/FJxES+W2uwcNkxGAV97U6sYhKLmkabL/usVL9gJwybMlWFKUlVptlDV/FZgnWOBLbFjLM0L0FGvh48WgeAe+K0edPGUxp3R1D8XUnf5aNCo3pI+zy8s5SvlRtcdiFfmWIIAIds2MSqzpuBjY2VybSCi1UT/oEeQghJEJt9xAW1A49rWRcJDglDV/FZgnWOBLbFjLM0L0FGvh48WgeAe+K0edPGUxp3R1D8XUnf5aNCo3pI+zy8s5SvlRtcdiFfmWIIAIds2MSqzpuBjY2VybSCi1UT/oEeQIlepDIFg0pKIzbG+JEb+nouHgmKCBARSMDvPQvnae4oCLmfIM/UTQI52DSEcWN0i+dEk1VgbrDnbppuYYqr1RRxHLifkb0sG3HJKFUTLr7pkV2RKeFDdt3IStq4WjC5mT+QyoSnr4KnhhQd5G/Xq5OYiqiWWtCZq+eQysX0BZBAs4ysnxcsBMVFS9otoLAYqjpdVcb50H527cHGcmccaLbdTi1x3mcIYkNEPMoCb13r55DKxfQFkEGFgp7Y6JEPfKlZqAGRNlUZ6c9O0Bg63VviwHveeTMqmzQS+GzP8/Ib67pZhSX17SNzu3ZOWHk4ienPTtAYOt1b4sB73nkzKps0Evhsz/PyGRvgfyGsBOHg0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek59v5hMcRL/0UDj2tZFwkOCQkP1FgSCfe/2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTIQAniHUP618BLT4On/TbjigXcylQpMNl0vZwDlzKIgxJoEOBo+KxnyhByivyDfY+Gff6IxV3Ch90qqoZSserD0QIaAy+tSTHE37Nk97b+6rpR9IvpCAgNMWmgBv7vT+q0hVGVzBgcX5kydOY4cCap9NaQ+/yt3IYuAbAWZCTK1uA/XOJfyF1XDY3sCEo28Fct8J/VrU9hea2suxKHYfDbF4SSlnUTC2Qiwb5BE4LPl1j8BqKRjeRUOwxYPtu7JX5m/EUKWXiWm56g18ZZFxsrf00TkGxtLRi7oRaHkFnZ2UNHTcO8NQp4B/VTovGr0QLodpjwl5w1JKcCYA2LhiYf9AXuICwaRr40sdNfLhY75zro+eR8FJ+6DQuDohD/SGc44L8BEXYczgByea7edLQgPGGu+3/L5gB3eDp2hARUqOwfKI7NfIIfCTUzukOvUyXZAhoDL61JMcYZD0YxFx+drndNQ2VtlEPSzpuBjY2VybSgkp2OQPbYJKVP553NK9K4T8UWWALyUfAKOglD3i92FGsnjlPKS68UaIwUHZLJLX4uHgmKCBARSVHpQye/BwYSEHKK/IN9j4Z9/ojFXcKH3Y01o7JXoJ47eDCLqVi0uMxI26MsU3OoL50K2YSXp6+2P8JOOoHD8kpoEOBo+KxnyhByivyDfY+E/AaikY3kVDuUBJlfGrw1yTQ0Qz8SsAz5aaAG/u9P6rawdFhuzas+MB8ojs18gh8J54P6wCA7h4MxBPmd3IyJnUzZu75YUdPUhYsLPBXpdbBI26MsU3OoLGiMFB2SyS1+Lh4JiggQEUkBVDninNkj/2K6hMdSPTRzvQl6N7+AIWFpoAb+70/qt5H38VJ1uWmY1pD7/K3chi6g18ZZFxsrf1i5t3ireDk/AWCwd+65pMPiwHveeTMqm55w9mue2arfggR+hzBPyxC8HZEGoTxCDAEpUG6CU5b5rHszq1lh4ri9+I38gCk0sKVP553NK9K4T8UWWALyUfFG5mylj9mW/PwGopGN5FQ6fmmS/7b21AJoEOBo+KxnyhByivyDfY+E/AaikY3kVDklaAgaR8PUc0BiPpbsi2brIGhYz4H/XH0Te3KALTTmko42SHFIoxvsCCPIM8UbzZVheXH98JSKsJ3t9Rawit/k0MGESyPyxPMnCozbEA5VC3hPusilpRTvvT1jAzmCmG3RpJoOd+hYUUlljQ/M39j08tc3YQOrzznyA/Cw3lzwqPmHr4Xr1T07lvTUuxDoeVIj6CHAwAzlcSvXkPabCstYwY9lPn2PW+ChEWmK+out6IygrQlXVWifeDp2hARUqOwfKI7NfIIfCY01o7JXoJ47ib9EZFcK1pj3qSB/xtszijXexUUVT4fKXz5rmDyTTKOrUwTkaCc0JwiO2pvYsFV8ue7H9bpqx5szqgSIDgZBXVMz8s7lE/N1HNCb/bE0kL7c0KWFdl5zghAcs6LblPoHPLW92kYge6Llg5fuBTrJozLLyP+34SHDixNqL4K6K+81rIRWQdyFCBrunOcy3DdEYa77f8vmAHb23f9HiueSywFgsHfuuaTDN2Y5/xWj+4eulPEJ+kyZjKlZqAGRNlUZ6c9O0Bg63Vr2rBUoGQrMw43YVY774KSEQ9BMUbPYIW3cMKmb+s8su+LAe955MyqbNBL4bM/z8hvrulmFJfXtIZi0w1agfHwKPkgBJUwhBsj7bQ/5ABJDjnwDziWeYZMy+MQYhrirnU82rIsZ2j1EyrE7zYZJyS7nI6AyniWV02a7Qi0pdUr5P0dNw7w1CngGoNfGWRcbK35PiRyc+G/jB3T3qOLnPAV2Gha5pqfgj8OajaoonzT2+4SSlnUTC2QgvfiN/IApNLClT+edzSvSuv8rU/J3S9L7qhC1ytIRZtCVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3/iwHveeTMqmJd5QDLgzV7rpo0tqMGKr4Vd5WV8gU76CcPeNm59NMYEMK41UJTu/SvnkMrF9AWQQYWCntjokQ9/0vMmB34y6UFR6UMnvwcGEhByivyDfY+E/AaikY3kVDsMWD7buyV+ZvxFCll4lpueoNfGWRcbK3/iwHveeTMqmJd5QDLgzV7rpo0tqMGKr4ZDsBdiaM3mLEjboyxTc6gvGIKB8BZXcQZ4r/tYjUq1/qN6SPs8vLOUA3xzinps+BFiCACHbNjEqGStneg1J7JoSNujLFNzqC8YgoHwFldxBniv+1iNSrX+o3pI+zy8s5QBPucmAm2lOkNEPMoCb13phZozdt25vcB+pBQUd/IzhvoiGCRllu1SRftjjGWJHTSzO2ClnTF0RWmgBv7vT+q1NOMIRwaIAjk5RPjL/18fI8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWX3Vlu5j6fqPJ90+HsrJq8NEnaLgnzfE3FrnL9KIepPJY1OkWGc8TNyuiL0XHn2AGrnh05PBA/u5JpEbzArGXUPI+VNfkKUW5QOwhoVlMlYUGkNmRqWznUdbhic2k5kLJaAQxxMFtWwN3y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8f9tScKmf5jihyqqIMZwKRKjfX96yewauUWAEeYJanWVWw046j9A4ZopU/nnc0r0rmjtGGoGbXhVGrSgLn7jD9B9v5hMcRL/0XVOxSw+bqJR2SQjd+5XpjIUX0HwUOirfFpoAb+70/qtYIQmwql9MYncmeZty2DsZ0lu4sES4sFVGGu+3/L5gB2+l82Ja+sw7c+iNdzv2+sDdlJuDLhMxCAP6iquqF8CPT8ciI7ukbXTeHz/QmRw5TYYa77f8vmAHXRP+ExMXcQ/ZYUGnAY7VRG5X0wq7M2fG6g18ZZFxsrfGaF4BwRend3yvbc3fCjCTH5+suu9eKcHZZEDGKzNUgIYa77f8vmAHTUFTNzDDw80N1fFlTmBkmcnn/eRhT9SxTUFTNzDDw80N1fFlTmBkmczw6Pe4cRH+1JrntLiRahq0Kur71o/fuioNfGWRcbK32A8dKC/IiZKWqTz3+mLoAi/3bzWigGMNjveSImX13A0X+xkqAgzksGXIk1JlZdjcqlT71QxNftDlhjpoPRdHjMovJ2PA2gz5AL0kEjdIIoXqDXxlkXGyt8S1F+P0jKq1cMd2hdfixOdv2yzTKfz+4wSNujLFNzqC4+SAElTCEGydyY3poxtDYxi7mYxX0WepD8BqKRjeRUOQ6vtJYI0ZE755DKxfQFkECzjKyfFywExUVL2i2gsBipm/Ryw5q+bkL/dvNaKAYw2lXeHI7I2QVsQ0gqCcU6w2pTUiD3/70rdzQS+GzP8/IY+MX0v/+FrLag18ZZFxsrfEtRfj9IyqtWKC7l9yZOqSPnkMrF9AWQQLOMrJ8XLATGkmn8ia1Gt/Bhrvt/y+YAdSLLlIdizBExC2906JuabGs1F4WizKZmEwFgsHfuuaTD+J3a3ILgRbPmQvJ/Gtg5qGEH0Ukw8qFRA49rWRcJDgojEpQP5hfCVbb/ntHEx/iioNfGWRcbK39z0JJUew4U+X6maz8Mf8VyU1Ig9/+9K3c0Evhsz/PyGmQ6dLF8thXH9bDxuZ9h+2Kg18ZZFxsrf3PQklR7DhT66JCkbq6Njm5TUiD3/70rdzQS+GzP8/IaZDp0sXy2FceFY229t0wAcqDXxlkXGyt+80fPVDUTOTZSmz4/fohxpo4Z43lAweeNaaAG/u9P6rcakeqz9p8Db5gYYMSvBWb6EHKK/IN9j4TmXVBfK4hJZ7WC2R9AtZVoYa77f8vmAHXTSnCmLL8pXMW1IP+hPk/wG3SJPCawg3py20QfQAbjTvlkP4vG3jtSioOnn/o5+efQQ3bGrJfI2xNmtH0x0CeuuHu+KzBdRsZSytehtpQqkGGu+3/L5gB22PMS5HBgUOVpoAb+70/qtPBRehIFeP5Bsq+4FytlE1umg+n6Xvr+whByivyDfY+EyuJC6xJTy1YiT/fnSNp5fKqLBu3yOMdroi9Fx59gBq6ShZNjR8iw55sC5Eqj1cJ5jeLHAlxQcW80hhN5Hi/ZjauayXcdn5O5Zb/h0F1jGImgGynhwCG/d0372ExX2DzzNIYTeR4v2Y2rmsl3HZ+TuIrFPH/HX6kEIsJMAqh2q1ajekj7PLyzlIdWHn/tImo2tu7YHRjGV2cBYLB37rmkw7uXDF6EZYDcpU/nnc0r0rqPBMYH68KDQF0rQ9eQCMCW2PMS5HBgUOVpoAb+70/qtPBRehIFeP5Dy53saRsV9hRhrvt/y+YAdtjzEuRwYFDlaaAG/u9P6re2UrLQHGtliCLCTAKodqtWo3pI+zy8s5YpE722OMBL4f2KOYefqesb5O8c1/X7uIKFQLu0n4T7W4m/RGRXCtaZMdANqS7ySiPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln5Ojh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2Zdiv2/PARSMOjFi3elKSewCnxs3xDrAxMJSOY+FYv+NyeGBjZGr56nWRmgyOnuynTKvJ+ar2PdBgUQpVDhBElXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOys1ZhDP6lMJ8XdUn5A3p2tkCA4GEI6PiEHKK/IN9j4ceT9DJ48gRZ/FJxES+W2uwcNkxGAV97U6sYhKLmkabL/usVL9gJwya1VGZro4U2EfjmLM+CtmyQ8nCmN7WTh3B9FhpMRFotQjWUlYtzEPb4xQJJ/9T3GuxibOrlFWKCRhuYozLwMEAyqNXzXd6GrG1kuCAfLW8/UhDZzHb92co053Yfl0Bwi1KDqpuYQqeSUXCpaDK8/CB0TXJM6ss//ElQfJSpzdhoA2S4IB8tbz9SENnMdv3ZyjRHOVhkZTSo+toL6RuXGpJAbUXfYiX6zhQh7ZqYKCFRvdB7Nm3y+0xcOZdUF8riElnib9EZFcK1pmX73LCg88ocVMz8s7lE/N0JrXE3nd7zlm1F32Il+s4U0kfhGIVJ+sp4LB8SnYnkWJuhHwoq8y0TY59MtPd72sG5YOX7gU6yaPocAm/gB5F1oPq8dYvXBDgfO5O88P9+afaqByDZ6jU0w5PI0uBw12RAhoDL61JMceRAr9Y3JhT7GmM340wuvpEcntMtpfiKIltDQX4ZtjgNKUC9UwPEUwFaaAG/u9P6rbB71lKJpE7gQIaAy+tSTHE37Nk97b+6rvjkhFrTpNh599W9as+3kQgrS38jQRJ5Rh3YiDdIyMUtNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOUh8uL99ptz2T/vBO++dtBrWG/RF1RFWNZDpqtZrfo5tourMmZ+Ww9Je3XicDJZZfQ1pFmvl22ruVzBspFARCWZacAGSF9jAb2K6hMdSPTRztJ1HzQxcqySjQuTfvCGgs+tPbMB1+uxzGEhMtEeNCkTpHZex+pcjKVNHUjdCULt68LoCjszcV0TNLGvQY48Ou9o1CgVlT1Yt8gPwsN5c8KtAN033DIpkTNtL5kgYrcA1E8BIVMYCVsfoMNWA7OOFaYc9V/ti4K/jFAkn/1Pca7M9eRGH9JQIcat0yLaDXGVElX26L3zEeg4h4BdF8CI0lZL+814w1rJaskPxLL+8gfZ7e8AKsiYpZBExjoZrrAHE4URe+RmtTaeJv0RkVwrWmNtKYg6sxuYOUTihxtJuHuJGMZSUNb0n0ck3AdF3nbDFqYiJJoX74IfKcrn+p14eKnrgr/BC+fs59x0PG2ahCSsBYLB37rmkwNZz0yFbviGag+rx1i9cEOKvHRLLjwvH15krfjBhZlP+7cHGcmccaLbdTi1x3mcIYkNEPMoCb13qdF1VrLELAopaiq4GeSeVvo/9ZldjJzl027GxhwPSxHExILR/FcFeqWmgBv7vT+q3GpHqs/afA22AxCKm4g/0KkNEPMoCb13pYa18FP5By6aFOWhvQIMdbYc9V/ti4K/jFAkn/1Pca7OVBwPRP57szGsnjlPKS68VkuCAfLW8/UhDZzHb92co00OmLBnNSH0gVi5VOCjCxWHCpaDK8/CB0TXJM6ss//EmyIDqErtreOlAPHiuHcPVLtwlgYrweSq9E8BIVMYCVsRyYmvUe+fd246ktm+MiKXYLfxkNwHUMMkbEgTYkUrdlmewN5sq8lH745izPgrZskPJwpje1k4dwcZinTM8Sur24S5g4i6k1Lxhrvt/y+YAd6SQqlZ/JIaqb6ghZnPxkKxfKw4ezGVzRGXYtUHZTjauoNfGWRcbK30TimM6oX3TUiGd8RVhhBBpWc2yTwbGGAuVyYA4EPBH7H4df574TJBtGKrnC3xFW8MUCSf/U9xrs5UHA9E/nuzMNVvWYccNDUaexfRDVq1G/UBp2wuvWpinAWCwd+65pMMBYLB37rmkwwFgsHfuuaTDAWCwd+65pMMBYLB37rmkwROKYzqhfdNSIZ3xFWGEEGlZzbJPBsYYC5XJgDgQ8EfvCoi58W3k997jsCuE8sbFl7Gfhw9lEZpuWIfqIs0eBJ6g18ZZFxsrf8xB7sp62pU2Q0Q8ygJvXes5NFSdNE6Z/jjLY3TEgHJGg8qFx7Ja/oBIvzOToHmTOlqKrgZ5J5W+j/1mV2MnOXWi9zQOX4tiG8K6qKDjiEwmg+rx1i9cEODz2v7UjS7DT2EGCqic1bmpr0IpCVjxOwuPlFyDCCNCFG1o37w1NpGBjEInwZUrqv7jc9VUHC9J3u4DzqoPiSyqVR5tB0yz9EcLNjnDogolaWrOWAxcwF8IpBW9ja8TZKKD6vHWL1wQ466l6hW7w/uhkuCAfLW8/UhDZzHb92co0uoHAqDJ8P1uThs5VrqkgMrIsYSM3OD0sK0t/I0ESeUYXXYD60WhEt9l9mvxruCGXqDXxlkXGyt+yLGEjNzg9LCtLfyNBEnlGHdiIN0jIxS1J425X6IfQozmXVBfK4hJZ4m/RGRXCtabZry6oinSCWZ8A84lnmGTM/vkPv/j5JwkMTZLQ9KzysMI7BDzRop/hzEE+Z3cjImfkLJZTSD5dJ2iHGsHzyqm5KVP553NK9K6flnPNJGYGKQzCwsjkVgCQqN6SPs8vLOVqf8YwCKLlL7lg5fuBTrJo4nDV/XrVdcc5l1QXyuISWeJv0RkVwrWmOPSbREx505hK4mvv3bsTwrZAgOBhCOj4hByivyDfY+H2j8PLQ1ycrmo5HDNB0yTFkNEPMoCb13rKVsPgxIwZHRlIdIFPDLEZWF5cf3wlIqxAdXnF4vjGJ+BdNO9ICE4+78gdgX4Vse5yjK7bCojOzxE7nNp8sszc5iKqJZa0JmpSHy4v32m3PZP+8E77520GtYb9EXVEVY0Gu6c5zLcN0ZflSbQ/7r+gNv1C5IcM116oNfGWRcbK31e6vxd6pfubDE2S0PSs8rBdzNiK5tOvPILQ04Y/0qyIniiGxY+UbgiiNsT6HltXTfZpsnAOPbse2Y8Wvq1zX4Ectas+oPi1vMq6NwyUzhs7EITvjH0B+aBdvRQ8e32aQhYQj1oUlAuZeCwfEp2J5FglqHv5TQrPwMnQZz73tRXfWQ8wxwY07XtXmAeYqCVGIMBYLB37rmkwEMkGQcEF6B0pBW9ja8TZKKD6vHWL1wQ49qoHINnqNTQT1zWClEYtH4XLjiOTjsUyqmsDxRVIPaKbj4OjJVMgFS/8NCuN60H4rn5Bj1eqyVZ6c9O0Bg63Vmo5HDNB0yTFBEzlrdCgbpw2/ULkhwzXXn36paaXJ0Fmq7BLCzMzdrmfF3VJ+QN6drZAgOBhCOj4hByivyDfY+HEkHluyjAW/fL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4Ull/LbH3nTSWXO1VYueuMIv1lt9pH2UAMIof7YWL0Jm4gU1dpumijwrqooOOITCajekj7PLyzlC1AURgVlqV20K7dSLPo5jykFb2NrxNkooPq8dYvXBDjOHsCLHOM4tffVvWrPt5EIK0t/I0ESeUYd2Ig3SMjFLdQVSQhFDqgEKUC9UwPEUwFaaAG/u9P6rfd9ZMWWJaTvP0fx17GOb03lOa7q651sZQ3iJkx7P6IXxFgICoR2R1vlOa7q651sZbHeljEya47LMj1EomkBOXDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8SuBpslhHO/IAe3n5GVz+k8CcNDsxKchWETwEhUxgJWxiMSa8TaHjr/8Mp19nPPxvkqc9BrDxsBIaa55jybRIvPprHEWwLJVJqsMWM4iqNh8OiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHKdbLFa/i38RW923dpWjeNa5oyoIXeJbFuwNu9pJr5KepciTUmVl2NyDcWDzbxYwjogotVE/6BHkK4Jk1m5wAEi/RR3NYigAxwNZJfX4cOWpG2iGP2HJykBWIIAIds2MSqzpuBjY2VybSCi1UT/oEeQrgmTWbnAASJCQ/UWBIJ97w1kl9fhw5akbaIY/YcnKQFYggAh2zYxKgo8IZFs7BM+DQUFJSyD4MVNhDOo5YPnV/ML3EO/WvzNjhwIGUocy7GoNfGWRcbK3yyfk7bHUbWe/XMQlPCamgy7cHGcmccaLau89FjbHlF3E9c1gpRGLR+OL9z0IaBXzLNEZ2s85WcBOWzy0Nx5asG+c8SO015jYlEJZt5I6hoNu3BxnJnHGi23U4tcd5nCGLOm4GNjZXJtOuIYo/f2D8D0x/AFB8GuKzSc3R/HQ5ndOSHV1ZqHYJlRCWbeSOoaDbQLbwE2vp5pEelJFGUuidkAAzdkf+JEEUC2V7cGw93mJV9ui98xHoOIeAXRfAiNJWS/vNeMNayWrJD8Sy/vIH1hzmCobOs//F06Zj0VaX9G8erlt9uTitJs/P9zr8kn/SVfbovfMR6DCZrVxtmjyhmQ0Q8ygJvXemcCPgVyqAsAtUopYyW03RY0OvP90zT1HixfGI9/oyonbPz/c6/JJ/0zJ/bYDVRTMKnDRjqcd8g4lB46/ONT5Pup8akuHxFzA0CGgMvrUkxx5ECv1jcmFPsaYzfjTC6+kejS7z5XwI5G8FPB8WT8BcdxGNS3NEnkZfaqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+qDXxlkXGyt8sn5O2x1G1nqnxqS4fEXMDQIaAy+tSTHE37Nk97b+6rhHpSRRlLonZAAM3ZH/iRBG+c8SO015jYlEJZt5I6hoN5iRnMMMFpPtmPJKZ4to+ygwdk2R1rKY9X85afUIPTVlRCWbeSOoaDeYkZzDDBaT7ZjySmeLaPsoMHZNkdaymPb5zxI7TXmNiUQlm3kjqGg3mJGcwwwWk+/cYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaKLw7qSoagOKtSPxfNwhGtQN6HOf6eUJHOuuIdRQ6Vdr/ermcXqbL2CubR49MEXXgzoxYt3pSkns+eQysX0BZBAxxwgOBF9AQUr15D2mwrLWLJ+TtsdRtZ68197s23yhybtwcZyZxxotq7z0WNseUXcT1zWClEYtH44v3PQhoFfMUAbSjVcAROkaTiTc6HMjoIrMhDJ8h7hkJV9ui98xHoOIeAXRfAiNJWS/vNeMNayWrJD8Sy/vIH0GY0NzhgYSbFnX8J/7J+1OtNo6E8jNFVL50STVWBusOdumm5hiqvVFHEcuJ+RvSwaqYHsggBJYRylT+edzSvSuqORYhzctgv6LAPxMv4f68ZDRDzKAm9d6rgmTWbnAASJCQ/UWBIJ975w2v10+o7b1WmgBv7vT+q0SwdBnDRh8I4IV+C9cfNIRExmDq+mjjShA49rWRcJDgonGPW0VL9kXY1/Vvk9ipkSoNfGWRcbK31smN4Cmq5n888vf6HForg7Hb7/tgU5nI0WAEeYJanWVkmqvYw2pqFkYa77f8vmAHWcCPgVyqAsAIXUEftJzC69y+5nx1JzUfOQLa7W/39OS/RR3NYigAxx4mg03TqOyIGoW0hepgRpQjT7YRXs13sfKXoCJJkzFhD9Loy1Fye11MosEwBjbwnKzRGdrPOVnATls8tDceWrBoxbIYYYZI5dPCt6o+mKBDxpOJNzocyOgJ49htbU7sqhdCK6l1VZK0fIfFKmnxE42Wdfwn/sn7U4anoR4ukg4akpRE9bVBTiel+VJtD/uv6CWIfqIs0eBJ6g18ZZFxsrfWyY3gKarmfwvbzyP4J4wwMdvv+2BTmcjRYAR5glqdZXa8c+urmLThMBYLB37rmkwLJ+TtsdRtZ4YLWCdPoMjEax3W73WWWwNLJ+TtsdRtZ50xHBCMc9xpqN00gN/fwqKvM0y+qTZnmY5bPLQ3HlqwQKEatuyvBzgFKbZMim8lWrAWCwd+65pMCyfk7bHUbWedsWyTYA6Fn2sd1u91llsDSyfk7bHUbWeSRvvAIaurpqjdNIDf38KirzNMvqk2Z5mOWzy0Nx5asE/E47R+9NyiRSm2TIpvJVqgypL2PvmW8Fx9OgdnkHJZ58A84lnmGTMRQJdpHPz088WhIKst6Ucs+kkKpWfySGq1U7FWimi4hrgvCfaSCNbt5G7d8H0C1ozAAM3ZH/iRBHH63RapyqEfFJN4YGgcwFhAAM3ZH/iRBE9KRPnA/eNbXWKGz+IMlYeuGK2oLWF5eUzz8ckyViae4hlyCo6vB2MI/GItrN3/2GRu3fB9AtaMwADN2R/4kQR91Xu478vyb9STeGBoHMBYQADN2R/4kQRhr5P+o7uo2R1ihs/iDJWHrhitqC1heXlU8KHB8LdGdEjQEe3g79GrSPxiLazd/9hAEpUG6CU5b4S7mzIwwp3t0Te3KALTTmk6bd6C8lsyVGoNfGWRcbK35cRiFXk5lH5SRcwuxVrjWUDDmo0qbnltqnDRjqcd8g4lB46/ONT5PuYcy1ZK3Lw3y2DKeo4lUXhHG40MeyrO4+UdWnKTbNzRSrjAtGKgOknwwRHov9SjG1KyAq4xL1ZkYnWoxG+KHzW5DB/53FFOOupw0Y6nHfIOJQeOvzjU+T7clgztW/oj4ctgynqOJVF4RxuNDHsqzuPuQQjd77NM5wq4wLRioDpJ8MER6L/UoxtpR7P75WRAiiJ1qMRvih81uQwf+dxRTjrvasFSgZCszCikJkdr3478ZGMZSUNb0n0EhdVi+uglwQR6UkUZS6J2QADN2R/4kQRKJ260MqesqOfmrunKoCvE7X0tdsL0YqR5ShB7+sCnNK8zTL6pNmeZjSYw9OBUUsbI6m2Cz5AsZ+zpuBjY2VybTriGKP39g/Al5GKzXDYP+G8zTL6pNmeZjSYw9OBUUsbKspCdHVX+9VqFtIXqYEaUCyfk7bHUbWepzh5T7FbTPKg0kTih4RM6J8A84lnmGTMLOsY+8PgSBkx6+h860tqEzQ5gleVGHfehbTaIcVNlmQJxq30VWVdbtz0JJUew4U+F5TvcqXOBv0S5s2AtQKcMYC/TgNN6yBU2ORIAnEKnqtQDRJ+hzGH7YTMyZvURocbZjySmeLaPsoMHZNkdaymPV7YQver1v2FAwl+HhDg0Wgsn5O2x1G1ns0kS0LQjlWTQtcDhLsU+Gj/NwFwC9cbSGo5HDNB0yTFogIjR7OGoDeFf1lN6qbqazkVHpC/m8bxHUv3Ydkkxqby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+RlB3leja3rfS3cdS8o8J0QJKWePQB2wkLSCXgofxdjQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Ltx5v2R/2i7QW6cR3ugt84yOSikUR84Jm6vt7lh6NPTEyIl9tcDvIrKwQFMBrptmFt2FocRTvBr2+YkbIMZ8A+du/y3mwoDlqvnujeI7UaGwAyrlX0gor6g1ND+mU4+mNmtmwwjkh/Y9RlZG9GFHxP4sGwRjmsKH3H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LE6S3a9z1k0WeUUQ57P2dZ/D0yVYSr1ZqQun+fadIqySUzsVX+qjJ2VWvn3zt+a+vNGzsQ7/B5p9Qw2GSyqIWv4kAEDsXn9JOtWHT9AV0+9AxkL91+oXh1Fsnph1GMPMA55MjocTbh2KxrN3wl7KRmuqTrZEeUCO655MjocTbh2Llj6Q9piTVVjNvcaGxFOTatfJjinfBJCHC/Akftdwe1xaMwmyDRPwoI2z39yYmxkvSgIrk3Duj8dZJwV5YQzzoz+C1ZKBRVxZ532mKjRs8AuQ9zsKk8AIidXQoFv1vZWBTV1Ow46mucuqTrZEeUCO655MjocTbh2Jg/CBO8Fj5vgm5qCV94BibIqrp3xKIxtCCeBlNilgh9mH8ArqPJQ+xztb79FklI5yiNFH2NtD6fq56w8vceuNoiaE4iAwtsipB6pIgDSrKgNJCZTW10xy+0kpBS5r4LY4+/8gGLek9mqHD/F1KTXj6wFgsHfuuaTAM9uQHNB2YXirPy6PIIrxXlLgB9YwaOIMXjIUSRp5iLFeQAiCPHqhvdE/4TExdxD8SZIflFwKTGFwNT4Su+gmAeIEWMn685D7yw56ELXbOTEbZ8+ehSgh6+tPbMB1+uxykab8tyNYGPy43GWN7xBKzbRVR2f+S08jvLBREZBsyKSznCTT1KMwTyb6gok+TsLX6/g+/xi8vHplDjbyGAKq+rdL18Y53nrBLdx1LyjwnRDHHCCEMf6C8CHiFB3ZQysfoi9Fx59gBq54dOTwQP7uSFdF9sNL77K4g83LAMYyQZCNbCVwY4RKuGACxZueQsta8iFN/SvSSe8TMVETQRPgsk9zh58NNPNRyKPh5FXIC6YQcor8g32PhILyEafY/TT+z8BLoTp1oq8m+oKJPk7C1Sw7CfIe0Fl3609swHX67HKB+4jtXrPJVhvy908q9WblUKWfrZ1reWCalmxDBvT6ycV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/m6EfCirzLRNmAmFR3LKaecIKQH9xapKWakY/FF8AzWg8tc3YQOrzzlzGchwav//MwV5kUMSlBLg/AaikY3kVDupsnDhTV7KDMCAsaLkc9sMgi9P5Q05ExJV3hyOyNkFbQFI6n/GhQcXJUIcMHf+R7A+w5CPuIzPya9CKQlY8TsIdg1suZ9E6/9AYj6W7Itm6cnxbdbZhAlZ1YKbw3tpRShxHLifkb0sGc8rFJQKPIgNIsuUh2LMETELb3Tom5psazUXhaLMpmYRhfQeIFI3IYjxStOXLI6x8jdJIW7Xv4pYl6D6ITEIyuQGrw5g00TiR3PQklR7DhT71sjhE51GMawcIiTMCV9H8MZPML60V2LXsY21T3uRMTUdn1ZhMqr1TtlnOaLA8gPP3IEJC81H1gTGFM4H4efwuTkGSJu/s69jC4OEyxUpTD4LF9nAZbW1Ml6r3CSjbOX5Z5YAumi6YjO6gnuh/ZnB5QhQaHWyXaE8BYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h1nlgC6aLpiMcij4eRVyAumEHKK/IN9j4eJY8MeStEN8nrgr/BC+fs6ia3IMTTWunlRWHJYQ/HeHWeWALpoumIyGL9tNOi/9KGehIcSq8HwlG+n1s+QzRGCeuCv8EL5+zk5Bkibv7OvYwuDhMsVKUw8Vw4+YPdbWBvCuqig44hMJqN6SPs8vLOXFqyrM77/6z7Hlx5s8YLHMr5EQVKqlJmfsY21T3uRMTUdn1ZhMqr1T85aPd7bXLue2QIDgYQjo+IQcor8g32Ph4ljwx5K0Q3yeuCv8EL5+zqJrcgxNNa6eVFYclhD8d4e7y7P5cV3Ptj3bNc5h58Js4sTai+Cuivsb6fWz5DNEYJTOxVf6qMnZwWFEse2vnPagOdmIOZ5ujGV+ciC9trJa8/TVDKwR8YQk4Feq0u3fy2YCYVHcspp5wgpAf3FqkpYfhcE4/+Cy30JedmLj8OTYD3EWbs3/qzbxdN+hDEejVpTOxVf6qMnZwWFEse2vnPZ+b81YoZuWE08MDQF/7jEYsHhv35Z6JybnS3neikNixGfnQvQKDKkh+JjqRdkszjkQXGMka48tj4tJFi57rHJCupmkdEVpLFttRd9iJfrOFMFOlKqDpMwoCmSzK+vxonKKso8+c3aOkCspC8S1AlPqD7DkI+4jM/Jr0IpCVjxOwh2DWy5n0Tr/8DR9AAKR4cASNujLFNzqC5YlHfB/zqZz/zdjE2h1RvcRaygtE5naOViCACHbNjEqs6bgY2Nlcm3u5cMXoRlgNylT+edzSvSuo8ExgfrwoNAwol3FYOBavzAgLGi5HPbDIIvT+UNORMTmoETK2hidRqjekj7PLyzlIdWHn/tImo2pFRTU3iAjTh3bcYOqDhgjKJnyGPmNyWbhwyaAxLfQPZucCMu1RG6NzSGE3keL9mNq5rJdx2fk7vo3Ivj0zua65Ld3OxyR92yUzsVX+qjJ2cFhRLHtr5z27uXDF6EZYDcpU/nnc0r0rsev3EEsczW5BggfoHS0qym3N2ItPs9tfuxjbVPe5ExN4UHRF2FP0mzG7Ce+W2HfcWXMSV2r0LxpkTk+9SxN4FUNfP/1CBud8VW7inPYRzEOc1E1Q2lqdtHRMgNHSLmAHm3gjXOEok0SFaxWXSQHf9Gev1XJ64vHB4bvWnk0VbzsrHEBNYVWkOfyB7SGLKppNxF/mjKMTrUtO8RlGCmkrig6D3w6o/XX1/J6/nou/PGxwwLI6PaEiG1VIEMkaX/hZYlZunU3QS6K61O2EiKeVXXnSv/rNmDxCdt8viD2Pcbo46FnwlZdCSjUrYBXlMQtxGvQikJWPE7CK+TC2YUt5PaW6tXGgD6qoibEf4pPKYQ6fobjCkrKLXpYggAh2zYxKvJMoiRRwIwd3YblGLjJTNr+auMVYDwYlNEMoXwrc0LWwgpAf3FqkpYUiOnUM637J/c3V6cwb0nT6Jzm+JTZIoGeuCv8EL5+zk5Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCfrQWiUhv22gv+7HiQZWY1Q1Zicz6VVMhCi+G04JfRlAVFYclhD8d4dBboDWT8dzI94u8CKO4j3DkdJtHh2KlbySh6M44dDkoyiZ8hj5jclm4cMmgMS30D35mIpPSMlFC8nghxtgSf/dGKbyRacrtkKidpiAqLWn+YtJFi57rHJCupmkdEVpLFttRd9iJfrOFKcnp15/O3TdQ48Klkl6qB9bBxKCjXZ6EEHI9aDL4/wTD7DkI+4jM/Jr0IpCVjxOwivkwtmFLeT2pxCxH/LdU6O9Oa2fH/gDQSzsCQRQzh7UEWsoLROZ2jlYggAh2zYxKvJMoiRRwIwdAn9N8Zep1WVNUDUdFl7g5564K/wQvn7OTkGSJu/s69jC4OEyxUpTD+dK/+s2YPEJESTztMuEgrtp0Bwxp8a5ixFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHQJ/TfGXqdVlZSaWnvZe2NwwO89C+dp7iiCL0/lDTkTEQW6A1k/HcyPheHRWukdGMtEMoXwrc0LWwgpAf3FqkpYUiOnUM637J9dl0GZ/leaoCn3e4CrK/cxByPWgy+P8Ew+w5CPuIzPya9CKQlY8TsIr5MLZhS3k9rjT6VyuHQayOfQe2WVEi0i+ZoMV+OHM4TGTzC+tFdi17GNtU97kTE2caiSB0pwUU0SII6Iyryq1SsGn4U4m6JCUzsVX+qjJ2ToUI3EUh97186rFGeIZsTb7uc8DbJ8+8AbPrROeGUVt/f5gSXwmQ0mlaqHQ6HYhZedK/+s2YPEJPmAsMHb7AOrheHRWukdGMtEMoXwrc0LWwgpAf3FqkpYUiOnUM637J0eCyXGTMbc/vTmtnx/4A0Es7AkEUM4e1BFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHTj/fUMiCbFK3skA2C1ljiO1BRYdoPVBonVgpvDe2lFKHEcuJ+RvSwaFVSD1FKcXtFFv6Bi0afoq6mjAnMsfNv+/psQaoFtOIAXI4jeSkqH8KuRaK+ZZ/5nhwyaAxLfQPRSI6dQzrfsn6wgfmtTePWsuIzQREW/iCLyshTI4z82i8hSSR3ajaK0cRy4n5G9LBoVVIPUUpxe0UW/oGLRp+irqaMCcyx82/4JdLh0g0PtQ1ociu3VKxwXObbBmchPkx+HDJoDEt9A9FIjp1DOt+ydxZFYEK2F249NWS4XzWpI5+QTvuMLqRE6dGlESu52O3gGTsNaRYYomHEcuJ+RvSwZFXGCifSifHBJrJJfgyQ/1nYrBGuqPwNaym6TZ+4ZAL5TOxVf6qMnZI4vTKyHBGc8YlCRV3OBRxIJ4fh36Dqz5QW6A1k/HcyM59B7ZZUSLSJPxWtMzAgGoSX1eYZ5oBk2JbNXR2Y2XTvEae5HQ/VvXXiu5UQV8FEPl2OZPzP4kvv5q4xVgPBiU0QyhfCtzQtbCCkB/cWqSlhSI6dQzrfsndasJ1vGB6X4NzJ6Ef67+O6+HjxaB4B74AavDmDTROJGnJ6defzt03V1RJNlAAqHwMJp9vrRWXeMxk8wvrRXYtexjbVPe5ExNnGokgdKcFFOUBi/Cc2FCyhknl1KpJK/kwgg/EGv40FBOQZIm7+zr2MLg4TLFSlMP50r/6zZg8QlDbzX4/bSz1O5mtt+2oBA9i0kWLnusckIJrXE3nd7zlm1F32Il+s4UDVFdmoI6PBjVpEbPMriWNT0toaJ1zhYvFLE6gy+KXP1YggAh2zYxKvJMoiRRwIwdOP99QyIJsUp8uP8B73xPpMIIPxBr+NBQ/JM0QwbobnXC4OEyxUpTD+dK/+s2YPEJSj3qncdyBmFVPWW+qKhb7InQe5Uf6V63WIIAIds2MSryTKIkUcCMHTj/fUMiCbFKejrVpkRaG8nCCD8Qa/jQUPyTNEMG6G51wuDhMsVKUw/nSv/rNmDxCcCUIkFv5qe3q0oMMMiW2kn5BO+4wupETp0aURK7nY7e4lliQR6AqWLDAsjo9oSIbWivf22M5pDn8Rp7kdD9W9cr5MLZhS3k9hm7SZ7t+P9vEOWA9WExwic1epxaUq4HuJtc8GpGHxkVpWqh0Oh2IWXnSv/rNmDxCVD692bx4iGyaTX623ZVV89mQxzABC1dbXVgpvDe2lFKHEcuJ+RvSwaFVSD1FKcXtJ165aKmwYoweddT3rsrfc7QGI+luyLZumO6ppjjBwmOD7DkI+4jM/Jr0IpCVjxOwivkwtmFLeT24x8dtCp3i6cD7xDjEan8Ur0/byzNr6MKMDvPQvnae4oCLmfIM/UTQI52DSEcWN0iKVP553NK9K5gx0wYE6lyMyX4TG+j1VUfgnh+HfoOrPlBboDWT8dzIxM3e7aqgMa4z8pNw5JTrIWym6TZ+4ZAL5TOxVf6qMnZI4vTKyHBGc9V+uoLYyB2AP1buDDf9fDntwa1lNNbSWacaiSB0pwUU6UlehN3zjnisU0/oJHfp/qM2tL6TG3QtAFg0CdygaSDnGokgdKcFFOVPC/DhPfjabZZzmiwPIDzozWXR791Zi+sPWg6FSenyHeAIBdpfm+xaCVUTx0Ldul3yGQ3+1v8dTQ7e1k80Qpni0kWLnusckKBxl0y+KwUu21F32Il+s4UyNuIjjJNURjVpEbPMriWNYB2QMhvPCeJNWYnM+lVTITu+49+N5j8NVRWHJYQ/HeHQW6A1k/HcyMMHZNkdaymPepsnDhTV7KDlM7FV/qoydmdE8lMvwJei2lAqlLKErBpxtd7T1IVlmTCCD8Qa/jQUE5Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCS7E9Q3b7xJCPS2honXOFi8RaygtE5naOViCACHbNjEqQLw4iiueoOJe/3IFH7+KMBJXgTipY6mor4ePFoHgHvitHnTxlMad0alyDWxEiU8Ja9CKQlY8TsIr5MLZhS3k9sav0b7CzNyrB+CZbzfAuFIBYNAncoGkg5LFaicXcUrcKL4bTgl9GUArBOhIF3Yy4kW3/xjgeN4byJMDPf58wFvfcf1Mf9P6Y52ZIevvosDuafAXapYNs5udCClQjtkLmsZEXwGx4BMOLuUM26rs8NvTVkuF81qSOdBGcNUDt/muS1VycFim3gqgczzEVznGKWXbI1w74mecNIPm9GswZnPhmswq3yY3WPgDySmSIpuEspuk2fuGQC9bGWYXNRwVq0stOds0J+YKRbf/GOB43hvIkwM9/nzAWw7hziso5mEtwJQiQW/mp7erSgwwyJbaSdBGcNUDt/muS1VycFim3gprfNWVWWYHSwEuZ0tVGH/EW9UgCDHWybhoNxvyQ8QW1lMD6O1jZsT2beCNc4SiTRK2Vj2rFF1UatEpX0cGoCbUtJHeYJF3ambng0BEe+B2qsLkHuGMG8HWB6zWvc54nLnHuhOXTeaFEQQTKhkCMCgM0RRoVXO6yLIKDTzY6X5jNHgu5ycM1HwOn+mkvPPHNolRCWbeSOoaDeYkZzDDBaT7d7n4+DSADDqur7lLJxgHGECGgMvrUkxxXLnjWymgEA46OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZH4k6FkaOzap8HO34+GtPOSAXGxzsd1P18v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTrFqZvIrlnE0JDduZ1NMfBJT1dzNIy08oHb9NaCTHvtVf96I/NeAv+XjSXWVvU5e0SKwVTJiCn7hBkx4VDCBbkp64K/wQvn7OdyRahjnpyC9f9W5MXt61N41gaYmce4gS7qCe6H9mcHmrRIuP3VR7r9WZoiiFN4qHOH0DzTrgtIp7VNiIJufxuJTOxVf6qMnZI4vTKyHBGc9CeMf2ZD1BIa4ff7MeCeGX8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCThSWX8tsfedNxKePCQssKMQR+XeTW+bH5HdiIN0jIxS0aPgrfiNL0tQj8I4DemQQwcij4eRVyAumEHKK/IN9j4bGc+sKfn6v3cPcMxRz91r92OEtofaIWDtvOLjyFka1VLE2o2qgPPbdUzPyzuUT83eiL0XHn2AGrnh05PBA/u5LjLG13HMSmXEC8OIornqDi8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEcTcvWuScXwr5PNZHjv92QfOnQHfseN1W1qiB6FwN50jc4x0IDx4VGcW5cYTe7mmfzTEd3DDWG8PqVUjlT2vocabNpSdunsHtby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOys1ZhDP6lMAUhrQL6c92nD79vTvHnOBKhYWAR161KjWdq6q+4iv7MalCoso7qGU4npv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWsElqjsKdbEtk6dAd+x43VbYjgSlc8ZhlVJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfIWmLqwovHZNc6J/fnZFbjvaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMvcaLydpsQM0S7519g7oX491FiiUOkfRs6a35DOqZ0CrvxFCll4lpueoNfGWRcbK3875+cDYpCPB5Gom/sLQz7BxQ5vTCrbMcTp0B37HjdVt3bOolX2jUIkSWqOwp1sS2S8jKhI7hEwpBq1t35MuvqXYmsSLNW+dTZ7+ehYbqhzmCjS7FrK8+zNqORwzQdMkxaICI0ezhqA3hX9ZTeqm6mtu5GsWQ+CTZqHhk7xaWUw1OiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHIyPUSiaQE5cPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxbTEslmXbaye3Sy3SdjZglTPCqYb32VRZKLRL53Na22IUyEIXbwbQeyx9dqYb1Nuq+SxVxujKQl1b/9Rz8nqbgyjsXgfB9luyZjUCWr/7OvcO9fka5oBwypdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmxtE/f/rL1MJjjt+45IBYuc0c4NDhG9giCyJ7naQr5WKsJZRsOPth+6bOTF1KWT1qhSYDdhWR8SaeExe6S/Vo23f+zZLf8Byc20UfxrAW9Z5oMcDzmvmwmRop3chTVXMBy1CEuOjaPZswlJ/5IYLwyXCv1OkUuFpEDqFeXIjVfUOP4r3tD8ykX0WyOTE2UwNchBdE73GNEXhycn0fczLPWCqiwbt8jjHafiqJ59OKOgAfILcYi00x4gezedDC0hirpdntYsoL4Pt+jzavHUBG/+eguvYqw5bJvsAljwu8TvWfAPOJZ5hkzCCDlfeLskX4x86/zhbm2TJoLj9s86Pjly+595hQ5cfij5IASVMIQbIFPGYARHVhHBUEU0INUM9Q/WlvQsu1ocWzxO7EBtu+KD8BqKRjeRUOKm0doPtSltcTGOzkkr8idoiT/fnSNp5fEtRfj9IyqtWKC7l9yZOqSGxHoMmoJRXKsvaYC65zKmiRjGUlDW9J9FHHyTQ0RZGMPc+PV/SsXAYzIeBJvgb5eKcLcQrv4Vv8e66BPmKRG8X4wIj090880/Sw9+g0AZxzv/lyBVcVHa1hfQeIFI3IYkLAf/WhvSmzns4pDZQYZm35vpcb49WAxr/dvNaKAYw2jfuoxOiR3gtM22n8LpeRSAiT6BkE7RX1uMZj34FAwSb/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk1vBvlGgaYRlOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHLsfhr90QTvmICDwKpv1gLAvdp5OfbAB/U+lhRsedS7VK0bXFy6oCg0Gl4td5t+6ERVof3mR9INtFP8SsxxMaGWWQAybzo+wjE1o60Sey2JFvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHpCXuUDj1M3e4DHJqmgAUTYV/WU3qpupr7Z36IFzy/QUfILcYi00x4iL+1Q2ZS9vlk7EXRx5S7nqmPID/4sxHvwpEyFXdzsvjMDvPQvnae4ogi9P5Q05ExOb98+AaJaEDsG+QROCz5dYaeSEc5Yud15hSJ4nVh6Bl2K6hMdSPTRxgPbjk1W9cL705rZ8f+ANBOuf5rG3jMzNs/P9zr8kn/aI9EAkCE4YeoeXPho84c/VwN86OhftVULtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXehEk87TLhIK7TVP9cq4atqRAhoDL61JMcTfs2T3tv7qu+OSEWtOk2Hn2dnAt9eOvpimyvrBUS1oHenPTtAYOt1ZPpqlrbjAIlxF1PLIfOqGMSc+YnhH5GrQW0lrq3fnd/b05rZ8f+ANBOuf5rG3jMzNs/P9zr8kn/aI9EAkCE4YeQfuxd1nIsVGXIuFzLk77WYE34qu09ArhJV9ui98xHoMwwgxUJiDsGag18ZZFxsrfPtbVLvDFqH1AaanXkj+vLpDRDzKAm9d6Ex/DHjOXLPZD59ZaIHdAtPHq5bfbk4rSbPz/c6/JJ/2iPRAJAhOGHqHlz4aPOHP1ZSaWnvZe2NxSQiTI9fxSyrtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXep1l2L8fMII8vT9vLM2vowr2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTLicNX9etV1x/lFtrqO89VPldmD65voKkpAhoDL61JMceRAr9Y3JhT7GmM340wuvpHo0u8+V8CORvGED6cYfjdoNrlzvRZ41imTysGfIDZrZ5jY2T67Es+9y5PpLEgYovSzxO7EBtu+KMb/fvZt05gScUkvEivHQvspCbjHIfzrNblg5fuBTrJo2T4abTESre5O92/6SVl4I7t45WpLXas5uKe9qMUrryjMQT5ndyMiZ/rQWiUhv22ggp3Y617rI1An9JP/q4MDx/ZRd3MobK1f2K6hMdSPTRzsZ+HD2URmm5/b4tAt7nSQcDfOjoX7VVD60FolIb9toCZK83EfNGpxJ/ST/6uDA8dWa7dVyjYxIhhrvt/y+YAdvbd/0eK55LLAWCwd+65pMB8/qeuN/AYlCn3e4CrK/cw0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4ASlQboJTlvsmhdMzPTwDOwFgsHfuuaTA8RlE6A/zVs3kaD45+EkxlnfeNVOspMYZwBcg577jo3opyfhf7Xtw1n9vi0C3udJCo6wAAYY8/oWRLHfzhdxa0b9A8hLrZ8fbYrqEx1I9NHLWNgoQIUVY//gpMCV1TPwcObZP0l+6/KC9nAOXMoiDE7Gfhw9lEZpv+BYdEK+bzarWNgoQIUVY//gpMCV1TPwcObZP0l+6/KBaWMcaIPh6m7Gfhw9lEZps2/ULkhwzXXsBYLB37rmkwj/IJGvCKUf7zIrLTmUKVoiAPT3ILvlS1MaDWF6xEKeaotdUHbRtfyYHjdxOtHWIkfXyJ8er5k6/1Ol2csmiILqg18ZZFxsrf85GvHtroOzHV6NZ9F+QyuC95usJthyqkwx0QCIlGggvg58T+baN4J4OiZaR9YS1rGLnstruChpHkv6JOVIQSsgR95u3QdqexiEYTVcFR9JeYUieJ1YegZdiuoTHUj00cYu5mMV9FnqSOKVDYIywfwQp93uAqyv3MK5mbRf1Nl1HL3gN/E+8VZhqWmfBNaDlHGGu+3/L5gB2h5c+Gjzhz9XA3zo6F+1VQu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6XsYktZ/dqBb3vCospftKNPHq5bfbk4rSbPz/c6/JJ/2iPRAJAhOGHsBYLB37rmkwUh8uL99ptz26UnSdgjFlR3aoYn9Prc44wFgsHfuuaTDWLm3eKt4OT8BYLB37rmkw4nDV/XrVdcd1RQe+066x64ncRifUhYOBFY4XHLxU9YHAWCwd+65pMOJw1f161XXHBAOTJZ275B4AEQbubAvX2/e8Kiyl+0o0UQDEX4lGWKzAWCwd+65pMMk3RwiFK+SuCjN+ccGCmnJw942bn00xgexn4cPZRGabNv1C5IcM117AWCwd+65pMKl8+09yWfa4wFgsHfuuaTAuIzQREW/iCPaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMsBYLB37rmkwOfQe2WVEi0iG2fVKV4V35FEJZt5I6hoN5iRnMMMFpPvAWCwd+65pMPNR81GeG0jIOB9tRAMrmtovZwDlzKIgxOxn4cPZRGabNv1C5IcM116oNfGWRcbK3wJGDnxjoTzECn3e4CrK/cw3Y+bdMpFTIL05rZ8f+ANB96NuItgiCOy/9heHH+03YLcwOH4Kkxp7gTfiq7T0CuHEHpF47UElc6icXrE9H7kEwFgsHfuuaTCJ3EYn1IWDgd922jJLw6ALbzk2LaqHvSwWzCjPOR9fRwhDyp/i7I/XzlVa6Adits3VViQb2qETk6MLY53ZGrdk0ZwJ4FzgqooVI6lt9WkL82o5HDNB0yTFkNEPMoCb13qdZdi/HzCCPAkrX9Ipxjl389ha9R5KfBsVPSuPbkJVcKHlz4aPOHP1ZSaWnvZe2NxSQiTI9fxSyj+4RV4ocmfrpHPm4OFi6edELo9K1Oj4YdNWS4XzWpI5bEhe84m7giw44KuW0tEdOkUHsyc6qooMBs+tE54ZRW3wgwHSOitc6E+mqWtuMAiXCnfuWxyzru9cIHqHcYjGZ01GQlQ7x8nzqFW/4BpViMlNRkJUO8fJ89yo2T6rEYhgNp+ipJFgnO+pCrrM9MGLIuF4dFa6R0Yy0xf1dm3aO3xSHy4v32m3PaDvKer7J+NhH6UHr+EZrBL4A8kpkiKbhJqfRNn5NMkn+APJKZIim4QWu86DM8FPLkGK0kCQb+z+JuArOjbYDxERJPO0y4SCuwhDyp/i7I/XajkcM0HTJMWiAiNHs4agN4V/WU3qpuprpCXuUDj1M3fTjp23SIQxVXAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsRzbA+B/t55XRRobWH6VNQ/E5DPjfwAWCBxuAgy4CNz0QRiZ8n2LLuNBfcgXPscSDtjQ+OWJ1YcqfzM/L46PZoeGFZZ+GnoozRdMvIJxLDCvDYb5zzBKjDG2506y/qPHd9xMJBBkE5JakLtuuCCc/3YQmSNOGFhTFALe6ECZWxlPpUbHuSKRXZTT1hwxVxj8l9PszoAcSSMB5Spz0GsPGwEgkpUa0mRHmH+mscRbAslUmqwxYziKo2Hw6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcnr4JqZBK6Oxv5PRIfaiLNt6Hu9O0DpjbPxScREvltrsHDZMRgFfe1OrGISi5pGmyw0neMfwQeBXHXH094QtKfntBS8LUiOBRSvMDcMPc5Bzqc63Np+FCsZNz7Ynn829T+7bZH2Wd7diX8r03BfIlYzeEIT8M8Gz9hFrKC0Tmdo5WIIAIds2MSqqTY2OIIr/yJ64K/wQvn7Op1hm7sqpRdFOUVnURYOp/yHtmpgoIVG9U7E7IfkUp+TjoWfCVl0JKI+ECzyoDEkO7GNtU97kTE0wdEqJVaiuG5lbwafy9kL9zFuDkwf6hjieuCv8EL5+zm/3UNnM6eLtwuDhMsVKUw/+6xUv2AnDJrOC5IBC2t+/VNsBhRtRIdUPeo34RK7Ax0HI9aDL4/wT4kwCqvEXDadr0IpCVjxOwtfzyeLG5RUgyTR+UIzCD2jV1nSmtbA90OzKeOakhOUTV5gHmKglRiAPARHWGN+GBmbCA1sizVO4cDfOjoX7VVC7cHGcmccaLbdTi1x3mcIYkNEPMoCb13qmB88yZ8LF9p/nWosf9rdvWbtMVWHMD2ds/P9zr8kn/SVfbovfMR6DCZrVxtmjyhmQ0Q8ygJvXeqYHzzJnwsX2n+daix/2t2+jkLKJG78SCWz8/3OvySf9JV9ui98xHoMJmtXG2aPKGZDRDzKAm9d6pgfPMmfCxfaf51qLH/a3b+ZWkZ9EnW+RbPz/c6/JJ/0lX26L3zEegwma1cbZo8oZBEzlrdCgbpySd3s1ClEDb2bN+cK+lOT1uF0OMqX8TPtwRVC+ZmzhmHEK95r9tEWskYxlJQ1vSfRdl4xEjYpVQuOpLZvjIil2VEL8UzMFA/pakulguSmx75ROKHG0m4e4pskNHrHn6gJSbiREETFkpFEJZt5I6hoN5iRnMMMFpPvAWCwd+65pMFYtoEX3NnZou3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6Jb53+keb6tQKdjFwWrwCr3s1hFdmshbkwkjCKPByRQdXmAeYqCVGIMBYLB37rmkwine8xpRL6xHIcjNxEaH/YrqpoQeYQ83uf+fyJyBGnkPsZ+HD2URmmzb9QuSHDNdewFgsHfuuaTAYpj7jys4vT6hCFy47j5uqjlXzZ0RjLO7R1M4N0EZvj3EK95r9tEWswFgsHfuuaTAUvdOMZEde/FB5OylphKT7sey7tg7gVLzv7TWr3ksuSmdfGMBniQifJyOB5VW4JdsASlQboJTlvmsezOrWWHiuDwER1hjfhgbqaMCcyx82/5AvGO1bWzIOByfEHQZfYcqbaCOWQUBWqXhYonbMS0/WVEbpeCnAPqBm1/WBNgQD84LF9nAZbW1Ml5cNmVcIcNL5BeWi7b7m3mL6OwOWFQ/LtFQ7L+vXBuddkINk58cbd3adfSxPiwNnZoFDoESkUlqTV5/uZYAeSFJN4YGgcwFhVNsBhRtRIdV2d0CcBisGtGsmhhMUx8fjpblPvi6KqMaZPeMX2uEKY92aBHyVNoymvTmtnx/4A0EB6LXa4V0EZApRfPLel7n725zi01rOKui9qwVKBkKzMKKQmR2vfjvxkYxlJQ1vSfSJGdz1w3KKxeOpLZvjIil2VEL8UzMFA/oSsyb8d0JLzpROKHG0m4e4KPoO14y1vBbi9lxYgYM1oEND/Oxo/JAorHdbvdZZbA0VjRbT63SkCtxGcCM++o8U3sTWKS3USPBagr3DD2lSFRmSTqVZ9OqIvuUXC7cjHv1mgUOgRKRSWjF++kU5VwnNlnJsWw88qtMNPn4+iTsdlABKVBuglOW+Eu5syMMKd7dE3tygC005pOm3egvJbMlRqDXxlkXGyt8P998TN28thi4jNBERb+IIu3qP1jQmgn4Vz7LnaIdlhi4jNBERb+IIhe22Uz90kSz8Te8XHFbWTxmSTqVZ9OqIvuUXC7cjHv1mgUOgRKRSWtrPoYvvAOhYwP4nrX1JisGQ0Q8ygJvXej5gLDB2+wDqLiM0ERFv4ghtbpVwn8q4oEHXZxRfPv1Q8GJCPoFXPAGf51qLH/a3b0oaPDy1uhLWTlFZ1EWDqf9qORwzQdMkxaICI0ezhqA3hX9ZTeqm6msa0nPZ2637dAV61D9XOMstWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM3JDd1Pv6qG5CPi6SkxdPs1WqPK795RV7gkMbjpKZoMJ5DdTUDjCgNzXy+MnH6dilHARJR6d6+b5+FAT4miU/DKI9jy5HpVciDwc5oBu9e0U1GQlQ7x8nzBxzeiB2SpbBKUOL+0EvdUTn0HtllRItIriVdHoWpqrH4A8kpkiKbhF4exXekNcaRrHEBNYVWkOfy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8W0xLJZl22snt0st0nY2YJUzwqmG99lUWSi0S+dzWtti/FArTAx6F7nLzMZVsHV+5Zdo9Zg//h1mW//Uc/J6m4Mo7F4HwfZbsmY1Alq/+zr3DvX5GuaAcMqXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZvwETEEAloPSFPO6jTFHBOHiQE4QSVh1bFxL+NLuJ8HVjXyMnfXingwGPFzb0e5Y6CfYmJTxiaHl/mX464GuAKfJwVstakVQ4kc5WGRlNKj6p25nh5KDIkCaAPwKVQZqQstGE+AYWW3n0Kur71o/fuioNfGWRcbK31i37jT+RQlYZ/nY7DOAj22zxO7EBtu+KBp5IRzli53X16l9QXE9fX6XlUsPHnitQS+595hQ5cfiWfoJvbUlc1mpolYzQEyQ2sGFSAxSUcbxK+lIboRweD9klm0yLGFEkCi0S+dzWttiDTln+TF5QhjeHv5fPyuFQWxHoMmoJRXK0vg5DvH2KTHkJbkeFXcf5KRtPgDOvscadyY3poxtDYxPWdlcJT28jf0UdzWIoAMcJ2dx1hmkvRVZeqAJEIMTLQ/sY/XEoa46BTwkza6/GlQB/WwMvpibSmVsn5R87rmOpINNJnnuT797cj+2fk46peZGjNYvuNYD/0+nXrAtOe44+QiFIudvQtPQ6howGw4vBbZmuQwQxEKoNfGWRcbK306vW1/XoWKnAcnFhpoXtIfudg7xw+/ONPPNhAEaBOj/kYxlJQ1vSfRRx8k0NEWRjJg5sFTclD0tUi9P2PWKL3A1X02QnciBzIjEpQP5hfCVBTxmAER1YRwbP7hNr+TAqYHgowb2FukwZjySmeLaPsoMHZNkdaymPUhesE66N7zGkjQig8puC3y/3bzWigGMNo37qMTokd4LU3gmErADo4QCyMmm6rvrZ3wYaSML+e4il2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGaju/ZUaNXKlk4xqMc6PPHEZSaWnvZe2Nxka3tvVLY8+YiDHudU55GC2v8Dx/FZSdBAxDl9RRXHVBrSc9nbrft0SclRXmW9paKhwLnsNEwlkpTXsonjQxQzwyg2J8Q7XtACyMmm6rvrZ75i1OBd28aLxDHH9Jv0G4DTVkuF81qSOdz+Xi3QFxjJOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2epCRbrACC7P6TAEs4vVOtOEHKK/IN9j4cQIFmzGG3lmrU2BNkJQdEYEbtc4Cer+/+Jv0RkVwrWmih+P8o/iH/kLvrgjgyEqJI9abCHFWZwAA+JaQRaY4r/q8NAhXGsEW/zF7w80FpKLkbV1of0WE6by/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPNjLuoLq6wnClT+edzSvSuw+6jiTXJfafiQE4QSVh1bEIGrHQECPGvKVP553NK9K42W2bbM2+wP3PpFBtQkSMfqcJVNzczxRKoNfGWRcbK3+NYGn9arYQvNO8PoE4fuf9PkJK4xKvxsL6J+dnhIo92AsbzO9w5pLhZ0VuuOp2LleUu1YUUUsC4XKvnN+4Vo9KnCpKqW9tmuVyr5zfuFaPS4Z1fPxEEO5UQrhvVTDYoK4Qcor8g32PhWAQtwjZy4eUwKaBFOCzwfIQcor8g32Ph9+jA7gNDJq2oNfGWRcbK31sNOOo/QOGaKVP553NK9K4KNED49oYyYtGg2WvKXcaQoPq8dYvXBDhpI8Lldtyg/C3dEWgk/3CQA+Oc1Npth69RY+fnLq7F/D1N9d+fX7PwqDXxlkXGyt+XIk1JlZdjcpMRkOQ5VOTcOtykQczYjX+fAPOJZ5hkzGdAD0Fzenj9s/fOdT+1++tQgnJmgVSSnpV3hyOyNkFbNXqcWlKuB7gN0RoZzEHli/5q4xVgPBiUYk+ciHfVdO6Vd4cjsjZBW1FS9otoLAYq8+YE5l+/3k1QYnf51uKnMH68/cyYin/plXeHI7I2QVsQ0gqCcU6w2qaBP0a9CkKPSx9WdznYh99PWdlcJT28jUJD9RYEgn3vmqbDPMFPyRnTakiY08pStZ8A84lnmGTMZ0APQXN6eP0nHJK7K5aHeyPL/CaaqnEGYX0HiBSNyGLUjJvBEBrO879ss0yn8/uM4Mf5Yij3Wry/3bzWigGMNo37qMTokd4LU3gmErADo4RDbzX4/bSz1HPis7cGEN7FRN7coAtNOaTV4cqecEQZ52DUy0bAGUzIWrOWAxcwF8IpBW9ja8TZKKD6vHWL1wQ4wwHBeGASTdzwrqooOOITCajekj7PLyzlCu2jGFHUMC5mPJKZ4to+yhDJBkHBBegdKQVvY2vE2Sig+rx1i9cEOERkx4hZcdy0Z+Qk3vLsY1yzkW7aevE694D0Wo4hwj4LYNTLRsAZTMgsTRZXXNZPMunbFRHGwnEJnQd8okuZsQkZN1rwBvr+l5P+8E77520GDtRhguZjYj+oNfGWRcbK36A52Yg5nm6MZX5yIL22slpLN+9GTIBSiQldkCFjwDorSNVuMZCqb1nE2a0fTHQJ6z++2+kUKePdRbI5MTZTA1xCXnZi4/Dk2A9xFm7N/6s21g9KUkAYliMlqHv5TQrPwMnQZz73tRXfEnTynOBleyuxiUHlBXT88IrOej0JtLplcDrRmuZdabT1qhHaBp+6N9N+9hMV9g88zSGE3keL9mNq5rJdx2fk7hB+VaJBV3EICLCTAKodqtWo3pI+zy8s5SHVh5/7SJqNqrSHE67+NZ4vufeYUOXH4vA0fQACkeHAEjboyxTc6guWJR3wf86mc0PyMJF0IG0S6aD6fpe+v7CEHKK/IN9j4TK4kLrElPLV8TA3ARFSATrTfvYTFfYPPM0hhN5Hi/ZjauayXcdn5O4isU8f8dfqQQiwkwCqHarVqN6SPs8vLOUh1Yef+0iaja27tgdGMZXZL7n3mFDlx+LwNH0AApHhwBI26MsU3OoLq7g57ipYIslD8jCRdCBtEumg+n6Xvr+whByivyDfY+EqEHNKcJDhm5FOuR6qT7CN0372ExX2DzzNIYTeR4v2Y+rUwTkaCc0Jb3XN+LvwPDrpoPp+l76/sIQcor8g32PhCG6FkUkT0GhwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk5ObRzSM0cQs8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEdb/9Rz8nqbg5zJSvLqzXH7BmPR6RYdZvt1xV2rE5Sg6fhlVPQXF3VPrnL9KIepPJY1OkWGc8TNyuiL0XHn2AGrnh05PBA/u5IJcarNM6m7nhpeLXebfuhEVaH95kfSDbTgDbOBdz1WIGY1Alq/+zr3DvX5GuaAcMqXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZrG4+lrpL6mzdX3J46S/MonjIZ9VzMT1rmApWcMElBKnN1mGDPIL1xBVof3mR9INtDXQWSJFOFAMAOv+cluy8gB3viIW9OFg6+8yDQTOUE5rWQAybzo+wjGZo7e4vutliQwetxTVmz/0TgzDPyV9mV4mXmk/7/DktWDwz9c8cX2oM3yHCRp5cv16eTMFa3S0m9JH4RiFSfrKeCwfEp2J5FiboR8KKvMtE2OfTLT3e9rBuWDl+4FOsmjdWUBMlkrk3tgXt3jDMxaMJV9ui98xHoMwwgxUJiDsGYBsBZkJMrW4D9c4l/IXVcNjewISjbwVy3wn9WtT2F5ray7Eodh8NsXhJKWdRMLZCDF+zS5Me/CUtItpLbTffbWMroHGyZS6tU2OEcWuUO7eFQRTQg1Qz1AXgCM814Ju2Wo5HDNB0yTFogIjR7OGoDeFf1lN6qbqawwetxTVmz/0w/wlsSVTGqeRlO8QHS5xexxxThBinnoikcsTidIjTYvR8WdJFTO+nXRTC31QlktNWAlvFpTYnxx3/s2S3/AcnNtFH8awFvWeaDHA85r5sJmUdCICoMN3FOMW1YAL+x3KicBM2G+IVyFTPPE6t6HRhOi3XtNp/A2H6IvRcefYAaueHTk8ED+7kglxqs0zqbue1QJ2bjeTfs6v+/CmGCc2TWgxwPOa+bCZYDx0oL8iJkpapPPf6YugCL/dvNaKAYw2HyC3GItNMeIffdSuUY3eUAIEa+1M42FMqDXxlkXGyt8VBFNCDVDPUMVCgDEWvRH5hkPRjEXH52vDHdoXX4sTnb/dvNaKAYw2bEegyaglFcpK1bSrLvw9FUwk/7pFIUSvqDXxlkXGyt/+J3a3ILgRbAvrURMFnh5wBPkJgn3q0jx7RlSkO6Ao/0YdhE8XYM7t7SgeXXuAMM0/G8MS9PnKJIG2zufW9P1rBC+80CRl4tJZGp/c0A8lBm2IZAJuaxDkRtVIfZAaxOKTsLP4PzWzu2f8qC/LW0llmMEu+JWkoYB2NTaPghKcHuPQpabB3ToEPfUIhdLbIHB06DpwrCGE2MtGE+AYWW3n0Kur71o/fuioNfGWRcbK31i37jT+RQlYZ/nY7DOAj22zxO7EBtu+KBp5IRzli53X16l9QXE9fX6XlUsPHnitQS+595hQ5cfitUglP28Ri19zg1LbqfhpobWX7IGEZzgnNV9NkJ3IgcwylYfWFh4AQHODUtup+Gmhyz5KDMtsMC1KUOL+0EvdUcHqcCthirvYRvgfyGsBOHjvuK/wRHveq3vQrd0mj4FkHEcuJ+RvSwZNbr6WMYdVBZQbQlB/29fgPwGopGN5FQ5BeIMKod3jqZevSiaXBfrG/JM0QwbobnVfIcjFMbaWmnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR1v/1HPyepuDU/KBFi3pm70UO9zbFzv8pTuH59hwIt/0T7V6GhwcixwL8XbTEN/l19ZxZQyZcXiXHc0dz7Wr5DWVe4rPFKp5N78nV9fJNxz9QgjmsVHNyn6AGrWzzjTqT4VUy7W+Ais8Pidopf7gsC8K01dMM4NIcTwvuFIuNWOKxVjc6Uj/cvHiD7GLyyFzLlfPF4Iq9iGx58NLjUi7Tdc99FpVoGdKsvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHDB63FNWbP/S8YqKDKfFsWsiYmsHgeVfiIPEEOOs5sYJFhs+T6mvC3Bp5IRzli53X5CRqz7/gFKofUxVuCXS5Y32Pkite4rtGKQ9XKZKOL02NVcWq422EsmFcV6pKQIgYBUpe48G8Uie9P28sza+jCvaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMvcaLydpsQM0S7519g7oX491FiiUOkfRs6a35DOqZ0CrvxFCll4lpueoNfGWRcbK34+SAElTCEGyCnfuWxyzru+j1LPZE6uc4jV6nFpSrge4FXzu693lZFQFSl7jwbxSJ70/byzNr6MKWhfB7jTkExej9a4NkQvW6dOL9h5nT1XI+u6WYUl9e0jTF/V2bdo7fGFmjN23bm9wM1ILnQKCFfPmjKghd4lsW6qF0jQ4DNTTMHiwATbD+KjDPI4Y22ZnyfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln52hlMwyRSeWoQ5YD1YTHCJzV6nFpSrge4iUiQ9QcZfDg1epxaUq4HuKKdQxa98qI6hdcP5rXzimU0hwqTZwXP5FnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZcH53YEX2q4K3exMfZSOej1QEpaRNSjkmB4gaeQMtWMLncL9tHUV5V6tP/8iyWTRRNb/9Rz8nqbg0pNePUEsCYGWQAybzo+wjE1o60Sey2JFvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHphePuqkHOmSYN1s6Sk8tYYV/WU3qpupr7Z36IFzy/QUfILcYi00x4udtI/0UeRgdZFdkSnhQ3bdyErauFowuZk/kMqEp6+Cp4YUHeRv16uTmIqollrQmauNZNOv2MOqRPFK05csjrHwW4s7HGeisBS8HZEGoTxCD9bWzbnugrBgMHZNkdaymPV/OWn1CD01ZUQlm3kjqGg3mJGcwwwWk+9jEzvSCEnoJd8hkN/tb/HUee83d/nVokbtwcZyZxxott1OLXHeZwhgETOWt0KBunJJ3ezUKUQNvZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYcQr3mv20Ray8iRQVfy8GYy20xkzWGDMO+ZC8n8a2DmpnhE/Ldsm2hBDlgPVhMcInNXqcWlKuB7i4eRyaWfFBYMA900UoGRKm2yooR3rR3bG71+pmN5dPwjqQZJOAjFEmaTX623ZVV8+CDEqk4KN3Coc9ERpnV/PIUPgVZBSMS11AODvAcOIFprOm4GNjZXJtwD3TRSgZEqaVhqsillAnUrutRDCvk7ipOpBkk4CMUSZpNfrbdlVXz6kL/+Pr3Ch+hz0RGmdX88hQ+BVkFIxLXStS3T/7WIGWs6bgY2Nlcm2tMg/TH8AwMJuwpfyRpuHUTMzqNaAeQE1lwStUaipM/JdXVEUhgA60l2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkzn2Cf6wkDYmIU6DqJ9JVmvWmnH9BH2l4KhyurFjgufo8ge0hiyqaTekVMR49ZXf1XlwIK+2YqHXBm/tDoEW3H3y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTQxvlIRzAKu4T7L7qo2pqAaFf1lN6qbqa+2d+iBc8v0FHyC3GItNMeLnbSP9FHkYHWRXZEp4UN23chK2rhaMLmZP5DKhKevgqeGFB3kb9erk5iKqJZa0JmouxPUN2+8SQsMqztNYZUr1dqhif0+tzjihKlCAG3SxEtSMm8EQGs7z9qoHINnqNTQT1zWClEYtH4XLjiOTjsUyMZzec4NYb6YoIKa6daczlDQ68/3TNPUeGmM340wuvpGzpuBjY2VybfOoYXf/L/aGpxk0KAaU9eZuCUJl+r1Ko6+dhSVvWRZXV5gHmKglRiChKlCAG3SxEjxStOXLI6x8NdbDn1NlOuTVpEbPMriWNSKcIW0S4ke4uHkcmlnxQWBgrcIThxdfFwib78JuTJdWF5GQDUhGqxiByiCpLrgl/tsqKEd60d2xmTZNdyfyGW5hXFeqSkCIGJWGqyKWUCdS6W7ldRrs11NZCgVqQqiccNWkRs8yuJY1RIxvErpswl9OUVnURYOp/2o5HDNB0yTFogIjR7OGoDeFf1lN6qbqa4BwIV4xUvMsOlu5v9spQ1T/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyPXyMGM0AOB/id2tyC4EWz5kLyfxrYOakb9FmBzmM2bD//YU7iEetlWTPX5i8iVPtsqKEd60d2xo9Sz2ROrnOLCxkfGYxEhttDnumNqBSSRHNYQoPY+k1ez8hPZk9AeGbReBOnbSegyOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2Scckrsrlod7htsEJq8gOaX2qFdVP8L/mHkDSvrx2tRcC9/atjq3bzHy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8U65bNWSRgdXfBIDRqGKAPpPOv9kGa7RsEsHmd1FUYed0JXvIVeIyaSy20T5+B+osGgKKyLBBcfgpH+iYXN2p5bgUVVy1alynwh8gkp9XXDmoi1Hn//j9/A68tJl60JPbzUqggyLD3Y9J3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb4VBFNCDVDPUBiU/p0DOgML7uCOwCkqMmV1X8bCTYx+03E8RO4Xfrw+CQ2AdkZql9BwfFE3jEDu6zdFhZVMWKsl6dGM3GzqJngwHeFlQlDk6dAYj6W7Itm6BdRCVefspm6jwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+yerg4Gueif9EJD9RYEgn3vC9UxHq3ksia6oe5ZwWKZz2bW3QOh4GysKsEgrZrautUsRcaZ+A7Ms4S5RxUgSUbFlfBDV8O6w2tafV9lbSLkiWAhKDvfFWaU+b6XG+PVgMa8Dy7ngtmVyvhoiL8D6lHOMZaJukqSckHL8ElX1S2IiWIE1XX73ux6cJHkeyCHV6+4ugDXg6fOP3NRNUNpanbR6ihOEYXlsHFldhL9taLl2nARTTIGopTtq2c5LF+tfNvSJD/qZn2kQVN82YRSaoyBjrhFco9P5yAua5OgYUwrP8vJyVyAn9P4q4j0S+aVfp5Lek8xFmzmIlJTuU3JkJFImN40pX576szdHCWTaRlZArT9KQ3pbn9G0JXvIVeIyaSy20T5+B+osGgumaGAZYcj0ohBiw0TNk7gUVVy1alynwh8gkp9XXDmoi1Hn//j9/CHfONQ67SkrkO+3ASB3K3ySp7agx0oPXIpUXp5yCcn5nSDCgXY/oNQTW6+ljGHVQW6oe5ZwWKZz2bW3QOh4GysL4tf+y80onMVVXQXeypM9IS5RxUgSUbFlfBDV8O6w2tafV9lbSLkiURSFihkcs+fT3rSKy8BbrDLyclcgJ/T+KuI9EvmlX6eggQgvlkfYpW0/SkN6W5/RtCV7yFXiMmksttE+fgfqLA+onDamL7IHtKIQYsNEzZO4FFVctWpcp8IfIJKfV1w5qItR5//4/fw1+eLFBUSCKVxtmIHGMoxHBuoeql1QGPUL5jRi1VXD1ApUXp5yCcn5nSDCgXY/oNQTW6+ljGHVQW6oe5ZwWKZz2bW3QOh4GysOAbGlV5h170VVXQXeypM9IS5RxUgSUbFlfBDV8O6w2tafV9lbSLkiVwK/SzxUqqtbDWNQylDsBgDByv9ndSrsjQEm3q+H0Yvo8DxcgTS24wpoifs1g0sYtzpl+SIzDkjFjQQ2ZXZpMatoa1lDJPN9PggHRm1WjZXXh44Eru+G2/DFdE/EjAVqFrVGulmlxBWtVFsxpT1HcQRvFg8OY9A3cWJVfx3H+Pdy8nJXICf0/iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUjv7TWr3ksuSlHl+9yKWTJZ5up/OZQTrX9Hb5ySiowbTfg+Md4A1ysMsOW9w8BUFblrS1TXObGJThhg/XGD5XiftlY9qxRdVGoo1DQgBUbZZPgDySmSIpuEvA8u54LZlcr4aIi/A+pRzjGWibpKknJBy/BJV9UtiIl+rIoi9GbuAebcn0Z4Qa4iYAcQM8A6degxtR3Q+abawLc5BJnnohG7M7kKG2fKh0coKmVcgLNIxVbTORy73wEzzrogeifzvRR8jRLnCqHAbj5gLDB2+wDqLiM0ERFv4gi8Dy7ngtmVyvhoiL8D6lHOMZaJukqSckHL8ElX1S2IidSjzaTTxMv4vTmtnx/4A0FR5fvcilkyWebqfzmUE61/R2+ckoqMG03e8fXyb78Qq7DlvcPAVBW5a0tU1zmxiU4YYP1xg+V4n7ZWPasUXVRqdBxwy5bBKlCSNCKDym4LfLwPLueC2ZXK+GiIvwPqUc4xlom6SpJyQcvwSVfVLYiJvSO24h1WXGr3gklsGh3IcWAHEDPAOnXoMbUd0Pmm2sC3OQSZ56IRu2ZY65kZm/ZcKCplXICzSMVW0zkcu98BM866IHon870UfI0S5wqhwG4CyMmm6rvrZ72qHWF7qOUAo8DxcgTS24wpoifs1g0sYgvlmBdWPHvsKRJhnplZbC+WJhxp7A9QBcMVHSMhCB3Emxzv3OMGq/q858KL7Pjc9sL+svkxfSHxNRMLgAVFn+dM17FUngeMAWzl9rDa49LyoQzo+xFDDesNjqHLZaF1TvVnxGpsSXtNc20Eq1oO6lop9Wi3byhVE8vJyVyAn9P4q4j0S+aVfp6CBCC+WR9ilXTxKxSkSzc8yLXF7GE8qgRFMyLAKz0jJARMY6Ga6wBxOFEXvkZrU2nib9EZFcK1pnnD5FlFAUS75SYuCB4yNtkAFjRhzGDuItCV7yFXiMmksttE+fgfqLBgJ3I4+djqhl4eOBK7vhtvwxXRPxIwFaha1RrpZpcQVrVRbMaU9R3E1rrLcksw1OnRON1SZ/eXZZ3cS8KvkPuHlIyGaEtDN/foXtjLQPXKgLU+dvifs+5uvA8u54LZlcr4aIi/A+pRzn7e4xvVnKJTmVAOLjyeJllnjIuUFYZHg+N9bq2d/DkWb09PynwLIq7o0u8+V8CORhY0ENmV2aTGraGtZQyTzfQ5M57ySSiSNMbhvgkPW9unpH+iYXN2p5bgUVVy1alynwh8gkp9XXDmoi1Hn//j9/DZEmj/kKluE440Uyxw0ygVfHm6Mz5irVCRC3g4juBGEeB38mpuzrnD53NMrwVe76uZYzuyDub2ki2nfLt+ZNl18ssgR/LIf8TO1vv0WSUjnGB3XgZZNAPjMBfWnVGZDT7WSWAw8/wUNAAWNGHMYO4i0JXvIVeIyaSy20T5+B+osPI7fLeAu06nXh44Eru+G2/DFdE/EjAVqFrVGulmlxBWtVFsxpT1HcT4T753QHw88fPJTjsgBIGZHa6914cfPfrWmH0QnDKBijzdrqjwcFWlYw1QmDWJm2knenpDSLhBEHcgbE5tYw5FEpvLiZo19zyo3pI+zy8s5U3EN4He1lQFb09PynwLIq7o0u8+V8CORhY0ENmV2aTGraGtZQyTzfQ5M57ySSiSNMdajQNPKKATpH+iYXN2p5bgUVVy1alynwh8gkp9XXDmoi1Hn//j9/A4HlizuWTCiurb5xHV4PaABForUTxmQ5bKs7f1SokZXzG9fqsAOHIUiUL0t/Mo4NQ+3wUp4AHlaZpBVhazntdDClTOQ4fmgDyEHKK/IN9j4TAX1p1RmQ0+1klgMPP8FDQAFjRhzGDuItCV7yFXiMmksttE+fgfqLD+NpmSBJn7m14eOBK7vhtvwxXRPxIwFaha1RrpZpcQVrVRbMaU9R3EZPtg6tBd+CQvPwrAjHHIVpSMhmhLQzf36F7Yy0D1yoC1Pnb4n7PubrwPLueC2ZXK+GiIvwPqUc5+3uMb1ZyiU5lQDi48niZZpKFk2NHyLDko4jTCFjRv+NZJYDDz/BQ0jl5YD7ZmhyYIMEmt5aG1PeAwa8Ni+6HHG6CItCHO0RQWNBDZldmkxq2hrWUMk830S8PFom1+yV0Efl3k1vmx+bJKxY3R/6JnInGe6JgvBcI1EwuABUWf50zXsVSeB4wBbOX2sNrj0vKhDOj7EUMN653Y4ycS9bm2rWz420kd3WDrxuw4ifj+2w/IYWiIqjyhXlB9PcWZIkk/XWJqccLGSmAHEDPAOnXoMbUd0Pmm2sCbUmNyJGMmv3Io+HkVcgLphByivyDfY+GYFx+lJCXDALDlvcPAVBW5a0tU1zmxiU4YYP1xg+V4n7ZWPasUXVRq0Mu6t40wzZNNd8JeP4StuSxcOq7ltmx0y8nJXICf0/iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUg0eO9Xo6RFKVNzngGgdFHYuLoA14Onzj9zUTVDaWp20eooThGF5bBxWw046j9A4ZopU/nnc0r0rqVbInNIQl/LXh44Eru+G2/DFdE/EjAVqFrVGulmlxBWtVFsxpT1HcRv8dLjRA9o3OZKPmxb5g/j6tvnEdXg9oC8Dy7ngtmVyvhoiL8D6lHOMZaJukqSckHL8ElX1S2IiYPrOdjFKeWSf0VZZq3eQ6e0/SkN6W5/RtCV7yFXiMmksttE+fgfqLCcNr9dPqO29VpoAb+70/qtp8974Fqk7GwACBDauxhAM3B8UTeMQO7rN0WFlUxYqyXp0YzcbOomeDAd4WVCUOTpr5Tvb3fE+wJ/rmtZlAA7yilRennIJyfmdIMKBdj+g1C7ZNdaujmE8tSUW6vUOi3IEOWA9WExwieNOQJDgAgCarT9KQ3pbn9G0JXvIVeIyaSy20T5+B+osJw2v10+o7b1WmgBv7vT+q3BPf2YkVSMqgAIENq7GEAzcHxRN4xA7us3RYWVTFirJenRjNxs6iZ4MB3hZUJQ5OnBgOZj5nk3XX+ua1mUADvKKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTy1JRbq9Q6LcgQ5YD1YTHCJ/9ADaGcPqDstP0pDeluf0bQle8hV4jJpLLbRPn4H6iwnDa/XT6jtvVaaAG/u9P6rYaHfrTu9+b+AAgQ2rsYQDNwfFE3jEDu6zdFhZVMWKsl6dGM3GzqJngwHeFlQlDk6UTCiOB3QGOGPGoMTr9MUY4+3wUp4AHlaZpBVhazntdDFXX9LD/Bi695zs5PRIUJliwfVEDW7E8KtP0pDeluf0bQle8hV4jJpLLbRPn4H6iwnDa/XT6jtvVaaAG/u9P6rTTMCo0+Vrj5AAgQ2rsYQDNwfFE3jEDu6zdFhZVMWKsl6dGM3GzqJngwHeFlQlDk6fdMSzxFLz3rPGoMTr9MUY4+3wUp4AHlaZpBVhazntdDFXX9LD/Bi695zs5PRIUJlqwbTrb/HNEQrHEBNYVWkOfHuhOXTeaFEQQTKhkCMCgM0RRoVXO6yLJwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwyKEsl0DET5ohz+Pg21Gw+w0zB9aWHlcmao00x1enIKFJVOS/zOfjAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctBWUqh8ccsm2utZi+wc2cjOx7LgKysZ1ioEByRFu5q/m9ftHBTauKeUesELTuRK270nmAeVpWqKqvgwI9x/utdQxQ/1o3LCLDdI9OVRdvOOQbCAZ+BPqfjm2T/oMotMcsB8o8UlyNZhmfKdOuCiuosGwRjmsKH3H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LE6S3a9z1k0WeUUQ57P2dZ/D0yVYSr1ZqQun+fadIqySUzsVX+qjJ2VWvn3zt+a+vNGzsQ7/B5p9Qw2GSyqIWv4kAEDsXn9JOtWHT9AV0+9AxkL91+oXh1Fsnph1GMPMA55MjocTbh2KxrN3wl7KRmuqTrZEeUCO655MjocTbh2JRJUM6pmF0UCCJTZ0WDcFxND5/1YD7AQ8v94TlSlGhCWL0YIzvLQ8VIqrp3xKIxtCCeBlNilgh9jJakekrNK1qG0skx/+6q3EjbPf3JibGS9KAiuTcO6PxjmJuTaztkfoSNujLFNzqC1NXU7Djqa5y6pOtkR5QI7oqjDr0IxGcVHHFDMsSomWTTMoZ70muRJpP32Qsz4x1ZmgxwPOa+bCZBAGEBFqQcFrvLBREZBsyKfMRCa9OZHwqG+fEe+nYDkKUuAH1jBo4gxeMhRJGnmIsV5ACII8eqG90T/hMTF3EP0mVALdrAqT407ZvP/PYbvG01EeehbpGDTfZ+KJDEY0ENVoVs56o14VLl81jhiXDQbiORkZlhxbX8+u7wWiuaDC+cPQZxIfoJABvQxf6LC66EgnnfcfbgkxZYgTtv5fy/vUTMJsCpZTYgxI5jQR7b3bUo8zBLpmHGjNje+Ce4Yw3uAXmsIu8x3NUKWfrZ1reWCalmxDBvT6ycV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/m6EfCirzLRNmAmFR3LKaecIKQH9xapKWp3F2/KZDZS0FSl7jwbxSJ1xLzhnLPbnBrD1oOhUnp8hO7JRb/x7EOGxHoMmoJRXKqQ9E78HC2+We89mzNgf3y2/3UNnM6eLtwuDhMsVKUw8B/WwMvpibSmVsn5R87rmOi32YOSX61aiPhAs8qAxJDuxjbVPe5ExNR2fVmEyqvVO2Wc5osDyA86M1l0e/dWYvYqUN4zQ2F0vCCkB/cWqSlvj10qKusZM22yooR3rR3bEb6fWz5DNEYItJFi57rHJCupmkdEVpLFttRd9iJfrOFNz0JJUew4U+gHZAyG88J4kHCIkzAlfR/DGTzC+tFdi17GNtU97kTE2foAOLnMoIH5YTxDsJ4TeBwNj1ICFNcO9UzPyzuUT83Si+G04JfRlAVFYclhD8d4c2PkIZHX1pOctExGHgI65b+PLhl1syijoxk8wvrRXYtexjbVPe5ExN4UHRF2FP0mzG7Ce+W2HfcW5PdQuqMv4NkTk+9SxN4FUNfP/1CBud8VW7inPYRzEOizw8Fsbag5INs+RMmCND0gS0SN/g8i75+u6WYUl9e0ggLWZKS10MIK+HjxaB4B74rR508ZTGndHM+H/iUy3h7vEae5HQ/VvXK+TC2YUt5PaH/7UNU58jTmZDHMAELV1tUtKXf0qA26scRy4n5G9LBoVVIPUUpxe0BLRI3+DyLvllbJ+UfO65jsIIPxBr+NBQb/dQ2czp4u3C4OEyxUpTD+dK/+s2YPEJzWsAdRETu3xjBfVosytm4ymKbl2BmuF0a9CKQlY8TsIr5MLZhS3k9pW8RIof/QllPS2honXOFi8UsTqDL4pc/ViCACHbNjEq8kyiJFHAjB1pQKpSyhKwaWMSvbi5o+Y3koejOOHQ5KPIlqyTjvEGuOHDJoDEt9A9FIjp1DOt+yeysXhkHKmrsPr4MdQxzMMEi0kWLnusckKBxl0y+KwUu21F32Il+s4UC8g1E4M0/TbNpa3ulvgHiwsyjBhW1qfXHEcuJ+RvSwaFVSD1FKcXtLVuaovWGxGbZnbbokUPDio4jPCkSyLcEViCACHbNjEq8kyiJFHAjB3FTczZP+QykJB6Fx0PxWyUKX6FkM9GFm4BgJmCwtDu5m1F32Il+s4UpyenXn87dN3f3rwpcvsKaMIIPxBr+NBQ1hAIlb2xXDLC4OEyxUpTD+dK/+s2YPEJu7xPZGzdaLQ1Zicz6VVMhKuMjhEadZ2SVFYclhD8d4dBboDWT8dzI21GcBp30haZkoejOOHQ5KMsK+jXre5gqOHDJoDEt9A9FIjp1DOt+yePkgwKL7hwuSXl9AvMcPsPNWYnM+lVTITUYceLkRH/QUfw4xTZ2SU17GNtU97kTE2caiSB0pwUU+7zJ4//EO7L6OpIWaTfNinCCD8Qa/jQUE5Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCT6ovuNWQ2fyTn7El89PXU91YKbw3tpRShxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnNPi6uk0GLKYwgg/EGv40FBOQZIm7+zr2MLg4TLFSlMP50r/6zZg8Qne2+IB6jW2q/3QKvhcCLHPMZPML60V2LXsY21T3uRMTW9zv0N7Jz4/1SRKyncGKZvy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Jhvg2ORkfDDZs/fOdT+1++vFEjVycPxU7PL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx0wTryAGe+6t928nvhV/4hyZeaT/v8OS1YPDP1zxxfagzfIcJGnly/Xp5MwVrdLSb0kfhGIVJ+sp4LB8SnYnkWJuhHwoq8y0TY59MtPd72sG5YOX7gU6yaNboZH+dJQSkMHiwATbD+KiV2YPrm+gqSkCGgMvrUkxxN+zZPe2/uq5hXFeqSkCIGP0UdzWIoAMc9qoHINnqNTQT1zWClEYtH4XLjiOTjsUyMZzec4NYb6Z9HcjokmCrV7twcZyZxxott1OLXHeZwhiQ0Q8ygJvXes1rAHURE7t88erlt9uTitJs/P9zr8kn/aI9EAkCE4YeDCuNVCU7v0plzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZqwJQiQW/mp7fukZUgm5l+TxMY7OSSvyJ2UQDEX4lGWKzW6GR/nSUEpCdRbueM7dJ7PwGopGN5FQ6yNcfwmy5SoVdhM5+RokiElpxU0j/k+QlLIwQy0msMzlkIQXZ/yiQaUjFYObx+9iWoNfGWRcbK34+SAElTCEGyCnfuWxyzru+j1LPZE6uc4jV6nFpSrge4FXzu693lZFQFSl7jwbxSJ70/byzNr6MKWhfB7jTkExej9a4NkQvW6dOL9h5nT1XI+u6WYUl9e0jTF/V2bdo7fGFmjN23bm9wM1ILnQKCFfPmjKghd4lsW9ME68gBnvurPXCvfBe3t3VZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk0MSw/dqK9HHl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGbqQ6X+shkHMeNUxfXBXYbMmV9Txacs2bug7TSb/dl8EHMki6J0QlCAbwUqEt4rQwe5MpoukXyeLmhV9xGVcXRVXQsGJxv3izAosMKZ2Jht7/B3px1I6lodPvkv3kOGiSnrXvk5qWty4JT87VPGePaFX6/m8gwCuzxkUXjwUTdvy/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHFQxf91Swmnm49eKqao4hlmVCiKiiXiKDw5GeydvR+LBu3IDn6lmkA+UmLggeMjbZVee9VOtSicmFwEJscIKK6qoLH7uFVaIihX9ZTeqm6mvtnfogXPL9BR8gtxiLTTHiIv7VDZlL2+Xm/fPgGiWhA8xBPmd3IyJnHyC3GItNMeLGLXITHOJplHEK95r9tEWskbt3wfQLWjObbwVYsPoY/zSc3R/HQ5ndZL+814w1rJYvxMuc4I56TgwrjVQlO79KZcxmz9AAC0ynxG91hzMy4FFj5+cursX8ETuc2nyyzNzmIqollrQmaldhM5+RokiElkBxnmLWvZNLIwQy0msMzlkIQXZ/yiQa0M7cUjtjT+moNfGWRcbK360yD9MfwDAwgz5oQLaYuGaFf1lN6qbqazGsmlPuyBhn/1N3sL/wjOA9kqpak07eS/k7xzX9fu4goVAu7SfhPtbB19WHuPejwuxQILc3cqlTzR/2Q4FWAB56SX2VhG97q2VCiKiiXiKDw5GeydvR+LAo73sTQOvsWz3wXqYfXsKtdp19LE+LA2dxDs/sYIBriSVfbovfMR6DMMIMVCYg7BkzUgudAoIV82UNpLBUAVv7h6N3qfsu4mVVzrtOR+/2cFnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTQxLD92or0ceXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZgsZAZgJDrkq+8BExJlLKEiBv4yF6xOLjvyC0hAnOffNPfO4a3aC/XQ94OhrzgOLfAJxW6TTM4W9fKyQYqm1/u9aoP+zE5GtlH/LBJJt900o8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTsrNWYQz+pTCyL91jI3Rw5eaMqCF3iWxbLKorACqS2fQnpv7XU6I3MQAaS5MeA3kgZcxmz9AAC0ynxG91hzMy4FFj5+cursX8ETuc2nyyzNzmIqollrQmasKoTt+qWcx+rfa8gq17JyA9SVUBaqrPg5XEitdKzVpQLtuuCCc/3YSJvNcwrG43Q8ffPy3ykWGRwx3aF1+LE52Gha5pqfgj8JacAGSF9jAb2K6hMdSPTRySoGtWHrMQoGMSvbi5o+Y3s/IT2ZPQHhlZt+SqJtO2gMBYLB37rmkw0BiPpbsi2bpThMqz5WPAU0JD9RYEgn3vkNEPMoCb13rskbMZwXu+eQVKXuPBvFInvT9vLM2vowpU5uizxpm6iVeYB5ioJUYgwFgsHfuuaTATGOzkkr8idg56ROpl9LPnQkP1FgSCfe+fmmS/7b21AJKga1YesxCgi57bcuegZJqz8hPZk9AeGTSNAh98z+tTqDXxlkXGyt+tMg/TH8AwMKZhREc2ssOTyz9Mojq2luCT1+R2gqRopKg18ZZFxsrfZ2eOMjMuho3AlCJBb+ant/xBnBX6pjn76uobMYIPNeSoNfGWRcbK30l671M8yflSwJQiQW/mp7drz/tPb3CQNR+EuPHdEZ91qDXxlkXGyt//E3P0C6tcADT1yjnxEkSvfituwZjT2jzhrEhB5K5JwTpYHflG6tYT5Kj/ZRoAgVDMQT5ndyMiZ8CUIkFv5qe3q0oMMMiW2kldFVsT0GpUWb8RQpZeJabnqDXxlkXGyt9nm/HbccBj+s/eQWe2Kgu5mkR55UAY78q6z/Acd5Ia+eHcdQqbL6zZqDXxlkXGyt+pfPtPcln2uPiPZQgtJ4XXSEOEe6b9Y4sb1j7cjHuy3+wNykNFPTcGG0valbzf4elKXBKO9XCukL2rBUoGQrMw43YVY774KSGTcePKG9wAs0hDhHum/WOLa5pyonMfqRvkPfWwECyyiL2rBUoGQrMwvnE5wKNaMBRiCjv/vpJYcJMF7ANKa+yJPlzmJopa7f7y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPFpbEnY3Ckt1nKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZfLbMWGDxvDKK+/YdeoACsnnV3Mce/w92fy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPJ+a4mRx7Kdet07PxdIyzOjbLqxK00IOWFf1lN6qbqa+2d+iBc8v0FHyC3GItNMeLnbSP9FHkYHWRXZEp4UN23chK2rhaMLmZP5DKhKevgqeGFB3kb9erk5iKqJZa0Jmp/1uAcjxO4n1gXWJF3SUPYu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6lGsFPNI15xUWr4hOtznGViVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3z1fALIrSJM0qfGpLh8RcwNAhoDL61JMcTfs2T3tv7quVVtw4ikZM8KBvmiZ5/gwsvaqByDZ6jU0E9c1gpRGLR+Fy44jk47FMgD16ny9fmk7HUb7o88XwSK7cHGcmccaLbdTi1x3mcIYkNEPMoCb13qN+6jE6JHeCw//2FO4hHrZjRBmQQXz8GWoNfGWRcbK3/4ndrcguBFsCJvvwm5Ml1YlX26L3zEegzDCDFQmIOwZqDXxlkXGyt/+J3a3ILgRbJ3j9Df7gZDzJV9ui98xHoMwwgxUJiDsGYBsBZkJMrW4D9c4l/IXVcNjewISjbwVy3wn9WtT2F5ray7Eodh8NsXhJKWdRMLZCEWDixS+Zk+wNN4j7JAuqQoJ9wpaONExHbz5wJKYI9cX6LBBjaQcy+X/nXd1gCviNJDRDzKAm9d6lGsFPNI15xUWr4hOtznGVrSkkB3ZsLwyBfbMsDNHeAQDebtNyiW2lttbv+xeLKxwQvZOoeWO9V+PkgBJUwhBsgp37lscs67vJQrzcTNzDzjLk+ksSBii9Bhrvt/y+YAdPqi+41ZDZ/IMd8dMfgkJA4+sD0v8t3QaPC7n3244wpn3GKSbJQo2s2qObKHokHBEMHiwATbD+KjNfxxZYVhC6BE7nNp8sszc5iKqJZa0Jmq/Db78aSN4/Qib78JuTJdWPV8AsitIkzQXgCM814Ju2ZHHobpjcJk1s6G/BDHDNQC91ZxjHmU+SLyPmdspFBHYl+VJtD/uv6A2/ULkhwzXXqg18ZZFxsrf/id2tyC4EWz5kLyfxrYOapJIJff7NywdvGKigynxbFo4IDZyRuYUTJDRDzKAm9d6jfuoxOiR3guQhsMj3WeLXN7b4gHqNbarn5pkv+29tQCnC3EK7+Fb/ExXPmRW2GhfjrxshDSOUUXQxjvZI/ggvxD0ExRs9ghbLNKtkJNGg+W4EkG4xCRtzP05XZUYVPrNR07EIzlhgQNEretmpTjbSPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4mNcckY+0YJ6t2BRUdrOABUBKPN3GUEFpf7seS2ir8i0ruTV91SZC4fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwuJKt7Kze/qfEg2GBGWdp6+ba4tYSGGu76g6WVlzc1l0pOTpOcBgaCoXHACojHgtWWxd7lNh/wwskDvGcVrJOJStW35N7S1tYN/XtlbBqfF9Pa2rh3gftwJ/AYG4VS7mGU62YvjZ5yzqWypkCG8hA/837uhci3nvipW9EiFfraz+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/SOUqXqc4IdsI6Op4SZut/nDzHsULEgQUFnNNo97vtp0uXiEffkxxqc/Jhw+MxWm4J4GU2KWCH2o7IgfUbYao66E0Ypsh6pbTKbtlqu6/gxKow69CMRnFRYhtkfcJFp3rb/uHctfBfgiyv7FCOOlfGHY0vEVzVeKfPxUuxmn4rWFjocVPi77H2HKqogxnApEgz25Ac0HZheKs/Lo8givFfRRK2AynbnX57b4zPPKA4pOKemJYYxr9/CkKMGaZiAxdd4nH42vs1UalGkJ+i79qGimZzjQEhc7cBYLB37rmkwXCjyJM9eBPPUqcS18oLPlSH/Az7EINaUyCsc6J41TV1CVpf0fc8K4MPxbAaJM4pXVASjzdxlBBZG93gikoryXwjqK/Yt6Um04m/RGRXCtaaKH4/yj+If+bHqvjDwRwgsIPNywDGMkGQMHQwXOl2lGNHz0brRV14uvIhTf0r0kntd73vksJ/7u4MQLhpxmxu6MPenqpFMMafoi9Fx59gBq54dOTwQP7uSlPGwF7a1yULWmH0QnDKBilVIIBmEB/f+AEUrsNWzMJPCkKMGaZiAxQHvIXKjGBPsLm7hilQTdnbkL7++j2RmPV64AFrmEp/GEjboyxTc6gu+f8CkopUc+Qz25Ac0HZheKs/Lo8givFe2GBR+Tp587aMMNbS4MtVXJLVlnCRieQ1bhom0J0WqgJeXDZlXCHDSLwL0gn1AbsspU/nnc0r0rmDHTBgTqXIz3sjlPbKKDcLixS0fZB1znzdEspXdWi8xgt08FGkSxVbR03DvDUKeAZkQelFZ/eLjI94KHVBpBFUI6iv2LelJtNGg2WvKXcaQoPq8dYvXBDgOdnVdkll0qSDzcsAxjJBkI1sJXBjhEq4YALFm55Cy1ryIU39K9JJ7Xe975LCf+7uDEC4acZsbujD3p6qRTDGnWw046j9A4ZopU/nnc0r0rpr33IXWN3AE1ph9EJwygYqbHW3sedOO/ToxYt3pSknswpCjBmmYgMUB7yFyoxgT7C5u4YpUE3Z25C+/vo9kZj0aKd3IU1VzAeJv0RkVwrWmZUrld5ojtCkM9uQHNB2YXirPy6PIIrxXs/44G2kt1zGjDDW0uDLVVyS1ZZwkYnkNW4aJtCdFqoCXlw2ZVwhw0i8C9IJ9QG7L+dEk1VgbrDkUoNgNHZ4w5TCfeTM9uG9xq80jmz7Dkh4Ouoxb7ZIcKe9O9cyzyc+00dNw7w1CngGZEHpRWf3i4yPeCh1QaQRVad+WbYZY/O1oMcDzmvmwmbl9wsIcAO/aMCAsaLkc9sMgi9P5Q05ExDveSImX13A0+XS6JX6v8WPBH6ab6nFM+gGrw5g00TiR6vwdSZBVz3vBD69SO8F2PM1F4WizKZmEAf1sDL6Ym0r67pZhSX17SGJu0vDWy4qIlM7FV/qoydnBYUSx7a+c9hUEU0INUM9QL8StHlHjq9o1Zicz6VVMhO77j343mPw1VFYclhD8d4eVd4cjsjZBW+98B1Mj5z6UyVCHDB3/kezqfUNT01XmRmvQikJWPE7CNuF9Szb8bc8riyPp1ahjhlHHyTQ0RZGMUIJyZoFUkp6N+6jE6JHeCw//2FO4hHrZQhQaHWyXaE8BYNAncoGkg0dn1ZhMqr1TtlnOaLA8gPNZ36WaPk0oGzGFM4H4efwuTkGSJu/s69jC4OEyxUpTD2F9B4gUjchiHNYQoPY+k1dCFBodbJdoT3VgpvDe2lFKHEcuJ+RvSwZzysUlAo8iA21uXnOUL/ia+GpcnNosxo5UVEqmjG+nLiNsOatI3HtJj2idcEsQWxrNzaJy93Vs0RfzvLOuA1LyupmkdEVpLFttRd9iJfrOFHD3DMUc/da/lDjcrSCMxzFTShjDmBWSJpTOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMPgyUd5QEQvBBdHSO3AsZMsD2CflnpM83/Jeg+iExCMrmtHnTxlMad0alyDWxEiU8Ja9CKQlY8TsI6Sgfx+TritnNRNUNpanbRBA5piQpUwawgZH/Prfb6w9WZoiiFN4qHr1AgXgzKfvVYggAh2zYxKrOm4GNjZXJtz/8OLwI9o17eUT4w4RllRI9onXBLEFsazc2icvd1bNEX87yzrgNS8rqZpHRFaSxbbUXfYiX6zhRw9wzFHP3Wv9Gg2WvKXcaQoPq8dYvXBDiWQWQEl4HgvFM2bu+WFHT1uZimT2kQX2DC4OEyxUpTD4MlHeUBELwQXm6MfsYWaQcpU/nnc0r0rksrShcjbgOejMV4TVdqFIrQcUkDek10aWvQikJWPE7COkoH8fk64rbmapvu8GTtFeJv0RkVwrWmzod+smLGbBgdVC1tgFiwjjlmsLGCk0KdWIIAIds2MSqzpuBjY2VybVppo2+UjsoY+dEk1VgbrDkUoNgNHZ4w5V7yAeG6jn8jVMz8s7lE/N0JrXE3nd7zlm1F32Il+s4UcPcMxRz91r92OEtofaIWDtvOLjyFka1VlkFkBJeB4LxTNm7vlhR09SiZ8hj5jclm4cMmgMS30D025av4RRNNKF0t3pJwKv8bbesCLgYotUO9treNY1Gz8rHlx5s8YLHMEWsoLROZ2jlYggAh2zYxKrOm4GNjZXJtWmmjb5SOyhj44oIh9mYzmI/n1WAt1gjCXvIB4bqOfyNUzPyzuUT83Si+G04JfRlAVFYclhD8d4dZ5YAumi6YjIYv2006L/0oZ6EhxKrwfCXdZkCex15AMUngnZslNY0/D7DkI+4jM/Jr0IpCVjxOwjpKB/H5OuK25mqb7vBk7RW9w0HqmYWYM+u7zzFRyYwpXvIB4bqOfyNUzPyzuUT83QmtcTed3vOWbUXfYiX6zhRw9wzFHP3WvyKxJWMbtP+K4g6XAIaM8hh0yXRb4WLJTYzFeE1XahSK0HFJA3pNdGlr0IpCVjxOwjpKB/H5OuK25mqb7vBk7RW9w0HqmYWYM2BRqRBAIijhXvIB4bqOfyNUzPyzuUT83QmtcTed3vOWbUXfYiX6zhRw9wzFHP3WvyKxJWMbtP+K4g6XAIaM8hiKXxtxSeI/e4zFeE1XahSK0HFJA3pNdGlr0IpCVjxOwjpKB/H5OuK2TnsJf44REAdUVGGFf1TOxTmXVBfK4hJZU0oYw5gVkiaeuCv8EL5+zqJrcgxNNa6eVFYclhD8d4dZ5YAumi6YjPOWj3e21y7nnPvrzUAkMW0VQYzcy9jpIh1ULW2AWLCOOWawsYKTQp1YggAh2zYxKrOm4GNjZXJtGjM89qAA/CGheTGTzEMSDxULXnWGb3lIe2KKAI0yLWZJ4J2bJTWNP+eSNGl1cCaS4cMmgMS30D025av4RRNNKGvu6TVpIgPAvcNB6pmFmDO23HsUbuuAtV7yAeG6jn8jVMz8s7lE/N0JrXE3nd7zlm1F32Il+s4UcPcMxRz91r+4NYWZC3rCCyS+Rcv2KmnOpGgIylgTbd1ipQ3jNDYXS8IKQH9xapKWNuWr+EUTTSh76HVCkFwS1MKRtQL/KaalkuNUFu+C5a63Nv7ImqW0oJTOxVf6qMnZwWFEse2vnPbaPWCFUspSOtnTBVNxD3DLXxLt6MFIZvhEQj3KOxUlhHHO1gemEq84IIvT+UNORMRZ5YAumi6YjDpOP/sHbWg2WtEXmuBxTQnDpKy+48LpC49onXBLEFsaUzMxN3ZVssA24X1LNvxtz2gLnMoJSJnyHYNbLmfROv8nD1iWiaJSnwldkCFjwDorJ1AqBPke3MEBYNAncoGkg5+gA4ucyggfAOcFxSNMQtsEujim6sxPX3ojKMgrgmb8cV9sX9MGuKJTMzE3dlWywGTF6WjHxqxiHZRXYx8mS6cf3i5JiFZy84LQ04Y/0qyIHYNbLmfROv/BJGktlrWsO1DFSZ18At2ob5a18IBpPj1mAmFR3LKaecIKQH9xapKWm5wIy7VEbo3CHTnGJiwHXcTZrR9MdAnrgzDpmo9++/BeCQMHKUbNsKVqodDodiFlKqLBu3yOMdoAQnJ+BiGA7qKg6ef+jn553ngGDIv8iOAwICxouRz2wyCL0/lDTkTE5qBEytoYnUYkicNNMWhMwGXf8k5ctsyC6bkVwIZBuuLBH6ab6nFM+gGrw5g00TiRwU6UqoOkzCiGv/s16QMD+iRYufMz54BS7dGZTVLjMkd865Y4/YCsNgFg0CdygaSDn6ADi5zKCB+I8Fr57XLiYm5jMyU+AnNu/nLahDZxASg0vdnlEABTMF4JAwcpRs2wpWqh0Oh2IWUqosG7fI4x2raOQZwLKZ7xMA6OixUw6rRBUf+h5bl0QriYA3FRomsprD1oOhUnp8hO7JRb/x7EONmzID3ndQXqo5b2Gfh6SO6ZzxjF9EhfAwDqg32YtJMacV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/wSRpLZa1rDsYpvJFpyu2QscqZyX+NEWS+PLhl1syijoxk8wvrRXYtexjbVPe5ExNn6ADi5zKCB+I8Fr57XLiYjp0B37HjdVtEUl1Jfxf3nwGCB+gdLSrKRFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybdD0jPoHAd0i0PpIV6W3I+BWbq1chxCvXPG7E3QxTiCgdWCm8N7aUUocRy4n5G9LBnPKxSUCjyID2bMgPed1BepwG3LBXMR64fX4OJH6BGbpEFxjJGuPLY+LSRYue6xyQrqZpHRFaSxbbUXfYiX6zhTBTpSqg6TMKMRMPKQaiwwWXOif352RW45OVry/zlmQLp64K/wQvn7OTkGSJu/s69jC4OEyxUpTDyqiwbt8jjHakex5NYkW0nHL3gN/E+8VZtppLLjPaU8vKykLxLUCU+oPsOQj7iMz8mvQikJWPE7CHYNbLmfROv/BJGktlrWsOwpksyvr8aJypRouHe/cyEIGCB+gdLSrKRFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybdD0jPoHAd0iFtoNCfe/cTf1+DiR+gRm6RBcYyRrjy2Pi0kWLnusckK6maR0RWksW21F32Il+s4UwU6UqoOkzCjI7HXAdufalxI26MsU3OoLAiiPL9wuI3BSlJxu09djeYtJFi57rHJCupmkdEVpLFttRd9iJfrOFMFOlKqDpMwoyOx1wHbn2pcSNujLFNzqCwIojy/cLiNwMKJdxWDgWr8wICxouRz2wyCL0/lDTkTE5qBEytoYnUb49sHv18Hvs4Qcor8g32PhNYegUgJZ4PnO2tIEHj2/xDVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3h+agRMraGJ1G+PbB79fB77OEHKK/IN9j4TWHoFICWeD5cDCyOjc4bvZeCQMHKUbNsKVqodDodiFlKqLBu3yOMdrzkgYjmawpSilT+edzSvSuo8ExgfrwoNDkR5TJwQr3X57z2bM2B/fLTkGSJu/s69jC4OEyxUpTDyqiwbt8jjHa85IGI5msKUopU/nnc0r0rqPBMYH68KDQCp4MBTDNz7JmAmFR3LKaecIKQH9xapKWm5wIy7VEbo3MU4UVpv+iFFpoAb+70/qtPBRehIFeP5DBoLT4HQsX6R3bcYOqDhgjKJnyGPmNyWbhwyaAxLfQPZucCMu1RG6NzFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QS05+7CbzaKhxX2xf0wa4olMzMTd2VbLAHYNbLmfROv/BJGktlrWsO+Jv0RkVwrWmWnw//gC8XDqxz7VxwyLzm8lQhwwd/5HsD7DkI+4jM/Jr0IpCVjxOwh2DWy5n0Tr/wSRpLZa1rDvib9EZFcK1plp8P/4AvFw6pqCNPdiDPh3BNg3LDLX2ZQFg0CdygaSDn6ADi5zKCB+I8Fr57XLiYqjekj7PLyzlIdWHn/tImo3XwFxU+jQytot9mDkl+tWoMZPML60V2LXsY21T3uRMTZ+gA4ucyggfiPBa+e1y4mKo3pI+zy8s5SHVh5/7SJqNegl7nWhT+1Xkt3c7HJH3bJTOxVf6qMnZwWFEse2vnPbQ9Iz6BwHdIgGAQX2IpawmpKFk2NHyLDmtduay5T/uc/83YxNodUb3EWsoLROZ2jlYggAh2zYxKrOm4GNjZXJt0PSM+gcB3SIBgEF9iKWsJqShZNjR8iw5rXbmsuU/7nMpa8rPfcFPWKw9aDoVJ6fITuyUW/8exDjZsyA953UF6l0t3pJwKv8bauayXcdn5O75ewgZKQep5HJ8W3W2YQJWdWCm8N7aUUocRy4n5G9LBnPKxSUCjyID2bMgPed1BepdLd6ScCr/G2rmsl3HZ+Tu+XsIGSkHqeTFibXPSil278EfppvqcUz6AavDmDTROJHBTpSqg6TMKMjsdcB259qXEjboyxTc6gua+78znw3ikgYIH6B0tKsptzdiLT7PbX7sY21T3uRMTZ+gA4ucyggfiPBa+e1y4mKo3pI+zy8s5YpE722OMBL4i195SnhsyJJTNm7vlhR09f4yfXr78HOawuDhMsVKUw8qosG7fI4x2vOSBiOZrClKKVP553NK9K7+yGWVnr85YBBcYyRrjy2PmLeeZbuMJ5EcRy4n5G9LBnPKxSUCjyID2bMgPed1BepdLd6ScCr/G+rUwTkaCc0JARLWdPclGxz48uGXWzKKOtStgFeUxC3Ea9CKQlY8TsIdg1suZ9E6/8EkaS2Wtaw7GiMFB2SyS1/sN4y5hqAjrPG7E3QxTiCgdWCm8N7aUUocRy4n5G9LBnPKxSUCjyID2bMgPed1BepsoM5fG8CZ7UcmUejfS7U0c4SNAPWFs2eeuCv8EL5+zk5Bkibv7OvYwuDhMsVKUw8qosG7fI4x2sQzp20SDb8DjmenhxlvRnhqGJn+CLQNDwYIH6B0tKspEWsoLROZ2jlYggAh2zYxKrOm4GNjZXJt0PSM+gcB3SKo5FiHNy2C/kK3RJ5lwuL0c4SNAPWFs2eeuCv8EL5+zk5Bkibv7OvYcdmIiNk4jAj63I2TU/dOmyKkk5GRrj0RE8vBtvg9T9aGp+J6yuY9aCX0ErQyxUNNVjW1fM47WbvRafQqGpk4qbBQFOQvZ3yiVjW1fM47WbtJi8mo3u4XzqNUbehcOlfX6pOtkR5QI7rnkyOhxNuHYvuKiazyQ07CygDEbahTo5m18mOKd8EkIcL8CR+13B7XLlk89pyoh1QKcIdUpPLmJTRs7EO/weafO0+iUPoaTRHN/jys/Hw1bLBQFOQvZ3yiVjW1fM47WbunY+wI9aowrgC6kcQC+v+PygDEbahTo5m18mOKd8EkIcL8CR+13B7XJw9YlomiUp/3eNoOgk516O0bWTRss2SZohz+Pg21Gw+w0zB9aWHlcmHOrclVvQBaPLXN2EDq885+jvPiRLJcaPJ6/nou/PGxVFQf51dFuyer73Isr9tVv8EKigEo1SnubAQcOy7/A7Tyev56LvzxseJv0RkVwrWmih+P8o/iH/miw3Dru/3KHpDAAUFNMy/LJSOpD5+0nMrVWOhARem1g3GYp0zPErq9tFb89eU5ixYCcOf8sCcKkzApoEU4LPB8hByivyDfY+FV+A+aShy2QWuRZTUMPC0ZGhu9DEhD27haaAG/u9P6rcpFAKM9WD4wo6yNCesxp30bNCLazsctMajekj7PLyzlJfqPbVbhADJEHLmJDbWEScHJ0md63CjkNQVM3MMPDzQ3V8WVOYGSZ8wTi0PUtsv/e0ZUpDugKP9t4I1zhKJNEgJWu7877GJiKVP553NK9K4ktiaH4ymtPpDAAUFNMy/LJSOpD5+0nMrVWOhARem1g3GYp0zPErq9tFb89eU5ixYCcOf8sCcKkxo38GtLH1LwqN6SPs8vLOUxB6XM5gvvY/+UZCFbJzU/Gjfwa0sfUvCo3pI+zy8s5f/KIfQMqp/GOd1pjOAzV28aN/BrSx9S8Kjekj7PLyzljNYvwaFo+DXl3YAfgxxM6xo38GtLH1LwqN6SPs8vLOWYXcqqnIjNYinBQ55mE3EBx/9BN7g4CcpdHSO3AsZMsIHXJhT1FXpFzMVeOF5AAi1ny4xNyhR4rNVR5Rj0dqq/OV2xrpK/nDrsY21T3uRMTZxqJIHSnBRTlvEgkQyUjhvRoNlryl3GkKD6vHWL1wQ4jFH6xbEADBZD7yxSCyuYmNVY6EBF6bWDcZinTM8Sur0w0mP3skyStFRWHJYQ/HeHQW6A1k/HcyPI7HXAdufal4KLY1BA6bZNt/AppCGSgkCuq5RgVyJXFSJPUwU+QGUkT80g3hJAfBjuIY+Fii8a7liCACHbNjEq8kyiJFHAjB14eK2+BZCIEsCTsqSLk1SmXslGlDKq0rZw3LSn03UDPvXzClMVnPUWsJcLQ3VyEwFFy1NiCVwoZNhBgqonNW5qa9CKQlY8TsIr5MLZhS3k9kPvduJuB2FTTQbM7YMtlDbiDpcAhozyGMeVdu0BwjeR/e33G6k5A2eOZSgChCE4twePxLG2o3WY1NJEJFqXK1rhwyaAxLfQPRSI6dQzrfsn2Hdq+FKLGKzZ0wVTcQ9wy18S7ejBSGb4G9N4biOT1vadGlESu52O3uJZYkEegKlijmUoAoQhOLcHj8SxtqN1mNTSRCRalyta4cMmgMS30D0UiOnUM637J6URBhW0GSXt0e+vGXgoG48k4Feq0u3fy6+HjxaB4B74rR508ZTGndEiMvY6Q2mATs6MQApuBRE7MFN9ua4dqTc44KuW0tEdOm1F32Il+s4UpyenXn87dN0N0mWZqCU3HxQjWoieQyMsVtfM3gqBsEzA9XGWsKHPdJ0aURK7nY7e4lliQR6AqWKOZSgChCE4twePxLG2o3WY1NJEJFqXK1rhwyaAxLfQPRSI6dQzrfsnpREGFbQZJe3Q+khXpbcj4Lv8Ik5kGtKer6XAk0olsDge0pn32vN1miXoFeEwmnw1FXNBKZaZmVIcRy4n5G9LBoVVIPUUpxe0xvZrfAFJ45yR7Hk1iRbSccveA38T7xVmQrzB1j/N0PEEAcndc3eVqrCXC0N1chMBRctTYglcKGTYQYKqJzVuamvQikJWPE7CK+TC2YUt5PY4ikiSAZSiTl0t3pJwKv8bauayXcdn5O4QflWiQVdxCEl9XmGeaAZNQ+8sUgsrmJjVWOhARem1g3GYp0zPErq9MNJj97JMkrRUVhyWEPx3h0FugNZPx3MjwSRpLZa1rDvib9EZFcK1plp8P/4AvFw6/ZQRZKzLOf+vh48WgeAe+K0edPGUxp3RIjL2OkNpgE7OjEAKbgUROzBTfbmuHak3OOCrltLRHTptRd9iJfrOFKcnp15/O3TdzFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QNYOnexOTNWJjr71WCqHSa2fLjE3KFHis1VHlGPR2qr85XbGukr+cOuxjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3cjsdcB259qXEjboyxTc6guruDnuKlgiySAvZetnnrzMzc2icvd1bNHavFdz3pmbF7CXC0N1chMBRctTYglcKGTYQYKqJzVuamvQikJWPE7CK+TC2YUt5PY4ikiSAZSiTl0t3pJwKv8b6tTBORoJzQkbGoFqhta0ZnL55H3lE1PUsJcLQ3VyEwFFy1NiCVwoZNhBgqonNW5qa9CKQlY8TsJeK7lRBXwUQ3h4rb4FkIgSEjboyxTc6guwT8X/oXxNlaw9aDoVJ6fI6m3ZnKEGKjwe0pn32vN1miXoFeEwmnw1FXNBKZaZmVIcRy4n5G9LBoVVIPUUpxe06aoy1WiNitY4Zk4WCpxifqKg6ef+jn55haKKk2mq+JbNzaJy93Vs0dq8V3PemZsXsJcLQ3VyEwFFy1NiCVwoZNhBgqonNW5qa9CKQlY8TsIr5MLZhS3k9nDHjp3AnvIdFCNaiJ5DIyxW18zeCoGwTMD1cZawoc90nRpRErudjt7iWWJBHoCpYo5lKAKEITi3B4/EsbajdZjU0kQkWpcrWuHDJoDEt9A9FIjp1DOt+ye0f2eHNSWQfvThJyXFBSaVZMUPkuV6iZFUQxceJ6Vh5ZTOxVf6qMnZI4vTKyHBGc8iT1MFPkBlJE/NIN4SQHwY7iGPhYovGu5YggAh2zYxKvJMoiRRwIwdeHitvgWQiBLgx/liKPdavMpTUhlIxK14Enga0CwyceEiT1MFPkBlJE/NIN4SQHwYQEECCmIQDytr0IpCVjxOwivkwtmFLeT2uVDOITUIvshcCRC82HZbeUtK5BBW2zMUBAHJ3XN3laqwlwtDdXITAUXLU2IJXChkXkpPsZ+dnSHC4OEyxUpTD+dK/+s2YPEJZax0spYeFH138AitcHVEIfJuIsHCp9sTzc2icvd1bNHavFdz3pmbF7CXC0N1chMBRctTYglcKGReSk+xn52dIcLg4TLFSlMPK+TC2YUt5PanboegnGsd/mhmECt9KzkIfobjCkrKLXpYggAh2zYxKvJMoiRRwIwdhAslpYUxBtsh3lUHYet7OFTM/LO5RPzdgcZdMvisFLttRd9iJfrOFPOqxRniGbE2BXZXUrs81rD67pZhSX17SNEMoXwrc0LWwgpAf3FqkpYUiOnUM637J0eCyXGTMbc/PwGopGN5FQ5/rmlOCs+pkTGTzC+tFdi17GNtU97kTE2caiSB0pwUU0ibB9nx8EYwCrUNkWofJ48tji7xe9XGUHVgpvDe2lFKHEcuJ+RvSwaFVSD1FKcXtMf/QTe4OAnKqORYhzctgv75kLyfxrYOaq+HjxaB4B74AavDmDTROJHbA8chY5Tt3Ign5UWLR4Y6NDt7WTzRCmeLSRYue6xyQoHGXTL4rBS7bUXfYiX6zhTbA8chY5Tt3Ign5UWLR4Y6MdwO7xcwqNuLSRYue6xyQoHGXTL4rBS7bUXfYiX6zhRvsIoaBB34idsqKEd60d2xYwX1aLMrZuMPsOQj7iMz8mvQikJWPE7CK+TC2YUt5Pb9rNQ9pMjFpzHcDu8XMKjbi0kWLnusckK6maR0RWksW21F32Il+s4UXv9yBR+/ijDTgI+gsDxqVTA7z0L52nuKAh7GJdVdRXcRgZf3KU7i+Xe5+Pg0gAw6gkXTrB5PTrHmnWkGLugJ85dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmaR5kMQ01CIuNBOIwVCPkWKOrWInZKBWSl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZPJbAL9tHLEGWHX6YEdj0Tnrgr/BC+fs6yXzekylNbvuME3AWcNJDTFzIuTzuQM1ZUVB/nV0W7Jxo+Ct+I0vS1KgE7/Wg2oF9HK1m18oZigrf/TaIogyMjIs0vThxS1XzH7B0bn4S9DqtEi4/dVHuv1ZmiKIU3ioc4fQPNOuC0intU2Igm5/G4lM7FV/qoydkji9MrIcEZz0J4x/ZkPUEhrh9/sx4J4Zfy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNsAfu4fjqbOnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTiqYUd+1+I9sNsLj8+1LArYp2Esb2xo32WR5b28YUL+LQBh6HFoi6KbpBVE/12+GrTlQmC8P+3GDyeFxINQuuL5u0JJVmBOW7l2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZw9wzFHP3Wv5Q43K0gjMcxFKnq6h8DmkfuoJ7of2Zweb/gSNtnTmQLz/8OLwI9o17Y4QQJqbO87tTp7U2MqFK2kg1GqmGzqDZamgl93Gvh5nNRNUNpanbRbal1u1efLIS9plC+cyyDYQf4Yh9NJGhzEnA+qtoY84NdHSO3AsZMsIIKjfLl3ZbED/XfrYjohNzYWjo6O8Jhu3D3DMUc/da/0aDZa8pdxpCg+rx1i9cEOEXb67T6dm4QXm6MfsYWaQcpU/nnc0r0rgiJpNbV7ZkHcPcMxRz91r/RoNlryl3GkKD6vHWL1wQ4rRZfsWcdGPFebox+xhZpBylT+edzSvSuTqWbBXWJIWxw9wzFHP3Wv9Gg2WvKXcaQoPq8dYvXBDiV7rIXypR8MF5ujH7GFmkHKVP553NK9K6CKtHVZIlUm3D3DMUc/da/0aDZa8pdxpCg+rx1i9cEOFIzKO1ujFZYXm6MfsYWaQcpU/nnc0r0rj8UyvNSeFV+cPcMxRz91r92OEtofaIWDtvOLjyFka1VRdvrtPp2bhDC1/fCupsoFA9aq6MBhUYU9UMyDf3LSmlw9wzFHP3Wv3Y4S2h9ohYO284uPIWRrVWtFl+xZx0Y8cLX98K6mygUD1qrowGFRhQjfjxbQlFzMnD3DMUc/da/djhLaH2iFg7bzi48hZGtVZXushfKlHwwwtf3wrqbKBQPWqujAYVGFFhQAKZZMa31cPcMxRz91r92OEtofaIWDtvOLjyFka1VUjMo7W6MVljC1/fCupsoFA9aq6MBhUYUAcdlHw6AJJxw9wzFHP3WvyKxJWMbtP+K4g6XAIaM8hh7HeNG+/pX0eZqm+7wZO0VvcNB6pmFmDMAPSxBKWuLGVqaCX3ca+Hm5mqb7vBk7RW9w0HqmYWYMxjo7G2zTl3RZQL/oMAG4rIisSVjG7T/iuIOlwCGjPIYXRiYuK/YXftw9wzFHP3WvyKxJWMbtP+K4g6XAIaM8hifbR3T5TM1fuZqm+7wZO0VvcNB6pmFmDPszcMp6FdHelqaCX3ca+Hm5mqb7vBk7RW9w0HqmYWYM7bcexRu64C1ZQL/oMAG4rIisSVjG7T/iuIOlwCGjPIYu9izdxs229Vw9wzFHP3Wvxj+FmzHJW3ZXslGlDKq0rYQ5jOphMVE0JKo6qB5+p5fLDw1gsxVpXifsyT7eXUhjb/gSNtnTmQLGjM89qAA/CGheTGTzEMSDxULXnWGb3lIP43hjlhA7a5r7uk1aSIDwL3DQeqZhZgzwb8M+BjJYjxamgl93Gvh5k57CX+OERAHVFRhhX9UzsU5l1QXyuISWaFj858ehtyw85aPd7bXLuec++vNQCQxbVcXFEpHJjI8EnA+qtoY84MB0rdEwIGjwTToHlm2V76QdwrrbERPHvmjaT1pKeBddU0GzO2DLZQ24g6XAIaM8hi72LN3Gzbb1XD3DMUc/da/uDWFmQt6wgskvkXL9ippzsFMGP+lkylBFsGuEV+tOYXZ0wVTcQ9wy18S7ejBSGb4OMX4bxb2E4Nw9wzFHP3Wv7g1hZkLesILJL5Fy/Yqac6D3IXdjMVoXhbBrhFfrTmF2dMFU3EPcMtfEu3owUhm+HthVJtZqBcVcPcMxRz91r+4NYWZC3rCCyS+Rcv2KmnOBgIQovxrrHoWwa4RX605hdnTBVNxD3DLXxLt6MFIZviULlnJ8sZq83D3DMUc/da/uDWFmQt6wgskvkXL9ippznFPDK6sKqVmFsGuEV+tOYXZ0wVTcQ9wy18S7ejBSGb4zLJsoAVoLpoZgbHqdcpCwycPWJaJolKfCV2QIWPAOiv2rx8kyeqwrYEaJL2thns32bMgPed1BerO1vv0WSUjnN096ji5zwFdxGPe4bucB96aMf1rE3LnacEkaS2Wtaw7UMVJnXwC3ajHEXkGqj0LkTndaYzgM1dvCLCTAKodqtUkicNNMWhMwGXf8k5ctsyCEpUeUcyxK2rp/R9h5DelodD0jPoHAd0i0e+vGXgoG4/5bcPIy81zPTNifuT+9HiUDdJlmaglNx8UI1qInkMjLFbXzN4KgbBMn3U1q5CRms3RbTL2mz8el07gS1r63R5Dhr/7NekDA/okWLnzM+eAUu3RmU1S4zJHa5FlNQw8LRmIW1OMeqk9JA3SZZmoJTcfFCNaiJ5DIyxW18zeCoGwTFKYFNfUmR3VD+tV1YrzprXQ9Iz6BwHdIvThJyXFBSaVZMUPkuV6iZEpTZ/GXPlL4+XdgB+DHEzrCLCTAKodqtUA5wXFI0xC2wS6OKbqzE9feiMoyCuCZvwJf95veuyARMEkaS2Wtaw7GKbyRacrtkKWD2l6Al3TxAJw5/ywJwqTCLCTAKodqtVEYxRziOLSXPiY6kXZLM45xGPe4bucB96aMf1rE3LnacEkaS2Wtaw7GKbyRacrtkJEvwRMaTUJvVSrUnJRST3i2bMgPed1BepwG3LBXMR64YHgfTkjpAjIf5ZqjnBY+ivXqX1BcT19flLmp3lPgRYv8EsjfGHwQ4UZxHiQkh1RvanpXNyAmjLPLyMqEjuETCkGrW3fky6+pWgxwPOa+bCZ74UOEKx29rSoTXC84ul14Z7+ehYbqhzmWkbI1I1Mu6vPDah99te57dmzID3ndQXqOS2bMRXLafiImZoORXXgsf8C2SZVmDNdHQRRoJw/+2KoTXC84ul14Z7+ehYbqhzmibs4d/4+CUrBydJnetwo5NmzID3ndQXqOS2bMRXLafiImZoORXXgsTNifuT+9HiUzFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QqfGpLh8RcwMCcOf8sCcKkwiwkwCqHarV+PbB79fB77OEHKK/IN9j4TWHoFICWeD5UHLSet2GzjeiAvTc3UWxu4jwWvntcuJiqN6SPs8vLOUh1Yef+0iajQ3LW5cIdQCfOd1pjOAzV28IsJMAqh2q1fj2we/Xwe+zhByivyDfY+Gwfo+h/zyUvFBy0nrdhs43Qy8gpr1ISwCI8Fr57XLiYqjekj7PLyzlIdWHn/tImo2cUbIJ9ys9Q26ZmKiPu09v+PbB79fB77OEHKK/IN9j4TK4kLrElPLVDAko/mYmeUU0fsXS7rLoRNepfUFxPX1+85IGI5msKUopU/nnc0r0rqPBMYH68KDQlWJnz9w9Q/f/lGQhWyc1PwiwkwCqHarV+PbB79fB77OEHKK/IN9j4funjUNO/1cljnsh4VZhZLFYguOSuVUdG07gS1r63R5DyOx1wHbn2pcSNujLFNzqC1eag1PUkG54Drn8EXq+wzfBydJnetwo5NmzID3ndQXqXS3eknAq/xtq5rJdx2fk7s+54arRnuKX5hp1Z5nFx6IEWaoAMA0T8gGAQX2IpawmpKFk2NHyLDmjtxhuLD/JGORaK+jVTVinA+mvjg8B7HHBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDqK+J6TvRaiS8ZVeGkwOQRWTuBLWvrdHkPI7HXAdufalxI26MsU3OoL68EzLdZBncHwXT4A2AnSw/OjOFmORVMKwSRpLZa1rDvib9EZFcK1plp8P/4AvFw6TAHKhhX0wKCYYhw+sxYl1U7gS1r63R5DyOx1wHbn2pcSNujLFNzqCxjxHcXQS7GBmBtactbH9s7BJGktlrWsO+Jv0RkVwrWmWnw//gC8XDpqp+dU65i0NUxe50z1V+NAAy0e5wgwXMeI8Fr57XLiYqjekj7PLyzlIdWHn/tImo3AMozU4es7PGgGynhwCG/dmjH9axNy52nBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDo/lLhk/ggMrjcgfXEg9tLEHQRRoJw/+2LMU4UVpv+iFFpoAb+70/qtPBRehIFeP5DXD3ogJOY4CX+Wao5wWPor16l9QXE9fX7zkgYjmawpSilT+edzSvSuo8ExgfrwoNCTgGroNfcMyW6ZmKiPu09v+PbB79fB77OEHKK/IN9j4Uctn+VEzmHLaDHA85r5sJnvhQ4QrHb2tMxThRWm/6IUWmgBv7vT+q31WfcG33pX/WuRZTUMPC0ZiFtTjHqpPSTMU4UVpv+iFFpoAb+70/qt9Vn3Bt96V/3/AtkmVZgzXR0EUaCcP/tizFOFFab/ohRaaAG/u9P6rfVZ9wbfelf9icBM2G+IVyGG7IQi1d1TJcxThRWm/6IUWmgBv7vT+q31WfcG33pX/TkUV1TzDakf8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWXtiCIHQOiIcf92dte6LcbG51dzHHv8Pdn8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTT0qKIjqzbVXZaLveUM2A9tkkI3fuV6YyMpwzPoRrUBT+Q5PGEIXMOHf+zZLf8Byc20UfxrAW9Z5oMcDzmvmwmeQ7B9SHnHTb2dV1iQFiJw/ZdRQqYcqcO9i0SXWMoC19waFJ//MVAarvJsseUX7QBpF/KGBLAuOctnmc0Gr44Jfa1Zni5uVvKw6OyG6bnoLJL7n3mFDlx+KMyy9ofvlbCVlMoCCcErT30372ExX2DzxP5DKhKevgqTMG/erWsTnq8/TnSPPDjO4B/WwMvpibSvrulmFJfXtIi5hjbLWrggWPkgBJUwhBsncmN6aMbQ2MT1nZXCU9vI39FHc1iKADHCY9EvBAEIvmPjF9L//hay2oNfGWRcbK3xUEU0INUM9Q5WOgwK0Z78M/AaikY3kVDvBdPgDYCdLDpwtxCu/hW/x7roE+YpEbxS1CIIGS1geuFEB+jvEgReE1epxaUq4HuJ7JkW377qQR3PQklR7DhT5fqZrPwx/xXADJtPfo94m8PwGopGN5FQ5TPAJSXOY2s6cLcQrv4Vv8TFc+ZFbYaF/kJbkeFXcf5BMx80za+64H/xzTeVt3aPdLEFGrHS4RpNCE00JDV6wsTuBLWvrdHkPIAIyXWxsyLm8Oxz8TxEynUHLSet2GzjdLEFGrHS4RpNU9GlAiXdw0TuBLWvrdHkPIAIyXWxsyLm8Oxz8TxEynfBhpIwv57iKXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZmLGnFFoQhegCCluMxN3mEGNGYX60UQYBlKUJySrmw1K14XBKVwYCguyJ1lgfqDrBwX94OU4e/c4Jw9YlomiUp8JXZAhY8A6K/Hq5bfbk4rSbPz/c6/JJ/0MIhaGFMINVqKg6ef+jn55Da6ygPY6P1OOnHt02tNEKxI26MsU3OoLwH2wOq/fkXNsclhcoUcxl6Kg6ef+jn55tZxbj4yjxprBJGktlrWsO1DFSZ18At2oSu3dJh+2uVHS3x7mk9U6EzAOjosVMOq0QVH/oeW5dELDcD+9R55FOGz8/3OvySf9QDmp5qMwprkwDo6LFTDqtEFR/6HluXRCCjbg08w1myqJ8kfQ6OJ29hQjWoieQyMsVtfM3gqBsEz/zuT3TJ9/u/ThJyXFBSaVZMUPkuV6iZFts67pJvAzdKnpXNyAmjLPbmMzJT4Cc27+ctqENnEBKBog9ZIDYXsTcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJP0e81vVW9ueNK3XnZ6aCuj/FQNkXvsMHapwriAGCcPo4FEKVQ4QRJV8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9kbOaaK9y6QkotDm2SkoC7mOyBttLSJ8lhTO/1HjlsfWmWsdLKWHhR9uYIrU+CZte1y5IhhzLqwUwV2V1K7PNawh/iCN3JOYzFwY1qZHZMRiB/QlkiN+pvxHVlyws4S8Ogabgj936CNHj8BqKRjeRUOYcajpA7YTTJTPnMuafyLILZ1IJx1aJgMzgsFth785LLk434FxrlvywVKXuPBvFInoOMOuKvU1GdZVoBpsL9UIp6qxLjRfEbxRRd3vfRmFATpJCqVn8khqrcsyY3m+q2rsJcLQ3VyEwFFy1NiCVwoZGCMihUaWmCYPfBeph9ewq379D1fVRwVwHNRNUNpanbRlE0THxm4EUDRoNlryl3GkKD6vHWL1wQ4hZCi6HuH59VlDaSwVAFb+6g18ZZFxsrfc1E1Q2lqdtELInudpCvlYqwllGw4+2H74V5ngPiPCPRRhkt8ygaKBHPpFBtQkSMfqcJVNzczxRKoNfGWRcbK3z7/yAYt6T2aeHz/QmRw5TYYa77f8vmAHd40NK133aiQD8bmdyp4oyTDkZ7J29H4sKP2hmw1RuLwxzqio0ZomnfAWCwd+65pMBmheAcEXp3d8r23N3wowkx+frLrvXinB2WRAxiszVICGGu+3/L5gB0QrhvVTDYoK4Qcor8g32PhWAQtwjZy4eUuOo/ZGolPU4Qcor8g32PhEP5I66euI4tudwpRJStzjw/qKq6oXwI9cij4eRVyAumEHKK/IN9j4ZeXVQaR/+/mBH5d5Nb5sfn3gA+/forxpujJU5N1wcZpJqSHugx1dPEj8G3eo7Q9Chhrvt/y+YAdJqWbEMG9PrK6WFEGdh5P7HhjxeqVii0rL7n3mFDlx+KboR8KKvMtE6xlrn6QXuemiccdViuS2KDAWCwd+65pMEiy5SHYswRMpVSOVPa+hxq0//yLJZNFE8BYLB37rmkwbEegyaglFcrS+DkO8fYpMdDPkCN5inJnRpo1VzgallqqDBY2SeSwS7/dvNaKAYw2T1nZXCU9vI39FHc1iKADHCZty4Gc+RblZOkwYzLjVEvtYLZH0C1lWhhrvt/y+YAdlXeHI7I2QVs9UeFmpYZozIXISCx2JoVzQH1USW7XdDdeI2hxaq/IasBYLB37rmkwSLLlIdizBExC2906JuabGs1F4WizKZmEwFgsHfuuaTDc9CSVHsOFPiKcIW0S4ke4OCuvmV197yxjkZpwmQhR3CNlpIV43hTC6lLszuAb+/3AWCwd+65pMI37qMTokd4L8/U06gnCF+plrHSylh4UfbmCK1PgmbXtRhdXxtZM3mDAWCwd+65pMNz0JJUew4U+uiQpG6ujY5uFyEgsdiaFc0B9VElu13Q372G4nAulXUcYa77f8vmAHSB6N9AruewH3hw/17fmDLfAWCwd+65pMM//Di8CPaNefHWjXjdtXbu9plC+cyyDYYndsK8141KEqDXxlkXGyt+DJR3lARC8EF5ujH7GFmkHKVP553NK9K6yaI1w6RUvUF5ujH7GFmkHKVP553NK9K5SO5Pj113PdMBYLB37rmkwcPcMxRz91r92OEtofaIWDtvOLjyFka1VJm3LgZz5FuV2OEtofaIWDtvOLjyFka1V8jHUuAsZ7HHAWCwd+65pMCqfI5t3Vcm+tkCA4GEI6PiEHKK/IN9j4RHzPb5732p1wJOypIuTVKZeyUaUMqrStvDc+JKlN8rLGGu+3/L5gB27y7P5cV3PtgzCwsjkVgCQqN6SPs8vLOWelHy5kyLF2JKo6qB5+p5fLDw1gsxVpXifsyT7eXUhjfIx1LgLGexxwFgsHfuuaTA/R/HXsY5vTeU5rurrnWxlJwTt36MkGCLl5Q+Fxn3tJ9nTBVNxD3DLXxLt6MFIZvjuuVyPS98a+8BYLB37rmkwJGTiO4QTk9YF/eDlOHv3OMBYLB37rmkw8/TVDKwR8YQk4Feq0u3fy8omqXrMYYjkztb79FklI5zdPeo4uc8BXfIx1LgLGexxwFgsHfuuaTDGNJ2E3BZ7kqrSNGlab0YqnQd8okuZsQmOnHt02tNEK25jMyU+AnNu/nLahDZxASgeRraBm+NxYag18ZZFxsrfsYlB5QV0/PCKzno9CbS6ZXA60ZrmXWm09aoR2gafujfAWCwd+65pMNmzID3ndQXqfpRLPm1xe9x7goybPfp5F1Lmp3lPgRYv8EsjfGHwQ4UP3RgCupB5GMBYLB37rmkw2JrEizVvnU2e/noWG6oc5pEIU61qlpNhqE1wvOLpdeGe/noWG6oc5rXLNo6q0aQFGGu+3/L5gB3moETK2hidRqjekj7PLyzlIdWHn/tImo2AFp01VCBqdanpXNyAmjLPqN6SPs8vLOUh1Yef+0iajdMr+bwGkQLzv9281ooBjDbTfvYTFfYPPM0hhN5Hi/ZjauayXcdn5O5Zb/h0F1jGIiVgifm0v68T85IGI5msKUopU/nnc0r0rqPBMYH68KDQSs/OJpfR7FK/3bzWigGMNtN+9hMV9g88zSGE3keL9mNq5rJdx2fk7iKxTx/x1+pBnUDnH/Z9p7BdLd6ScCr/G2rmsl3HZ+TuA3vtrwnv1wFudwpRJStzj2LuZjFfRZ6k6aD6fpe+v7CEHKK/IN9j4SoQc0pwkOGbXNJuUrHz0jzBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDrg8MxZ7cKwom53ClElK3OPYu5mMV9FnqTpoPp+l76/sIQcor8g32PhTnxwVNaDwL6p6VzcgJoyz6jekj7PLyzlikTvbY4wEvgCXevWbRfP072rBUoGQrMwZQ2ksFQBW/uRAexMN6ip3oxXewkyAg4wWRqf3NAPJQY5ZkjAZ4zkc9KYxRqvtbJh24vKAAoVQKao3pI+zy8s5f4vCzo7OmVVO/PlKCabzkU98F6mH17CrUTe3KALTTmkK4sj6dWoY4ZRx8k0NEWRjFCCcmaBVJKeJGWEAM+2tg9GmjVXOBqWWqfhlhZiQhmejgciMNIBQ7dN9HZDM4oFzZiq+gKZgdxdVE7wPsYqY/FKefk00o3M3WTpMGMy41RLUn5U1efqLMFlAv+gwAbismTpMGMy41RLf2OhbxKR9MsbfKdF9AnQ9lM+cy5p/Isg1yWChz5Wi46rnLKW4/Y621M+cy5p/Isg1yWChz5Wi46zpuBjY2VybbzR89UNRM5NlKbPj9+iHGkSV4srYgD9OpoknK+VQWdeRKf2+Y4zEZhs/P9zr8kn/aI9EAkCE4Ye91QBIb/AHapyKPh5FXIC6YQcor8g32PhXVOFvdGwRWAlX26L3zEegzDCDFQmIOwZqDXxlkXGyt/I7HXAdufal4KLY1BA6bZNZJICK8Y3x500nN0fx0OZ3WS/vNeMNayWL8TLnOCOek606ysuXeyLqrZ3Gf53ZAxHFQtedYZveUiCnzLOGTzsjiVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3057CX+OERAHVFRhhX9UzsWQBAlbjgszgl8bfd3tzkA4UQlm3kjqGg3mJGcwwwWk+wOmtfJ0DasJjdqez8K2Jjg5XH+13tvMxO+GSEmE4yxfrk4jl4Pq8hgETOWt0KBunPk7xzX9fu4goVAu7SfhPtbj4pgeTCL138McM+486ro2QmYYXfngN8oBF5x/e4AMjdCV7yFXiMmkyaMHFiW8g4zkXWvrW8eZ8au57+H51PXiWh+Ir3l0H4jcVMA06ZdvmF5SPkMfiTL99wRyp4eWjoqIJ+VFi0eGOpCGwyPdZ4tcXe8xLkcBDI3gx/liKPdavBQCZy5IKBAj/Z8wu79Zx3dHOVhkZTSo+r/C0CFEbDEncGNamR2TEYgMHZNkdaymPWUKiXmsnCgJQIUQutbmvtBAfVRJbtd0Nx7Smffa83WaJegV4TCafDV+8wZPt7z+wH/n8icgRp5DZax0spYeFH17roE+YpEbxQAEJIX02sNFTfR2QzOKBc2YqvoCmYHcXSJPUwU+QGUkT80g3hJAfBhAYBhMVsCNOHAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTk5tHNIzRxCzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR48BR4cfHsJrm63jaaqNovEtWoZ7GLFEjzokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRySfIcbFARtTalhVaSdINj+T8bwxL0+cokgbbO59b0/WuHLjVt4S72X9yZ5m3LYOxnSW7iwRLiwVVPkJK4xKvxsAYGsMjn6WTZ/wLZJlWYM13z8VLsZp+K1hfzVCER8IC8v9281ooBjDbFgJrZJIg0xre89BhN90ZAAJxQckar1N6a4B0zYio8JEbVSH2QGsTiJqWbEMG9PrK6WFEGdh5P7HhjxeqVii0r0oMS3RldC8LQNO+VCg0OpRp5IRzli53Xv9281ooBjDZsR6DJqCUVytL4OQ7x9ikx0M+QI3mKcmeIxKUD+YXwlXcmN6aMbQ2MT1nZXCU9vI39FHc1iKADHCZty4Gc+RblDB2TZHWspj1TPAJSXOY2s5V3hyOyNkFbPVHhZqWGaMyFyEgsdiaFcxzWEKD2PpNXv9281ooBjDaN+6jE6JHeCw//2FO4hHrZ3j/2W3Zfci88UrTlyyOsfL/5cgVXFR2tYX0HiBSNyGLUjJvBEBrO8y9flAtC7R090PufJx7egIZg1MtGwBlMyLZZzmiwPIDz/Qz5Qa/K3RmVhqsillAnUkLQhhfkIQJ624FvBU8HXOF8r2bXyX8exdD0jPoHAd0iqORYhzctgv5Ct0SeZcLi9FM8AlJc5jazNj5CGR19aTlLSJUhbBPaWtmzID3ndQXqiCflRYtHhjqaILl5KLQ9RnwYaSML+e4il2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGY1ydMezGn0OINFfR0AhOV367gLJ+CTSRXQ57pjagUkkdSMm8EQGs7zs/IT2ZPQHhnxiaFR/tfzL9OZgk+wyD5DTFc+ZFbYaF9G/RZgc5jNm2Z2JKG1Ab8BWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFl08nQc4jWEmxEWirsvf/0zOLt7Yp1VWFUIJjubSHeqZ2fPFJUI4vifHy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2Jse6E5dN5oURBBMqGQIwKAyj+ihftNPNpri6ANeDp84/5ON+Bca5b8v9FHc1iKADHCE2/WqAu5XREiBKXmipad4FdldSuzzWsAY3NfbQXckUtP0pDeluf0YTN37P7AYMo9AYj6W7Itm6TmhUq/u91EUvQ0Ibh4iZvuTjfgXGuW/LQkP1FgSCfe/DFR0jIQgdxMQzp20SDb8D3rwQ4EgH2Homh0qIRSq++lJTuU3JkJFIUbU2r04p2Km5gitT4Jm17Y76QwT80CFfFjQQ2ZXZpMa2Wc5osDyA8wCCdGm07ksPFXX9LD/Bi69SpEv0kiDL7x/QlkiN+pvxB/c5jI49Xd+4ugDXg6fOP8gAjJdbGzIuB46OGl9UjUghNv1qgLuV0cFtbmSFg2wqUz5zLmn8iyBEN8vP0viDygvVMR6t5LImmOQCVyLExfmcDpwBd7YCYn4VAc3Gw6WPy/BJV9UtiInOm8J0daJArEB9VElu13Q3LNAKhBsU0yvu4I7AKSoyZajkWIc3LYL+1GLtMtfemLua/sbTdmm9xUmHqaw2YBBL4Mf5Yij3WryxJ/zTbrmU9LT9KQ3pbn9GA0RlPktigXsAxRL+EobTHk5oVKv7vdRFL0NCG4eImb7IAIyXWxsyLmsAXV4TO5kHu+CC4E3dooPjMCCJDBx2Wyj9qJndmR6SkIbDI91ni1wVdf0sP8GLr3nOzk9EhQmWxKIrZ0cOdru4ugDXg6fOP+TjfgXGuW/LlYarIpZQJ1JOaFSr+73URS9DQhuHiJm+DB2TZHWspj2yKpeMOS2Hre7gjsApKjJlGHO+d2kpQcwzuQobZ8qHRygqZVyAs0jFdGXt2euF0xZ9CajtNeobhTUqggyLD3Y9D8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDAqplN3cVEzU/AaikY3kVDt4Mvp02gP+vFjQQ2ZXZpMa80cUcUuQRFgAIENq7GEAzcHxRN4xA7uuqCw5z8R7caan7NglYj85b2RvGzODhFquZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4tAYj6W7Itm6YOS3/iuq/EPm6n85lBOtf+7qdMFrMieHXh44Eru+G2/DFdE/EjAVqOxz/UmTPfDTPmAsMHb7AOoTGOzkkr8idl2C69wHVd1PPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuvnSlOlW8OGOQKtQ2Rah8nj6N0AVPk9YbPYAcQM8A6dejxQzZkyNkLl+F939GPE/8icBFNMgailO2rZzksX6182328zjnKGYrICrUNkWofJ48C5UN1XAKxCA/IYWiIqjyhXlB9PcWZIklyA8lDag+GgxIgSl5oqWneBXZXUrs81rDrVedGrotX28MVHSMhCB3Ey2sfGRJ5U5hZv4+itd+NICxFxpn4DsyzhLlHFSBJRsW0PhT6PCGD/Ygn5UWLR4Y6usYanHoofj0nenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvsgAjJdbGzIuLB9UQNbsTwq0/SkN6W5/RkU+G0HYj8smWUxf0x6bokll5iu8XGxV40zXsVSeB4wBmRpCIh+h4iuo5FiHNy2C/j/pKbRms9PqD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDwW1uZIWDbCqIJ+VFi0eGOuDhEHI21dy0uLoA14Onzj9iy0p0pBKJy9dzQNyGLarrpH+iYXN2p5bgUVVy1alyn3FelMlJmN9AwJOypIuTVKZeyUaUMqrStp4qm8TJ5PDQQZl+0QKwT4iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUid06uLbciJmlRUYYV/VM7FkAQJW44LM4KEupzfsB0UvhY0ENmV2aTGqQbOd+pLH44ACBDauxhAM3B8UTeMQO7rqgsOc/Ee3GkMp+iHD/Ja4dA83omXDZzLn7Mk+3l1IY0yt8V/NMhP4JljO7IO5vaSLad8u35k2XXFUlVUTWKaM6hDsuOwxl0dYdN2pxK1+dCc++vNQCQxbeOaIADZIsHLwxUdIyEIHcTLax8ZEnlTmEN31FYMp4zFLEXGmfgOzLOEuUcVIElGxbQ+FPo8IYP9S6QSDAWWgag06B5Ztle+kFtTAVlKRRsBbHL4xeW2cKkpUXp5yCcn5nSDCgXY/oNQu2TXWro5hPL6EvIt0EqAX7Z3Gf53ZAxHFQtedYZveUgomSlT17GGkGAHEDPAOnXo8UM2ZMjZC5fAbWV8y0btFXARTTIGopTtq2c5LF+tfNvehJoGpiOY5CKxJWMbtP+K4g6XAIaM8hjWob9UV7T7YSd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+5mqb7vBk7RW9w0HqmYWYM0trmsNOkbajHJ7TLaX4iiLm6n85lBOtf97Qrs+EB8Q1AAgQ2rsYQDNwfFE3jEDu66oLDnPxHtxpFBfeuvmDgd54XgLSZRtKdQ/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8EmZGuEoHlf2yooR3rR3bHY3vUVTnX3mObqfzmUE61/DZ47GUbdnKIACBDauxhAM3B8UTeMQO7rqgsOc/Ee3GkUF966+YOB3j/pKbRms9PqD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDwSZka4SgeV+VhqsillAnUmDkt/4rqvxD5up/OZQTrX8go2OQ5IRqTgAIENq7GEAzcHxRN4xA7uuqCw5z8R7caa0dVe7iTaogHwvZ3bgc7cmAvOCwHeTjbQ/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8FtbmSFg2wqUz5zLmn8iyBG4hg2iglMPxye0y2l+Ioi5up/OZQTrX9Bze3Pj1d4bAAIENq7GEAzcHxRN4xA7uuqCw5z8R7caa0dVe7iTaogQH1USW7XdDeAvOCwHeTjbQ/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8FtbmSFg2wqUz5zLmn8iyBTk7ZpUvB1nxye0y2l+Ioi5up/OZQTrX/kfgIrz95PZAAIENq7GEAzcHxRN4xA7uuqCw5z8R7caa0dVe7iTaogHwvZ3bgc7cnvcCYkII9qFg/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8FtbmSFg2wqUz5zLmn8iyBEN8vP0viDyhye0y2l+Ioi5up/OZQTrX+qPBzu2I66tQAIENq7GEAzcHxRN4xA7uuqCw5z8R7caa0dVe7iTaogQH1USW7XdDfvcCYkII9qFg/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8FtbmSFg2wqUz5zLmn8iyAvcq7oNwtxcdUr6WdxQVzP7uCOwCkqMmXKA4kX//DraZwf0M1gFFqmZeYrvFxsVeOHXjnEs5qlO/UWDsIJp/5JautoXujtsnmH860fPQD/v/hoiL8D6lHOMZaJukqSckHL8ElX1S2IiXxpZJSDjlAnCoMDdDSaWK64ugDXg6fOP0DeFbQdyaYIUZng4HY3Blyw5b3DwFQVuWtLVNc5sYlOVHhwVSfQjW7QGI+luyLZunKktKCfYgnyPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuvmNJa65VppwDrVedGrotX28MVHSMhCB3E4HupafghKjhKg5+1vcC/pAkNgHZGapfQcHxRN4xA7utKRHJCBL7wHdxP4sBiSHxpPHrYr99U5d+ZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4sEkaS2Wtaw7GiMFB2SyS1+Eyb4ko77PQ8MVHSMhCB3E4HupafghKjh5ARjasmhIPwkNgHZGapfQcHxRN4xA7utKRHJCBL7wHdxP4sBiSHxpgYxcyYN63+yZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4sEkaS2Wtaw7GiMFB2SyS1+cd7Yk5eqV08MVHSMhCB3E4HupafghKjidZ92yqwN24AkNgHZGapfQcHxRN4xA7utKRHJCBL7wHbQYaWirHqtbCYQ7e2dQXkaZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjMqwkCXMsFjnRRAfo7xIEXhjTkCQ4AIAmq0/SkN6W5/Rlj5ABPnt5iWPkgOcaYXn+9eHjgSu74bb8MV0T8SMBWoFn1HcPHcOkYuxPUN2+8SQr2qHWF7qOUAo8DxcgTS24wpoifs1g0sYgvlmBdWPHvspoNZZH35B2+hDShfbp0ofwgRSgFujcDCMeez4Wyv2dPge6lp+CEqOMsDfwwWR/EJW+PLWHJwcdsoKmVcgLNIxWW7fUGWdFS/4uHChJQoK4Wh+6WYAleXJyd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+yACMl1sbMi4sH1RA1uxPCrT9KQ3pbn9GWPkAE+e3mJZ3FMN4gK4+dwkNgHZGapfQcHxRN4xA7uuTJ7waA9Pt9F/pozoqkiE/AuVDdVwCsQgPyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoPBbW5khYNsKogn5UWLR4Y64OEQcjbV3LS4ugDXg6fOP0DeFbQdyaYIVdbS25li+vxeHjgSu74bb8MV0T8SMBWoE1isglIQbUtI95ulwcX+qTx62K/fVOXfmWM7sg7m9pItp3y7fmTZdcVSVVRNYpozshsyfOCZT+LBJGktlrWsOwwdk2R1rKY9LgCPmYBxuk8L1TEereSyJoonk1nQhv9VzjUPwX1Br9BldhL9taLl2nARTTIGopTtCaezB0BxP6JnZbl/TR7oCeYja5QdxnwhQZl+0QKwT4iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUjBSInkgkznPogn5UWLR4Y6miC5eSi0PUbnRtsmIhkLd+7gjsApKjJlULsX8fby+WxInpw+XUcVHixFxpn4DsyzuENd/xwlui/SZ4vGg75zhwwdk2R1rKY9e9DNL0JiEfk+3wUp4AHlaZpBVhazntdDFXX9LD/Bi695zs5PRIUJliwfVEDW7E8KtP0pDeluf0ZY+QAT57eYljFt1Uh+k/jvCQ2AdkZql9BwfFE3jEDu65MnvBoD0+30PCmsD21LywkIqzJr0O6rZQ/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8EmZGuEoHlflYarIpZQJ1JYLfnqC3KLi+7gjsApKjJl0e+vGXgoG49ICcjYAhxhTubqfzmUE61/zlUcE/kMgsPm6n85lBOtf88TcoFBIGQ1gL4h8L7dc5TAWCwd+65pMMBYLB37rmkwibqvoBhHy2oxtR3Q+abawFIMZZvCIRTZ5SPM+hJzjW3ib9EZFcK1pq+HyfyXV4dpCUY4f0NlNxXAWCwd+65pMMBYLB37rmkw/1U4QQ+VIc+6oe5ZwWKZz/6nD7KtPrUjpy9c5V1y28LRoNlryl3GkKD6vHWL1wQ4UcgSq20hpbaAviHwvt1zlMBYLB37rmkwwFgsHfuuaTCJuq+gGEfLajG1HdD5ptrAebJzwzT13SLlI8z6EnONbeJv0RkVwrWmCKIPZGb6AdkJRjh/Q2U3FcBYLB37rmkwwFgsHfuuaTD/VThBD5Uhz7qh7lnBYpnPeY4UkN+WwXenL1zlXXLbwtGg2WvKXcaQoPq8dYvXBDgPcesR+JIAFIC+IfC+3XOUwFgsHfuuaTDAWCwd+65pMIm6r6AYR8tqfMbopcIV/2AEm5ZiMMicMSSJw00xaEzAiTDnoEFFNUGDuQfuaEzh6AEuZ0tVGH/EW9UgCDHWybhoNxvyQ8QW1ibI4OU01kkG8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTiY1xyRj7Rgnq3YFFR2s4AFQEo83cZQQWl/ux5LaKvyLSu5NX3VJkLh+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC4kq3srN7+p8SDYYEZZ2nr5tri1hIYa7vqDpZWXNzWXSk5Ok5wGBoKhccAKiMeC1ZbF3uU2H/DCyQO8ZxWsk4lK1bfk3tLW1g39e2VsGp8X0SHMr6Lrz5MSI6TSiGsXwH7B4b9+WeicmI/iWZAKMPakcoEm6npVGk1zyng9+sV+MVvRIhX62s/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv0jlKl6nOCHbCOjqeEmbrf5w8x7FCxIEFBZzTaPe77adLl4hH35McanPyYcPjMVpvtG1k0bLNkme26DEPZAh35c1E1Q2lqdtFazGz0g/SmcE8IhG/YUbO4zZK7g4ampf7WKXzNyqi3M+gY5Vv5jPDWw6PQKP4NFnHYJGrtkz11nH6O8+JEslxo8nr+ei788bEm5qj0sPQYIO6gnuh/ZnB5wFgsHfuuaTDAWCwd+65pMDawSr20lhs4g5NPl9WzoWZahzYZ9tJ0oM221Vos8FzOxE/4L/XDFvWlN+pvRdTl2l4QwmYzlPiZHOIUBjz17Vj6nY9cDso9N79X4crs+u5RewPNu32f/eGjfpLEgKvDGxXShtQxdP0CeKH7lgMGsxjyev56LvzxsSbmqPSw9BggOnQHfseN1W2iJey38Y+ojMBYLB37rmkwNrBKvbSWGziDk0+X1bOhZtIlAvFZUXkZV6tt62a8zsPET/gv9cMW9aU36m9F1OXaExWZul1JXMYBsayBXPyLMICT2Jt4VBR2v1fhyuz67lF7A827fZ/94fRreCzFsdSbFdKG1DF0/QJ4ofuWAwazGPJ6/nou/PGxJuao9LD0GCDIZBJy55F5B2PfHdw3b2XBwFgsHfuuaTA2sEq9tJYbOIOTT5fVs6FmZZuZtM1PHBRXq23rZrzOw8RP+C/1wxb1pTfqb0XU5dr49sHv18Hvs4Qcor8g32PhKhBzSnCQ4Zvmt36QlX0Q+XsDzbt9n/3h/FBdnSjlYy2l7bduICzwyHih+5YDBrMY8nr+ei788bEm5qj0sPQYIKjekj7PLyzlIdWHn/tImo1S7PdmcHtQkDawSr20lhs4g5NPl9WzoWbqDrFSP5gmhrwm8cgZNBLlxE/4L/XDFvWlN+pvRdTl2vj2we/Xwe+zhByivyDfY+FFfhon9Z63XL9X4crs+u5RewPNu32f/eHjQMkG2uqQeRXShtQxdP0CFVx6xUxL6WLyev56LvzxsSbmqPSw9BggLyMqEjuETCk+6l4HoFkDusBYLB37rmkwNrBKvbSWGziDk0+X1bOhZtkXVyocKJ+FAsZgPlJkaEzORTQOSZQ9adb6GFURAaIfDululkiFa5lB2HI455bXqbQPXlvw1m1bKgczd/8Z9mfI/BNjjA+uCOqHnTxe7YG788PibVjkjOCZtOaV3rbA4yDSP9OTl9aL+OKCIfZmM5iLqUS1T6hWSAW+NPo/SQQpc09lhEMC2PECca2Mr6/QFWJponaqEc2oUH1h3alkV9BwdEvRp/kjAajekj7PLyzlfOKrunFvcMnWmH0QnDKBioTGSR7/wOaPupmkdEVpLFv1vofQevc2tmuiOljGxGW0fpRLPm1xe9wElSR0X5ynT/GwAIE0kyRp1Zhhgo82CzXkaib+wtDPsEodg7Lws3CNS+NUGOoRoh/JeV/VJ1seV+WKUQGTYMurzZK7g4ampf4KZLMr6/GicuTWdIsLxu3YmbTmld62wONHnAPdOL3wfsveA38T7xVm+hcwU+8igCxoGTNZWuj7uC09xTeuFeweEWC7FcyAyxdixpxRaEIXoGvu6TVpIgPAGYgIHXcSjdM9xXRXH+EVT/GwAIE0kyRp5mqb7vBk7RW9w0HqmYWYMwbuk8DkJFmvBb40+j9JBClzT2WEQwLY8QGAmYLC0O7mYmmidqoRzahQfWHdqWRX0BMVmbpdSVzGLDw1gsxVpXifsyT7eXUhjVCtKGqLmpTaWPCrRU0PtFrRyiDpp7quVMoWlcOw4K3IOMKA1BJV2ZNCTfkjIiJ1ezpOP/sHbWg2WtEXmuBxTQnbSmVqwiEmDr90/v0Oz005t1gwaU1AuTsMK9t+o8D0dchkEnLnkXkHYDiOqM/SkqczbXroVfCi1iTBylNvINu0vFOYt1VUKzQq7g44yy4ZF8fUFAOJ9pO0Yg7sjBccnaQRYLsVzIDLF2LGnFFoQhegXS3eknAq/xtq5rJdx2fk7kWfVdjHDYIfmbTmld62wOMg0j/Tk5fWiylT+edzSvSu+LMsTVxkkjRKHYOy8LNwjUvjVBjqEaIfyXlf1SdbHlflilEBk2DLq82Su4OGpqX+4m/RGRXCtaauhT3ZL8d6DtRipjlsWqciMlkMGSopX0EBgEF9iKWsJiZ5YxE26THe//uvj0VI3s9oGTNZWuj7uOHXq/nAzeXBHLvdloCY0mzz0K/G13USSXU6W6ipCpMtD/XfrYjohNxU7sH0ORZZlalY9muNMqqWUMc8eAUmMqAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsAyrlX0gor6tVKtg7aPDoVB3ByGK/VBOniK3a0yLM5mRQQDm0+FyW5cCrRrGz4N4rFPwThf4xO935KcFXXGVwNLFN64LgH5CMAyrlX0gor6oXOWdKa6EuwDk8imoV7y6D307+4oPX6k7Qzy7YJtQYj2jmz4lCH4bEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsvZXzvFjDk/E8jCmrTA34ECueWGoonK3GY9BCSCKyXy1idipxlUuI0S33hUU5oIdEEWH4+LwrdSY1qeF/3xLYVZd6RBKNM6Eip9JBxvAjUF5wM/7WNDT+Ht3Ho6t/zr3ksoGaY57rssvI/lEFVd2N1YsywZ1gXwb6mbVrC4uDyJdep2m4JtoMoFA6vM2qPhqpzUTVDaWp20VjtB2TEMtvNad+WbYZY/O1oMcDzmvmwmbl9wsIcAO/aMCAsaLkc9sMgi9P5Q05ExDveSImX13A0+XS6JX6v8WPBH6ab6nFM+gGrw5g00TiRSPnsHct0Z2uGhC8xWXi+vkB1ecXi+MYnJCA3jbO26lYwICxouRz2wyCL0/lDTkTEPbEZ6naIcP6yJ7wgeFyU0wFg0CdygaSDn6ADi5zKCB+ti4k5ZgE8lTAgLGi5HPbDAi5nyDP1E0AcKEGREeUMHmvQikJWPE7CHYNbLmfROv/hVAuScmh6714JAwcpRs2w1ZmiKIU3ioevUCBeDMp+9ViCACHbNjEqs6bgY2Nlcm1I9kKMFmdfDUIUGh1sl2hPAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4eKGpOrlOiEVxvp9bPkM0RglM7FV/qoydnBYUSx7a+c9gGOw6IbIHiyW7JZH99t+/fV4cqecEQZ5x+FwTj/4LLfD/XfrYjohNxibtLw1suKiJTOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMPKnNj3pkyIuRebox+xhZpBylT+edzSvSu/vtmPKIB8DWUzsVX+qjJ2SOL0yshwRnPGJQkVdzgUcRUVhyWEPx3h366FIYjonHOhi/bTTov/ShnoSHEqvB8JSdQKgT5HtzBAWDQJ3KBpIOSxWonF3FK3AJxrYyvr9AVbUXfYiX6zhStTa3BCpnBViKxJWMbtP+K4g6XAIaM8hjt2GEi72SQ8pTOxVf6qMnZI4vTKyHBGc8YlCRV3OBRxFRWHJYQ/HeHfroUhiOicc7zlo93ttcu55z7681AJDFt8O9AYQKqaGTBH6ab6nFM+q0edPGUxp3R1VqsDAgUsejhwyaAxLfQPR+FwTj/4LLfe+h1QpBcEtTCkbUC/ymmpWapAtUxcGjDZgJhUdyymnnCCkB/cWqSlh+FwTj/4LLfXS3eknAq/xvq1ME5GgnNCY7krx2Hekt1rD1oOhUnp8jqbdmcoQYqPHRC9BQrQSJ4wuDhMsVKUw+HosDvcT/uYYrOej0JtLplmNyYxOvt3Dj1qhHaBp+6NwY9SJR7MwFURGMUc4ji0lz4mOpF2SzOOUIUGh1sl2hPAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4cGPUiUezMBVOXOd1VVqUVwW5cYTe7mmfxMF+YwSIF2OpTOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMPsUJYN6b3gXuhiWHG0TehoZLFsfdigeEoDrmenQuEMZasPWg6FSenyOpt2ZyhBio8A6iWb6ni9GLC4OEyxUpTD7FCWDem94F785IGI5msKUopU/nnc0r0rqPBMYH68KDQgJnn4ZpykqCsPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPXVkydSh8I56zFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QCHQmrIhRtd9ipQ3jNDYXS8IKQH9xapKWdWTJ1KHwjnrMU4UVpv+iFFpoAb+70/qtPBRehIFeP5D3IEJC81H1gSXoPohMQjK5rR508ZTGndGpcg1sRIlPCWvQikJWPE7COkoH8fk64rbBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDpqp+dU65i0NY9onXBLEFsaUzMxN3ZVssA6Sgfx+TritsEkaS2Wtaw74m/RGRXCtaauhT3ZL8d6DkIUGh1sl2hPAWDQJ3KBpIOSxWonF3FK3IHGXTL4rBS7bUXfYiX6zhRcF9VXEWYWH8jsdcB259qXEjboyxTc6gtBTMhRiSfbJo9onXBLEFsaeTCTjlA57Y34SW4WqIeN74mhOIgMLbIqYsywZ1gXwb4XS1JnD+2owaIc/j4NtRsPsNMwfWlh5XJhzq3JVb0AWgteLEy/ay1AaMSTESCu1grAk8yfFtp1eSgaRNLNiI+VNz3gAPE1y+XnSv/rNmDxCR+lFIzyhXH2NcLAKWIy4N3VmaIohTeKhyUGtg9pP9WQ7GNtU97kTE2caiSB0pwUU4Ke3RH6KbgnPB33uCU9gsmdGlESu52O3qWv15BBneM3HEcuJ+RvSwaFVSD1FKcXtBMFz68YcXSzNGERh5UHqB+laqHQ6HYhZedK/+s2YPEJC4aCMXedht5TMzE3dlWywCvkwtmFLeT2MLHXl0A1q5CUzsVX+qjJ2ToUI3EUh971pyenXn87dN0ZpIVGa7hueH6USz5tcXvcImO2CPc/mOydGlESu52O3qWv15BBneM3HEcuJ+RvSwaFVSD1FKcXtMb2a3wBSeOckex5NYkW0nHL3gN/E+8VZiJjtgj3P5jsnRpRErudjt6lr9eQQZ3jNxxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnKGJYcbRN6GhksWx92KB4Sj1p3wp7+lMkZ0aURK7nY7e2zczD3UmsM1YggAh2zYxKvJMoiRRwIwd7tFfp7RZlEH49sHv18Hvs4Qcor8g32PhMriQusSU8tU9zQjfrwajONWZoiiFN4qHr1AgXgzKfvVYggAh2zYxKvJMoiRRwIwd7tFfp7RZlEH49sHv18Hvs4Qcor8g32PhKhBzSnCQ4ZvthTHR3gweKdWZoiiFN4qHr1AgXgzKfvVYggAh2zYxKh4IBUHNephVBRR3UE83WBLy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR01H72YelCd0zaFhFdGDGyYF/eDlOHv3OPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHhjKp2FzSqRcFPFe6/fnC3eJAThBJWHVsO0+iUPoaTRGUjOdoYvdN1E4TwpSzHp6Ar/vwphgnNk1oMcDzmvmwmWA8dKC/IiZKWqTz3+mLoAi/3bzWigGMNh8gtxiLTTHiH33UrlGN3lACBGvtTONhTKg18ZZFxsrfHF34gAZl5q3pCgYVS10ee6g18ZZFxsrf9FxOwknxBjDmj3izMDWou7PE7sQG274o/OTSx5nBfjoZQxDboJX1nKg18ZZFxsrf3McuJTQciynLTjWqmsp8bL/dvNaKAYw2xPY/UBscfahTwKEe72PazyL4/FnHICy/ZjySmeLaPspsru3Y1NZombakuKnTOGrNnwDziWeYZMwT4zO4pj1qZBEDngQVB3aKK5CNUm9ffMgJtl20oOO+OlebVLa/4c/QYNTLRsAZTMjCqXKmYipQJp7JkW377qQRQ2VMWsqE7wX2pmJ83qD0Bi5HanjcYjPwrudjzAtOtIQx8+fSCxlRIGxst5+uOWZi/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMj18jBjNADgTct4uUjQIxzu2TXWro5hPKgST972Z2KoUf9IYEvNtEtBgcBPwf5Ux46OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZWeKdmTkEiU0T1OYMshcsCf5/znXpc+s3cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMk632GcagQymWr0q4Z/j5AJl5pP+/w5LVg8M/XPHF9qDN8hwkaeXL9enkzBWt0tJvSR+EYhUn6yngsHxKdieRYm6EfCirzLRNjn0y093vawblg5fuBTrJoBFmqADANE/LQ+khXpbcj4Aatbd+TLr6lu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6qelc3ICaMs8vIyoSO4RMKQatbd+TLr6lu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6qelc3ICaMs/IZBJy55F5B1trLI1DCBJku3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6qelc3ICaMs+o3pI+zy8s5SHVh5/7SJqNieFpP4FWKPa7cHGcmccaLbdTi1x3mcIYkNEPMoCb13rs5bybePbTw10t3pJwKv8bauayXcdn5O5Zb/h0F1jGIpZWH16/+TeYenPTtAYOt1YEWaoAMA0T8gGAQX2IpawmpKFk2NHyLDmjtxhuLD/JGDQ68/3TNPUeGmM340wuvpGzpuBjY2VybVwX1VcRZhYfyOx1wHbn2pcSNujLFNzqC6u4Oe4qWCLJNeiLyn7WySUvB2RBqE8QgwY9SJR7MwFU+PbB79fB77OEHKK/IN9j4Uctn+VEzmHLu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d67OW8m3j208NdLd6ScCr/G+rUwTkaCc0JHbOaRAXT0K52qGJ/T63OOPcYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaFwX1VcRZhYfyOx1wHbn2pcSNujLFNzqC5YlHfB/zqZzNeiLyn7WySUvB2RBqE8QgwY9SJR7MwFU+PbB79fB77OEHKK/IN9j4SoQc0pwkOGbpWNWXJa/ayhJz5ieEfkatLFCWDem94F785IGI5msKUopU/nnc0r0ro1AyzbeWK2KesjGH/xN4DeQ0Q8ygJvXehgAssjGryytETuc2nyyzNzmIqollrQmapy3rp3QMllqb2xHjiFyDfwYa77f8vmAHXg7KXxLmSbKvg4z4i8XZ59wG3LBXMR64XT3wXUszLSfSMGkaYCErkSC9TX5sAYwGhmkhUZruG54fpRLPm1xe9wG4YpXUZXOeKzkHOTCS30lcBtywVzEeuHoK2LoobfvSqg18ZZFxsrfeYj6+rMrrz2pkEbAltJTXcRMPKQaiwwWXOif352RW45oVOelkqJIZ8BYLB37rmkwqelc3ICaMs8vIyoSO4RMKQatbd+TLr6lbi+kv3mC/7NHnAPdOL3wfsveA38T7xVmhGZrIqJy0orAWCwd+65pMP9YOIVlvcdJyPwTY4wPrgjjBbh5aeA0wLTNVOuBc+aOGGu+3/L5gB0SWqOwp1sS2da701axnPDWKfaITWj4BHx4kcummI9H4FqAH25hGVE6o8ExgfrwoNDZfZr8a7ghl6g18ZZFxsrfeYj6+rMrrz2pkEbAltJTXcjsdcB259qXEjboyxTc6guWJR3wf86mc2hU56WSokhnwFgsHfuuaTDs5bybePbTw10t3pJwKv8bauayXcdn5O5Zb/h0F1jGIhyniG+FtOw2enPTtAYOt1bAWCwd+65pMMEkaS2Wtaw74m/RGRXCtaZafD/+ALxcOu9+5wueZjvPYKWMQYJDY4X49sHv18Hvs4Qcor8g32PhNyyZzWckHYGoNfGWRcbK33mI+vqzK689qZBGwJbSU13I7HXAdufalxI26MsU3OoLq7g57ipYIsloVOelkqJIZ8BYLB37rmkw7OW8m3j208NdLd6ScCr/G2rmsl3HZ+Tu+jci+PTO5rocp4hvhbTsNnpz07QGDrdWwFgsHfuuaTDBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDpXKYJnDCCQGWCljEGCQ2OF+PbB79fB77OEHKK/IN9j4Tcsmc1nJB2BqDXxlkXGyt95iPr6syuvPamQRsCW0lNdyOx1wHbn2pcSNujLFNzqCxVg51sseBcXGGu+3/L5gB2DVgVGxEJLFsxThRWm/6IUWmgBv7vT+q3tlKy0BxrZYqLFi/scuo1Mkez6ymeMObzib9EZFcK1pq6FPdkvx3oOs6bgY2Nlcm3AWCwd+65pMJWtQOXMvcI5AYBBfYilrCYmeWMRNukx3rgAR1pFKyWsFpYxxog+HqbAWCwd+65pMKplFao/xeJqWsZICMKqI68Ya77f8vmAHZoEOBo+KxnymlYqV8JzNNS9qwVKBkKzMMFs0X7NnVetAEpUG6CU5b5rHszq1lh4rmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqayqeX/Rm8uL/8yH9OclHsqCXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiYrwj6/ble3V8b2J4ODUGYe/n/Odelz6zdwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyTrfYZxqBDKPvyh0RNWxkOFf1lN6qbqa+2d+iBc8v0FHyC3GItNMeLnbSP9FHkYHWRXZEp4UN23chK2rhaMLmZP5DKhKevgqeGFB3kb9erk5iKqJZa0JmrYMn+n/hOve+0xGyrcuuIebPz/c6/JJ/2iPRAJAhOGHgwrjVQlO79KZcxmz9AAC0ynxG91hzMy4FFj5+cursX8ETuc2nyyzNzmIqollrQmatgyf6f+E6977TEbKty64h5s/P9zr8kn/U/64RAvyEUwdS3Qs1O+kMtg5eK7mvUD1g/ausd1vV5GeeTDpjMk28+WnABkhfYwG9iuoTHUj00c2NMLgoDWiuxM0u5Yi2s55XyA/Cw3lzwqkYxlJQ1vSfRzUTVDaWp20ZJXSb5WtpQPWsvbF38YWeRrZ+Gtr7w0egZFOCT/k9dTfHWjXjdtXbuoNfGWRcbK32Y8kpni2j7K3OXkGArzLsPlwA+e7vpE+CZk7z5A4NNOqDXxlkXGyt95iPr6syuvPamQRsCW0lNdAl4sQ6AqDUYoKKuNvHGhBmhU56WSokhnwFgsHfuuaTDYMn+n/hOve5Hs+spnjDm8djhLaH2iFg7bzi48hZGtVXh3H4ZkRldnXS3eknAq/xtt6wIuBii1Qwa9J8dSovWewFgsHfuuaTB72cywEGpcnODXEbg5Anphcij4eRVyAumEHKK/IN9j4Rdv3p8ka1QY5mqb7vBk7RXib9EZFcK1pu7y7xKZUUK4wFgsHfuuaTDfm5UNID2G0ybmqPSw9BggOnQHfseN1W1Gb4vFzpjnLBhrvt/y+YAdg1YFRsRCSxapl7Nk+TGKVdWYYYKPNgs1PR1ZPkCG95H8Ug8BLyqKN9WYYYKPNgs15RaV/VNBYMuoNfGWRcbK33mI+vqzK689qZBGwJbSU13ETDykGosMFlzon9+dkVuOaFTnpZKiSGfAWCwd+65pMNgyf6f+E697kez6ymeMObwKZLMr6/GicvNfRUg6mxuUqelc3ICaMs8vIyoSO4RMKSSlAliNaL4KwFgsHfuuaTBF86nqKnwwoXiwRHgxhUbuo8ExgfrwoNDnoJXGukoD3EjBpGmAhK5EOvzm46oTw3GUUHQYVZ+36L3VzsCVlJsRksWx92KB4SgZk84juCgeRhmkhUZruG54vFOYt1VUKzQnbT1CXrelv8BYLB37rmkw/1g4hWW9x0nI/BNjjA+uCKhhBFMpp/+J6HR8CEQJtVdL/DLYQ9qk3MBYLB37rmkwSPZCjBZnXw2B/JGDlqdOXrZ3Gf53ZAxHFQtedYZveUjH+FnN8AkdWOZqm+7wZO0VvcNB6pmFmDNKA9y5nMGi/Rhrvt/y+YAdg1YFRsRCSxapl7Nk+TGKVU57CX+OERAHVFRhhX9UzsUyfGSk/TQONvbKzPqjkHxfAdK3RMCBo8E06B5Ztle+kCKxoq1FrDYswFgsHfuuaTB/SH/kfW8Kmry12QL5tbb2e+h1QpBcEtTCkbUC/ymmpTH4bUBAm8bq9srM+qOQfF+N2p7PwrYmODlcf7Xe28zEuS6pK8U6jEUYa77f8vmAHXg7KXxLmSbKvg4z4i8XZ59dLd6ScCr/G2rmsl3HZ+TuEH5VokFXcQhL/DLYQ9qk3MBYLB37rmkwSPZCjBZnXw2B/JGDlqdOXlpoAb+70/qtPBRehIFeP5BfWADTFbkpBPj2we/Xwe+zhByivyDfY+EyuJC6xJTy1VEAxF+JRlisWsvbF38YWeRrZ+Gtr7w0eusFWlD/XbfQKVP553NK9K6jwTGB+vCg0JwAIm6voaaLwFgsHfuuaTCNmlGfQjyG1lqAH25hGVE6AYBBfYilrCakoWTY0fIsOWslaivClYdOwSRpLZa1rDvib9EZFcK1plp8P/4AvFw6aKW2sdGKPJvAWCwd+65pMN+blQ0gPYbTJuao9LD0GCCo3pI+zy8s5YpE722OMBL4/QaMRZ2eYTTAWCwd+65pMHvZzLAQalyc4NcRuDkCemGo3pI+zy8s5YpE722OMBL4pJekojrv4K3I7HXAdufalxI26MsU3OoLlRe277/u6FHAWCwd+65pMKplFao/xeJqWsZICMKqI68Ya77f8vmAHZoEOBo+KxnymlYqV8JzNNS9qwVKBkKzMMFs0X7NnVetAEpUG6CU5b5rHszq1lh4rmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa27kaxZD4JNmB6dMgmnMCSPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+XJ3oG7RzGOQRGMUc4ji0lz4mOpF2SzOOfxSDwEvKoo31Zhhgo82CzXlFpX9U0Fgy+zNictq7nhGkex5NYkW0nHL3gN/E+8VZo3M0rvEzQHukex5NYkW0nHL3gN/E+8VZqrn4HUfnwG0iPBa+e1y4mLIZBJy55F5B1trLI1DCBJkqelc3ICaMs/IZBJy55F5B0N1XstUC8zIXBfVVxFmFh/I7HXAdufalxI26MsU3OoLliUd8H/OpnP8Ug8BLyqKN8jsdcB259qXEjboyxTc6guWJR3wf86mcxmErH2aWvtpzFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QRnSNGW11ZNnMU4UVpv+iFFpoAb+70/qtPBRehIFeP5Cq953i5K6w+qDLoNsELlx7S3cdS8o8J0QJKWePQB2wkLSCXgofxdjQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Ltx5v2R/2i7QW6cR3ugt84yOSikUR84Jm6vt7lh6NPTEyIl9tcDvIrKwQFMBrptmFt2FocRTvBr2+YkbIMZ8A+du/y3mwoDlqvnujeI7UaGwAyrlX0gor6r2mUL5zLINh0xHdww1hvD787xs4Igtz+f5W5TAUTX/n5GZOfoZUdm+AK8wOanajkx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC8axWoQJD0/V8wrXqzAFqTpoOtXRJq6nKxoeVOYqyZ8qAWDQJ3KBpIN3BLsxLlj0rNKAiuTcO6Pxj5hK0qFhWSu9bIqll76wTNep2m4JtoMosI6Op4SZut82DRk4iUI12S/3hOVKUaEJ4V5ngPiPCPQv88qbGbLEZ7BQFOQvZ3yipgq0LWib304II7KNV4xCEDSCYyn8060xoSF3Q0r6i7ZbXClJvGx7XM6CrTtw71PvEK4b1Uw2KCuEHKK/IN9j4VgELcI2cuHlRg0eF18pdwGOls1gEoxGuzoxYt3pSknswpCjBmmYgMW1u7nMy4XTYxvwPBeGDe/SVCln62da3lgmpZsQwb0+snFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/5uhHwoq8y0TZgJhUdyymnnCCkB/cWqSlmpGPxRfAM1oyMokQ8Xzmo/R8jzVqDLOsZZruN9kNGOkcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/ruy3PTCzp+zBH6ab6nFM+gGrw5g00TiRDy0I+VfMnMZxX2xf0wa4os3NonL3dWzRV6fhQIgtprEcRy4n5G9LBnPKxSUCjyIDxPY/UBscfajVoAiB1/rvWAFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHjZpRn0I8htZCQfT0TITgDyXoPohMQjK5rR508ZTGndGpcg1sRIlPCWvQikJWPE7COkoH8fk64rbXRRoUldjjPXHO1gemEq84IIvT+UNORMQU6HCot6Ji8IacZmbQr1UlWl/Wb6CXunL4alyc2izGjh+9Z2GdoKbiz9+B5bv6EKgwICxouRz2wwIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTZ+gA4ucyggfcHRL0af5IwGo3pI+zy8s5cWrKszvv/rP+PLhl1syijpOYJTDnJE81WvQikJWPE7CHYNbLmfROv/I7HXAdufal4KLY1BA6bZNyFcFEqvNbKgrKQvEtQJT6v61wG12TAEF4cMmgMS30D0fhcE4/+Cy30ukEgwFloGoNOgeWbZXvpCEEQlJ7h2uIPjy4ZdbMoo6TmCUw5yRPNVr0IpCVjxOwh2DWy5n0Tr/TnsJf44REAdUVGGFf1TOxZ0JM8ktFmf88bsTdDFOIKACG93JMuWgEViCACHbNjEqs6bgY2Nlcm2oTNF0tV1F+dnTBVNxD3DLXxLt6MFIZvgcng7b/emm3JTOxVf6qMnZwWFEse2vnPbi4XgOVDPh/08MDQF/7jEYzasixnaPUTISW9VF0VD+74jwWvntcuJiOnQHfseN1W2us2AGBIuFmozFeE1XahSKMZPML60V2LXsY21T3uRMTUdn1ZhMqr1TiPBa+e1y4mIvIyoSO4RMKbv8Ik5kGtKeseXHmzxgscwRaygtE5naOViCACHbNjEqs6bgY2Nlcm2VrUDlzL3COaPBMYH68KDQ64PPJGXeuIlipQ3jNDYXS50aURK7nY7e2zczD3UmsM1YggAh2zYxKrOm4GNjZXJtla1A5cy9wjkBgEF9iKWsJqShZNjR8iw5oHRlQ8QWhbsHCIkzAlfR/DGTzC+tFdi17GNtU97kTE1HZ9WYTKq9U4jwWvntcuJiqN6SPs8vLOUh1Yef+0iajWb6dEN41M4dQhQaHWyXaE8BYNAncoGkg0dn1ZhMqr1TiPBa+e1y4mKo3pI+zy8s5SHVh5/7SJqNqRUU1N4gI04fSSbQfgTQYg+w5CPuIzPya9CKQlY8TsI6Sgfx+TritsEkaS2Wtaw74m/RGRXCtaZafD/+ALxcOmqn51TrmLQ1j2idcEsQWxpTMzE3dlWywDpKB/H5OuK2wSRpLZa1rDvib9EZFcK1pq6FPdkvx3oOXvIB4bqOfyNUzPyzuUT83YHGXTL4rBS77N9ax/BvGXN+TFSQ0YK9gCkijeLlTTJuZGbUJZXSqmMuc92gsVwEKq4Ga14AP/SQcyP8LAktKTF0U64xg9zGNqPzmJ8jav8gQVlWo4auvX0F7pVL7p7RG+7RX6e0WZRBRGMUc4ji0lz4mOpF2SzOOTA7z0L52nuKAi5nyDP1E0C7mVmb2+QTluxjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3cRMPKQaiwwWXOif352RW44wO89C+dp7igIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTZxqJIHSnBRTyeCHG2BJ/93I7HXAdufalxI26MsU3OoLliUd8H/OpnMwO89C+dp7igIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTZxqJIHSnBRTyeCHG2BJ/93I7HXAdufalxI26MsU3OoLq7g57ipYIskwO89C+dp7igIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTZxqJIHSnBRTyeCHG2BJ/93I7HXAdufalxI26MsU3OoLliUd8H/OpnMaqFZvLSpfoMIKQH9xapKWFIjp1DOt+yelEQYVtBkl7QGAQX2IpawmpKFk2NHyLDliI0tlVN5G8zlyP1CVms/HIIvT+UNORMRBboDWT8dzI8EkaS2Wtaw74m/RGRXCtaauhT3ZL8d6DjA7z0L52nuKAi5nyDP1E0BUWxYGrwGYr2vQikJWPE7CK+TC2YUt5PYG0dbeBYeZllpoAb+70/qt7ZSstAca2WJByPWgy+P8E4NxIMYhzmp74cMmgMS30D0UiOnUM637J6URBhW0GSXtAYBBfYilrCYmeWMRNukx3lAetOBgipkylM7FV/qoydmtIS3jmEoPV9Bi1HNIhaN5D/XfrYjohNyJUnCjx0TtPPBwnZcmTAaAjmJuTaztkfqj85ifI2r/IGIdbto7m/FTr/vwphgnNk1oMcDzmvmwmWA8dKC/IiZKWqTz3+mLoAi/3bzWigGMNh8gtxiLTTHiH33UrlGN3lACBGvtTONhTKg18ZZFxsrfHF34gAZl5q3pCgYVS10ee6g18ZZFxsrf9FxOwknxBjDmj3izMDWou7PE7sQG274o/OTSx5nBfjoZQxDboJX1nKg18ZZFxsrf3McuJTQciynLTjWqmsp8bL/dvNaKAYw2xPY/UBscfahTwKEe72PazyL4/FnHICy/ZjySmeLaPsqdTLLphyYjxEtOkCp1eAL5VOzOzyJ4+1+KGpOrlOiEV8iCHbceiYTstR99sDa+ZA8zXPk4u663XPfTv7ig9fqTQiO1mgCru3SUps+P36IcaX66FIYjonHO7qCe6H9mcHnk1R/0qxfD9V0dI7cCxkywnsmRbfvupBGtTa3BCpnBVtGg2WvKXcaQoPq8dYvXBDjhAiuoYSpfrNWZoiiFN4qH4/74IpolEUAhKQtkFpVbalpoAb+70/qt61ejeB7CfllFsjkxNlMDXF0t3pJwKv8bbesCLgYotUMlu6JFlLo2wgFg0CdygaSDksVqJxdxStycapXrT6wSxPjigiH2ZjOYXdwyg3Vvw+eoNfGWRcbK35xqletPrBLE0DzeiZcNnMufsyT7eXUhjeECK6hhKl+s1ZmiKIU3iofj/vgimiURQEukEgwFloGoNOgeWbZXvpAoFxQz+OPu27PE7sQG274oExWZul1JXMYsPDWCzFWleJ+zJPt5dSGN4QIrqGEqX6zVmaIohTeKh+P++CKaJRFAa+7pNWkiA8C9w0HqmYWYMz/zggxTgkvWqDXxlkXGyt+oTNF0tV1F+dnTBVNxD3DLXxLt6MFIZvgEZsiqy5mvqY5lKAKEITi3vcNB6pmFmDNLHKr89pLzx7/dvNaKAYw27UaAb8Cd6MNaaAG/u9P6re2UrLQHGtliuGU6IEifNW4CLmfIM/UTQDzeJ4w52xBf4m/RGRXCtaauhT3ZL8d6DivpSG6EcHg/5RdZpRNTfA3jES9EfGyAKJis8nXcgBlZsrgO018QId8GPUiUezMBVERjFHOI4tJc+JjqRdkszjmbvgjOrX4mndWYYYKPNgs18QOiFCwIqoOoNfGWRcbK35WtQOXMvcI5FtoNCfe/cTd098F1LMy0n+B4LDznFf8qFtoNCfe/cTcmkPvW1+PXu2DUy0bAGUzIiPBa+e1y4mKo3pI+zy8s5SHVh5/7SJqNgBadNVQganWp6VzcgJoyz6jekj7PLyzlIdWHn/tImo2qtIcTrv41nmY8kpni2j7KwSRpLZa1rDvib9EZFcK1plp8P/4AvFw6/ZQRZKzLOf+dQOcf9n2nsF0t3pJwKv8bauayXcdn5O5Zb/h0F1jGImgGynhwCG/dBj1IlHszAVT49sHv18Hvs4Qcor8g32PhKhBzSnCQ4ZvN+bs+aHRbQPj2we/Xwe+zhByivyDfY+EqEHNKcJDhm0LQhhfkIQJ6XBfVVxFmFh/I7HXAdufalxI26MsU3OoLq7g57ipYIsl0xfW9MHVL3MxThRWm/6IUWmgBv7vT+q08FF6EgV4/kPLnexpGxX2FYNTLRsAZTMiI8Fr57XLiYqjekj7PLyzlikTvbY4wEvgbcNzpKwLX1Pj2we/Xwe+zhByivyDfY+Ftxbng338D5GY8kpni2j7KwSRpLZa1rDvib9EZFcK1pq6FPdkvx3oOdMX1vTB1S9zMU4UVpv+iFFpoAb+70/qt9Vn3Bt96V/1VDUsmMpH18lwX1VcRZhYf1Zhhgo82CzXkaib+wtDPsBbu5R4EL2JM+hVxEg4lpobVmGGCjzYLNT0dWT5AhveRGYSsfZpa+2moTXC84ul14Z7+ehYbqhzmucyxB55ZqQ1UzPyzuUT83cEkaS2Wtaw7CmSzK+vxonKNpXOBHzA7JFwX1VcRZhYfyOx1wHbn2pcSNujLFNzqC5YlHfB/zqZzxAHZv+4XFSxHWVEWiH2ZXl0t3pJwKv8bauayXcdn5O4nh/4cr3gUyBmErH2aWvtpzFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QIdvHuI01VL7WXTbMqsvSyPOSBiOZrClKKVP553NK9K6jwTGB+vCg0JgbWnLWx/bOla1A5cy9wjkBgEF9iKWsJqShZNjR8iw55sC5Eqj1cJ6QPtliQjzua/j2we/Xwe+zhByivyDfY+EyuJC6xJTy1bdB5F7FgPPG7OW8m3j208NdLd6ScCr/G2rmsl3HZ+Tu+jci+PTO5rriIjjpLFg77POSBiOZrClKKVP553NK9K6jwTGB+vCg0Di9a2BL4IX/WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFlx2fsw7CTQN24Jza30sa+RMfJuig+e8Pw+eaWrVG2eRMhyqqIMZwKRK8INt7Oi9OUnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTEV9N6Vokm8MpU/nnc0r0rsev3EEsczW5hX9ZTeqm6mvtnfogXPL9BR8gtxiLTTHi520j/RR5GB1kV2RKeFDdt3IStq4WjC5mT+QyoSnr4KnhhQd5G/Xq5OYiqiWWtCZqw19njuDvH2SEHKK/IN9j4Uctn+VEzmHLu3BxnJnHGi23U4tcd5nCGARM5a3QoG6cknd7NQpRA29mzfnCvpTk9bhdDjKl/Ez7cEVQvmZs4ZhxCvea/bRFrEL2TqHljvVfwSRpLZa1rDvib9EZFcK1pq6FPdkvx3oO0z27FDTt2FFXmAeYqCVGIMBYLB37rmkwyOx1wHbn2pcSNujLFNzqCzct4uUjQIxznrgr/BC+fs7N4uOh+kDjVqjekj7PLyzlikTvbY4wEvh2cn2ZqVXC7gwrjVQlO79Kqelc3ICaMs+o3pI+zy8s5SHVh5/7SJqNZvp0Q3jUzh2WnABkhfYwG9iuoTHUj00ckYxlJQ1vSfRWqPPshXK/MS4c+pcu3MV+uU0nLMA4Q//EgSv2O5WLUMSy6S9fGYN/6xDC+wC+o9lC9k6h5Y71X8jsdcB259qXEjboyxTc6guxhjzBgynmHqjekj7PLyzlJfqPbVbhADLahIj4LKg2r7lg5fuBTrJoA6a18nQNqwkBgEF9iKWsJiZ5YxE26THe5VhNOXCTDXgBgEF9iKWsJiZ5YxE26THecDDJtkD/KOkYa77f8vmAHb23f9HiueSywFgsHfuuaTDDX2eO4O8fZIQcor8g32PhRy2f5UTOYcu7cHGcmccaLbdTi1x3mcIYkNEPMoCb13oQ9BMUbPYIW3cMKmb+s8suajkcM0HTJMUETOWt0KBunDb9QuSHDNdeffqlppcnQWarsEsLMzN2ueJv0RkVwrWmroU92S/Heg7/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyPXyMGM0AOBla1A5cy9wjkBgEF9iKWsJiZ5YxE26THe5VhNOXCTDXgBgEF9iKWsJiZ5YxE26THewLrm9EHO66/q3YFFR2s4AFQEo83cZQQWl/ux5LaKvyLSu5NX3VJkLh+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC4kq3srN7+p8SDYYEZZ2nr5tri1hIYa7vqDpZWXNzWXSk5Ok5wGBoKhccAKiMeC1ZbF3uU2H/DCyQO8ZxWsk4lK1bfk3tLW1g39e2VsGp8X0SHMr6Lrz5MTO1vv0WSUjnNcq85VK+8vIo2NRHqTm3DxjdOVZjr39Aa2zEUq06bqVnBZlDDWPRc0fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv19JhV0Bg8FAX8cYC1vw6ZInrSOdnQKWp0tGcGsxfg0omtQ797AIb1pn5zUaoL+FImERhWsm5kQl8+HpiKWFvZCqlntSoAU7ex9+KGCXaa2T5v2IOUDBbobJUDlhYm1sYnD1iWiaJSn5FduQCOCMXeIonZ3rfEKafU1D/3jySdSQ7pbpZIhWuZMCeBBE3ASyzziCaTcQUoHNf2bOmVI2lUx+wdG5+EvQ7AWCwd+65pMMBYLB37rmkwNrBKvbSWGziDk0+X1bOhZlqHNhn20nSgzbbVWizwXM7ET/gv9cMW9aU36m9F1OXaJInDTTFoTMB0M1RvfJwNe2aN6VPfbOypYbo5NtfjTJPGPbG4bYuGlpSGygbCZLb6jWzKGLj+tqCQt1DnHGtR+23gjXOEok0Svg4z4i8XZ5+jlvYZ+HpI7pnPGMX0SF8DVgs9h4+iTue/V+HK7PruUXsDzbt9n/3hg+v9BeenSyyl7bduICzwyHih+5YDBrMY8nr+ei788bEm5qj0sPQYID8BqKRjeRUOHeMzOwvuJqnAWCwd+65pMCR64g5RIKvAmo59SWkrRX4/L4nKw8/pwKHSBYNLJWQtMCeBBE3ASyzziCaTcQUoHE0/IayWTXHR5SjyIM1enMcsnYen9zEpFcBYLB37rmkwNrBKvbSWGziDk0+X1bOhZmWbmbTNTxwUAsZgPlJkaEzORTQOSZQ9adb6GFURAaIfDululkiFa5lB2HI455bXqdHvrxl4KBuPYsacUWhCF6DO1vv0WSUjnFf1cPx4P1yKl2V2DVOsVDhJoF+NBx45uM7W+/RZJSOcV/Vw/Hg/XIpF3UN4ScCf1FCtKGqLmpTaWPCrRU0PtFpOlXUImUS+qOWKUQGTYMurzZK7g4ampf5+2dxAkrjxp4GDntZqY3nMTSJFaI2CnfpQfWHdqWRX0ADnBcUjTELbv9BdAi47BxyQBAeMuZcUI2YV88QK4B2gk5n01VZXCAqo5SojrNIEZQwr236jwPR1PwGopGN5FQ6s6xl1MTEpqjNteuhV8KLWtzwGk+i//fL3U4yioDBJCyutjB7GXbSIx9QUA4n2k7TUJ0gEyB12uliCACHbNjEqTTtsYR1Ybc5lrHSylh4UfewcnqbgcQbs6szc2pk6r3HxsACBNJMkacgAjJdbGzIuWJ7/LE7Dk+j0ypEypYbPcWYV88QK4B2gjZNCqE6lQOEcu92WgJjSbPPQr8bXdRJJdTpbqKkKky3O1vv0WSUjnM3+PKz8fDVslTNqJ4OEiDvSu5NX3VJkLh+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC4kq3srN7+p8SDYYEZZ2nr5tri1hIYa7vqDpZWXNzWXSk5Ok5wGBoKhccAKiMeC1ZbF3uU2H/DCyQO8ZxWsk4lK1bfk3tLW1g39e2VsGp8X09rauHeB+3And51mwfGfVtZrZsMI5If2PUZWRvRhR8T+LBsEY5rCh9x+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCxOkt2vc9ZNFnlFEOez9nWfw9MlWEq9WakLp/n2nSKsklM7FV/qoydlVr5987fmvrzRs7EO/weafUMNhksqiFr+JABA7F5/STrVh0/QFdPvQMZC/dfqF4dRbJ6YdRjDzAOeTI6HE24diYPwgTvBY+b6x9+KGCXaa2Qpwh1Sk8uYlrnrDy9x642iJoTiIDC2yKtHvrxl4KBuPWO0HZMQy281p35Zthlj87WgxwPOa+bCZuX3CwhwA79owICxouRz2wyCL0/lDTkTEO95IiZfXcDT5dLolfq/xY8EfppvqcUz6AavDmDTROJFI+ewdy3Rna4aELzFZeL6+QHV5xeL4xickIDeNs7bqVjAgLGi5HPbDIIvT+UNORMQ9sRnqdohw/rInvCB4XJTTAWDQJ3KBpIOfoAOLnMoIH62LiTlmATyVMCAsaLkc9sMCLmfIM/UTQBwoQZER5Qwea9CKQlY8TsIdg1suZ9E6/+FUC5JyaHrvXgkDBylGzbDVmaIohTeKh69QIF4Myn71WIIAIds2MSqzpuBjY2VybUj2QowWZ18NQhQaHWyXaE8BYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h4oak6uU6IRXG+n1s+QzRGCUzsVX+qjJ2cFhRLHtr5z2AY7DohsgeLJbslkf323799Xhyp5wRBnnH4XBOP/gst/O1vv0WSUjnCAes/8zYB4fwR+mm+pxTPqtHnTxlMad0alyDWxEiU8Ja9CKQlY8TsI24X1LNvxtz/njf4QVSG0zJw0XpeH2hGtwgI33e8UC9nVkydSh8I56wh05xiYsB13E2a0fTHQJ6yRRWoYm3c8icc7WB6YSrzgCLmfIM/UTQBwoQZER5Qwea9CKQlY8TsI6Sgfx+TritsEkaS2Wtaw7ftncQJK48aeBg57WamN5zNesPyE/IoCsJeg+iExCMrmtHnTxlMad0UGWRiIb9KWh4cMmgMS30D11ZMnUofCOepuhl9Tp+p7Z91OMoqAwSQv0eng9sr0GPyXoPohMQjK5rR508ZTGndGpcg1sRIlPCWvQikJWPE7COkoH8fk64rbBJGktlrWsOwwdk2R1rKY9si/dYyN0cOUgZH/Prfb6w9WZoiiFN4qHr1AgXgzKfvVYggAh2zYxKhG4sbj7Agur8HCdlyZMBoAnD1iWiaJSn6s92FF+IubfkTk+9SxN4FUNfP/1CBud8VW7inPYRzEOJw9YlomiUp95EjyIu+UKAgXulUvuntEbgtH98El+k2k8U3XVh8LZrqpgPjy26nTK86rFGeIZsTbhagTmjDzRSq+HjxaB4B74rR508ZTGndFBlkYiG/SloeHDJoDEt9A9FIjp1DOt+yfCOUNz2J8cyzA7z0L52nuKAi5nyDP1E0C7mVmb2+QTluxjbVPe5ExNnGokgdKcFFOabbQl3mJc96w9aDoVJ6fId4AgF2l+b7H/QiY+QmZbGjA7z0L52nuKIIvT+UNORMRBboDWT8dzI8EkaS2Wtaw7UMVJnXwC3aifAo4nHH+TJ5TOxVf6qMnZI4vTKyHBGc8+7fMKTrRNy1RWHJYQ/HeHQW6A1k/HcyPBJGktlrWsOxojBQdksktfSMqPXgUslBwBYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h0FugNZPx3MjwSRpLZa1rDsMHZNkdaymPbIv3WMjdHDllM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw/m/fPgGiWhA1nKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZeweG/flnonJnT/O9OWBsaTWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPBRnQ4KXnZiDFYMcF+g/n5EC5cX7HhIOjcskGuRzF0LrkEA/9gIkb2ZSaj3fKNwBja1Zni5uVvKw6OyG6bnoLJL7n3mFDlx+KMyy9ofvlbCVlMoCCcErT30372ExX2DzxP5DKhKevgqTMG/erWsTnq8/TnSPPDjO5o+5jTK0ldzHSKnJYuzPGGK5CNUm9ffMjbvA1ZBHXQ+1R/FcXzcC8uthxzW1vQl1A9sRnqdohw/u8urnAR93nky6GUon86Ic9f2PIKNcBb966GG09whqBRLkdqeNxiM/C8qkyybZPDJjHz59ILGVEgxPY/UBscfai+i47LNHaWlyuV0j7hfrI3hbHLiLClnz4tpyoisIJaeLIiYXiAtFkBfqX5RZE0PwrpCgYVS10ee6g18ZZFxsrfmOjc0xlHvOtoBsp4cAhv3RiMMjZy3Mgwb6BlpaooVb1mPJKZ4to+ynvqzdifKM1tDn9W7ccooda/3bzWigGMNmEf31XJNKnei5AyVKShBF+XlGGeQD7iI5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmIy9snkq4jxghNv1qgLuV0Ybv14ozNnq5VMz8s7lE/N0Of1btxyih1t+3BFUyRUa0l2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZ5apJj9XwnyAOnomoLxLlodGypHfWQNvyzMdPeyZg5QvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxxoEDM4VuHcK2Kfzgyku+2yZ/SDtPy6KROZ2MLP56m91/Q3YtcqFzn9fzyeLG5RUgyTR+UIzCD2jV1nSmtbA90OzKeOakhOUTV5gHmKglRiCRx6G6Y3CZNQBCcn4GIYDuoqDp5/6Ofnnjg8yLWpBbekCGgMvrUkxxN+zZPe2/uq5g1MtGwBlMyIjwWvntcuJibmMzJT4Cc27+ctqENnEBKAbGmNFBNoZ4JV9ui98xHoMwwgxUJiDsGag18ZZFxsrfwSRpLZa1rDsaIwUHZLJLX+RI2+DeHKYLrYcHyJR4fckbXl1MfIIIXmS/vNeMNayWL8TLnOCOek6COCDSuabAYYgn5UWLR4Y6miC5eSi0PUbl4X/5vvZUwCQq5T3BDWXyQIaAy+tSTHE37Nk97b+6rmi6syZn5bD0l7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHAY9SJR7MwFUAOcFxSNMQtsEujim6sxPX3ojKMgrgmb89qoHINnqNTQT1zWClEYtH1owyMlfNJgd6fP2fXflSwoFTCo9XIB1AtOsNyE57QpRfmjkoPh4FxgpCbjHIfzrNblg5fuBTrJoLuoa7fVqDjdrKTa8ca0i6qg18ZZFxsrfaPuY0ytJXczO1vv0WSUjnBy1qz6g+LW8pAc/hVAOtpjJUu6i4j6R0SSJw00xaEzAdDNUb3ycDXt+Eapg313n/8BYLB37rmkwIfsv+SkPX9wnD1iWiaJSnwldkCFjwDorZ4xFh1OwKjpagB9uYRlROtHvrxl4KBuPjb9uZP+VgrrbqJEeVd5An5DRDzKAm9d6pAc/hVAOtpjJUu6i4j6R0QDnBcUjTELbBLo4purMT196IyjIK4Jm/GhU56WSokhnwFgsHfuuaTDs5bybePbTw6OW9hn4ekjumc8YxfRIXwMLHlWR+6Hi4VW7ozuVoOLI5resT2VruzSIgMCjrtOs7I2l56GsfE6lwFgsHfuuaTDfm5UNID2G0ybmqPSw9BggPwGopGN5FQ5ws3YfZ2+p/ag18ZZFxsrfkcehumNwmTXEM6dtEg2/A3yrdhzVneuzvzO5g2BtT8ms5Bzkwkt9JWygzl8bwJnt5ySYMBwNUZ2Q0Q8ygJvXeqQHP4VQDraYyVLuouI+kdEDRGU+S2KBe+wcnqbgcQbsrguWLun/rBjAWCwd+65pMII4INK5psBhiCflRYtHhjqaILl5KLQ9RojhdZV0IuFQ4NcRuDkCemG2Wc5osDyA89Wm2BoFmAgSqDXxlkXGyt95iPr6syuvPYtwiQQxAq/5S/wy2EPapNzAWCwd+65pMDW7sCrFExPH7Gfhw9lEZpvG4+SZ6/62xqg18ZZFxsrfrTIP0x/AMDCDPmhAtpi4ZmsezOrWWHiu9orqZYAgHpvG3NjDV3BgyxNha2VNWl81WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNDEsP3aivRx5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmeWqSY/V8J8jZ4JntdtcmueMdUqWV9McPyZ4JHOwzPVry/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTQZhnrV/LA+/iFN34nXB0lH8UnERL5ba7Bw2TEYBX3tTqxiEouaRpssvFfG+fBhu2ssCk5CiXq3flyJNSZWXY3L5W+rEb8XoruEkpZ1EwtkIf0h/5H1vCpqweSSCHUioFSVfbovfMR6DMMIMVCYg7BmAbAWZCTK1uA/XOJfyF1XDY3sCEo28Fct8J/VrU9hea2suxKHYfDbF4SSlnUTC2Qh/SH/kfW8KmrB5JIIdSKgVJV9ui98xHoMwwgxUJiDsGcBYLB37rmkwBAfW+eQstE79+JdC81Y+H25U37/HTypsQvZOoeWO9V/Gqsp9yJLieHEK95r9tEWsCjztA2FYcnwqgHrgP0Ys0NjTutw/wzMvRIoLn9egg/AqVmtebrbNeTBOxsWdPiRLwFgsHfuuaTD/WDiFZb3HScj8E2OMD64IRBmzYCl31FwICS8/dRweScBYLB37rmkwe9nMsBBqXJzTigpD6jq16icPWJaJolKfcbxZexuo4arAWCwd+65pMEXzqeoqfDCheLBEeDGFRu7R768ZeCgbj42/bmT/lYK6aFTnpZKiSGfAWCwd+65pMNgyf6f+E697kez6ymeMObxq5rJdx2fk7ipNh0o/ZvWTu1krzJFXQzM0j9Hpu0C8HtHvrxl4KBuPddPwtGtwIsaoNfGWRcbK33mI+vqzK689qZBGwJbSU13IAIyXWxsyLm8Oxz8TxEynaFTnpZKiSGfAWCwd+65pMNgyf6f+E697kez6ymeMObwaIwUHZLJLX5ff+lhffmvjqelc3ICaMs8/AaikY3kVDuxQILc3cqlTwFgsHfuuaTBF86nqKnwwoXiwRHgxhUbuqORYhzctgv7EGxY4F/U6Okv8MthD2qTcwFgsHfuuaTBI9kKMFmdfDVznD+IVNyZG5SjyIM1enMeX3/pYX35r46npXNyAmjLPtlnOaLA8gPP+yZdJ/bTTIBhrvt/y+YAdeDspfEuZJspAhoDL61JMcUjBpGmAhK5E70Jeje/gCFg4VEE7RIqMX4MqS9j75lvBO05LCnqgWo+X5Um0P+6/oDb9QuSHDNdevasFSgZCszC+cTnAo1owFGIKO/++klhwRvk1cis1RYS7iV9Wgf/ylzokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyA2f5OWNrScHCHTnGJiwHXcTZrR9MdAnrMTJa+vfBrITBJGktlrWsO1DFSZ18At2oSu3dJh+2uVFcF9VXEWYWH8gAjJdbGzIubw7HPxPETKf8Ug8BLyqKN8gAjJdbGzIubw7HPxPETKcZhKx9mlr7aZuhl9Tp+p7Z5SjyIM1enMfkSNvg3hymC8EkaS2Wtaw7DB2TZHWspj3sUCC3N3KpU9q++V6uymFYWuBI0G9+rQ7yJShURQtb/ADKuVfSCivqH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LmmFES8+Cm8cGkhh4DauPmQGCFICShv5G1xg+mXKd5vkWAwRWLohduWwWyFLGq9l95dHXktQENbxD23+ziOLLX21Ukx/l+oXSo4f+2AKQ/RJI9cV2ZZxh2/hkgu1LnWMCAulZItuVyRAfEiPPmAIvbWfWN+YokTjfdg9riVUbWNecFmUMNY9FzR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/X0mFXQGDwUBfxxgLW/DpkietI52dApanS0ZwazF+DSia1Dv3sAhvWmfnNRqgv4UiYRGFaybmRCQWc02j3u+2kOy44C5ZqFQCn5vz96kpWbarmDIzkr822b6s8qwQE970EPDmeXSehvjmJuTaztkfoSNujLFNzqC1TuwfQ5FlmVND5/1YD7AQ+uWC3qjmSkEdAi6bE66DeLahfsP1kIF7KhIXdDSvqLtmnflm2GWPztaDHA85r5sJm5fcLCHADv2jAgLGi5HPbDIIvT+UNORMQ73kiJl9dwNPl0uiV+r/FjwR+mm+pxTPoBq8OYNNE4kUj57B3LdGdrhoQvMVl4vr5AdXnF4vjGJyQgN42ztupWMCAsaLkc9sMgi9P5Q05ExD2xGep2iHD+sie8IHhclNMBYNAncoGkg5+gA4ucyggfrYuJOWYBPJUwICxouRz2wwIuZ8gz9RNAHChBkRHlDB5r0IpCVjxOwh2DWy5n0Tr/4VQLknJoeu9eCQMHKUbNsNWZoiiFN4qHr1AgXgzKfvVYggAh2zYxKrOm4GNjZXJtSPZCjBZnXw1CFBodbJdoTwFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHihqTq5TohFcb6fWz5DNEYJTOxVf6qMnZwWFEse2vnPYBjsOiGyB4sluyWR/fbfv31eHKnnBEGecfhcE4/+Cy387W+/RZJSOcIB6z/zNgHh/BH6ab6nFM+q0edPGUxp3RqXINbESJTwlr0IpCVjxOwjbhfUs2/G3P+eN/hBVIbTMnDRel4faEa3CAjfd7xQL2dWTJ1KHwjnrCHTnGJiwHXcTZrR9MdAnrJFFahibdzyJxztYHphKvOAIuZ8gz9RNAHChBkRHlDB5r0IpCVjxOwjpKB/H5OuK2wSRpLZa1rDt+2dxAkrjxp4GDntZqY3nM16w/IT8igKwl6D6ITEIyua0edPGUxp3RQZZGIhv0paHhwyaAxLfQPXVkydSh8I56m6GX1On6ntn3U4yioDBJC/R6eD2yvQY/SeCdmyU1jT8PsOQj7iMz8mvQikJWPE7COkoH8fk64rbBJGktlrWsOwwdk2R1rKY9si/dYyN0cOWx5cebPGCxzBFrKC0Tmdo5WIIAIds2MSoRuLG4+wILq/BwnZcmTAaAJw9YlomiUp+Be5ChltkEmi5z3aCxXAQqrgZrXgA/9JBzI/wsCS0pMXRTrjGD3MY2EjboyxTc6gvAV/O7+mBoutF2UR5TB5rH86rFGeIZsTb5NgNaBz9I4Gygzl8bwJntloSaBDig42+vh48WgeAe+K0edPGUxp3RqXINbESJTwlr0IpCVjxOwivkwtmFLeT2QG97gxmI8s2boZfU6fqe2eUo8iDNXpzHSMqPXgUslBwBYNAncoGkg5LFaicXcUrcKL4bTgl9GUDYbMNM9q7myBGBl/cpTuL53KSr8CnBu/mx9+KGCXaa2WXsI5auldge3LJBrkcxdC5g/CBO8Fj5vrH34oYJdprZ8FS4hpmCSp4t3RFoJP9wkAPjnNTabYevUWPn5y6uxfw9TfXfn1+z8Kg18ZZFxsrflyJNSZWXY3KTEZDkOVTk3DrcpEHM2I1/nwDziWeYZMyjlAeoYmWTQacnMu1L3SPEs8TuxAbbvii6qnClgm/kvfDb8ejw1EdjL7n3mFDlx+IrISzJ3vGu1uf3+BjnrrDts8TuxAbbvihOfHBU1oPAviwY41BfgizSqDXxlkXGyt9uef7bBxJu0qJeh5N3mxYoNk/hRZZ21vSDVgVGxEJLFspzTMIxSnr12DJ/p/4Tr3u+i47LNHaWlyuV0j7hfrI3hbHLiLClnz4tpyoisIJaeBTocKi3omLwhpxmZtCvVSVaX9ZvoJe6cvhqXJzaLMaOrU2twQqZwVZEGbNgKXfUXJeWqdvtSnOuztb79FklI5zUH4R7DCV4fpGMZSUNb0n05O7zh9Syxi0e9p3K6OuLN2xYNjq+U59gZjySmeLaPsrBJGktlrWsO1DFSZ18At2ob7wggUCVjBns5bybePbTw87W+/RZJSOc3T3qOLnPAV2/3bzWigGMNuzlvJt49tPDo5b2Gfh6SO6ZzxjF9EhfA9Fkk4qMsZDxvuT/A2beRxeGv/s16QMD+iRYufMz54BSK5Pj6mLQwSGoNfGWRcbK35WtQOXMvcI5E/FFlgC8lHwhX+8ZTcMudVoZOiOw4iUmxDOnbRINvwN8q3Yc1Z3rs1q4EdcFYjuQBj1IlHszAVQDRGU+S2KBe+wcnqbgcQbsTJBixh8s/y3jZ9RPG/9z46jkWIc3LYL+rJ7ifHHcmDxDBVGFhn0TYojwWvntcuJiPwGopGN5FQ6/Rq8lGp/drlM2bu+WFHT1H6vHHN4gzovEM6dtEg2/A3yrdhzVneuzuBYISOx1nyWVrUDlzL3COajkWIc3LYL+xBsWOBf1OjoW7uUeBC9iTEf9IYEvNtEtwSRpLZa1rDsMHZNkdaymPY1SkNEqcpXgRQKJqxTIEf9a4EjQb36tDvIlKFRFC1v8AMq5V9IKK+ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwuaYURLz4KbxwaSGHgNq4+ZAYIUgJKG/kbXGD6Zcp3m+RYDBFYuiF25bBbIUsar2X3l0deS1AQ1vEPbf7OI4stfbVSTH+X6hdKjh/7YApD9Ekj1xXZlnGHbLFOWKLFxHuyn6oRC5W3WdGjXSZfx/Vb6VIMPLFspXmrcD8Aw6xwPwwbdIk8JrCDe/VFj6JngMKINX3dpFlTAfTCgwNA5DqFb0WpJUrH6bOgM9CWfn8z6Hs7W+/RZJSOcTE/Lefq2tsuLBsEY5rCh9x+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCxOkt2vc9ZNFnlFEOez9nWfw9MlWEq9WakLp/n2nSKsklM7FV/qoydlVr5987fmvrzRs7EO/weafUMNhksqiFr+JABA7F5/STrVh0/QFdPvQrlgt6o5kpBHQIumxOug3i4hgNZFXKsgxi++Ryg5I4/jZ1hd+V95nkAjqK/Yt6Um0wdfVh7j3o8LQ9YEyzZAeJAz25Ac0HZheKs/Lo8givFfRRK2AynbnX57b4zPPKA4pOKemJYYxr9/CkKMGaZiAxdd4nH42vs1UalGkJ+i79qGimZzjQEhc7VwNT4Su+gmAeIEWMn685D7hJXEyD7bOjVO9d4D4TNSL6mJLQ5OSBi9iH6cJsNrRkFrgSNBvfq0OWs6WJnNpvEwi/t7H9yXqybUncqGOjeCSih+P8o/iH/mx6r4w8EcILCDzcsAxjJBkDB0MFzpdpRjR89G60VdeLryIU39K9JJ7Xe975LCf+7uDEC4acZsbujD3p6qRTDGn127eRuaxTwVgx0wYE6lyM4dhgLV3SWd44sUtH2Qdc583RLKV3VovMYLdPBRpEsVW0dNw7w1CngGZEHpRWf3i41AQcwlmn0BLCOor9i3pSbR8HzEiHkiY9L5/wKSilRz5DPbkBzQdmF4qz8ujyCK8V7YYFH5Onnztoww1tLgy1VcktWWcJGJ5DVuGibQnRaqAl5cNmVcIcNLAbMYyTtB81Z4dOTwQP7uSutJcpVWhHoTWmH0QnDKBilVIIBmEB/f+AEUrsNWzMJPCkKMGaZiAxQHvIXKjGBPsLm7hilQTdnbmQfBzoMgtaXJcC90fsIs2lcxFj+2+tzQOdnVdkll0qSDzcsAxjJBkI1sJXBjhEq4YALFm55Cy1ryIU39K9JJ7Xe975LCf+7uDEC4acZsbujD3p6qRTDGnqbVp/Vbhm851TsUsPm6iUTCfeTM9uG9x4sUtH2Qdc58Ouoxb7ZIcKe9O9cyzyc+00dNw7w1CngGZEHpRWf3i41AQcwlmn0BLCOor9i3pSbToUllVpvk3RCexByKrgu9EDPbkBzQdmF4qz8ujyCK8V7P+OBtpLdcxoww1tLgy1VcktWWcJGJ5DVuGibQnRaqAl5cNmVcIcNJEP98XS3m3N1TLv/vdm2QcGWdvkDp2qjDWmH0QnDKBihcgHd782XmkOjFi3elKSezCkKMGaZiAxQHvIXKjGBPsLm7hilQTdnbmQfBzoMgtaSqfjMxCeS3XDwbn6gg9H1jqqHUMB4nvSgFg0CdygaSDn6ADi5zKCB/yOT/aNSRZb3FfbF/TBriiUzMxN3ZVssAdg1suZ9E6/5uhHwoq8y0TZgJhUdyymnnCCkB/cWqSlpucCMu1RG6Nepwz2FlQUCsa+4JkKGk8XJTOxVf6qMnZwWFEse2vnPbpG4jXwUtOiPEZM0BP048II8v8JpqqcQYS1F+P0jKq1cMd2hdfixOdcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/Exjs5JK/InYnUCoE+R7cwVLSl39KgNurHEcuJ+RvSwZzysUlAo8iA2xHoMmoJRXK2SOt4epHEo6e89mzNgf3y2/3UNnM6eLtwuDhMsVKUw+WGOmg9F0eM8OHGDpqTVyGibWHIFPZElBHbf98+LjC3LZZzmiwPIDzozWXR791Zi9ipQ3jNDYXS8IKQH9xapKW+PXSoq6xkzbbKihHetHdsRvp9bPkM0Rgi0kWLnusckK6maR0RWksW21F32Il+s4U3PQklR7DhT6AdkDIbzwniQcIiTMCV9H8MZPML60V2LXsY21T3uRMTQg2TCPiayVf8momoKYW6Ig6Sgfx+Tritk57CX+OERAHi8jYpW4ftHFluY1BLHaQUWKlDeM0NhdLnRpRErudjt6Pa8hQIu2MdliCACHbNjEqs6bgY2Nlcm2gOdmIOZ5ujGV+ciC9trJaDCIWhhTCDVaioOnn/o5+eWUx5hnADsYsrD1oOhUnp8hO7JRb/x7EOPQAhe/j9717iIDAo67TrOzvnwCxWu6flKw9aDoVJ6fITuyUW/8exDgrmuyD7Mm4h85R7faEOK8e6vSPrYlMVDtbLZa7SqARxMEfppvqcUz6AavDmDTROJFM+L0EvCUbXHFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/1m4YvJ53MUiwR+mm+pxTPqtHnTxlMad0YafmkrDD/Fd4cMmgMS30D2QGNxLYmU7NhjnPh4lsF29MCAsaLkc9sMCLmfIM/UTQLuZWZvb5BOW7GNtU97kTE1HZ9WYTKq9U8LWAtdQboS1j2idcEsQWxrNzaJy93Vs0RfzvLOuA1LyupmkdEVpLFttRd9iJfrOFCuV0j7hfrI3QhQaHWyXaE8BYNAncoGkg+FB0RdhT9Jsxuwnvlth33HO1vv0WSUjnA9BPo42HcXYhqfiesrmPWgl9BK0MsVDTVY1tXzOO1m70Wn0KhqZOKmwUBTkL2d8olY1tXzOO1m7yvSCqDbzX+imbVrC4uDyJbXyY4p3wSQhwvwJH7XcHtcnD1iWiaJSn/d42g6CTnXo7RtZNGyzZJmiHP4+DbUbD7DTMH1pYeVyYc6tyVW9AFrrW/2UQz6Fya6lw5RRYKNdafAXapYNs5viF9Xide6Pi/aRpF30MQ+OfddPh5+IBq5fFCkwlJi+bY7Vcpa3x0Xt+VqsHKyV31TR9Jx8VJPO5ktesC9dZtwl1mJR8yO+TOMbnwqD6OZjkQaxiTNs8MaesefX11P3gmTqwor1v2bSEgGJyIKnSgwq9zmANLO/pMwt/IYHU0jtl03Ptiefzb1PRJKkskFDD1g3V8WVOYGSZxi+QVDl/tcYpmH7SyfPW5VV2yRFNNAe1bCXC0N1chMBRctTYglcKGSTD0HZA0t8reRaK+jVTVin1DSaIrWvd298HzEiHkiY9OmefjRHGgFZDB8DLSd8qcZFeaAI/husB54dOTwQP7uSzCHUZ+c2gb5YguOSuVUdGy/5ixeKIDk0ih+P8o/iH/l2COKGbcKew+n9H2HkN6Wh127eRuaxTwVgx0wYE6lyMyIIFfVzizs4OMKA1BJV2ZO0I436IX4GtKjekj7PLyzlxasqzO+/+s+mYftLJ89blVXbJEU00B7VsJcLQ3VyEwFFy1NiCVwoZJMPQdkDS3yt5For6NVNWKfUNJoita93b+hSWVWm+TdEkxnyX9Ry9hPGVXhpMDkEVsj4juCraZfMlcxFj+2+tzT/BIbpgYV/EBhPdpg7lzno6FJZVab5N0RahHd0l5xhjZhiHD6zFiXVyPiO4Ktpl8yVzEWP7b63NCIIFfVzizs4UaXl6z3PdmRMZ0lgI7F2m2LMsGdYF8G+/QxNMJDc60i80ZOBuPlToAAB4LgJfBifbkDvGpU7n2GOZSgChCE4twePxLG2o3WYXJiFjy+Rl6hoMcDzmvmwmZ7q/YtCGrHjD/XfrYjohNyrVs3e8Ho22QCGN6OvDnnfDB8DLSd8qcZO9wCLXegEbW/78RTI7wwQNYuQn2dDgkv6KaXfbhyt5DndaYzgM1dvNzsef3WTV7qwazyVpQizNU3f5glWk8xyhYpYGyxjb0KYYhw+sxYl1X39UlipstLL9TJH5edPkyWAPeXNQ8AQrB4FDevtDiVU+ZiKT0jJRQu60Os6y0eYhvCLlv6ah2eUzc2icvd1bNHavFdz3pmbF9CV7yFXiMmkU5vxeJL2a6p52q2LL6b32V5rWeBxOwLWGq/Ze9PU2kdm6N03kOe76YA95c1DwBCsHgUN6+0OJVQUiOnUM637J+EE5k82EFMYHKEKG9O+lS7CCkB/cWqSlhSI6dQzrfsnxN4slmapfj6wOsBc4HaQqJ0aURK7nY7ej2vIUCLtjHZYggAh2zYxKvJMoiRRwIwdYaIkjItxTX6lqmFVgZ1MPq+HjxaB4B74rR508ZTGndGpcg1sRIlPCWvQikJWPE7CK+TC2YUt5PbhKsp+f+SqUvYMAb28qXNflM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCXAV1p2bf4sLPc0I368GozilaqHQ6HYhZedK/+s2YPEJ0CLpsTroN4sr/woLldCAyDwd97glPYLJnRpRErudjt6lr9eQQZ3jNxxHLifkb0sGhVUg9RSnF7TH/0E3uDgJytHvrxl4KBuPo4ORZXvKFCKUzsVX+qjJ2Z0TyUy/Al6LeHitvgWQiBKyfJP0mpuVkaRxskdtCCx90LQQDfTTMUQNAvY4w9le2M6MQApuBRE7MFN9ua4dqTc44KuW0tEdOm1F32Il+s4U2wPHIWOU7dwP9d+tiOiE3OBHGN2nvuNhAWDQJ3KBpIOSxWonF3FK3GfLjE3KFHis1VHlGPR2qr85XbGukr+cOuxjbVPe5ExNKcFDnmYTcQHH/0E3uDgJytHvrxl4KBuP1XgPaO0Wi4rNzaJy93Vs0RfzvLOuA1LyupmkdEVpLFttRd9iJfrOFNsDxyFjlO3cD/XfrYjohNx9rMO+sJK4viG+kpyK5fDDIk9TBT5AZSRPzSDeEkB8GO4hj4WKLxruWIIAIds2MSryTKIkUcCMHXh4rb4FkIgScij4eRVyAumEHKK/IN9j4Xr8dNEVzMoBFAJnLkgoECP9nzC7v1nHd0c5WGRlNKj6QeNlthsd/EfC4OEyxUpTD+dK/+s2YPEJw19njuDvH2QBvITLBMC2tpNA/lE5ubxrr6XAk0olsDge0pn32vN1miXoFeEwmnw1FXNBKZaZmVIcRy4n5G9LBoVVIPUUpxe0x/9BN7g4Ccph03anErX50Jz7681AJDFtfLTDrNY9w1j9rDa4Sx3haGfLjE3KFHis1VHlGPR2qr85XbGukr+cOuxjbVPe5ExNnGokgdKcFFOW8SCRDJSOGxj+FmzHJW3ZXslGlDKq0rZw3LSn03UDPvXzClMVnPUWsJcLQ3VyEwFFy1NiCVwoZNhBgqonNW5qa9CKQlY8TsIr5MLZhS3k9kPvduJuB2FTi3hQ1IL/NyPSeiz8JRNVSJtc8GpGHxkV1ZmiKIU3iodeO3r38NXwdf2fMLu/Wcd3RzlYZGU0qPpB42W2Gx38R8Lg4TLFSlMP50r/6zZg8Qmp6VzcgJoyzxI26MsU3OoLsE/F/6F8TZWsPWg6FSenyOpt2ZyhBio8HtKZ99rzdZol6BXhMJp8NRVzQSmWmZlSHEcuJ+RvSwaFVSD1FKcXtMb2a3wBSeOcto5BnAspnvEGGCY8M4nxuMD1cZawoc90nRpRErudjt7iWWJBHoCpYo5lKAKEITi3B4/EsbajdZjU0kQkWpcrWuHDJoDEt9A9FIjp1DOt+yelEQYVtBkl7dD6SFeltyPgu/wiTmQa0p6vpcCTSiWwOB7Smffa83WaJegV4TCafDUVc0EplpmZUhxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnJHseTWJFtJxy94DfxPvFWZCvMHWP83Q8QQByd1zd5WqsJcLQ3VyEwFFy1NiCVwoZNhBgqonNW5qa9CKQlY8TsIr5MLZhS3k9jiKSJIBlKJOXS3eknAq/xtq5rJdx2fk7hB+VaJBV3EISX1eYZ5oBk1D7yxSCyuYmNVY6EBF6bWDcZinTM8Sur0w0mP3skyStFRWHJYQ/HeHQW6A1k/HcyPBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDr9lBFkrMs5/6+HjxaB4B74rR508ZTGndEiMvY6Q2mATs6MQApuBRE7MFN9ua4dqTc44KuW0tEdOm1F32Il+s4UpyenXn87dN3MU4UVpv+iFFpoAb+70/qtPBRehIFeP5A1g6d7E5M1YmOvvVYKodJrZ8uMTcoUeKzVUeUY9Haqvzldsa6Sv5w67GNtU97kTE2caiSB0pwUU8nghxtgSf/dyOx1wHbn2pcSNujLFNzqC6u4Oe4qWCLJIC9l62eevMzNzaJy93Vs0dq8V3PemZsXsJcLQ3VyEwFFy1NiCVwoZNhBgqonNW5qa9CKQlY8TsIr5MLZhS3k9jiKSJIBlKJOXS3eknAq/xvq1ME5GgnNCRsagWqG1rRmcvnkfeUTU9SwlwtDdXITAUXLU2IJXChk2EGCqic1bmpr0IpCVjxOwivkwtmFLeT2OIpIkgGUok5soM5fG8CZ7UcmUejfS7U0gwY6DoEkbIN1YKbw3tpRShxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnMQzp20SDb8DfKt2HNWd67PLRMRh4COuW564K/wQvn7OTkGSJu/s69jC4OEyxUpTD+dK/+s2YPEJqelc3ICaMs+2Wc5osDyA85YTxDsJ4TeBIXPT22KgGxYRaygtE5naOViCACHbNjEq8kyiJFHAjB3u0V+ntFmUQQNEZT5LYoF77ByepuBxBuzLRMRh4COuW564K/wQvn7OTkGSJu/s69jC4OEyxUpTD2nwF2qWDbObuxqzJmOoTNGWDiOzQ76WJCFxvwzLWr+n0GaT9Geh3N1lyJ/wR/kzpycPWJaJolKfJlVY4v7eh3ToJn7x5wSUwJzvYl3hDcdLunFppJC6tyycCepFjS3OmdAi6bE66DeLWASWAIiDjww/G8MS9PnKJIG2zufW9P1rbMIOY/UGBGcYKYvSvC3NekNqfLrFo1S0A+Oc1Npth690T/hMTF3EPygt4LMVYyCGieOJLs8eaqrHJt0jCwEnmbWuptDHGlcHSxsgrKJQ93C/BE6xYdQGmHFRSNmbJEr2x3NEmM5ATahxUUjZmyRK9r/dvNaKAYw2NQVM3MMPDzQ3V8WVOYGSZ2OKzqjfS+L0JSOB5TEcRGwl+o9tVuEAMngcf74frgB55S7VhRRSwLjib9EZFcK1poofj/KP4h/52X232+bN80nXbt5G5rFPBWDHTBgTqXIz/wSG6YGFfxAQrhvVTDYoK4Qcor8g32PhVfgPmkoctkHxdcCSAV0m5TdXxZU5gZJnHZLfJEkuMDioNfGWRcbK3+iL0XHn2AGrnh05PBA/u5JZ+7778PWMpi/5ixeKIDk0ih+P8o/iH/n8OQW0PfoyysnBWy1qRVDiBH5d5Nb5sfmOMtjdMSAckdUqsUUNv80Y0gmGylV8dZlaiDSZ909GE+Uu1YUUUsC40aDZa8pdxpCg+rx1i9cEOKyoIuqkNvzn6FJZVab5N0SMm1vl7CFg0k+QkrjEq/Gwcij4eRVyAumEHKK/IN9j4ZuhE7RCxKJELWcgwekdLnEa/9EEFAyBeag18ZZFxsrfWw046j9A4ZopU/nnc0r0rk+p6KubcHQVqbVp/Vbhm85wR4EH4t53KWkjwuV23KD8Ld0RaCT/cJAD45zU2m2Hr1Fj5+cursX8PU31359fs/CoNfGWRcbK35ciTUmVl2NykxGQ5DlU5Nw63KRBzNiNf58A84lnmGTMZ0APQXN6eP2z9851P7X761CCcmaBVJKelXeHI7I2QVs1epxaUq4HuL3bzv+4iPWpBUpe48G8Uie/+XIFVxUdrQH9bAy+mJtKRvgfyGsBOHgWzGQMJTUEZaYzax1MSndms8TuxAbbvig/AaikY3kVDhSt7apcRCOK0BiPpbsi2bpC0IYX5CECeur8HUmQVc97hbTaIcVNlmRy5MK0fr/EkmDUy0bAGUzItlnOaLA8gPPFQoAxFr0R+W1WnmoxFkAxIpwhbRLiR7ieyZFt++6kEdz0JJUew4U+X6maz8Mf8VxtVp5qMRZAMdD7nyce3oCGYNTLRsAZTMi2Wc5osDyA80Aop8gQS747tlnOaLA8gPP/HNN5W3do94LF9nAZbW1Ml6r3CSjbOX6B5vN6lMor7M7W+/RZJSOcQECr9go5854nD1iWiaJSn6e1SpNNt9qkZjySmeLaPspzUTVDaWp20Tp2J9kSzb9qvaZQvnMsg2EadyxsJyh3lag18ZZFxsrfz/8OLwI9o17Y4QQJqbO87iqTZPV2VoXJkg1GqmGzqDYr6UhuhHB4P3D3DMUc/da/lDjcrSCMxzFGsh9bzCKSx+6gnuh/ZnB596RMIaTRtG+DJR3lARC8EF0dI7cCxkywpcJf/1ZBiW0P9d+tiOiE3LNppDBVzKAyZjySmeLaPsrmapvu8GTtFeJv0RkVwrWmKFBN76mDcskugNuttMl1fPnRJNVYG6w5A9dE52dTkJYr6UhuhHB4P3D3DMUc/da/0aDZa8pdxpCg+rx1i9cEOMnQloDIKK4JXm6MfsYWaQcpU/nnc0r0rrB9mdwKcpOwZjySmeLaPsrmapvu8GTtFeJv0RkVwrWmmzex8mhFdxougNuttMl1fPnRJNVYG6w5hD/C9tAnC3Qr6UhuhHB4P3D3DMUc/da/0aDZa8pdxpCg+rx1i9cEOD4Ri9crbmFAXm6MfsYWaQcpU/nnc0r0rnai66J660EJZjySmeLaPsrI7HXAdufal4KLY1BA6bZNV65xPiNw594ugNuttMl1fPjigiH2ZjOY2AtciUXIvXkr6UhuhHB4P3D3DMUc/da/djhLaH2iFg7bzi48hZGtVcnQloDIKK4Jwtf3wrqbKBQPWqujAYVGFP2aJGFV3NlpZjySmeLaPsrI7HXAdufal4KLY1BA6bZNteLxNCsLfYougNuttMl1fPjigiH2ZjOYYJbkOrQdkPMr6UhuhHB4P3D3DMUc/da/djhLaH2iFg7bzi48hZGtVT4Ri9crbmFAwtf3wrqbKBQPWqujAYVGFGEQaDGu3LvFZjySmeLaPsrmapvu8GTtFb3DQeqZhZgz67vPMVHJjCkmbcuBnPkW5SKxJWMbtP+K4g6XAIaM8hioQPXDgYLHx2Y8kpni2j7K5mqb7vBk7RW9w0HqmYWYMxjo7G2zTl3RJm3LgZz5FuUisSVjG7T/iuIOlwCGjPIYDdRmmnX9NtJmPJKZ4to+yuZqm+7wZO0VvcNB6pmFmDNgUakQQCIo4SZty4Gc+RblIrElYxu0/4riDpcAhozyGPjR9GAgWVvSZjySmeLaPsrmapvu8GTtFb3DQeqZhZgzttx7FG7rgLUmbcuBnPkW5SKxJWMbtP+K4g6XAIaM8hgSjMzO3mSihWY8kpni2j7KTnsJf44REAdUVGGFf1TOxTmXVBfK4hJZ6H/pG1S+2BXzlo93ttcu55z7681AJDFtM+d9VQNM0QuoNfGWRcbK3xozPPagAPwhoXkxk8xDEg8VC151hm95SFhzrN3cXobJa+7pNWkiA8C9w0HqmYWYM8G/DPgYyWI8K+lIboRweD9w9wzFHP3Wvxj+FmzHJW3ZXslGlDKq0rbWNWMGXryoGpKo6qB5+p5fLDw1gsxVpXifsyT7eXUhjfekTCGk0bRvgyUd5QEQvBAB0rdEwIGjwTToHlm2V76QdwrrbERPHvneAnkkG3cpnk0GzO2DLZQ24g6XAIaM8hgSjMzO3mSihWY8kpni2j7KjmUoAoQhOLe9w0HqmYWYM0scqvz2kvPHXOIfOx19r32/yRcdIlPKOF9n59S+kdLXPhNrs29cLVyoNfGWRcbK39o9YIVSylI62dMFU3EPcMtfEu3owUhm+PEZGxamF3wBTnsJf44REAeLyNilbh+0cXEHM4QD7mjxK+lIboRweD9w9wzFHP3Wv7g1hZkLesILJL5Fy/Yqac6LjDNuryK+GXTdGv7jL5CeDJp/pQZKDeJxCbuKBT0CTvekTCGk0bRvgyUd5QEQvBCN2p7PwrYmODlcf7Xe28zEN//SSiT+uscmbcuBnPkW5TVeXi0DFZS+tUuDEvz2ZIIo00iRIc+N/0Te3KALTTmkaAucyglImfKoNfGWRcbK3wwiFoYUwg1WoqDp5/6OfnniY6/zAGiYviSJw00xaEzAZd/yTly2zIJauBHXBWI7kH66FIYjonHObmMzJT4Cc27+ctqENnEBKD+XRXK82DJ0QDmp5qMwprkGGCY8M4nxuDvrS6VLqEMHsYlB5QV0/PCKzno9CbS6ZZjcmMTr7dw49aoR2gafujfTfvYTFfYPPMIdOcYmLAddxNmtH0x0CetNrztQyWMZVuB4LDznFf8q0e+vGXgoG4+b65afJWPMNxew4YYQevj+5qBEytoYnUYkicNNMWhMwGXf8k5ctsyCxyGXcS2GWl7BJGktlrWsO1DFSZ18At2o8Hy9I/URyxm/3bzWigGMNtmzID3ndQXqztb79FklI5zdPeo4uc8BXZ9akvex6qX5AEJyfgYhgO6ioOnn/o5+eX/LWRejNmiYs8TuxAbbviiI8Fr57XLiYhI26MsU3OoLuA4w2eAvm+KbvgjOrX4mnScPWJaJolKfCV2QIWPAOiuJ3z8IcZPX7dN+9hMV9g88DdJlmaglNx8UI1qInkMjLFbXzN4KgbBMHlpQ9GLg1X3BJGktlrWsO10ZgVxXJY21ldaA3MM7bhioNfGWRcbK39D0jPoHAd0i9OEnJcUFJpVkxQ+S5XqJkYJ21nAmxqHjnUDnH/Z9p7CjlvYZ+HpI7tVumz2A9tWGo22LrPJSog7moETK2hidRgDnBcUjTELbBLo4purMT196IyjIK4Jm/J9akvex6qX5to5BnAspnvEGGCY8M4nxuDxoUHU4zF3xL7n3mFDlx+LBJGktlrWsO37Z3ECSuPGngYOe1mpjeczpse661rgrPKnpXNyAmjLP5qr7N0RfswIZtfdKdtWR6b/dvNaKAYw22bMgPed1BepwG3LBXMR64cCRFbjeoE9Bm74Izq1+Jp3VmGGCjzYLNRP2XjZRKC+vF7DhhhB6+P7moETK2hidRkRjFHOI4tJc+JjqRdkszjlcHBGCgN2fU1Lmp3lPgRYv8EsjfGHwQ4W7bhuOJgVUj9N+9hMV9g88GaSFRmu4bnh+lEs+bXF73FL16ZTemMj7wSRpLZa1rDsYpvJFpyu2Qsq0xlHe7Gdrs8TuxAbbviiI8Fr57XLiYjp0B37HjdVtcJXQCKOgLXbgeCw85xX/KtD6SFeltyPgSYewBNcyWO6/3bzWigGMNtmzID3ndQXqOS2bMRXLafiImZoORXXgsRsUVFiaUZmM5c53VVWpRXBblxhN7uaZ/NCptC7KY+qD0372ExX2DzyoTXC84ul14Z7+ehYbqhzmqsZksc8FV8yp6VzcgJoyzy8jKhI7hEwpOvnqAzq55s6/3bzWigGMNtmzID3ndQXqOS2bMRXLafiImZoORXXgsS07SZiCkrBK5c53VVWpRXBblxhN7uaZ/KYpXmMJbs230372ExX2DzyoTXC84ul14Z7+ehYbqhzmynnnnDdutt+p6VzcgJoyzy8jKhI7hEwpSYewBNcyWO6/3bzWigGMNtmzID3ndQXqXS3eknAq/xtq5rJdx2fk7sN/AaPOJhdkA0r/wpDl56b49sHv18Hvs4Qcor8g32PhMriQusSU8tXhuIxkA+nXs9N+9hMV9g88zFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QhToi7N3L6cebvgjOrX4mncjsdcB259qXEjboyxTc6guWJR3wf86mc1b7lQsvEPggs8TuxAbbviiI8Fr57XLiYqjekj7PLyzlIdWHn/tImo3BMiQUSEgOwp1A5x/2faewXS3eknAq/xtq5rJdx2fk7gN77a8J79cBF7DhhhB6+P7moETK2hidRvj2we/Xwe+zhByivyDfY+E1h6BSAlng+ev0mOS1Mikc4HgsPOcV/yoBgEF9iKWsJqShZNjR8iw5YiNLZVTeRvPc3PVmIdA7btN+9hMV9g88zFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QefSDKMKaSJip6VzcgJoyz6jekj7PLyzlIdWHn/tImo0oARQ3vGeKNL/dvNaKAYw22bMgPed1BepdLd6ScCr/G2rmsl3HZ+Tu4Sbk8sMeY9qGgTiL5XJ6z8EkaS2Wtaw74m/RGRXCtaZafD/+ALxcOljkoRbCtXm9o22LrPJSog7moETK2hidRvj2we/Xwe+zhByivyDfY+H7p41DTv9XJVqfcSqHhFX8zFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QdvYmcQLH37mzxO7EBtu+KIjwWvntcuJiqN6SPs8vLOUh1Yef+0iajfynYmlTs0SdJWCJ+bS/rxPzkgYjmawpSilT+edzSvSuo8ExgfrwoND9dbI6EhB4E7/dvNaKAYw22bMgPed1BepdLd6ScCr/G2rmsl3HZ+Tu9IsVOoq1jUoDSv/CkOXnpvj2we/Xwe+zhByivyDfY+EyuJC6xJTy1bTIR5HcsFfa0372ExX2DzzMU4UVpv+iFFpoAb+70/qtPBRehIFeP5A+rTKOcwEyiZu+CM6tfiadyOx1wHbn2pcSNujLFNzqC5YlHfB/zqZzjEHRYwBDgHmzxO7EBtu+KIjwWvntcuJiqN6SPs8vLOUh1Yef+0iajdfAXFT6NDK2nUDnH/Z9p7BdLd6ScCr/G2rmsl3HZ+TuA3vtrwnv1wFrnrPtxDHxGOagRMraGJ1G+PbB79fB77OEHKK/IN9j4bB+j6H/PJS86/SY5LUyKRzgeCw85xX/KgGAQX2IpawmpKFk2NHyLDliI0tlVN5G82BG9ubztjpy0372ExX2DzzMU4UVpv+iFFpoAb+70/qtPBRehIFeP5DPtY2mfAlLnqnpXNyAmjLPqN6SPs8vLOUh1Yef+0iajSwyPKCUOXjwv9281ooBjDbZsyA953UF6l0t3pJwKv8bauayXcdn5O7PueGq0Z7il4aBOIvlcnrPwSRpLZa1rDvib9EZFcK1plp8P/4AvFw6WOShFsK1eb1dBi8ahMoUJeagRMraGJ1G+PbB79fB77OEHKK/IN9j4TI+iCSmW2b1Wp9xKoeEVfzMU4UVpv+iFFpoAb+70/qtPBRehIFeP5CeMM6VNn4/97PE7sQG274oiPBa+e1y4mKo3pI+zy8s5SHVh5/7SJqN302IdSH7Uv0lYIn5tL+vE/OSBiOZrClKKVP553NK9K6jwTGB+vCg0Bni0MK1vMvfv9281ooBjDbZsyA953UF6l0t3pJwKv8b6tTBORoJzQk/jBupACPSs6npXNyAmjLPqN6SPs8vLOWKRO9tjjAS+Nzc9WYh0Dtu0372ExX2DzzMU4UVpv+iFFpoAb+70/qt9Vn3Bt96V/1b9NcEpVQwPfj2we/Xwe+zhByivyDfY+GKtuXTM6+LKr/dvNaKAYw22bMgPed1BepdLd6ScCr/G+rUwTkaCc0J7W0fD8hWIxGp6VzcgJoyz6jekj7PLyzlikTvbY4wEvhgRvbm87Y6ctN+9hMV9g88zFOFFab/ohRaaAG/u9P6rfVZ9wbfelf9kn+588BSThr49sHv18Hvs4Qcor8g32PhXK+hUwMhxAy/3bzWigGMNtmzID3ndQXqbKDOXxvAme1HJlHo30u1NPvGlyy9XUBGxDOnbRINvwN8q3Yc1Z3rs0pIZmZpsMAhL7n3mFDlx+LBJGktlrWsOxojBQdksktfm28FWLD6GP+dQOcf9n2nsGygzl8bwJntRyZR6N9LtTTwXT4A2AnSw+agRMraGJ1GA0RlPktigXvsHJ6m4HEG7KalkM7yHxFmqelc3ICaMs+2Wc5osDyA85YTxDsJ4TeBiJP9+dI2nl/BTpSqg6TMKMgAjJdbGzIuWJ7/LE7Dk+iqfAtLY6eGvcEkaS2Wtaw7DB2TZHWspj3tSdBKbbWyQEC8OIornqDiGjM89qAA/CEMmn+lBkoN4nEJu4oFPQJOZQL/oMAG4rI1Xl4tAxWUvrVLgxL89mSCcOM9LbLRcpAZiCCGOFXW6yreBqO2mrOeK7v8TeBT4K3cskGuRzF0Lg+Gs8cao2oYPJ4+RyNocYHdKnc/75K1rKPrf0CC1QVuj+K97Q/MpF9BrZawyDg53+oq3t2cELoXV3ThbjCmjuR9/VJYqbLSy2bo3TeQ57vpgD3lzUPAEKxjhrsRW0Xh8+Uu1YUUUsC4hX9l0fm8U4VXdOFuMKaO5H39UlipstLL9TJH5edPkyWAPeXNQ8AQrBlmfcHmfdp72tWZ4ublbysOjshum56CyS+595hQ5cfihcv+0GNHQXI3TTckh4etg+dQJe3e58jCDwbn6gg9H1jZ3G1z13uk5Gf52OwzgI9ts8TuxAbbviiOvroGNV3EmEz2f6eex8n9oQpAMATGjcohbxV3AF2ZFtN+9hMV9g88oSfncoHHiH4ffdSuUY3eUAIEa+1M42FMqDXxlkXGyt+20VeWcjSa+IaELzFZeL6+QHV5xeL4xifX9aRAVbJI9dinGeNkVH4E5o94szA1qLuzxO7EBtu+KF2rl2PEELc7G4jp3h8J04jcaUoX8x86ri+595hQ5cfiS2mR7DTFg0yuhhtPcIagUS5HanjcYjPwRbI5MTZTA1xWW3LJDaclYBWme4zwVejCMMhEA1p0AaOoNfGWRcbK3/539MkHDITCnUyy6YcmI8RLTpAqdXgC+VTszs8iePtfd3/YqMorY/pdEuMAhwI2YeZayS/+pXGLiJP9+dI2nl/8AHUmsrXqVx/lW72eqcDi0fI81agyzrGB5vN6lMor7KioecrDQoAy1jPO+7s8jK/JEKU4QhXiLIHm83qUyivsTTib+DQieApUSO5DZHH5Riwt+ugE7hVKYNTLRsAZTMj05bZ6Zmo/f3vqzdifKM1tCSIDT+JAzFO/3bzWigGMNmETpzZc2/VMlvAmEYi0AhLTo69b5g0SgJpb1tIBC0VVs8TuxAbbvij05bZ6Zmo/f51MsumHJiPEuOjSDrviT6w2T+FFlnbW9EWyOTE2UwNcIoYxmfYA5WpCmbSxslgqltjDxy6ReLZik5tHNIzRxCwnD1iWiaJSn4F7kKGW2QSadLYrCn4++jjwcJ2XJkwGgI5ibk2s7ZH6EjboyxTc6gvAV/O7+mBouvQElGAQng4bLd0RaCT/cJAD45zU2m2Hr1Fj5+cursX8PU31359fs/CoNfGWRcbK35ciTUmVl2NykxGQ5DlU5Nw63KRBzNiNf58A84lnmGTMo5QHqGJlk0GnJzLtS90jxLPE7sQG274ouqpwpYJv5L3hAcO6G5IPMJheVxIlN1kTsffihgl2mtkHrOB+WKftPDLfOCduQDKyvKpMsm2Twybv4KVLFCXqhNoy/XBfDCQeqDXxlkXGyt/cxy4lNByLKaAQJUTq4jM6AjdJ0MTSjNbZKyAna4xzwjlewXUoPBy8hvsRWHNpsjC+i47LNHaWl3vZzLAQalycyOO9ITgLdD/R768ZeCgbj7ZmjHDNp2DBqDXxlkXGyt/NVaB58sH37UWy6sQtA6V7vXCs8C1s9IqIk/350jaeX3lqkmP1fCfIrDpW/ay1R5/kx6dJJwY9BnyA/Cw3lzwqMpcev8pQg+zH7B0bn4S9DiZty4Gc+RblRBmzYCl31FyeyZFt++6kEeUXWaUTU3wN4xEvRHxsgCiYrPJ13IAZWbK4DtNfECHfBj1IlHszAVQkicNNMWhMwGXf8k5ctsyCOWkn1mupLPsAQnJ+BiGA7qKg6ef+jn55NRjP9Z260P2xQlg3pveBe7aOQZwLKZ7xMA6OixUw6rRBUf+h5bl0Qo5BonJZZYOiAOcFxSNMQtu/0F0CLjsHHIBKh+Dvf72/XBfVVxFmFh/IAIyXWxsyLm8Oxz8TxEynm74Izq1+Jp3IAIyXWxsyLm8Oxz8TxEynUHLSet2GzjexQlg3pveBe8Qzp20SDb8DjmenhxlvRnjUaZEGNKkA25uhl9Tp+p7Z5SjyIM1enMeEyb4ko77PQ/Vx9YCrqc3Wm6GX1On6ntn3U4yioDBJC2qtoMUtTNPcNDrz/dM09R4aYzfjTC6+kRadgV3/8ZHoxDOnbRINvwOOZ6eHGW9GeGqtoMUtTNPcNDrz/dM09R4aYzfjTC6+kUC8OIornqDihiD2MFpMCzQLXixMv2stQOAZ2a7dXuH6MO1bv9UEx+1GxIE2JFK3ZS/SJds6FEw1T80g3hJAfBjuIY+Fii8a7mUNpLBUAVv7WRqf3NAPJQZycrCMUqm+FxkewXbZtiYycij4eRVyAumEHKK/IN9j4Yx1ndaINLPZj6GcPLJb1P6xHXReuN0pRL2mUL5zLINh40HwhHQp/DoLfWXEKHgzLT8bwxL0+cokgbbO59b0/WsLXixMv2stQAMX+GNx09+7wFgsHfuuaTCj639AgtUFbo/ive0PzKRfwFgsHfuuaTA1BUzcww8PNDdXxZU5gZJnJ5/3kYU/UsVEkqSyQUMPWDdXxZU5gZJn+UJxygjglB2kpXQ2AbQsVBgAsWbnkLLWvIhTf0r0knvEzFRE0ET4LHyA/Cw3lzwqDqFeXIjVfUOP4r3tD8ykX8BYLB37rmkwUWPn5y6uxfw9TfXfn1+z8Kg18ZZFxsrfKqLBu3yOMdp+Konn04o6AB8gtxiLTTHiB7N50MLSGKtEiguf16CD8KOUB6hiZZNBpycy7UvdI8QYa77f8vmAHZZruN9kNGOk06OvW+YNEoAE05v+Y2j2qmLMsGdYF8G+/QxNMJDc60iC3dJHqUQJO7/dvNaKAYw2vKpMsm2Twybv4KVLFCXqhNoy/XBfDCQeqDXxlkXGyt9f2PIKNcBb97sHEWsuDrnZdKqv2TzOuH8Ya77f8vmAHdkrICdrjHPCOV7BdSg8HLyG+xFYc2myML6Ljss0dpaXZjySmeLaPsqdTLLphyYjxBhYmoNdd33ypNl2Y1QdyI2SZ2KQNe8fTcBYLB37rmkwdUxkXl+Y/lAqk2T1dlaFydB5qlrIavmx8jHUuAsZ7HHAWCwd+65pMAGOw6IbIHiyW7JZH99t+/fV4cqecEQZ5xhrvt/y+YAdfroUhiOicc7uoJ7of2ZweSZty4Gc+Rbl6v/pubIgulBudwpRJStzj2LuZjFfRZ6kcHRL0af5IwGo3pI+zy8s5Z6UfLmTIsXYYLkXeRIMPlWo3pI+zy8s5f4vCzo7OmVVGJQkVdzgUcTjKIp8U6MtZcBYLB37rmkw7UaAb8Cd6MPTi7+sobmlE8Z50MirKYEM3h/L7CuRxlfTi7+sobmlE/VMKjyMdEa731D7mhcnSaRvRvZllj142Bhrvt/y+YAdfroUhiOicc7Ak7Kki5NUpl7JRpQyqtK2dLJAdWC5kppLpBIMBZaBqDToHlm2V76QWLV4z/KBWpsYlCRV3OBRxOMoinxToy1lwFgsHfuuaTAdro/YE+cGjk0GzO2DLZQ24g6XAIaM8hg3gRrBM8WwsAHSt0TAgaPBNOgeWbZXvpBYtXjP8oFamxiUJFXc4FHE4yiKfFOjLWXAWCwd+65pMPTT+tHNEkYQRnk7RsJSIrnXUAxLKr8IiwhTBvOkeoUqa+7pNWkiA8AiYgpI24Kok4yr9CVEQsIAv9281ooBjDaRjGUlDW9J9OTu84fUssYtHvadyujrizdsWDY6vlOfYMBYLB37rmkwXBfVVxFmFh/VmGGCjzYLNeRqJv7C0M+wnUDnH/Z9p7BwG3LBXMR64W8b1fRALXv9K+lIboRweD9mPJKZ4to+ysEkaS2Wtaw7CmSzK+vxonKnsCtZxsN3yMEkaS2Wtaw7CmSzK+vxonLW6sLKKFp5U6g18ZZFxsrfsUJYN6b3gXuhiWHG0TehoZLFsfdigeEodJ3YXRnViWwbVtTey9i1nGd5bEFp01puHZ+zDsJNA3ZS+4j3QfMqEzFtSD/oT5P8dflakqN+CvsYa77f8vmAHQY9SJR7MwFU+PbB79fB77OEHKK/IN9j4TK4kLrElPLVA0r/wpDl56b49sHv18Hvs4Qcor8g32PhMriQusSU8tVVKNcQPx/WQsBYLB37rmkw7OW8m3j208NdLd6ScCr/G2rmsl3HZ+TuWW/4dBdYxiIlYIn5tL+vE/OSBiOZrClKKVP553NK9K6jwTGB+vCg0ErPziaX0exSv9281ooBjDaDVgVGxEJLFsxThRWm/6IUWmgBv7vT+q08FF6EgV4/kFqfcSqHhFX8zFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QVA93oL05NlAYa77f8vmAHQY9SJR7MwFU+PbB79fB77OEHKK/IN9j4SoQc0pwkOGbXNJuUrHz0jzBJGktlrWsO+Jv0RkVwrWmWnw//gC8XDrg8MxZ7cKwom53ClElK3OPOvzm46oTw3GI8Fr57XLiYqjekj7PLyzlikTvbY4wEvgbcNzpKwLX1Pj2we/Xwe+zhByivyDfY+EotmZGFL4eU7Om4GNjZXJtQmYYXfngN8oBF5x/e4AMjXdDWff4sP2OAoHnaArgPt120QnqtGlOZLaNbDMil5XTOqbyDCZjC/oEfl3k1vmx+feAD79+ivGmjriYL1OXFoZlDaSwVAFb+6g18ZZFxsrfmtJYAprcY+KW3J1Cbc1Ieun7yTUhBQDieb4k4i+3XNSZrZx7SJki4hezEX+45eHjwxNh6hxU3Refha+Ff/1Yd2aoaHqckevDibUDgDdIncjg58T+baN4J154Ce/HkQvFl9WcS3HRv6SFf1lN6qbqa+2d+iBc8v0FHyC3GItNMeIi/tUNmUvb5SfMwToEKp96qDXxlkXGyt9yErauFowuZk/kMqEp6+Cp4YUHeRv16uTmIqollrQmavdUASG/wB2qWc0gvZzBA3Q2RPNnJNz0by9nAOXMoiDE7Gfhw9lEZpuSd3s1ClEDb2bN+cK+lOT1uF0OMqX8TPtwRVC+ZmzhmHEK95r9tEWswFgsHfuuaTC9plC+cyyDYWlWiHyrgMLnUn7vOTOrLz+46nwRN+G67A/1362I6ITch+scPhRacN65QhknzOiP9rOm4GNjZXJtvasFSgZCszDjdhVjvvgpIQ6OiSF92RA4TMzqNaAeQE1OWrilswXNRH2GK9U0xZSOG3ynRfQJ0PYP9d+tiOiE3LHpjTru+7rFRKf2+Y4zEZhs/P9zr8kn/aI9EAkCE4YeElqjsKdbEtlEYxRziOLSXPiY6kXZLM45poh/rkOrnydAhoDL61JMcTfs2T3tv7quVVtw4ikZM8KoTXC84ul14Z7+ehYbqhzm/zwVBKWDvkg0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm0EWaoAMA0T8gGAQX2IpawmpKFk2NHyLDkgc41TU8KUS0Sn9vmOMxGYbPz/c6/JJ/2iPRAJAhOGHhJao7CnWxLZ+PbB79fB77OEHKK/IN9j4TK4kLrElPLVuBj0pP+MawlkOmq1mt+jm1VbcOIpGTPCzFOFFab/ohRaaAG/u9P6rTwUXoSBXj+QclgztW/oj4c0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm0EWaoAMA0T8gGAQX2IpawmpKFk2NHyLDliI0tlVN5G84NQRtKjncDcSc+YnhH5GrSf5g/iCtxkFSVHGXsjrdkzI2qbkA28RZcdhWHV7FD6VZ/mD+IK3GQVJUcZeyOt2TMa2OhQcHTLNC6SngbgjHbf6dUjba9BfC1yukvJ0+dhsP7fZmiWx8wIdIGwmce3wWL5HWC7eO+D8il4RWdivyT34RDm32/AKyGtjIEIu5IRbZ2gSwAcBie18JHGTsBB+CadF75WlC6PsTaMWyOJnvaY0g0kBjBle0Zm6N03kOe76auml5LZ2vyZD/XfrYjohNwvpJbXVC3PbScPWJaJolKfs6ySRYK1mG29plC+cyyDYad3/ccu/yA8G5ijMvAwQDKo1fNd3oasbdl1B2mzxk7JrD1oOhUnp8jqbdmcoQYqPHPT6yNUvnsS4cMmgMS30D0bmKMy8DBAMqjV813ehqxt4EcY3ae+42EBYNAncoGkgzFNXd2820FOH1MVbgl0uWOwCjrchNdOcdDbt2mQ2CjrZujdN5Dnu+m34Pjhcb2TzaPUHKcLuUJsGLJlWAlYXuXR768ZeCgbj1Gxj+pBQPcqnt7wAqyJilkETGOhmusAcRqv2XvT1NpHJegV4TCafDUVc0EplpmZUuC8J9pII1u3f1vKEWhJUvxw9OtOuL2H+j7YuDL6tJDjKU4zRAOAPRCyfJP0mpuVkTh07YyEg/zPqDXxlkXGyt/N4LG/1tUNgoX537xg0LLElUAdu6kpU9ECslbJEJZVpObnpuYEUwCUVEbpeCnAPqBm1/WBNgQD86x9HHMqRXLGsHkkgh1IqBWwCjrchNdOccct6g70ZoLXt9Tx1KQXcUhfBMBGq+HXdHQe+Y7GMjhvuBJBuMQkbczzkgZxSxkdwd13GeSeB0+X89ghTu5aRdlqbuITBtwgaw18//UIG53xSobEgpG71M9wukwNlc6T+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3eCMgS2aQYlSf8lVN2ZZgfoxCFMy3ABQrty9SLWj9MahDVHhRSEtqXSdRsYz5JZBMnmvXHN8NcKUL5H3JR+gnQZvxh72Y6FA+VPnyoAOCdrJtrrWYvsHNlUFh09Ch4hbk83FaAXWxGqILsq4ZGa6SjvtQTrroWfUQDKuVfSCivq03NQQFCgtDwfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctPT/IbYgO2uVnwg/IMu6/6X3GFc3FY3ZPv+ggUqaEPvXOGXMNJvXM3NonL3dWzRS56qn3s1umWWSlHcguKCnO5t7uAJKNEdEjboyxTc6gup/ne6FLBzRS7MoYZt3WznxE/4L/XDFvUbzNeVTltYXrWuptDHGlcH654JAdfiHMHTtm8/89hu8fA+ZerL0IEUN9n4okMRjQQ6+TMg31DiDriORkZlhxbXmM8y5mijaut+jvPiRLJcaPJ6/nou/PGxXKvnN+4Vo9Kbe8A1xv5IgAz25Ac0HZheuDbewZkqGhrhJXEyD7bOjVO9d4D4TNSL6mJLQ5OSBi9iH6cJsNrRkFrgSNBvfq0OWs6WJnNpvEwi/t7H9yXqyU3Ptiefzb1PWhloO57RoIvKRQCjPVg+MNMicrSChxLT8xEJr05kfCo9zz90/pxAjH/MKC66+P0LtNbwRSh+Hr4y+nXuWVoO3E2Cc4UcsrspMCeBBE3ASyx1udby7Mm0Qp4dOTwQP7uSlPGwF7a1yULWmH0QnDKBiqj2y3sG2TVRsIre1k7L1jguz9XP6j8B0FPOYmcs5Ok1gxAuGnGbG7qaoNxzKr28XxuofeqqBDYtlcxFj+2+tzRV+A+aShy2QUJ0mQcCaCCcuWnmWQMqdNIsxt5FnVxi4i+jCiFH9NVpPLXN2EDq886YWZZFop59sBOprLWAi8DBxE/4L/XDFvVmigA2sxfh3Yofj/KP4h/5qI1SbY5FM1fTtm8/89hu8RnxL5R7FWBiJBSBA5x57C5AqGGvXIwvo1EZBRFscI+cI94KHVBpBFWMw98LvuzZjwH/qNNQ4/XU0gmGylV8dZnvYig7y1TEsEYNHhdfKXcBBg/6c8R0Jjo+W1W6qWY55hXxsg3wq/hvXe975LCf+7uDEC4acZsbunsFvKzrLv6jG6h96qoENi0tZyDB6R0ucXP5I5WTGaeaXCjyJM9eBPPrITzA4MsxVEu2rphJr3+lX9Wqq8GrCpkB7yFyoxgT7C5u4YpUE3Z25C+/vo9kZj1Nz7Ynn829T0Uq+igkh6EqfB8xIh5ImPTK/HC4WETPVvMRCa9OZHwqR4f9j1IyzojA4UP3yB2G0eEyOT6Jg5gwmFmWRaKefbATqay1gIvAwcRP+C/1wxb1OQr/jvQrWkiVzEWP7b63NBhLotClKDpo07ZvP/PYbvFfb0r6eTF4DZR23nvqFVJSHdiIN0jIxS1bhom0J0WqgHGrboavNCi07LOXWm4/mIO0WCK5EQkod9Hvrxl4KBuPn9J2qUUeSCYTS9z5yesqt7SCXgofxdjQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Ltx5v2R/2i7QW6cR3ugt84yOSikUR84Jm6vt7lh6NPTEyIl9tcDvIrKwQFMBrptmFt2FocRTvBr2+YkbIMZ8A+du/y3mwoDlqvnujeI7UaGwAyrlX0gor6g1ND+mU4+mNYKajqXaHTllZ29fen32sg5wWZQw1j0XNH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8L9fSYVdAYPBQF/HGAtb8OmSJ60jnZ0ClqdLRnBrMX4NKJrUO/ewCG9aZ+c1GqC/hSJhEYVrJuZEKuWC3qjmSkEdAi6bE66DeL87iiQsvbGCFSbaDc4Qlm51h5E0gkpomTYDx0oL8iJkrAWCwd+65pMMBYLB37rmkwnbRqRLVzwSvpqQ6UP5ANaSCL0/lDTkTEJqWbEMG9PrK6BPW1+WiwP8BYLB37rmkwXA1PhK76CYDpNxToeEza06VqodDodiFlKqLBu3yOMdqroMFZmDjoqcBYLB37rmkwYbo5NtfjTJOD4b2SkwbVy8IKQH9xapKWm5wIy7VEbo16nDPYWVBQK9z/bGhnHqdawFgsHfuuaTCrNegB7BAwelMzMTd2VbLANuF9Szb8bc8riyPp1ahjhotDm2SkoC7m+fu3S3MoLDAVBFNCDVDPUGQFnj/A3sElwFgsHfuuaTDKvnlKNQJDCqw9aDoVJ6fITuyUW/8exDhsR6DJqCUVyvUyOYQ7zCgdwFgsHfuuaTDvLBREZBsyKW3MGdQoK7o5rR508ZTGndEKPItwc6DyW2vQikJWPE7CHYNbLmfROv/QGI+luyLZulcjp01RZXdDwFgsHfuuaTAvGoUUDSu+fwFg0CdygaSDksVqJxdxStzu+49+N5j8NVRWHJYQ/HeH0eLVINCmTFb/wfD5J7MibwL0kEjdIIoXOkoH8fk64rYMHZNkdaymPUtKhzFRaSADwFgsHfuuaTBCFBodbJdoTwFg0CdygaSDR2fVmEyqvVO2Wc5osDyA89R7j6mvjT7PwFgsHfuuaTAd9k0kAgIZXZTOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMPYX0HiBSNyGIc1hCg9j6TV8BYLB37rmkwYbo5NtfjTJNipQ3jNDYXS50aURK7nY7epa/XkEGd4zccRy4n5G9LBnPKxSUCjyIDbW5ec5Qv+Jr4alyc2izGjhozPPagAPwhDJp/pQZKDeJxCbuKBT0CTkIUGh1sl2hPAWDQJ3KBpIOSxWonF3FK3DgddvbdX6MFbUXfYiX6zhQkZOI7hBOT1gX94OU4e/c4rU2twQqZwVZQxUmdfALdqO3DhHxxYjAQnbRqRLVzwSvpqQ6UP5ANaSCL0/lDTkTEfroUhiOicc7mqvs3RF+zAve9HXWBATytXA1PhK76CYDpNxToeEza06VqodDodiFlaPuY0ytJXcx0ipyWLszxhiuQjVJvX3zIMVN4UCyUmVbAWCwd+65pMMBYLB37rmkwnbRqRLVzwSvpqQ6UP5ANaSCL0/lDTkTEPbEZ6naIcP6kGqMpcrzT6MBYLB37rmkwXA1PhK76CYDpNxToeEza06VqodDodiFlX9jyCjXAW/dS22145xhhF8BYLB37rmkwYbo5NtfjTJOD4b2SkwbVy50aURK7nY7ebu/xo9Qn2EBYggAh2zYxKrOm4GNjZXJtbnn+2wcSbtLAWCwd+65pMMBYLB37rmkwyr55SjUCQwqsPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPXVkydSh8I561GC34m3nhGPAWCwd+65pMMBYLB37rmkwj2idcEsQWxrNzaJy93Vs0RfzvLOuA1LyupmkdEVpLFttRd9iJfrOFCuV0j7hfrI3wFgsHfuuaTDAWCwd+65pMFjkF5+MYWA6cc7WB6YSrzjrhFTlXHuZ/8NSDFCecw87hfV/AzQi7unqCBQ6NPcb47fjfPd89LlknlFEOez9nWfw9MlWEq9WakLp/n2nSKskbTggdaVT/2CFXu+JyennczGQv3X6heHUWyemHUYw8wDnkyOhxNuHYmD8IE7wWPm+8HjL2Qw43bAjbPf3JibGS4qSAAlznYzJvt0W25erGIQD9tcnMj9RLv/u2T0BZF4r8HjL2Qw43bAuzKGGbd1s5+Aq0sbJ7EcEy+PRN4Wv4VEWI7P9oUS0PSjGEerW18uQc+kUG1CRIx+HY0vEVzVeKThU6TM2OsLJ4BgaHzW/UhEZ/SvsYPMGAjCfeTM9uG9x4sUtH2Qdc5+y0vYnS1liCqxnm9rCo0OvctZ8wH2tsNPhCXA+0K6+P5y20QfQAbjTGaF4BwRend3gw6vhm4hincBYLB37rmkwDPbkBzQdmF4qz8ujyCK8V7P+OBtpLdcxl8NC30BFnA+XwhesyV2dPD/9IbdeOigRPIDqj4g/TL7xrGoQHSNmnE+QkrjEq/GwlcxFj+2+tzRV+A+aShy2QRJuGFWCOxHAeIEWMn685D6Df/7fl+hYvqF4IVEXXnu7Ae8hcqMYE+wubuGKVBN2doLaZudjLGm9wGzGMk7QfNWeHTk8ED+7kssRUvpwEF58MJ95Mz24b3HixS0fZB1znyQUgQOceewuQKhhr1yML6OrcdiTQEM57g29rVwWCkjb6F+0TU7SlHPq6av9CaIXlspFAKM9WD4wmfbEXZ4OyxVGDR4XXyl3Aabc1GFAXQMAL6MKIUf01Wkd2Ig3SMjFLVuGibQnRaqAl5cNmVcIcNLlLtWFFFLAuHwfMSIeSJj09CJCGkzeYACdtGpEtXPBKyDzcsAxjJBksIre1k7L1jguz9XP6j8B0MVz29t1PvyY0Zhqz3Ki6p8hmrqfHLJrsXUw75byfRaj3O3Hu/jZuBCTKnwj09WqoFwo8iTPXgTz1KnEtfKCz5WSJje8E/l2/rTW8EUofh6+mRB6UVn94uMibxF1ACdn9qg18ZZFxsrfqbVp/Vbhm851TsUsPm6iUWG6OTbX40yT1ph9EJwygYqsxWZyIrthGsDhQ/fIHYbR4TI5PomDmDCYWZZFop59sM14CqWbAaVLV69Uh7cU7ObSCYbKVXx1mZIRsIPvxNC97ywURGQbMiks5wk09SjMEz5bVbqpZjnmFfGyDfCr+G9d73vksJ/7u4MQLhpxmxu6L288j+CeMMByXAvdH7CLNpXMRY/tvrc0rKY5gEPljOsM9uQHNB2YXuxDndysk4Yh5ynGMp9bSSleoXvjTFbluTL6de5ZWg7ciRnc9cNyisUK3OJbrgocAvcUFVcuet2FJqWbEMG9PrLAWCwd+65pMMBYLB37rmkwXA1PhK76CYDpNxToeEza06VqodDodiFlL7n3mFDlx+KIQuHkK1LeTcBYLB37rmkwwFgsHfuuaTAvGoUUDSu+fwFg0CdygaSDkNEPMoCb13ofILcYi00x4tz/bGhnHqdawFgsHfuuaTDvLBREZBsyKW3MGdQoK7o5AavDmDTROJEqosG7fI4x2oMeYwbJbELEpBqjKXK80+hhujk21+NMk4PhvZKTBtXLwgpAf3FqkpafAPOJZ5hkzGdAD0Fzenj9s/fOdT+1++tQgnJmgVSSnpV3hyOyNkFbNXqcWlKuB7gc62LjIBAnGVwNT4Su+gmA6TcU6HhM2tOlaqHQ6HYhZS+595hQ5cfiExjs5JK/InZt5HwYZgixkcBYLB37rmkwLxqFFA0rvn9S0pd/SoDbqxxHLifkb0sGc8rFJQKPIgOVd4cjsjZBW/Z2WS5WM+OVwFgsHfuuaTBcDU+ErvoJgNe4F6gSImz76n1DU9NV5kZr0IpCVjxOwqg18ZZFxsrf6RuI18FLToiYAIPUc68MBrT//Islk0UTNV9NkJ3IgcyIxKUD+YXwlUcyp1o8bE8jwFgsHfuuaTCPaJ1wSxBbGlMzMTd2VbLAqDXxlkXGyt/+J3a3ILgRbOmW1XMCUUAjwFgsHfuuaTDctJ2zoa1XsjVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3hzVfTZCdyIHMlYarIpZQJ1JXI6dNUWV3Q8BYLB37rmkwTCIv7ttHc24RaygtE5naOViCACHbNjEqs6bgY2Nlcm280fPVDUTOTZSmz4/fohxpWeWALpoumIxBLOrL1RTB3/IbLJzd1XoBp6QZr6kNSXQgZH/Prfb6w9WZoiiFN4qHJQa2D2k/1ZDsY21T3uRMTZDRDzKAm9d6cUdnVqQv4Njs2BhB3bcYhX66FIYjonHOEjboyxTc6gtH3qg3UeDtZ1wNT4Su+gmA6TcU6HhM2tOlaqHQ6HYhZS+595hQ5cfihr/7NekDA/riROEB4O4qE8BYLB37rmkwLxqFFA0rvn8BYNAncoGkg5DRDzKAm9d6K5rsg+zJuIfOUe32hDivHrEddF643SlEGehG8pYEvlXAWCwd+65pMMBYLB37rmkw7ywURGQbMiltzBnUKCu6OQGrw5g00TiRyvZhKluyThnYLfAGSBhjU8BYLB37rmkwYbo5NtfjTJOD4b2SkwbVy8IKQH9xapKWs8TuxAbbvihFfhon9Z63XMBYLB37rmkwwFgsHfuuaTA00uTno9W5oZTOxVf6qMnZI4vTKyHBGc+ZVQRIwsVmhFRWHJYQ/HeHvKpMsm2TwyZ7HSNLCCxOFMBYLB37rmkwwFgsHfuuaTCrNegB7BAwes3NonL3dWzRF/O8s64DUvK6maR0RWksW21F32Il+s4Uf0h/5H1vCppZXxwJEPmTbsBYLB37rmkwYbo5NtfjTJNipQ3jNDYXS50aURK7nY7epa/XkEGd4zccRy4n5G9LBnPKxSUCjyIDihqTq5TohFdt5HwYZgixkcBYLB37rmkwXA1PhK76CYAgZH/Prfb6w68voH2jFdgaudmwWraDKuRj0OQYfJiMxNAi6bE66DeLiGA1kVcqyDEpwUOeZhNxAQS0SN/g8i751IybwRAazvPAWCwd+65pMFwNT4Su+gmAi0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+ImVhqsillAnUlcjp01RZXdDYbo5NtfjTJM1Zicz6VVMhCi+G04JfRlAKwToSBd2MuIKDTzY6X5jNHBjWpkdkxGI61v9lEM+hckLfWXEKHgzLScPWJaJolKf6uHFVqmNRsN3/s2S3/AcnNtFH8awFvWeaDHA85r5sJnz8VLsZp+K1rWuptDHGlcHcMgfVzBp7zfn23xFCVteleAYGh81v1IRxzqio0ZomnflLtWFFFLAuFyr5zfuFaPSm3vANcb+SIBU1ib0s4ZGzPuDKsVH32k5GolaQle9y6BY9Gu8ZUOPfDdXxZU5gZJnY4rOqN9L4vSS/HKuP8Rf2JXMRY/tvrc0VfgPmkoctkFrkWU1DDwtGbUncqGOjeCSih+P8o/iH/nvRN+cuCvVtwWVRSIVqJFZnh05PBA/u5LMIdRn5zaBvk+QkrjEq/GwlcxFj+2+tzRV+A+aShy2QahIxMPOep9JWhloO57RoIvKRQCjPVg+MN+8KwEmJSepwGzGMk7QfNWeHTk8ED+7kg0VMIwNVlvF+pcWgyPqzV58HzEiHkiY9PQiQhpM3mAAv9281ooBjDYRKro5GXzlN3wfMSIeSJj0xP174gDGwo/UiE2L08vMT9ztx7v42bgQ3ZaB0sL4BOJEP98XS3m3N1TLv/vdm2Qcm2jRuQt1TYH6lxaDI+rNXuhSWVWm+TdEjJtb5ewhYNJPkJK4xKvxsC1nIMHpHS5xR5vU75Io8uRN4Zj44qxiRkUq+igkh6EqfB8xIh5ImPSJwEzYb4hXIXJcC90fsIs2lcxFj+2+tzSspjmAQ+WM6xBjqS0++rYBVMu/+92bZBxCvCFOhwrV5w6hXlyI1X1Dj+K97Q/MpF9FsjkxNlMDXKmbQ7J8vHK8wFgsHfuuaTDAWCwd+65pMFqk89/pi6AIv9281ooBjDZIT4nit6q+tLRmW10L0ixywFgsHfuuaTC+g8bgsU36svI5P9o1JFlvv9281ooBjDYfILcYi00x4tz/bGhnHqdawFgsHfuuaTC+g8bgsU36shp5IRzli53Xv9281ooBjDYfILcYi00x4qmyYXQd5shOwFgsHfuuaTC+g8bgsU36sqEKQDAExo3KIW8VdwBdmRaRjGUlDW9J9Dy1zdhA6vPOXMZyHBq//8yKPVGY51VV1mxHoMmoJRXK0vg5DvH2KTHAWCwd+65pML6DxuCxTfqyPwGopGN5FQ6B4KMG9hbpMC+595hQ5cfiExjs5JK/InZt5HwYZgixkcBYLB37rmkwJ2dx1hmkvRVDywnIQkQ36v5xjx8wY2LPqDXxlkXGyt8VBFNCDVDPUJ4DsouCSOckwFgsHfuuaTBYQzOZRDCbithksuNh+cYAQkP1FgSCfe8r6UhuhHB4P+r8HUmQVc97hbTaIcVNlmRy5MK0fr/EkmDUy0bAGUzItlnOaLA8gPNkBZ4/wN7BJcBYLB37rmkwNFav2H0sXKqIxKUD+YXwlXcmN6aMbQ2MNV9NkJ3IgczbKihHetHdsW3kfBhmCLGRwFgsHfuuaTBieCBrHGhoxmrWX8axLz2GZjySmeLaPsoMHZNkdaymPc882PM8gf4rwFgsHfuuaTAvX5QLQu0dPZoF4z28LONpnwDziWeYZMzyaiagphboiKg18ZZFxsrfGjM89qAA/CEMmn+lBkoN4nEJu4oFPQJO68byGCBOYAO/yRcdIlPKOF9n59S+kdLXHX3JOQsHU+CRjGUlDW9J9AuxizP2bUcBs8TuxAbbvigkicNNMWhMwGXf8k5ctsyCZdrYrgIKmgvD81KSt20OEc7W+/RZJSOc3T3qOLnPAV2/3bzWigGMNvQAhe/j9717iIDAo67TrOwuehH7LzbnwL6DxuCxTfqyAOcFxSNMQtu/0F0CLjsHHIBKh+Dvf72/SPnsHct0Z2uGhC8xWXi+vkB1ecXi+MYnMVN4UCyUmVbAWCwd+65pMMBYLB37rmkwVNYm9LOGRszw2/Ho8NRHYy+595hQ5cfiyW20jIkTGnjAWCwd+65pMMBYLB37rmkwol6Hk3ebFijBBL+fRwJ4RShRdHogOf/cfUqjpxOJssrAWCwd+65pME3hmPjirGJGLBjjUF+CLNKoNfGWRcbK3255/tsHEm7SwFgsHfuuaTDAWCwd+65pMKF0dwMb5l1FmlvW0gELRVVg1MtGwBlMyMLWAtdQboS1wFgsHfuuaTDAWCwd+65pMAQJ6tvIhfjtw1rgTYtyBHxmPJKZ4to+yjFsdm7TBDCCwFgsHfuuaTDAWCwd+65pMIWxy4iwpZ8+8CY83mAYs6Tc9CSVHsOFPheU73Klzgb9zlTaFc8J/TStHnTxlMad0QVL5kzZncwYjzeDdEvx55bTmYJPsMg+Q0xXPmRW2GhfEARN0oZ7PF0CLmfIM/UTQP+U1FahioRxHo78dc8FoAwMihLJdAxE+aIc/j4NtRsPsNMwfWlh5XISp9suVyXdDSJ60jnZ0ClqdLRnBrMX4NKJrUO/ewCG9aZ+c1GqC/hSJhEYVrJuZEKuWC3qjmSkEdAi6bE66DeLC83rqPbCSzqQEery/c4fRFQpZ+tnWt5YJqWbEMG9PrJxX2xf0wa4olMzMTd2VbLAHYNbLmfROv+IQuHkK1LeTWYCYVHcspp5wgpAf3FqkpabnAjLtURuje0g+Lz8kbCgXgkDBylGzbClaqHQ6HYhZSqiwbt8jjHagx5jBslsQsSyJ7wgeFyU0wFg0CdygaSDCDZMI+JrJV9nQA9Bc3p4/bP3znU/tfvrUIJyZoFUkp5sR6DJqCUVytL4OQ7x9ikxZgJhUdyymnnCCkB/cWqSlqdxdvymQ2Ut/RR3NYigAxxxX2xf0wa4os3NonL3dWzRF/O8s64DUvKBxl0y+KwUu21F32Il+s4UEtRfj9IyqtXPgXetxsYfRTAgLGi5HPbDAi5nyDP1E0A7LBFakgTSF+xjbVPe5ExNCDZMI+JrJV9nQA9Bc3p4/Scckrsrlod7I8v8JpqqcQbc9CSVHsOFPiKcIW0S4ke4j7GeEBde/DuUzsVX+qjJ2cFhRLHtr5z2/id2tyC4EWx0t5l/KSVXDHHO1gemEq84Ai5nyDP1E0C7mVmb2+QTluxjbVPe5ExNR2fVmEyqvVO2Wc5osDyA8/cgQkLzUfWBJeg+iExCMrmtHnTxlMad0alyDWxEiU8Ja9CKQlY8TsI24X1LNvxtz9Xhyp5wRBnnNuWr+EUTTShr7uk1aSIDwCJiCkjbgqiTQyf4c5CixD8gZH/Prfb6w9WZoiiFN4qHJQa2D2k/1ZDsY21T3uRMTQg2TCPiayVfl2dZHauNLhiAHFK8SMRXrSSJw00xaEzAZd/yTly2zIK79c/TOjO0vZTOxVf6qMnZwWFEse2vnPZAOanmozCmuQYYJjwzifG49+zcW/tqmGeUzsVX+qjJ2cFhRLHtr5z2HF34gAZl5q3pCgYVS10eex2DWy5n0Tr/RU5OGMXZ4nysPWg6FSenyE7slFv/HsQ4Y/3FFXKQO95mAmFR3LKaecIKQH9xapKWixdRZESkTMKO5K8dh3pLdaw9aDoVJ6fI6m3ZnKEGKjzy/5ZoxbazucLg4TLFSlMPyvZhKluyThlNbFwOWiv+X8EfppvqcUz6rR508ZTGndGpcg1sRIlPCWvQikJWPE7COkoH8fk64rbZdQdps8ZOyWKlDeM0NhdLnRpRErudjt6lr9eQQZ3jNxxHLifkb0sGc8rFJQKPIgN1TGReX5j+UI9onXBLEFsaeTCTjlA57Y34SW4WqIeN74mhOIgMLbIq0e+vGXgoG48JvFAzQiLcx+SOCFwaOINhKN+o8Y3Bzwt1Q22CFKYv69Hvrxl4KBuPdE7kIVyHArAr5MLZhS3k9of/tQ1TnyNO0vg5DvH2KTGvh48WgeAe+AGrw5g00TiRb7CKGgQd+In9FHc1iKADHDA7z0L52nuKAi5nyDP1E0A7LBFakgTSF+xjbVPe5ExNnGokgdKcFFMEqBWW0JLx7s+Bd63Gxh9FlM7FV/qoydkji9MrIcEZz2/3UNnM6eLtwuDhMsVKUw/nSv/rNmDxCQWqkBy0jfPtwx3aF1+LE50wO89C+dp7iiCL0/lDTkTEQW6A1k/HcyPfBZW1/xX+hmZDHMAELV1tAWDQJ3KBpIOSxWonF3FK3O77j343mPw1VFYclhD8d4dBboDWT8dzI98FlbX/Ff6GLY4u8XvVxlABYNAncoGkg5LFaicXcUrc7vuPfjeY/DVUVhyWEPx3h0FugNZPx3MjvJCpmQlowYGIgMCjrtOs7BWq1hd8bcVLUzMxN3ZVssCbhlmvWfHeKcOcPsm7HRZy4Cxv9dxY9YWhzggIVuBuTGlAqlLKErBpe66BPmKRG8XRDKF8K3NC1sIKQH9xapKWFIjp1DOt+yfdv7czRvnKL97Wo1mKhDIgAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4dBboDWT8dzIwwdk2R1rKY9rW1P/AYE4pGdGlESu52O3qWv15BBneM3HEcuJ+RvSwaFVSD1FKcXtE9CnTVxY3vYtlnOaLA8gPOjNZdHv3VmL6w9aDoVJ6fId4AgF2l+b7FPQp01cWN72LZZzmiwPIDzRUKpi2fQRDXNzaJy93Vs0RfzvLOuA1LyupmkdEVpLFttRd9iJfrOFKcnp15/O3TdM7pWWtiRBLF25uOVPuyY8QFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHgehPADCJihRNIkVojYKd+sf/QTe4OAnKv8kXHSJTyjhfZ+fUvpHS1/I6C/BlP5D0AWDQJ3KBpIOSxWonF3FK3DgddvbdX6MFbUXfYiX6zhSnJ6defzt03b8+axcXccjnDJp/pQZKDeJxCbuKBT0CTjA7z0L52nuKAi5nyDP1E0AcKEGREeUMHmvQikJWPE7CYsacUWhCF6A77yCI4vDW4edK/+s2YPEJ0CLpsTroN4tl3/JOXLbMgnHqsG+fU83mr4ePFoHgHvitHnTxlMad0TtU9Hco4V/Z77ga/cJ2fpnH/0E3uDgJyvThJyXFBSaVPsSVUmfjib+sPWg6FSenyBl4xHnoc5F3o5QHqGJlk0GnJzLtS90jxBSI6dQzrfsn1ceqXdpBMS2UzsVX+qjJ2Z0TyUy/Al6L2yuopaJ3WbFe0loikmcP6KVqodDodiFl50r/6zZg8QmSyE1KaDflSJTOxVf6qMnZI4vTKyHBGc+ZVQRIwsVmhFRWHJYQ/HeHQW6A1k/HcyPhVAuScmh676w9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9FIjp1DOt+yd1KoutmKmK4jA7z0L52nuKIIvT+UNORMRBboDWT8dzI2TTzt4udd7Vr4ePFoHgHvgBq8OYNNE4kacnp15/O3TdbaghYXlpv6usPWg6FSenyOpt2ZyhBio88v+WaMW2s7nC4OEyxUpTD+dK/+s2YPEJ2bCj2fcQIXo8Hfe4JT2CyZ0aURK7nY7epa/XkEGd4zccRy4n5G9LBoVVIPUUpxe0/0ImPkJmWxr9dttIfq43CQFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHQW6A1k/HcyPgRxjdp77jYQFg0CdygaSDnGokgdKcFFOYsJ+3Ynti3vYMAb28qXNflM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCc29H8QfFoaYMDvPQvnae4qf1Ly4rVHjsEW3/xjgeN4byJMDPf58wFvfcf1Mf9P6Y52ZIevvosDuafAXapYNs5udCClQjtkLmsZEXwGx4BMO/+7ZPQFkXiuioOnn/o5+eWz+KYrx7nU/WXk+RRG5wTBmtRIae+35+uR19P3SUAiEK29pv2p2ZiwnD1iWiaJSny+wDNWT6NrP8FS4hpmCSp5UKWfrZ1reWEWyOTE2UwNcqZtDsny8crzAWCwd+65pMMBYLB37rmkwqzXoAewQMHpTMzE3dlWywKg18ZZFxsrfOGdD8dBHJYT6nY9cDso9N8BYLB37rmkwyr55SjUCQwqsPWg6FSenyE7slFv/HsQ4O95IiZfXcDRztK1HbwK788BYLB37rmkwXA1PhK76CYDpNxToeEza06VqodDodiFlL7n3mFDlx+KR2oL8nuFWz6HyHRQ0QKdRwFgsHfuuaTAvGoUUDSu+fwFg0CdygaSDkNEPMoCb13pIsuUh2LMETKVUjlT2vocatP/8iyWTRRNPWdlcJT28jQVKXuPBvFIn/87+eme0CV7AWCwd+65pMKs16AHsEDB6UzMxN3ZVssCoNfGWRcbK3xUEU0INUM9Q1HuPqa+NPs/AWCwd+65pMMq+eUo1AkMKrD1oOhUnp8jqbdmcoQYqPGt4HkPgqkJs4cMmgMS30D2zxO7EBtu+KD8BqKRjeRUOzzzY8zyB/ivAWCwd+65pMDTS5Oej1bmhlM7FV/qoydkji9MrIcEZz2/3UNnM6eLtwuDhMsVKUw9E3tygC005pCuLI+nVqGOGUcfJNDRFkYxQgnJmgVSSnqcLcQrv4Vv8e66BPmKRG8V7EtXq63l7iVwNT4Su+gmAIGR/z632+sOlaqHQ6HYhZWY8kpni2j7KDB2TZHWspj3RVKRms1ftdMBYLB37rmkwQhQaHWyXaE8BYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3hzVfTZCdyIHMlYarIpZQJ1JXI6dNUWV3Q8BYLB37rmkwj2idcEsQWxrNzaJy93Vs0RfzvLOuA1LyupmkdEVpLFttRd9iJfrOFILF9nAZbW1Ml6r3CSjbOX6B5vN6lMor7Gvu6TVpIgPAImIKSNuCqJP2pcAdaRKjvo9onXBLEFsazc2icvd1bNFXp+FAiC2msRxHLifkb0sGc8rFJQKPIgPtJ1HzQxcqyTFqDDBGqQLmRbI5MTZTA1zO1vv0WSUjnN096ji5zwFdwFgsHfuuaTCrNegB7BAwelMzMTd2VbLAqDXxlkXGyt9AOanmozCmuQYYJjwzifG4hoPjasusdD1tzBnUKCu6OQGrw5g00TiRaPuY0ytJXcx0ipyWLszxhiuQjVJvX3zI27wNWQR10PsxjHhxXS1Mv8BYLB37rmkwYbo5NtfjTJOD4b2SkwbVy8IKQH9xapKWs8TuxAbbvihb13wdrtS2ScBYLB37rmkwwFgsHfuuaTA00uTno9W5oZTOxVf6qMnZwWFEse2vnPYPLQj5V8ycxsBYLB37rmkwwFgsHfuuaTCdtGpEtXPBK+mpDpQ/kA1pAi5nyDP1E0DfF+j+J/HrZGvQikJWPE7CqDXxlkXGyt9uef7bBxJu0sBYLB37rmkwwFgsHfuuaTDKvnlKNQJDCqw9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9YNTLRsAZTMjC1gLXUG6EtcBYLB37rmkwwFgsHfuuaTAd9k0kAgIZXZTOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMPZjySmeLaPsoxbHZu0wQwgsBYLB37rmkwwFgsHfuuaTBCFBodbJdoTwFg0CdygaSDZmVQ/iwXbytr72NxY56leiYteRndDGLsaSOpSxNmlKmDeIyo7l2sXAUUd1BPN1gSJw9YlomiUp9hwZ/mRtOSotFDXlcnDT2Y6ggUOjT3G+P0BJRgEJ4OGy3dEWgk/3CQA+Oc1Npth69RY+fnLq7F/D1N9d+fX7PwqDXxlkXGyt84Z0Px0EclhOj39CSptuk74FEk8PLjGvyzxO7EBtu+KBp5IRzli53X16l9QXE9fX6XlUsPHnitQS+595hQ5cfikdqC/J7hVs/4nT3J0ViNpqEKQDAExo3KIW8VdwBdmRaRjGUlDW9J9Dy1zdhA6vPOXMZyHBq//8yKPVGY51VV1mxHoMmoJRXK0vg5DvH2KTEr0c/ovno5F/rulmFJfXtIYk+ciHfVdO6Vd4cjsjZBWxDSCoJxTrDaDxMzKqbEDxOmM2sdTEp3ZrPE7sQG274oPwGopGN5FQ5T6DMz1NlKVj8BqKRjeRUO8F0+ANgJ0sPR4tUg0KZMVv/B8PknsyJvAvSQSN0giheoNfGWRcbK3/4ndrcguBFs+ZC8n8a2DmpieCBrHGhoxg//2FO4hHrZv9281ooBjDaN+6jE6JHeC/P1NOoJwhfqLsT1DdvvEkJQctJ63YbON2F9B4gUjchiHNYQoPY+k1cvX5QLQu0dPZoF4z28LONpnwDziWeYZMzyaiagphboiKg18ZZFxsrfGjM89qAA/CEMmn+lBkoN4nEJu4oFPQJOJm3LgZz5FuU1Xl4tAxWUvrVLgxL89mSCnb35auPGcy/tJ1HzQxcqyTFqDDBGqQLmRbI5MTZTA1zO1vv0WSUjnN096ji5zwFdJm3LgZz5FuVQxUmdfALdqHRTvYezWROGaBA8TC5ucacvufeYUOXH4oa/+zXpAwP64kThAeDuKhMouFWb46jhYaOW9hn4ekjuK5Pj6mLQwSGoNfGWRcbK3xxd+IAGZeat6QoGFUtdHnuoNfGWRcbK3/RcTsJJ8QYw1RZw/FVGmt6oNfGWRcbK34mWRjIxk25wDvNDqSsIMaupU+9UMTX7Qw8tCPlXzJzGkqe3BprsTdHASdLvMqoB3cr2YSpbsk4Zk9kEG02JCz5DJKbZDHDaVL6Ljss0dpaXe9nMsBBqXJzZDxcApcmySDZP4UWWdtb0NV9NkJ3IgcxClJFtvcQ+6je6aDKv64egoHmzsNLB/HIyyS9tD8WULoV/WU3qpuprCJmH48QV0CPX88nixuUVIMk0flCMwg9o94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaGSWbTIsYUSQdZW6GV6T+u036mVZNAlLLNL4OQ7x9ikxfPBntcazikk1epxaUq4HuLh5HJpZ8UFg1uhkf50lBKRRuZspY/Zlvz8BqKRjeRUOn5pkv+29tQA36mVZNAlLLIJIoCLLjeYmFQRTQg1Qz1C4o+rELtG0r9ZbUSIgt1qhBUpe48G8Uidn7jRzMl7GhgVKXuPBvFInyIzN2gOlS4rWW1EiILdaof0UdzWIoAMcs/IT2ZPQHhlZt+SqJtO2gKOEbht4BwRyPwGopGN5FQ5JqWNRDiSJdGWxPwOOlMm6qDXxlkXGyt8nD1iWiaJSnwldkCFjwDorvW1uJ09i8hPlwA+e7vpE+FDFSZ18At2o7uoPzr5OQH4nD1iWiaJSnwldkCFjwDorq+4xvEoC5O/7l2JhySd9lVDFSZ18At2odFO9h7NZE4ZsSF7zibuCLCcjgeVVuCXbdeuKdsfJ7huIgMCjrtOs7JMmL3IRJNPCAOcFxSNMQtu/0F0CLjsHHPaPw8tDXJyuoksIRLPkiuPmqvs3RF+zAjdE0Tn2xtBRI5PzjVy2enW/0F0CLjsHHE8CrRFZfhfIXOLFD8ojL79U11gnm1y7wqOEbht4BwRytlnOaLA8gPPDKs7TWGVK9SbGr8YxPH9rMR68lVqQce2oNfGWRcbK34Z6ZIxqv/aCkIbDI91ni1wuxPUN2+8SQheAIzzXgm7Z1ltRIiC3WqGVhqsillAnUjRQAJFG6IIZ6bY4q+uA9AuoNfGWRcbK3/4ndrcguBFs+ZC8n8a2DmpXHTABR4KFlDxStOXLI6x8yIzN2gOlS4phfQeIFI3IYtSMm8EQGs7ztdyC87UfxxHbKihHetHdsVEAxF+JRlis3PQklR7DhT4oIKa6daczlF6Nd2t4XHpw6bY4q+uA9Avj5RcgwgjQhaJLCESz5IrjQSzqy9UUwd/yGyyc3dV6Ab1pLXHM4BUna+7pNWkiA8AiYgpI24Kok2LZ0RBkKj/BZjySmeLaPspOewl/jhEQB4vI2KVuH7RxL5J75j0HMuVaISAtYThB0kEs6svVFMHf8hssnN3VegFXWhNbHeE16Wo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa/+gtEFzV2Z5i2ivfD2nwYPBSay3l6556MeT9DJ48gRZ/FJxES+W2uy59GIrxYFC/Cem/tdTojcxABpLkx4DeSBIT4nit6q+tPsgv2m/uvmUuF0OMqX8TPs7nLtgj8wGuRE7nNp8sszc5iKqJZa0JmqvLLPxVFX1Ke0u0VsWSN4rtfBNeZpk/I2QaH0B0kLJFCpnBI0n/RJkMF5K3H8eP4rMin5pblEnIil9m5P6d5QorQbn/1U3SxXTigpD6jq16tPNwYjpCrYIVVtw4ikZM8LNfgAg5nDYHCSJ1f5MukVLX4CHGxF1gxO+aKF8/OgqHypnBI0n/RJkX4CHGxF1gxM3LeLlI0CMc5UXtu+/7uhRX4CHGxF1gxOk/f5AuYfuclW7ozuVoOLIAoHnaArgPt1uY62PEL53q7B5JIIdSKgV0nI2V/2B+1JVW3DiKRkzwiGVUf1Ew5nGt6BxeFxINmlg1MtGwBlMyMLWAtdQboS15A7V6S3r4tjVsVft9q2P1TVfTZCdyIHMQZUflK3iu1gekCAbLLKQJoM+aEC2mLhmax7M6tZYeK72iuplgCAem8bc2MNXcGDLZCaossf1EG/q3YFFR2s4AFQEo83cZQQWl/ux5LaKvyLSu5NX3VJkLh+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC4kq3srN7+p8SDYYEZZ2nr5tri1hIYa7vqDpZWXNzWXSk5Ok5wGBoKhccAKiMeC1ZbF3uU2H/DCyQO8ZxWsk4lK1bfk3tLW1g39e2VsGp8X0R5/Ln8SPrc/jUoqU3tzHnaFe+Y+2cTHgD3b6AdMxWsS0M8u2CbUGI9o5s+JQh+GxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LL2V87xYw5PxPIwpq0wN+BArnlhqKJytxmPQQkgisl8tYnYqcZVLiNEt94VFOaCHRBFh+Pi8K3UmNanhf98S2FWXekQSjTOhIqfSQcbwI1BecDP+1jQ0/h7dx6Orf8695LKBmmOe67LI7T6JQ+hpNEaI0UfY20Pp+NGzsQ7/B5p87T6JQ+hpNERX7BV54BMbzed9pio0bPALkPc7CpPACInV0KBb9b2VgVO7B9DkWWZU0Pn/VgPsBD65YLeqOZKQR2w6uZ3qRATcGJVGYi5tDsft2THkfDG77rBxXQD2wvp4fhcE4/+Cy3whKCCDytczOlM7FV/qoydnBYUSx7a+c9pciTUmVl2Nysie8IHhclNMBYNAncoGkgwg2TCPiayVfIIOV94uyRfgjy/wmmqpxBhLUX4/SMqrV8+pcdtwlFegnUCoE+R7cwQFg0CdygaSDn6ADi5zKCB8/AaikY3kVDlKUnG7T12N5i0kWLnusckK6maR0RWksW21F32Il+s4UEtRfj9IyqtXPgXetxsYfRR3bcYOqDhgjKJnyGPmNyWbhwyaAxLfQPWpGPxRfAM1oUcfJNDRFkYxQgnJmgVSSno37qMTokd4LD//YU7iEetlCFBodbJdoTwFg0CdygaSDR2fVmEyqvVO2Wc5osDyA81nfpZo+TSgbMYUzgfh5/C5OQZIm7+zr2MLg4TLFSlMPYX0HiBSNyGIc1hCg9j6TV0IUGh1sl2hPdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDbW5ec5Qv+Jr4alyc2izGjn5sQLuUwh4fz9+B5bv6EKggZH/Prfb6w9WZoiiFN4qHr1AgXgzKfvVYggAh2zYxKrOm4GNjZXJtgGzR/3QXaeRlfnIgvbayWqLIDNIzkHgxYUE3gRWQ3Uz/N2MTaHVG96+REFSqpSZn7GNtU97kTE3hQdEXYU/SbOVaJp8vfd5ys1KS/zkt0hvrArnGJXol6D0ppXEwM1yMWuBI0G9+rQ5l/XWxX8MRVEowBTBDTHuV5gu6cFolLo+2/7h3LXwX4DAngQRNwEssD4olhis9ms9nHy36d8LQTL90/v0Oz005sjkyE/EtHt4UiOnUM637JxA1EJ+0ThX/3hCE/DPBs/a3N2ItPs9tfuxjbVPe5ExNnGokgdKcFFPMrinkvOLhJf8UaSQ3aOtAmLeeZbuMJ5EcRy4n5G9LBsjzVMb2WergQW6A1k/HcyPfBZW1/xX+hmZDHMAELV1tdWCm8N7aUUocRy4n5G9LBoVVIPUUpxe02+OgMcAM3pyMJ/HmWrKilXVgpvDe2lFKHEcuJ+RvSwaFVSD1FKcXtNvjoDHADN6cSl8lpO6CT8J1YKbw3tpRShxHLifkb0sGhVUg9RSnF7ReFrBhJuZaJeY4NvWfIyqmr5EQVKqlJmfsY21T3uRMTZxqJIHSnBRTriz57x3bIHh0jTR7QpT+X9/4fk0LORRk8v+WaMW2s7nC4OEyxUpTD+dK/+s2YPEJRuNnSfU5OOqSh6M44dDko8iWrJOO8Qa44cMmgMS30D0UiOnUM637J6YJYDZ8Hf7io6Fxp5dO7pXqfUNT01XmRmvQikJWPE7CK+TC2YUt5PaArhUKTBgj6Ig2+XVXDrBit7g7hkhmqeQcRy4n5G9LBoVVIPUUpxe0+yQikIWbDVbQcyzlC4hPvvSJ52KAGWjkRgvHF21aQvfhwyaAxLfQPRSI6dQzrfsnIR/RIxbY8VKwYqGyCgiLHCpRMnkZNqxCWIIAIds2MSryTKIkUcCMHdnxLCf/5l/ispuk2fuGQC9w6ZSDkfj/lMfxg9KgCdBgwuDhMsVKUw/nSv/rNmDxCftxGgHUwF/pNWYnM+lVTIS66cbV/3KUkVRWHJYQ/HeHQW6A1k/HcyOEjH0DU2cbLItJFi57rHJC4LuegnKGAs5tRd9iJfrOFG+wihoEHfiJYPd032EYaYM3PfZF/mYRxBxHLifkb0sGhVUg9RSnF7Rqp7a0UEnGpI/+V7WO9DwLoJ8YWcJWsqBYggAh2zYxKvJMoiRRwIwdSGOfMlIPT3fndEVhlQFMsa7TLBTVr3Gn7GNtU97kTE2caiSB0pwUU4/XkN7KgPfFo6Fxp5dO7pWA82G8rECYlGvQikJWPE7CK+TC2YUt5Pac/7ZRIl/9F5KHozjh0OSjptAJInjr3WjhwyaAxLfQPRSI6dQzrfsnvj7JADSApbXCCD8Qa/jQUL72zT9rXnkBwuDhMsVKUw/nSv/rNmDxCeksM2xnQ3YLi0kWLnusckLgu56CcoYCzm1F32Il+s4UpyenXn87dN0PUWVBQl/1EKCfGFnCVrKgWIIAIds2MSryTKIkUcCMHW2ep0HnyKqht2m+24Kj1NiA82G8rECYlGvQikJWPE7CK+TC2YUt5PZaVaWYc7x7C8IIPxBr+NBQvvbNP2teeQHC4OEyxUpTD+dK/+s2YPEJbK2ONC6dtJaLSRYue6xyQuC7noJyhgLObUXfYiX6zhSnJ6defzt03fNb+NVshyXaoJ8YWcJWsqBYggAh2zYxKvJMoiRRwIwdjKao8w367t+3ab7bgqPU2IDzYbysQJiUa9CKQlY8TsIr5MLZhS3k9moKJRxejdqNwgg/EGv40FC+9s0/a155AcLg4TLFSlMP50r/6zZg8QmnVKlZ+8sNcotJFi57rHJC4LuegnKGAs5tRd9iJfrOFKcnp15/O3TdAgCoxve1S/qgnxhZwlayoFiCACHbNjEq8kyiJFHAjB0MVydUdWbMoXhP69nvk2w9gPNhvKxAmJRr0IpCVjxOwivkwtmFLeT2CtPeWFHOxJXCCD8Qa/jQUL72zT9rXnkBwuDhMsVKUw/nSv/rNmDxCS7ejH5im5+Oi0kWLnusckLgu56CcoYCzm1F32Il+s4UyhTlqu2FfIMRZ+JkkvOB5UTaP5SVi2/z7GNtU97kTE2caiSB0pwUU4asnNukj2n0wgg/EGv40FB+BeXeg9i3cMLg4TLFSlMP50r/6zZg8Qn/FYXkWkkpsBxUpe6e3KRVHEcuJ+RvSwaFVSD1FKcXtCiAf3Ssl7mBBcsOI3TA2xkJ5jCrQXuHN2vQikJWPE7CK+TC2YUt5PZazp58RsepyzVmJzPpVUyE85PQKcPDenBUVhyWEPx3h0FugNZPx3Mj5vFCdhpXMacwbjsaKEauTliCACHbNjEq8kyiJFHAjB2UIWNcob/9I5KHozjh0OSjptAJInjr3WjhwyaAxLfQPRSI6dQzrfsnATWN0qboxwaLSRYue6xyQuC7noJyhgLObUXfYiX6zhTzqsUZ4hmxNmaYQhqPazlYrtMsFNWvcafsY21T3uRMTZxqJIHSnBRTFYXcIqbiy2HCCD8Qa/jQUL72zT9rXnkBwuDhMsVKUw/nSv/rNmDxCcbh/Qa7+K8eo/fcjlASIKz1girRWgAdKW1F32Il+s4UvD90zBEMvO6dhOb2ajAi+Ilr6Ie+/QEHWIIAIds2MSryTKIkUcCMHZOIn24nSXdED/ah7JUhA8SLSRYue6xyQgJxrYyvr9AVbUXfYiX6zhTbA8chY5Tt3MIu8uYJO+XJkoejOOHQ5KMomfIY+Y3JZuHDJoDEt9A9FIjp1DOt+yekLhEkIVg6Ox4QPaaUFCn7NWYnM+lVTIQovhtOCX0ZQFRWHJYQ/HeHQW6A1k/HcyOlVhlfLVsZCjgQVfo6qdn1JlCbtD44IE/EgjECtmptXCvkwtmFLeT2JUkYfHnctoKINvl1Vw6wYgAuUmMNk8vBOOCrltLRHTrtN2GeUw+Ykqcnp15/O3TdqpiM1HANGtbFHvpbjrt36kQxQsi2xslRxIIxArZqbVwivd4MLtYJAf3RpbD7/vXm8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/H4oX+KSqn8nyTEqUDomNrlzmt2ko6MMbby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8dNERnB9b9x1Gj4K34jS9LUqATv9aDagXwapNs8kxEvP3QECkKWF9L9heAsGL4dJ1ibZ+QaY07vLr5jbKD008HRMVt+R5f9H03BNudsi2ngm0y500Sbu28OIt1VHmsDk5BTnIMVgLZ+azc2icvd1bNHavFdz3pmbF+so7nbu8mqBeNYYKjqEH6StHnTxlMad0Utl0MVy1OFL2NLBLzRFHMzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+To4dhv1qMaw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9m0jk95j5G3Djl4qRcMiLXxG7yRYmplVlNJOVcFLrQgnc2tM3AeNaPgzyjRpm453F8Ep6XLleL7hp3iUflwWpraOWDQJQVUMt3eAPW4ucvJ5YvyE3/NT4DnO/LoMT3gc3E1K0XyfF55kilXlysJTQHE8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/GqhdI0OAzU09rL7bLiQk9uIPEEOOs5sYJFhs+T6mvC3Bp5IRzli53X5CRqz7/gFKofUxVuCXS5Y32Pkite4rtGKQ9XKZKOL02NVcWq422EslVbcOIpGTPCH7mUaPtluaqp8akuHxFzA0CGgMvrUkxxN+zZPe2/uq5hXFeqSkCIGA4tHM49qAi1u3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6QiCqQNMvp2g0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek7/smYr+WTcY/aqByDZ6jU0E9c1gpRGLR+Fy44jk47FMpzdOt7KYglnKhicQBYJfeQ0OvP90zT1HixfGI9/oyonbPz/c6/JJ/0zJ/bYDVRTMPcYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaBq8gbPerYPmQjEwLog94FWMroHGyZS6tVm35Kom07aAqDXxlkXGyt+QnBWQZlybtarz/5Dft8cjQmBYsh6oM+lxCvea/bRFrP9VOEEPlSHPDi0czj2oCLUFqpActI3z7Vm35Kom07aAwFgsHfuuaTCxaXLnB01YPoyugcbJlLq1L5pREXvfxYMWnOIbR1Um54MoNZA6HRxHSUw1fI2054NTSeLqSGnLm9AYj6W7Itm6TKVS+fDCQUJJTDV8jbTng6yAfAZKDBVBPwGopGN5FQ6fmmS/7b21ABD0ExRs9ghb0uwTtBtpz0TkJ38aOfGtD/wfllR9T21BO2fS5qZhn/Fx8tfLfHJerbBvkETgs+XWPwGopGN5FQ5+jzavHUBG/xE7nNp8sszc5iKqJZa0Jmr/smYr+WTcY0/MTsEX+1QQUWSRcqjUbYTyAfioHpHTMABKVBuglOW+ax7M6tZYeK6c3TreymIJZyoYnEAWCX3k2yfH0gfyTVBMidbPXl/yrNwXpnpCDDozQPVHMmkNW9PGzEHVOiRgPB7MgvPaeKEq2Q0WC4t11ZOE7pvWpjzbDr2rBUoGQrMwvnE5wKNaMBRiCjv/vpJYcA/ZyqaUStSaOoYBtSmxCIpZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3NbD6g90SZWE75Z5C4k3E0fg/dxrdljanPNuZp8G1pywA9kMejUbeuaURoY3qwFw5PTtLOpVKj7it1xii0jXPYfg/dxrdljaoQQk1MP5XAxwA9kMejUbevwtQJaSuH+a2HY1KyzivUyl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGaBxI/NQhYrFtr4cyR+8KMm6637rD1jOjny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTSZHbeUSmYeJM5+MbNvSg0mFf1lN6qbqa+2d+iBc8v0FHyC3GItNMeLnbSP9FHkYHWRXZEp4UN23chK2rhaMLmZP5DKhKevgqeGFB3kb9erk5iKqJZa0JmraCO15ZLEyw/aqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+qDXxlkXGyt+/FMUSc15bz/aqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+qDXxlkXGyt9JbNI9vIjR2zSc3R/HQ5ndOSHV1ZqHYJlRCWbeSOoaDbQLbwE2vp5pYVxXqkpAiBhK8O6KdQYTdTSc3R/HQ5ndOSHV1ZqHYJlRCWbeSOoaDbQLbwE2vp5paLqzJmflsPSXt14nAyWWX0NaRZr5dtq7lcwbKRQEQlmWnABkhfYwG9iuoTHUj00cm9dfGYFWkf6p0CVakGWe4B4shfUOivwDFrvOgzPBTy5BitJAkG/s/lAbV/pq3+Q2jGFGQDlBT257Y7FX7V/uVH4rbsGY09o8L4kzwEdzQHap0CVakGWe4BNDewXXW1v2T3Da5cz11sxA9UcyaQ1b0+0aCqKW9N8dvxyMK0QSw6EDWKYzQStW/8yNickEs4ezYVxXqkpAiBibfY9fJAL2tRzlw8QLgf6PDsP/uGAygqusNWZ4XQCGlRxHLifkb0sGSFse/o5UMU+UMeN1MqFCHcWLKjNQnIjWYVxXqkpAiBhK8O6KdQYTdZFJPvOk2dplFk3/3O6iogfcqNk+qxGIYDafoqSRYJzvt4eh0QBo3jmMYUZAOUFPbgDeJ7DMa/1ZUD6VkhIFiC1hZozdt25vcDNSC50CghXz5oyoIXeJbFtTnYC1zg6kS07HqzFUYFswWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNzWw+oPdEmVkmnp9XyTwj+xXgMv8XbsER6pKzXpWco3+Qwf+dxRTjr8bJ6c7o0aB+q5cCftaVYON/b2c6WFk1d82+vD8TPOOJr+TQ2G7uft4Uu1Ox/A3YwS4E8kVDuIQsSQUD0/7Pgg5lcsn/5iRxxSmECqubyxfHoMJ1XyK/9Z0b2eEbbrcBUykV2MzVoLQzz8AAo9hhykyTEOaFTiP8bkc9j6lHIF20hfhDiZVaJh40J/yrMBaXLbvlJyn70jzBlcJ8QHSx2awILWXTpRYUCyPNUxvZZ6uBX9u6rppjieNfDpr+oqVdrhs5jgPWkfV1y+74S1KdbPI9GlJPpEKAkmcJi4MSY4v+XTf7IG0UNahJBQPT/s+CDR3NC44zcQ9+XYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZgLfEAoiKF8CDZQvE71G9cZx8tfLfHJerfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHwqpRVjxnz+XV+1ar9SbW7oV/WU3qpupr7Z36IFzy/QUfILcYi00x4udtI/0UeRgdZFdkSnhQ3bdyErauFowuZk/kMqEp6+Cp4YUHeRv16uTmIqollrQmavZnxI/YRvUtu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6HH26M3el8Lm7cHGcmccaLbdTi1x3mcIYkNEPMoCb13oWhrDdTVc4EbtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXen7C6VERnyqEu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6egLxgqlpcIa7cHGcmccaLbdTi1x3mcIYkNEPMoCb13q72zx0S+CpUbtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXemNoiI9rxRS5u3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6VJDf+bnxiA+7cHGcmccaLbdTi1x3mcIYkNEPMoCb13oYeJqLH5STV7twcZyZxxott1OLXHeZwhiQ0Q8ygJvXevavX0SI6HKwu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6mjzGbPQJprG7cHGcmccaLbdTi1x3mcIYkNEPMoCb13qdHBZXsVzIhrtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXettE4yxDB36Wu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6t5PabniS2WD2qgcg2eo1NMOTyNLgcNdkQIaAy+tSTHGq/E96ZInMfqg18ZZFxsrfpVYZXy1bGQo0nN0fx0OZ3Tkh1dWah2CZUQlm3kjqGg20C28BNr6eaVVbcOIpGTPC3GeZegu9qMA0OvP90zT1HixfGI9/oyonbPz/c6/JJ/0zJ/bYDVRTMPcYpJslCjaz94EbwpZrvjSQrFoNqx8+m2L9BnFMDbKCKQm4xyH86zW5YOX7gU6yaDa+4QU3RPr5rbqO8tJOiTKQ0Q8ygJvXehx9ujN3pfC5qM/i9JTSBWyWGyHcMQ926ccW3BFTTQE9ybzO1qijzjJZovcgxsRVrFA+lZISBYgtijwGMnDVvQE92mh43+POFHCI+NeFN0tn4+UXIMII0IUGyYLbgdNucnfLhJhjvyQjqDXxlkXGyt+Xv2AzoR1u+XNS5RuMthAaHeZQZbWslnpo+alAwUhAXef/LtKYD0xpOMqqLQrydnpv6qUwOF2sJJqvegb+vwowE38RzqEAvfKAyAaDCYq7K6ZhREc2ssOTGHiaix+Uk1ey6uqUkX/Ge1VbcOIpGTPCQGjay0D3SwdHR3ZB10wyPtvt+ZWcMqhVuZoWB3SbxCN5YdgOegMiMsVoUdGx2cTNAoHnaArgPt2fg+40vZfCqntTECW5LqsHkNEPMoCb13rbROMsQwd+lqqvbZuWL9SeqDXxlkXGyt+AcTFIOQiwIzLenxss480Pi7H5oT7MrPtsSF7zibuCLDjgq5bS0R06sLcbhRl9tGhYzMx0NX4VjQeLWEITgQr9cviWQ99kcYePpgSsO9diXBa7zoMzwU8uQYrSQJBv7P53PDtWMWrbTupsYkh//nQeD+Qk8tyMavlSQiTI9fxSyvpuwthAdXlK4rXWWhvuQDFaF8HuNOQTF6RZ1wRU88A+V5VAZbfi8jIETOWt0KBunDb9QuSHDNdeffqlppcnQWarsEsLMzN2uQtzbtkZ/ozUwzyOGNtmZ8ny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+To4dhv1qMaw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9lu1ZKE7sYMba3vAPCmghKL8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEd+eFCV/vUoIII4KkL9ljjxhX9ZTeqm6msImYfjxBXQI9fzyeLG5RUgyTR+UIzCD2j3gRvClmu+NJCsWg2rHz6bYv0GcUwNsoIpCbjHIfzrNblg5fuBTrJoDpfLb3L5qx9jZaaT0bMjLxkWlValnsrqGldaXEMdfttoc58c4jYggqg18ZZFxsrfTi6gfGLzQzukJBs2QFmbHV3gpLQ826asnpoklFeql65qmIG4MOpQxzV2e5LCFT4khSmClL5kJWeTM4jmqp4Bm21ulXCfyrigFG17LFGjQe5KF8s3dVvda4RvOWh7OfXVs6bgY2Nlcm1d6U6o4Q6KkYQv/6mTXR6UdeGEYCjOSTUR6UkUZS6J2cVrCVbbQ9EwqpovBFeobYyU/QqKXDzNFKg18ZZFxsrf0X13RW8YcN6Z1GKLhR6zPnSqrrkSenUWlHpmQ+2f7uLJAhsO7T73ov3mH94hRCpZCfcKWjjRMR2orxT2hF/XkbOm4GNjZXJtWEB+tFXdP69ESvNQK7C4eWT1PpA8T/PwTAHbaTlQplTpxKuOtozkusgWVo9TXx2AvasFSgZCszC+cTnAo1owFGIKO/++klhwV90mh/ov2/dXwcEAVytlqv+o6hWtmGM88v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTW8G+UaBphGU6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcooGN70S/xyynsGEu9vL+xIrJqxZuQaNK/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxH41nPGV3Y6TXEGxY4F/U6OiZeaT/v8OS1YPDP1zxxfagzfIcJGnly/Xp5MwVrdLSb0kfhGIVJ+sp4LB8SnYnkWJuhHwoq8y0TY59MtPd72sG5YOX7gU6yaIaGVqlPEEg8u3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6h2huW/yxIDAlX26L3zEegzDCDFQmIOwZqDXxlkXGyt9L02kUj9eSkTSc3R/HQ5ndZL+814w1rJYvxMuc4I56Tt0B4vwfYTemBHVUdwKRnS5AhoDL61JMcTfs2T3tv7quVVtw4ikZM8K6Vpuqv5jeaMrc4L476B1FUQlm3kjqGg3mJGcwwwWk+2Y8kpni2j7KDB2TZHWspj1HTf8B3+//fS9nAOXMoiDEDCuNVCU7v0plzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZqq4gRFTMbBZCmljTZ2svwcNrWBxWxo0xFiLgDLkBG7TKQ0Q8ygJvXeodoblv8sSAw1EUEp6zcjCy8mcWf19Umjt7qoTfcqOji0UHBZ03U44XM1AU01fCQeR9Vdz5tax2++xi3UxyMm4rBTB4wQehlNOOdoOv5H15gReQpWVmVuKa0pJAd2bC8MlRTbXhVlHrvqzUqO96X8MWjhG4beAcEcooVw963u0KFHXzGmSHaAL06JPml36ZtuWY8kpni2j7KDB2TZHWspj1HTf8B3+//fWxHoMmoJRXKUrlAD3ayx90ETOWt0KBunDb9QuSHDNdeffqlppcnQWarsEsLMzN2uRolwLWZ2eryk7O8kK2eOGaXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZtDnumNqBSSR1IybwRAazvN1CeY/Z888B9DtUqWtbIryjfuoxOiR3gsee83d/nVokYDPG5bJpjnpSOr6+KAx1wMZQd5Xo2t630t3HUvKPCdECSlnj0AdsJAAyrlX0gor6h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC5phREvPgpvHBpIYeA2rj5kBghSAkob+RtcYPplyneb5FgMEVi6IXblsFshSxqvZfeXR15LUBDW8Q9t/s4jiy19tVJMf5fqF0qOH/tgCkP0SSPXFdmWcYdu+YirjGbFRDuYLunBaJS6Paw2LgEagx0MgXkvOp3LB8dgkau2TPXWc77UE666Fn1EAyrlX0gor6tNzUEBQoLQ8H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3LT0/yG2IDtrlZ8IPyDLuv+l9xhXNxWN2T7/oIFKmhD71zhlzDSb1zNzaJy93Vs0Uueqp97NbpllkpR3ILigpxIbsUInXYeDrUSzfIrnC+zZujdN5Dnu+mmbVrC4uDyJS7MoYZt3WznxE/4L/XDFvWlN+pvRdTl2n0wxupMnKBKIimUWc526HfAWCwd+65pMGG6OTbX40yTxj2xuG2LhpaUhsoGwmS2+ixnwlnFDolDkLLT45GzH0Nt4I1zhKJNEvghM3C6Z1tas1KS/zkt0hv6LTgH+PaxEcBYLB37rmkwv1fhyuz67lF7A827fZ/94aN+ksSAq8MbFdKG1DF0/QImghdobMGAZk3v1XY3LF0RncT5vhWUMTUqWp6RM8rmH1B9Yd2pZFfQb/HBCwSJLTjLSGuYI5AJdsfUFAOJ9pO0Om5cZBqGn8kRYLsVzIDLFwyKEsl0DET57boMQ9kCHfkC7YKbRCnvybHkJ+pYPBZSzf48rPx8NWyVM2ong4SIO9K7k1fdUmQuH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LiSreys3v6nxINhgRlnaevm2uLWEhhru+oOllZc3NZdKTk6TnAYGgqFxwAqIx4LVlsXe5TYf8MLJA7xnFayTiUrVt+Te0tbWDf17ZWwanxfSfXLeUnYxOt1QUSEWiq+2JzasixnaPUTKGJVhXHVksriba61mL7BzZH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LsMN/64x7yBQ3jzhesRtAYfKcEnzPHlzUPUV6or0AJU/mm0Q/uaedKEGFwdQab4wcGpNPJuPUpAd0tGcGsxfg0gGLdQeyYI73q47DanIsQyPnq6oodTOP47oStch1nvBHnJbp6P6y4xa0Lg5DcbD+YLNSkv85LdIb6wK5xiV6JehazGz0g/SmcOqTrZEeUCO6Kow69CMRnFRJ9KMULFZWyifQD2F7fPktahfsP1kIF7KQEery/c4fRFQpZ+tnWt5YJqWbEMG9PrJxX2xf0wa4olMzMTd2VbLAHYNbLmfROv+boR8KKvMtE2YCYVHcspp5wgpAf3FqkpZqRj8UXwDNaMjKJEPF85qP0fI81agyzrGWa7jfZDRjpHFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/67stz0ws6fswR+mm+pxTPoBq8OYNNE4kQ8tCPlXzJzGcV9sX9MGuKLNzaJy93Vs0Ven4UCILaaxHEcuJ+RvSwZzysUlAo8iA8T2P1AbHH2o1aAIgdf671gBYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h42aUZ9CPIbWQkH09EyE4A8l6D6ITEIyua0edPGUxp3RqXINbESJTwlr0IpCVjxOwjpKB/H5OuK210UaFJXY4z1xztYHphKvOCCL0/lDTkTEFOhwqLeiYvCGnGZm0K9VJVpf1m+gl7py+GpcnNosxo7sjDe+J1h1K8/fgeW7+hCoMCAsaLkc9sMCLmfIM/UTQLuZWZvb5BOW7GNtU97kTE0INkwj4mslX2su/f6TMXUbH94uSYhWcvOC0NOGP9KsiDpKB/H5OuK2/8Qp1S2I2UD4x4bcEWBzamKlDeM0NhdLnRpRErudjt4tsSOtacc4ZViCACHbNjEqEbixuPsCC6vwcJ2XJkwGgALtgptEKe/JseQn6lg8FlL+bjS+7yrWXq2ZNt296QfyVASjzdxlBBYQmlo6ieCnxLNSkv85LdIb6wK5xiV6JehY7QdkxDLbzSvkwtmFLeT2pxNw5otIq1mr73Isr9tVvxvmUrx3I4a5Pox6NPSU9aWti4k5ZgE8lZTOxVf6qMnZI4vTKyHBGc8+7fMKTrRNy1RWHJYQ/HeHQW6A1k/HcyPhVAuScmh676w9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9FIjp1DOt+yfVx6pd2kExLZTOxVf6qMnZnRPJTL8CXos0Jma1PtADXa+HjxaB4B74AavDmDTROJGnJ6defzt03Ztc8GpGHxkVpWqh0Oh2IWUr5MLZhS3k9vyDTdTph4FFs1KS/zkt0hvHlp94FH+f6NWZoiiFN4qHANr2HJGcwW3sY21T3uRMTdRAJDJae6Vd/dGlsPv+9eby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8QGOw6IbIHiyJcnz0TqBjr8xMjtuZDR5RPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxttYk4SW206ZYK7ii7+OTifBwnZcmTAaA1knBXlhDPOgxWDHBfoP5+bK6DZlaWixPLd0RaCT/cJAD45zU2m2Hr1Fj5+cursX8PU31359fs/CoNfGWRcbK35ciTUmVl2NykxGQ5DlU5Nw63KRBzNiNf58A84lnmGTMo5QHqGJlk0GnJzLtS90jxLPE7sQG274ouqpwpYJv5L3w2/Ho8NRHYy+595hQ5cfiKyEsyd7xrtbn9/gY566w7bPE7sQG274oTnxwVNaDwL4sGONQX4Is0qg18ZZFxsrfbnn+2wcSbtKiXoeTd5sWKDZP4UWWdtb0NV9NkJ3Igcz8UBb5BLcpOmnqd8FFSwZKRN7coAtNOaQG3SJPCawg3j9P7Sa8Wdsuy1M00oFeww50BuqRu5sZqNd93JTxeLn3ZjySmeLaPsqHwix4uxzC7b/dvNaKAYw27lIRdvxVOvvsxQca/NBtNsBJ0u8yqgHdCbZdtKDjvjqT2QQbTYkLPiUUdJ7e6NcGWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPGIQAC7T4b2k2J1zdnhaUWy/BJV9UtiIlbiYvUXNVjIv1q6zn5PSsngV85hUIehQlZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWXsHhv35Z6JyaGok/J+yiliNHGil1XtixJOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHLBSay3l6556Av0V9AN/q/mhX9ZTeqm6mvtnfogXPL9BR8gtxiLTTHi520j/RR5GB1kV2RKeFDdt3IStq4WjC5mT+QyoSnr4KnhhQd5G/Xq5OYiqiWWtCZqX7uWKSzEUpgCTRwHEedg/jSc3R/HQ5ndZL+814w1rJYvxMuc4I56TvGED6cYfjdoNrlzvRZ41imTysGfIDZrZ5jY2T67Es+9y5PpLEgYovSzxO7EBtu+KO07JzE+BWFqy5PpLEgYovQYa77f8vmAHXVkJLM29GloBy84YDvii7/AWCwd+65pMN+blQ0gPYbTKrpOoRCUaq0CTRwHEedg/kv8MthD2qTcwFgsHfuuaTD/xCnVLYjZQKfYXtsj0+pWBBiKYaOep6UOZleiCh30xw0Diqs8KofUkNEPMoCb13qkBz+FUA62mJcRaHwDcIfmaFTnpZKiSGfAWCwd+65pMETWRiWthyW/wFgsHfuuaTCWE52Q8Bi5V5DRDzKAm9d6YWaM3bdub3AfqQUFHfyM4b6IhgkZZbtUkX7Y4xliR00vbnRpTpbAFgIH3KRS8JbE/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNbwb5RoGmEZTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyXgl1F8i6XpCizJKIF/dhGGCozPos+YeqszHT3smYOULy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8bQiwAhHKW1O59yCLLyZKVehYWAR161KjWdq6q+4iv7MalCoso7qGU4npv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWsg1YFRsRCSxYHbaHAM0lMvbtwcZyZxxott1OLXHeZwhgETOWt0KBunJJ3ezUKUQNvZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYcQr3mv20RayDVgVGxEJLFgdtocAzSUy9u3BxnJnHGi23U4tcd5nCGLmaVBt4pSEwrBDmgt5xZth6Mogp1C4PZLPE7sQG274oWGBGj/tq5A7Lk+ksSBii9Bhrvt/y+YAddWQkszb0aWgHLzhgO+KLv8BYLB37rmkw35uVDSA9htPejFaMipzgKu6gnuh/ZnB5aFTnpZKiSGfAWCwd+65pMNgyf6f+E697HN+FpcH/seWIt1VHmsDk5NMX9XZt2jt8HmWvyhCceuj0vBtD6T7gfQnbwKYcJeFtB59eXk9x5vGoNfGWRcbK32Y8kpni2j7KNmcKzFr+wOdv8cELBIktOGXAfejA8TZB/8Qp1S2I2UCYJfFIwDAaCxhrvt/y+YAdeDspfEuZJspAhoDL61JMcUjBpGmAhK5E70Jeje/gCFg4VEE7RIqMX4MqS9j75lvBO05LCnqgWo+X5Um0P+6/oDb9QuSHDNdevasFSgZCszC+cTnAo1owFGIKO/++klhwRvk1cis1RYS7iV9Wgf/ylzokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyA2f5OWNrScHuqzrUUL6jA2CdaBxFayITX7uWKSzEUphMla+A5Ics465fg2pGBtVhdmx6myoLZxRzI/wsCS0pMUKH1RpANeJ/UMc8eAUmMqAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsAyrlX0gor6tVKtg7aPDoVB3ByGK/VBOniK3a0yLM5mRQQDm0+FyW5cCrRrGz4N4rFPwThf4xO935KcFXXGVwNLFN64LgH5CMAyrlX0gor6lBEFqNi1+VNtRLN8iucL7MjXjWux6bcKvfTv7ig9fqTLy5d4EeqX6CLfN8pY7Efqto5s+JQh+GxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LL2V87xYw5PxPIwpq0wN+BArnlhqKJytxmPQQkgisl8tYnYqcZVLiNEt94VFOaCHRBFh+Pi8K3UmNanhf98S2FWXekQSjTOhIqfSQcbwI1BfvCv6L7me0zVphF1C8ucOotRLN8iucL7Nm6N03kOe76d4POnGkg9Q2kBHq8v3OH0RUKWfrZ1reWCalmxDBvT6ycV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/m6EfCirzLRNmAmFR3LKaecIKQH9xapKWakY/FF8AzWjIyiRDxfOaj9HyPNWoMs6xlmu432Q0Y6RxX2xf0wa4olMzMTd2VbLAHYNbLmfROv+u7Lc9MLOn7MEfppvqcUz6AavDmDTROJEPLQj5V8ycxnFfbF/TBriizc2icvd1bNFXp+FAiC2msRxHLifkb0sGc8rFJQKPIgPE9j9QGxx9qNWgCIHX+u9YAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4eNmlGfQjyG1kJB9PRMhOAPJeg+iExCMrmtHnTxlMad0alyDWxEiU8Ja9CKQlY8TsI6Sgfx+TrittdFGhSV2OM9cc7WB6YSrzggi9P5Q05ExBTocKi3omLwhpxmZtCvVSVaX9ZvoJe6cvhqXJzaLMaO7Iw3vidYdSvP34Hlu/oQqDAgLGi5HPbDAi5nyDP1E0C7mVmb2+QTluxjbVPe5ExNCDZMI+JrJV9rLv3+kzF1Gx/eLkmIVnLzgtDThj/SrIg6Sgfx+Tritv/EKdUtiNlA+MeG3BFgc2oHCIkzAlfR/NBxSQN6TXRproTqTSgJi7T4SW4WqIeN7w42NTAAd+hxYUE3gRWQ3UwSNujLFNzqC8BX87v6YGi6nBfQZErDltC+3Rbbl6sYhAP21ycyP1EuNICka9FATM8n0A9he3z5LWoX7D9ZCBeyoSF3Q0r6i7Yr5MLZhS3k9vyDTdTph4FFs1KS/zkt0hvHlp94FH+f6NWZoiiFN4qHANr2HJGcwW3sY21T3uRMTfrzcrVPrhZXcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JpfxAzn1X6OquP9Sg89xHJKnaWEOBQNVw+kKBhVLXR57WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJO01iiGhgjXSLUSzfIrnC+zZujdN5Dnu+mjYMORVM74DT8bwxL0+cok6FvmHqM4CDR6IINe9lwbyGkmZKZxGELEYh1u2jub8VOv+/CmGCc2TWgxwPOa+bCZYDx0oL8iJkpapPPf6YugCL/dvNaKAYw2HyC3GItNMeIffdSuUY3eUAIEa+1M42FMqDXxlkXGyt8cXfiABmXmrekKBhVLXR57qDXxlkXGyt/0XE7CSfEGMOaPeLMwNai7s8TuxAbbvij85NLHmcF+OhlDENuglfWcqDXxlkXGyt/cxy4lNByLKctONaqaynxsv9281ooBjDbE9j9QGxx9qFPAoR7vY9rPIvj8WccgLL9mPJKZ4to+yp1MsumHJiPES06QKnV4AvlU7M7PInj7X4oak6uU6IRXyIIdtx6JhOy1H32wNr5kDzNc+Ti7rrdc99O/uKD1+pNCI7WaAKu7dJSmz4/fohxpieGqWa41vavuoJ7of2ZweTPD8AnDqP83AaZdunTmJQCeyZFt++6kEeUXWaUTU3wN4xEvRHxsgCiYrPJ13IAZWbK4DtNfECHfBj1IlHszAVRv8cELBIktOKFMg/MyhvXb7qs61FC+owPhFKCN6NmkhXAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTRlvRND2F/BT/xCnVLYjZQKfYXtsj0+pWtNd3+Ny1F6zsUOZPthNsLw0Diqs8KofUQzAT0rgnVAh2bHqbKgtnFHMj/CwJLSkxQofVGkA14n9Qxzx4BSYyoB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCwDKuVfSCivq1Uq2Dto8OhUHcHIYr9UE6eIrdrTIszmZFBAObT4XJblwKtGsbPg3isU/BOF/jE73fkpwVdcZXA0sU3rguAfkIwDKuVfSCivq4e+mXVwCkdq6zmgS9boByIu06pKxhrEZkOQKfICwrxXKoosXlmGqZ9m0sv7LJtanH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LvOELWtFYaJAxkL91+oXh1AAHKLhj4L3RjWp4X/fEthWNsdqxvyc0pvvhO+I7b9wotfJjinfBJCFC6f59p0irJG04IHWlU/9ghV7vicnp53OmCrQtaJvfTshI/qd4jaqj5gu6cFolLo8P2j+cq1y7T072JKioWTdeKp+MzEJ5LdcPBufqCD0fWOqodQwHie9KAWDQJ3KBpIOfoAOLnMoIHxp5IRzli53XcV9sX9MGuKJTMzE3dlWywDbhfUs2/G3Ps/fOdT+1++tQgnJmgVSSnmxHoMmoJRXKUrlAD3ayx91xX2xf0wa4olMzMTd2VbLAHYNbLmfROv8TGOzkkr8ididQKgT5HtzBdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDbEegyaglFcrZI63h6kcSjp7z2bM2B/fLTkGSJu/s69jC4OEyxUpTD1zixQ/KIy+/4Cxv9dxY9YX5+7dLcygsMP4ndrcguBFs+ZC8n8a2DmqPaJ1wSxBbGlMzMTd2VbLAOkoH8fk64rYMHZNkdaymPYCZ5+GacpKgNWYnM+lVTIQovhtOCX0ZQFRWHJYQ/HeHpwtxCu/hW/xMVz5kVthoX0wiL+7bR3NuEWsoLROZ2jlYggAh2zYxKrOm4GNjZXJt7K2kkTNq4vgSW9VF0VD+730wxupMnKBKSDlUA99K1Y9xztYHphKvOAIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTQg2TCPiayVfOLXN0jA8St2AHFK8SMRXrSUbMK7NzAG1Ak0cBxHnYP6LfZg5JfrVqNBxSQN6TXRproTqTSgJi7T4SW4WqIeN7w42NTAAd+hxYUE3gRWQ3UwSNujLFNzqC8idZgcKx7PrrZk23b3pB/JUBKPN3GUEFhCaWjqJ4KfEs1KS/zkt0hvrArnGJXol6HRO5CFchwKwtgy5h9MV2thcxnIcGr//zE+8mKRcokneBKgVltCS8e7z6lx23CUV6D3NCN+vBqM4pWqh0Oh2IWXnSv/rNmDxCcCUIkFv5qe3f65pTgrPqZExk8wvrRXYtexjbVPe5ExNnGokgdKcFFMEqBWW0JLx7s+Bd63Gxh9Fi0kWLnusckK6maR0RWksW21F32Il+s4UpyenXn87dN3uqzrUUL6jA1kP0muh7dxwNrGMjGis1QocRy4n5G9LBoVVIPUUpxe0T0KdNXFje9g/AaikY3kVDrsFpaV05J+DrD1oOhUnp8h3gCAXaX5vsU9CnTVxY3vYPwGopGN5FQ5/rmlOCs+pkTGTzC+tFdi17GNtU97kTE2caiSB0pwUU/VvfHslr74/QkP1FgSCfe+Sh6M44dDkoyiZ8hj5jclm4cMmgMS30D0UiOnUM637J5d7pU18snElb/HBCwSJLTjmODb1nyMqpq+REFSqpSZn7GNtU97kTE2caiSB0pwUUxR3ay1jqFIXGiMFB2SyS1/iJpPr8J+9BpTOxVf6qMnZnRPJTL8CXouKEX310ujlTT8BqKRjeRUOf65pTgrPqZExk8wvrRXYtexjbVPe5ExNnGokgdKcFFMUd2stY6hSF9AYj6W7Itm6Y7qmmOMHCY4PsOQj7iMz8mvQikJWPE7CK+TC2YUt5PbTlS26HCAMYu6rOtRQvqMDWQ/Sa6Ht3HA2sYyMaKzVChxHLifkb0sGhVUg9RSnF7RPQp01cWN72JY8nIeo9EwrmzXE6Su/2aivh48WgeAe+AGrw5g00TiRpyenXn87dN3fBSoVCEvSwmZDHMAELV1tdWCm8N7aUUocRy4n5G9LBoVVIPUUpxe0T0KdNXFje9iWPJyHqPRMKz0toaJ1zhYvEWsoLROZ2jlYggAh2zYxKvJMoiRRwIwdeQhhy5rUwxglGzCuzcwBtQJNHAcR52D+wgg/EGv40FCia3IMTTWunisE6EgXdjLiUf7ZcmeleQOJtYcgU9kSUE+8mKRcokneBKgVltCS8e4inCFtEuJHuJtc8GpGHxkVpWqh0Oh2IWXnSv/rNmDxCS7E9Q3b7xJCDles2xfXwOkRaygtE5naOViCACHbNjEq8kyiJFHAjB1pQKpSyhKwaUxXPmRW2Ghfwgg/EGv40FBOQZIm7+zr2MLg4TLFSlMP50r/6zZg8QkXzj+PAVPP1DtJuh+udLyiAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4dBboDWT8dzI4Z6ZIxqv/aCD//YU7iEetkwO89C+dp7iiCL0/lDTkTEQW6A1k/HcyOGemSMar/2gjQ7e1k80Qpni0kWLnusckK6maR0RWksW21F32Il+s4UpyenXn87dN0zulZa2JEEsXbm45U+7JjxdWCm8N7aUUocRy4n5G9LBoVVIPUUpxe0T0KdNXFje9h9MMbqTJygSjtJuh+udLyiAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4dBboDWT8dzI/cQ3XBh/OkTIpwhbRLiR7ibXPBqRh8ZFaVqodDodiFl50r/6zZg8QljjBA/BPmXD8bXe09SFZZkwgg/EGv40FBOQZIm7+zr2MLg4TLFSlMP50r/6zZg8QljjBA/BPmXD0xXPmRW2Ghfwgg/EGv40FBOQZIm7+zr2MLg4TLFSlMP50r/6zZg8QlBPvuJe3pw6e6gnuh/ZnB5MDvPQvnae4oCLmfIM/UTQLuZWZvb5BOW7GNtU97kTE2caiSB0pwUU/dt1RS3EWPzDB2TZHWspj3qbJw4U1eyg5TOxVf6qMnZnRPJTL8CXot5CGHLmtTDGLZZzmiwPIDzDles2xfXwOkRaygtE5naOViCACHbNjEq8kyiJFHAjB15CGHLmtTDGLZZzmiwPIDzPS2honXOFi8RaygtE5naOViCACHbNjEq8kyiJFHAjB15CGHLmtTDGH0wxupMnKBKO0m6H650vKIBYNAncoGkg5LFaicXcUrcKL4bTgl9GUDYbMNM9q7myBGBl/cpTuL5+F6KSl+HPgUn0A9he3z5LQvN66j2wks6CyJ7naQr5WKsJZRsOPth+znUbnqIuKLPBiVRmIubQ7FghCbCqX0xia/78KYYJzZNaDHA85r5sJlgPHSgvyImSlqk89/pi6AIv9281ooBjDYfILcYi00x4h991K5Rjd5QAgRr7UzjYUyoNfGWRcbK38FJly3JZjP2tP/8iyWTRRNPWdlcJT28jVDV/FZgnWOB09ceU6iKyTYIP42M+bJ8nPPqXHbcJRXoiJP9+dI2nl8S1F+P0jKq1VBEW1jlzLTXAU3hE65nfiCmM2sdTEp3ZrPE7sQG274oPwGopGN5FQ5T6DMz1NlKVpY8nIeo9Ewr/xzTeVt3aPdc4sUPyiMvv+Asb/XcWPWF+fu3S3MoLDDc9CSVHsOFPiKcIW0S4ke40fa7AmikQJ57roE+YpEbxWJPnIh31XTupwtxCu/hW/zG13tPUhWWZGJ4IGscaGjGatZfxrEvPYZmPJKZ4to+ygwdk2R1rKY9hGm+ZkHUfsIc1hCg9j6TV7/dvNaKAYw2bW5ec5Qv+Jr4alyc2izGjgiey5VRr1Ja00RGcH1v3HXxBt16gomEmHpWtUmfjM5znwDziWeYZMw4tc3SMDxK3VGGS3zKBooEAI4m8KiSRp+zUpL/OS3SG+UnxRZ+MdRoJRswrs3MAbUNA4qrPCqH1IMDDq8nHSbJdvgvANcb9+3UUZDHTWmw2qFhYBHXrUqNToBSsmnJ7i/SR+EYhUn6yngsHxKdieRYpxk0KAaU9eZuCUJl+r1Ko6+dhSVvWRZXV5gHmKglRiBE3tygC005pKKbTsfrBcDdYVxXqkpAiBhQ1fxWYJ1jgXqvOorn9k/PFQRTQg1Qz1DQPTF9chW+26g18ZZFxsrfExjs5JK/InYsJuhlHhzK0f0UdzWIoAMckNEPMoCb13rAlCJBb+ant0laAgaR8PUc0BiPpbsi2bpMpVL58MJBQkplbS9NCfY4YUE3gRWQ3UxPzE7BF/tUEFFkkXKo1G2E8gH4qB6R0zBfgIcbEXWDExojBQdksktfzYpwOScyB0fAlCJBb+ant4bwjE+jHV/TVVtw4ikZM8IfuZRo+2W5qq2vWgBBQ/Dg/RR3NYigAxyQ0Q8ygJvXegWqkBy0jfPtfR3I6JJgq1fAlCJBb+ant7I1x/CbLlKhIqF1wiBCXpRRZJFyqNRthNuZrYWnCcPB/8Qp1S2I2UCYJfFIwDAaC1VbcOIpGTPCW1s0Cp8ioKFSuUAPdrLH3bXcgvO1H8cRUNX8VmCdY4H/j8B/1GqPK6mao6BFCvHjPwGopGN5FQ7JWTD4txlFzD8BqKRjeRUOn5pkv+29tQDcKzK7Cq19kkJD9RYEgn3vtdyC87UfxxFCQ/UWBIJ975DRDzKAm9d6c937kGh4ONVv8cELBIktOF0f8/aXBDxCqX92jxdeQxNhQTeBFZDdTJDRDzKAm9d6AU3hE65nfiCq8/+Q37fHI3xhZvJSZo0KVsN/yaMKepjQPTF9chW+26g18ZZFxsrfCD+NjPmyfJxigEUXHcYdrmOMED8E+ZcPLcJ6k6ujQLtVW3DiKRkzwt8FKhUIS9LCgkigIsuN5ib3EN1wYfzpEy+aURF738WDo4RuG3gHBHJT8pPAdJM0CmFBN4EVkN1MgqV532rriTf/xCnVLYjZQJgl8UjAMBoLpmFERzayw5NJABgwKu/lQHWVuhlek/rtcXiPEvUIKOM8UrTlyyOsfGfuNHMyXsaGiMSlA/mF8JUVPSuPbkJVcF+AhxsRdYMTDB2TZHWspj1XCGjpkLBfedSMm8EQGs7zkNEPMoCb13oFqpActI3z7Sggprp1pzOUJsavxjE8f2vQxjvZI/ggv1+AhxsRdYMTZbxRTpfpj+x7dU3MEAGKfoi3VUeawOTk0xf1dm3aO3zcKzK7Cq19kojEpQP5hfCVEXU8sh86oYyGemSMar/2gg//2FO4hHrZkNEPMoCb13pjjBA/BPmXD8bXe09SFZZkVx0wAUeChZTUjJvBEBrO85DRDzKAm9d6Y4wQPwT5lw9MVz5kVthoX1cdMAFHgoWUHNYQoPY+k1eQ0Q8ygJvXekE++4l7enDp7qCe6H9mcHljNu2DGegviIi3VUeawOTk0xf1dm3aO3zVT8d49oCi5YjEpQP5hfCVEXU8sh86oYz3EN1wYfzpEyKcIW0S4ke4uHkcmlnxQWDJ9wG+z6DDj9SMm8EQGs7zgqV532rriTcMHZNkdaymPZ+aZL/tvbUA1U/HePaAouWVhqsillAnUvrkcM9BqKDEtlnOaLA8gPO4o+rELtG0r003VqXieKUvZbxRTpfpj+yrznUoCTiNlBzo24/0a7klYNc2V0KXuZpg1MtGwBlMyLZZzmiwPIDzwyrO01hlSvW+juaFIJGf9DxStOXLI6x8yIzN2gOlS4phfQeIFI3IYtSMm8EQGs7zywL2NC3fIJkMHZNkdaymPZ+aZL/tvbUApwtxCu/hW/xMVz5kVthoX9apOpsHMQT+lYarIpZQJ1JMpVL58MJBQgiey5VRr1Ja00RGcH1v3HUcUZQb/mtqGoi3VUeawOTk0xf1dm3aO3xhZozdt25vcDNSC50CghXz5oyoIXeJbFsQGrK531WL7lCTZQJ1f8qvnHPfy+yGTjEo36jxjcHPC/eybMCLpGD5cLpMDZXOk/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwt3gjIEtmkGJUn/JVTdmWYH6MQhTMtwAUK7cvUi1o/TGoQ1R4UUhLal0nUbGM+SWQTJ5r1xzfDXClC+R9yUfoJ0Gb8Ye9mOhQPlT58qADgnayba61mL7BzZoS6qGHjVETaEuQchZ9jhZt7vdQRvfCbXYZnynTrgorqLBsEY5rCh9x+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCxOkt2vc9ZNFnlFEOez9nWfw9MlWEq9WakLp/n2nSKsklM7FV/qoydlVr5987fmvr0iU5SiHsM8OKw8fX1YgZ8q8C1sSUY9by0xnruitJTU5bJUDlhYm1saDEjmNBHtvdlku9oDySbAGrBlQhZxfpnorWK08TVYnHxkX0zvzhHvUnju9lZO76Zvyev56LvzxsdDHspvqm9uLB9zEEX+AOJA2sEq9tJYbONMBLSjtrpl+3eesf3VcPDKVXJAVg6/EOGTEH3p0tn8JRdsuwgPfbBPyKP/VZ589t+6BkjvuNtCbp9dHGgRGuxNq0b+1Nm6gITQAkbMcM7oIWieEcSnZ5R8zbXroVfCi1peR21pKYK0SiFNwRE7HuWjWmH0QnDKBiq+e/QMc4uhnHEcuJ+RvSwYPRixkXcRrrPGwAIE0kyRpvtk5SKcFdH8Remk6DZSIjWYV88QK4B2gXyFnNDgdSTS/Z4DvPop7lsGOdbJ9JQtTe0JhOR+lUna8C1sSUY9by+hHfjmtfNSBFatmMisMCcR0wn3TSYmobycIi9SsM9XnTXpXGOsNPQzXyJL+JiGIPs/PeAffmo0bBCWHW9TV9zImLJ4lIfX4RdaYfRCcMoGKhMZJHv/A5o84HXb23V+jBWJponaqEc2oUH1h3alkV9CPTG6BNO9Ckkodg7Lws3CNS+NUGOoRoh+Yfi1r5vHGG3M3DQj1aU0b48GcdeSei/mFZQgKai5debHNfQ6zw2yNaBkzWVro+7h3kId/dA1X4y6sBcF0uLJIMHkDY6adzjQo5XEdke9YbHfUZYz9bG/O1ph9EJwygYpr7aX3qJ0uG+C7noJyhgLOQ14+UEyrRVl7A65MVBcQL7XEk8ytQS//C3Nu2Rn+jNSVM2ong4SIO9K7k1fdUmQuH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LiSreys3v6nxINhgRlnaevm2uLWEhhru+oOllZc3NZdKTk6TnAYGgqFxwAqIx4LVlsXe5TYf8MLJA7xnFayTiUrVt+Te0tbWDf17ZWwanxfT56ae3iXlTjrwLWxJRj1vL1yrzlUr7y8ijY1EepObcPGN05VmOvf0BrbMRSrTpupWcFmUMNY9FzR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/X0mFXQGDwUBfxxgLW/DpkietI52dApanS0ZwazF+DSia1Dv3sAhvWmfnNRqgv4UiYRGFaybmRCXz4emIpYW9m3eLBqrjPtBbH34oYJdprZPm/Yg5QMFuiaaX7DoqNeJ0PVRIjpHmGpw17qXdPR0NQbqH3qqgQ2LS01RLgS3JOs6y3ZOsQka3gc62LjIBAnGcBYLB37rmkwSmIo5j8yCJGJWbp1N0Euijojjbuvm8H6yocNttbci0KMw98LvuzZj4G3eXrLjNqtT/ckQex2loBq5rJdx2fk7texpo4/tQWKwFgsHfuuaTB2Gzbvha9BMobvWnk0VbzsnahTAyYvWqD6AkhmLx3jRzjCgNQSVdmTE+lrgtFc1cp3bR4eTzIU92+0363IHGe1GgBTqhBvzYjAWCwd+65pMKvvciyv21W/bYiDHSwIOaylP4b2LdZ/hKYGTwol37VOTc+2J5/NvU+pkEbAltJTXapTfN5kPhN94Pegtv9cRAr8C4QBpeCSiFwNT4Su+gmAv3T+/Q7PTTm0LZ9wrayIZxYZ/vTCkqXK+3UCQ6/Os9obqH3qqgQ2LS01RLgS3JOsx3Ki6aiOBv2pCJ+J5hgaSDSxDyF80OIRSmIo5j8yCJGJWbp1N0EuiuXRJfQwnoTEag9o9V03daeMw98LvuzZj4G3eXrLjNqtT/ckQex2loDQx7Kb6pvbi8GNJjwzUNz/0VSkZrNX7XR2Gzbvha9BMobvWnk0VbzsJg4X2jwj/SP6AkhmLx3jRzjCgNQSVdmTE+lrgtFc1cp3bR4eTzIU92+0363IHGe1pf01i22B/oPAWCwd+65pMKvvciyv21W/bYiDHSwIOaz/pv6l3T5NQ6YGTwol37VOTc+2J5/NvU+pkEbAltJTXapTfN5kPhN94Pegtv9cRAq8cPVGWUIKGlwNT4Su+gmAv3T+/Q7PTTn4BDvHgvMMXRYZ/vTCkqXK+3UCQ6/Os9obqH3qqgQ2LS01RLgS3JOsvikGWcuEr9RJY1oJDRFNuMBYLB37rmkwSmIo5j8yCJGJWbp1N0EuiunyFXYn8eaxag9o9V03daeMw98LvuzZj4G3eXrLjNqtT/ckQex2loAqQrnO+n4kyMeWVQfKpR9bwFgsHfuuaTB2Gzbvha9BMobvWnk0VbzsAd3rTlIz+UH6AkhmLx3jR9r9NS/2J1eOxB0dI1EaCdwuxinGJGN236O79lRo1cqWltgMhxD5lKmFGLYQaJIhbiMDhSXtJ91ajb9uZP+VgrrUYqY5bFqnIkFU5NHvR+RnIwOFJe0n3VqNv25k/5WCuiTgV6rS7d/LSh2DsvCzcI1L41QY6hGiHyvkRTUBtiP4ucAvtnCyRGSZtOaV3rbA4xvNBLPWdLQgvcyFVQU3e6aYXXVd9VLHGwW+NPo/SQQpc09lhEMC2PHgu56CcoYCzit4gBb86Z2AaJ/jC0zHDQZvtN+tyBxntfo/jM6gzEKMM2166FXwotbiMt/zl0xLMu2Nhkx7Il6t3U2mo9otigsFvjT6P0kEKXNPZYRDAtjx9YIq0VoAHSkHMXRy7pTpvWif4wtMxw0Gb7TfrcgcZ7VrV+iazSP1ouPBnHXknov55oGai5KquwzQx7Kb6pvbi+Zk9oc9lVE3UK0oaoualNpY8KtFTQ+0WkbBRayCAgO/5YpRAZNgy6sO/D03hOUZEdDHspvqm9uL7X7SipdtZo6BhSuEFw+dszNteuhV8KLW4jLf85dMSzLtjYZMeyJerQtfmmDOkG/VBb40+j9JBClzT2WEQwLY8Si+G04JfRlAucAvtnCyRGTXv5KguLILW+2Nhkx7Il6t9fHb6vyOOIELcNA95PIA4Zm05pXetsDjkmSQ+YwOqlJvtN+tyBxntR4+JH6FN75a1ph9EJwygYqExkke/8DmjzgddvbdX6MFBzF0cu6U6b3693WYPdydBVfLc8kWuFtE8wHkuysYjDzxsACBNJMkaQXQltuMiEX2V8GFf2CafJBQrShqi5qU2ljwq0VND7RarCcYEYdtdGCo5SojrNIEZaG+LHmCEkmKyfBCfkcxo5TYGAPhUE5iyVB9Yd2pZFfQ0k2Sa0dUsXDEeHcz/uXwWUodg7Lws3CNS+NUGOoRoh8oq19RUhiKziwTHkGQLJGKewOuTFQXEC+1xJPMrUEv/2bo3TeQ57vppm1awuLg8iVmqNNMdXpyChSVTkv8zn4wH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3LQVlKofHHLJtrrWYvsHNnIzsey4CsrGdYqBAckRbuav5vX7RwU2rinlHrBC07kStu9J5gHlaVqiqr4MCPcf7rXUMUP9aNywiw3SPTlUXbzjkGwgGfgT6nJ8+Ic1EikCCNeNa7Hptwq99O/uKD1+pO0M8u2CbUGI9o5s+JQh+GxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LL2V87xYw5PxPIwpq0wN+BArnlhqKJytxmPQQkgisl8tYnYqcZVLiNEt94VFOaCHRBFh+Pi8K3UmNanhf98S2FWXekQSjTOhIqfSQcbwI1BecDP+1jQ0/h7dx6Orf8695LKBmmOe67LLXZxhq9dA2FyMDhSXtJ91aWsxs9IP0pnDqk62RHlAjuiqMOvQjEZxU3Y+Cc4beCfOx9+KGCXaa2WjEkxEgrtYKKp+MzEJ5LdcPBufqCD0fWOqodQwHie9KAWDQJ3KBpIOfoAOLnMoIHxp5IRzli53XcV9sX9MGuKJTMzE3dlWywDbhfUs2/G3PNORLbik88sawoLfxgcs7Ctu8DVkEddD7DGu0313so38BYNAncoGkg5+gA4ucyggfFUquKxLk0JQwICxouRz2wyCL0/lDTkTEKFF0eiA5/9zBNg3LDLX2ZQFg0CdygaSDksVqJxdxStw4HXb23V+jBW1F32Il+s4UUjkQ+6AMoW++eXiXuWvz15TOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMPf0h/5H1vCpr33vQVFlWnA3HO1gemEq84Ai5nyDP1E0C7mVmb2+QTluxjbVPe5ExNR2fVmEyqvVOjg5Fle8oUIiBkf8+t9vrDpWqh0Oh2IWUzXPk4u663XPfTv7ig9fqTQiO1mgCru3SUps+P36IcaalMB0zBvqsUFLZSiKZsDMReCQMHKUbNsNWZoiiFN4qHr1AgXgzKfvVYggAh2zYxKrOm4GNjZXJt/9ZUxD39Lv9vtN+tyBxntfH7ZVE6QP3vXgkDBylGzbDVmaIohTeKhwDa9hyRnMFt7GNtU97kTE0INkwj4mslX2su/f6TMXUbH94uSYhWcvOC0NOGP9KsiDpKB/H5OuK2LwcRUQo+Yt9QxUmdfALdqJ8Cjiccf5MnIGR/z632+sPVmaIohTeKhyUGtg9pP9WQ7GNtU97kTE1HZ9WYTKq9Ux3MlbIhFGnUN4hp1u2WpNvfkflPppAGqq62IOawTKQ9lM7FV/qoydkji9MrIcEZz+bV9EPoBEz3VFYclhD8d4cGPUiUezMBVAyUaO8yXW5oPeD4ApjS4JkDDeRSg0Zq8XHO1gemEq84Ai5nyDP1E0CVmcrNSWnKPmvQikJWPE7COkoH8fk64rYvBxFRCj5i39DHspvqm9uLesB/gtsbSATYLGbIXy7cnaw9aDoVJ6fITuyUW/8exDjL57bRgHBMzL8RVDUv1DzkQe0wZoVXbNsD5eTr4S7FDiBkf8+t9vrD1ZmiKIU3ioevUCBeDMp+9ViCACHbNjEqs6bgY2Nlcm114MgsNq16Rsdyoumojgb9qQifieYYGkjdmcWW1yV4t3HO1gemEq84Ai5nyDP1E0C7mVmb2+QTluxjbVPe5ExNR2fVmEyqvVMdzJWyIRRp1E3mPOZwD+gIiQsW5WB6RqxZ36WaPk0oGyXoPohMQjK5rR508ZTGndHwthhZvKXBo2vQikJWPE7COkoH8fk64rYvBxFRCj5i39DHspvqm9uLwY0mPDNQ3P8rKLIYC7rZmqw9aDoVJ6fI6m3ZnKEGKjxYGTbi9rEg4uHDJoDEt9A9dWTJ1KHwjnoU+ZOe7mk+Se2Nhkx7Il6t+0r1YM0jh2QgZH/Prfb6w6VqodDodiFlsUJYN6b3gXtij/6YhOIJtm+0363IHGe18ftlUTpA/e9ipQ3jNDYXS50aURK7nY7eLbEjrWnHOGVYggAh2zYxKrOm4GNjZXJtdeDILDatekbHcqLpqI4G/f1uL/13Vq6xUB604GCKmTIgZH/Prfb6w6VqodDodiFlsUJYN6b3gXvds74XZpNAelfLc8kWuFtEbCo3ZqFJh3qsPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPXVkydSh8I56i9PnsM5wBWqTaQ9m61ELmyw3ojjDp5pSlM7FV/qoydkji9MrIcEZz+bV9EPoBEz3THuAGfcsPKDDUgxQnnMPO8lGkbQ9GqeDaSZkpnEYQsTAC8/lj5kKjVrgSNBvfq0OZf11sV/DEVQB5z3GLRBwn2kmZKZxGELEKGElgcvbLTpBboDWT8dzIw5LqLGRo1LF9215oa1VU9wUiOnUM637J6s4z1+Qw2XUsDrAXOB2kKidGlESu52O3o9ryFAi7Yx2WIIAIds2MSryTKIkUcCMHQSb5EBsmCp8Q+o+Dva+e3vNzaJy93Vs0RfzvLOuA1LyupmkdEVpLFttRd9iJfrOFPOqxRniGbE2ImO2CPc/mOzCCkB/cWqSlhSI6dQzrfsns2nLIpNLN9YBYNAncoGkg5xqJIHSnBRTEE70Xf2PEt2sPWg6FSenyPx9q8/kPpTrQW6A1k/HcyMvBxFRCj5i31DFSZ18At2onwKOJxx/kyeUzsVX+qjJ2SOL0yshwRnPPu3zCk60TctUVhyWEPx3h0FugNZPx3MjLwcRUQo+Yt80p4gZf3LrG2KUtlXKCXQbMDvPQvnae4oCLmfIM/UTQNqTlZfCjsNca9CKQlY8TsIr5MLZhS3k9gZNgkwu7nTyvxFUNS/UPORkDlE+6f2friJjtgj3P5jsnRpRErudjt64TI2SdkRWqFiCACHbNjEq8kyiJFHAjB3u0V+ntFmUQQyUaO8yXW5oPeD4ApjS4Jmti4k5ZgE8lZTOxVf6qMnZI4vTKyHBGc+ia3IMTTWunlRWHJYQ/HeHQW6A1k/HcyMvBxFRCj5i39DHspvqm9uL7X7SipdtZo4AJstaZSYTn50aURK7nY7epa/XkEGd4zccRy4n5G9LBoVVIPUUpxe0xvZrfAFJ45xij/6YhOIJtm+0363IHGe1pf01i22B/oMwO89C+dp7igIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTZxqJIHSnBRTyeCHG2BJ/92qU3zeZD4TfeD3oLb/XEQKgUQtcBZ0XUOsPWg6FSenyOpt2ZyhBio8WBk24vaxIOLhwyaAxLfQPRSI6dQzrfsnyVJ1EdJtC7LHcqLpqI4G/fxoyKKxJMhHdubjlT7smPEBYNAncoGkg5LFaicXcUrcDhqdZrFVIZ1UVhyWEPx3h0FugNZPx3MjLwcRUQo+Yt/Qx7Kb6pvbi3rAf4LbG0gEDWM66eBU1m3CCkB/cWqSlhSI6dQzrfsnyVJ1EdJtC7K+KQZZy4Sv1FFUgFr5JEchrD1oOhUnp8jqbdmcoQYqPHPT6yNUvnsS4cMmgMS30D0UiOnUM637J8lSdRHSbQuyCcW7fYl+tp7SAARLZedAlAFg0CdygaSDksVqJxdxStw44KuW0tEdOm1F32Il+s4UpyenXn87dN0U+ZOe7mk+Se2Nhkx7Il6tjR8mHG6A3h8NYzrp4FTWbcIKQH9xapKWFIjp1DOt+yfJUnUR0m0Lssdyoumojgb9oAba6pFzewQwO89C+dp7iiCL0/lDTkTEMsZX46ljmMxwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyOYkaacOUfl99O/uKD1+pO98Sxv08jFm3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTaB4D329Ctmto3dJewHB6Xgsie52kK+VirCWUbDj7YfugqjQZKQWKCvdTx/dhpm0gDqFeXIjVfUOP4r3tD8ykX0WyOTE2UwNchBdE73GNEXhycn0fczLPWCqiwbt8jjHafiqJ59OKOgAfILcYi00x4gezedDC0hirGB6jBl007Ic8OcUvtKIUaMtTNNKBXsMOlmu432Q0Y6RVtzG8TrCT+OFRRTcQx2eSTPi9BLwlG1yiXoeTd5sWKMEEv59HAnhFKFF0eiA5/9yI4P51zuvVDcBJ0u8yqgHdyvZhKluyThmT2QQbTYkLPm55/tsHEm7Sv9281ooBjDZ1TGReX5j+UOZayS/+pXGLiJP9+dI2nl8aYZi93EU3gCGflt/b2E+Npycy7UvdI8Rg1MtGwBlMyPRyTtTkYoh2NyB9cSD20sTJRg+1OgVe9QxQWILR7ZC4LQaIu5snXiLTRVBzMyUZ+HskI+AeHuzXqDXxlkXGyt8o6rJBXJOT+UbY90Xs8kxeGNMqQk807ovy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+VJL61xzk7W6wm2ChLjB6jQIRdnHrv9Vhi6d0PiQFatWfA9bzqHAVIRAvDiKK56g4vL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHTUfvZh6UJ3Rt7Fd27J/y61jffj5tpBkjyZ4JHOwzPVry/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMgYSMGKOKkTQsteX/pLtfRFxhDJnfvPqGhYWAR161KjWdq6q+4iv7MalCoso7qGU4npv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWsElqjsKdbEtm7YSnN0T/tJmXf8k5ctsyCCKaqVvfQbO1RCWbeSOoaDeYkZzDDBaT7kcehumNwmTVS6d5Mkv2EXL3MhVUFN3umZKLh5o22mDQ0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm3LoB5kgu0i5cdyoumojgb956FUpyEGrT1sZx8IuFFF+Gz8/3OvySf9oj0QCQIThh6DVgVGxEJLFhT5k57uaT5J7Y2GTHsiXq3hSEvQqGknf3rIxh/8TeA3kNEPMoCb13oTI/0gR9Cjy03mPOZwD+gIr767Cqo0gKo+PtLIAl07z2z8/3OvySf9oj0QCQIThh6DVgVGxEJLFhT5k57uaT5J7Y2GTHsiXq2NHyYcboDeH5ZWH16/+TeYenPTtAYOt1bLoB5kgu0i5cdyoumojgb9qQifieYYGkgZQzX6IVoHLyVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3y8HEVEKPmLf0Meym+qb24vtftKKl21mjr5zxI7TXmNiUQlm3kjqGg3mJGcwwwWk+5HHobpjcJk1Yo/+mITiCbZvtN+tyBxntdcmVs73QfVL9qoHINnqNTQT1zWClEYtH4XLjiOTjsUyIfsv+SkPX9yqU3zeZD4TfeD3oLb/XEQK/pW/a4n9rIE0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm1cF9VXEWYWH6pTfN5kPhN94Pegtv9cRAqWVh9ev/k3mHpz07QGDrdWy6AeZILtIuW+KQZZy4Sv1DBAJnLgpg8d70gkrfDjVa74zSrs37+G7cugHmSC7SLlCcW7fYl+tp7bma2FpwnDwSVfbovfMR6DMMIMVCYg7BmAbAWZCTK1uA/XOJfyF1XDY3sCEo28Fct8J/VrU9hea2suxKHYfDbF4SSlnUTC2QixQlg3pveBe2KP/piE4gm2b7TfrcgcZ7V6W6opwjLgsHrIxh/8TeA3TawgfeifQ7oO6D5O6paRf+u4Cyfgk0kVqDXxlkXGyt914MgsNq16Rsdyoumojgb9oAba6pFzewSNEGZBBfPwZag18ZZFxsrfdeDILDatekbHcqLpqI4G/eehVKchBq09xZyvXGDW/ohJz5ieEfkatKHZ/hv0mGyKCmPOkKxcp2ThJKWdRMLZCC41I5xgCX1epxpVKQ/Ih0L6ujgmFGIVYFrL2xd/GFnka2fhra+8NHrFcK2ax6q2C1A+qUgeAqkYKv9M4v1MTEgYa77f8vmAHRJao7CnWxLZu2EpzdE/7SZl3/JOXLbMguRAcXxW0+nAYKWMQYJDY4W7YSnN0T/tJnQzVG98nA17S2XdYnk0cFi4FghI7HWfJcBYLB37rmkwy6AeZILtIuWCeh85CtM9nj7BHqWnJadcx2kL9IpC3wpgpYxBgkNjhUEttyJGw3pnW7MWQAosb2kWsoUu/xdHpBhrvt/y+YAdeDspfEuZJson4D6LlIe4eL8RVDUv1DzkZA5RPun9n64IcPWT5/CpcsBYLB37rmkwmoGd7aFyHqG/EVQ1L9Q85GQOUT7p/Z+uUpPs1aFBV0dgpYxBgkNjhQyUaO8yXW5oPeD4ApjS4JnzdVE5FdGTW8BYLB37rmkwsUJYN6b3gXtij/6YhOIJtm+0363IHGe1to/m2LQIDAM1pD7/K3chi6g18ZZFxsrfeYj6+rMrrz2pkEbAltJTXapTfN5kPhN94Pegtv9cRAoVYOdbLHgXFxhrvt/y+YAdElqjsKdbEtkMlGjvMl1uaD3g+AKY0uCZRy2f5UTOYcvE9j9QGxx9qLvgZd8LOYTD0Meym+qb24vmZPaHPZVRN7Om4GNjZXJtwFgsHfuuaTB14MgsNq16Rsdyoumojgb9/W4v/XdWrrG4AEdaRSslrBaWMcaIPh6mwFgsHfuuaTDfm5UNID2G04KtkKCkTL9oTeY85nAP6Ajp0e1fN6J/KDDNqeIX8uuxwFgsHfuuaTAh+y/5KQ9f3KpTfN5kPhN94Pegtv9cRAoL0kMNOVInXwQYimGjnqel40RjUDgKerVN5jzmcA/oCOnR7V83on8os6bgY2Nlcm1ay9sXfxhZ5Gtn4a2vvDR6d20eHk8yFPdvtN+tyBxntdcmVs73QfVLaFTnpZKiSGfAWCwd+65pMBMj/SBH0KPLTeY85nAP6AiJCxblYHpGrFG5mylj9mW/c9TRPet/+tSSZJD5jA6qUm+0363IHGe1Aqaz/qoHd1MYa77f8vmAHXg7KXxLmSbKJ+A+i5SHuHi/EVQ1L9Q85EHtMGaFV2zbYR5vFgB1R8KoNfGWRcbK35HHobpjcJk1Yo/+mITiCbZvtN+tyBxntaX9NYttgf6DAOV3wiTp0ctmWjhhCW9KLr8RVDUv1DzkQe0wZoVXbNslEGorDWkjPMBYLB37rmkw/1g4hWW9x0lP9yRB7HaWgNDHspvqm9uLwY0mPDNQ3P+cACJur6Gmi8BYLB37rmkwmoGd7aFyHqG/EVQ1L9Q85B5UBtqgp+AChfifdVlpUAbE9j9QGxx9qLvgZd8LOYTD0Meym+qb24tmjDZTQ1z/R5DRDzKAm9d6Ovzm46oTw3EdzJWyIRRp1E3mPOZwD+gIAtjXpwrEp0EGu6c5zLcN0Rhrvt/y+YAdeDspfEuZJson4D6LlIe4eAeEOBi+zsIg7wALy2dhRIlL/DLYQ9qk3MBYLB37rmkwLwcRUQo+Yt8khEjm/Hlc4gnEQQWLv3LMbnn+2wcSbtJPv6nUSjX1VnPeoGGTEiybCGbOvvwjvd7AWCwd+65pMN+blQ0gPYbTgq2QoKRMv2jJ8EJ+RzGjlKyAcjPH76sAwFgsHfuuaTAh+y/5KQ9f3Ertvcs0aR2sp9he2yPT6lYEGIpho56npeNEY1A4Cnq1yfBCfkcxo5Soezryhl+be8BYLB37rmkwqmUVqj/F4mpaxkgIwqojrxhrvt/y+YAdmgQ4Gj4rGfKaVipXwnM01L2rBUoGQrMwwWzRfs2dV60ASlQboJTlvmsezOrWWHiuajkcM0HTJMWiAiNHs4agN4V/WU3qpuprKp5f9Gby4v/zIf05yUeyoJdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JivCPr9uV7dXxvYng4NQZh7+f8516XPrN3AjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTJOt9hnGoEMo+/KHRE1bGQ4V/WU3qpupr7Z36IFzy/QUfILcYi00x4udtI/0UeRgdZFdkSnhQ3bdyErauFowuZk/kMqEp6+Cp4YUHeRv16uTmIqollrQmatgyf6f+E6977TEbKty64h5s/P9zr8kn/aI9EAkCE4YeDCuNVCU7v0plzGbP0AALTKfEb3WHMzLgUWPn5y6uxfwRO5zafLLM3OYiqiWWtCZq2DJ/p/4Tr3vtMRsq3LriHmz8/3OvySf9T/rhEC/IRTB1LdCzU76Qy2Dl4rua9QPWD9q6x3W9XkZ55MOmMyTbz5acAGSF9jAb2K6hMdSPTRzY0wuCgNaK7EzS7liLaznlfID8LDeXPCqkBz+FUA62mMlS7qLiPpHRtuoKi9MTT9jRTLU8Zxa8Cxhrvt/y+YAdg1YFRsRCSxYHbaHAM0lMvalMB0zBvqsUYNc2V0KXuZoYa77f8vmAHXg7KXxLmSbKJ+A+i5SHuHi8C1sSUY9by1f1cPx4P1yKAv459fq8YF/AWCwd+65pMHvZzLAQalyc40RjUDgKerUSNujLFNzqC6GKrG3ZkjsR/RaoyA1QnOeRk0NhlNeeXbwLWxJRj1vL3T3qOLnPAV2Q0Q8ygJvXejr85uOqE8NxlFB0GFWft+gbzQSz1nS0IL3MhVUFN3umqeXL7fv9V++Rk0NhlNeeXYYhBxte8o9jmkshN3mk+8L5XtoTGR/qvsBYLB37rmkw/1g4hWW9x0lP9yRB7HaWgNDHspvqm9uLJVc6h4vwlzNL/DLYQ9qk3MBYLB37rmkwSPZCjBZnXw14ctCNVy74yO2Nhkx7Il6tNgIPx54TCsyRk0NhlNeeXb8RVDUv1DzkZA5RPun9n66vZqxD/bSsix5lr8oQnHro9LwbQ+k+4H2TZF7KdNBLS+2Nhkx7Il6tWInLwkIK3qxL/DLYQ9qk3MBYLB37rmkwSPZCjBZnXw14ctCNVy74yO2Nhkx7Il6tHV/PMdNMKE8sIDAL8qWdv8dyoumojgb9/W4v/XdWrrHMj7olA8apYR5lr8oQnHro9LwbQ+k+4H2TZF7KdNBLS+2Nhkx7Il6t5DGaDvoF195LX71Z4PNWdMBYLB37rmkwe9nMsBBqXJzjRGNQOAp6tU3mPOZwD+gI6dHtXzeifyhfWADTFbkpBAyUaO8yXW5oPeD4ApjS4JmrK7S5UHe/g6g18ZZFxsrfeYj6+rMrrz2pkEbAltJTXapTfN5kPhN94Pegtv9cRAq0Og3dc5y96EjBpGmAhK5EOvzm46oTw3GUUHQYVZ+36JJkkPmMDqpSb7TfrcgcZ7XFZEjbsFrpcTMhzbqoZRtwx3Ki6aiOBv38aMiisSTIRzjIco5X68CHwFgsHfuuaTDfm5UNID2G04KtkKCkTL9oTeY85nAP6Ajp0e1fN6J/KObjL9dqhg2IwFgsHfuuaTB/SH/kfW8KmmZaOGEJb0ouvxFUNS/UPORB7TBmhVds24BtXQpidgShFPmTnu5pPkntjYZMeyJerRVacDS94VfdTKVS+fDCQUJay9sXfxhZ5Gtn4a2vvDR6d20eHk8yFPdvtN+tyBxntUW22TXrMSR6aFTnpZKiSGfAWCwd+65pMNgyf6f+E697u+Bl3ws5hMPQx7Kb6pvbi2aMNlNDXP9H/FIPAS8qijeqU3zeZD4TfeD3oLb/XEQKjHTsMp+AvS8Ya77f8vmAHXg7KXxLmSbKJ+A+i5SHuHgHhDgYvs7CIO8AC8tnYUSJS/wy2EPapNzAWCwd+65pMEj2QowWZ18NT7+p1Eo19VZz3qBhkxIsm3BfGLnKLtKWLwcRUQo+Yt8khEjm/Hlc4rHWVtharg3AwFgsHfuuaTDfm5UNID2G04KtkKCkTL9oyfBCfkcxo5SsgHIzx++rAMBYLB37rmkwf0h/5H1vCppmWjhhCW9KLlAyHSH9z2AQ69gUGto0sq0zIc26qGUbcAnFu32Jfrae8gH4qB6R0zDAWCwd+65pMKplFao/xeJqWsZICMKqI68Ya77f8vmAHZoEOBo+KxnymlYqV8JzNNS9qwVKBkKzMMFs0X7NnVetAEpUG6CU5b5rHszq1lh4rmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa27kaxZD4JNmB6dMgmnMCSPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdn+wichJZ+QNn+Tlja0nBBjpehuhoK9LE2a0fTHQJ6zEyWvr3wayELwcRUQo+Yt9QxUmdfALdqErt3SYftrlRXBfVVxFmFh/U1aiDD1ZpbuyLfjfLOY7bCIWowqdSWEEvBxFRCj5i3zSniBl/cusbYpS2VcoJdBsZhKx9mlr7aRT5k57uaT5J7Y2GTHsiXq0mwYphmOBmEjMhzbqoZRtwx3Ki6aiOBv3noVSnIQatPSiVgq1S7EspLwcRUQo+Yt/Qx7Kb6pvbi+Zk9oc9lVE3/FIPAS8qijeqU3zeZD4TfeD3oLb/XEQKlRe277/u6FHL57bRgHBMzL8RVDUv1DzkQe0wZoVXbNu4nAJq9UTZAhMj/SBH0KPLTeY85nAP6Ajp0e1fN6J/KBeAIzzXgm7ZdeDILDatekbHcqLpqI4G/akIn4nmGBpIQmJSyNHRScMvBxFRCj5i39DHspvqm9uL7X7SipdtZo6GiQDOZX86LR3MlbIhFGnUTeY85nAP6AiJCxblYHpGrC55r8llU0/ZFPmTnu5pPkntjYZMeyJerfXx2+r8jjiBCxfiU/ScNtovBxFRCj5i39DHspvqm9uLwY0mPDNQ3P8CTv6eBnWO22KP/piE4gm2b7TfrcgcZ7VFttk16zEkehmErH2aWvtpbN0KekdCEetz3qBhkxIsm+YrymY63GyybN0KekdCEetz3qBhkxIsm9p1curPH7kXdeDILDatekYJxbt9iX62ntuZrYWnCcPBLwcRUQo+Yt8qQrnO+n4kyB8aJLTW+dk0am7iEwbcIGsNfP/1CBud8UqGxIKRu9TPcLpMDZXOk/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwt3gjIEtmkGJUn/JVTdmWYH6MQhTMtwAUK7cvUi1o/TGoQ1R4UUhLal0nUbGM+SWQTJ5r1xzfDXClC+R9yUfoJ0Gb8Ye9mOhQPlT58qADgnayba61mL7BzZMT65WrDAzbyRXbkAjgjF3prZsMI5If2PhAev1DEE6KLrB3HOvAkqn4sGwRjmsKH3H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LE6S3a9z1k0WeUUQ57P2dZ/D0yVYSr1ZqQun+fadIqySUzsVX+qjJ2VWvn3zt+a+vNGzsQ7/B5p9Qw2GSyqIWv4kAEDsXn9JOtWHT9AV0+9AxkL91+oXh1Fsnph1GMPMA55MjocTbh2KCDdow07H8h7H34oYJdprZCnCHVKTy5iU0bOxDv8Hmn9dnGGr10DYXIwOFJe0n3VojbPf3JibGS+8K/ovuZ7TNohZyDHoAx1QSNujLFNzqC8BX87v6YGi60XZRHlMHmscqn4zMQnkt1w8G5+oIPR9Y6qh1DAeJ70oBYNAncoGkg5+gA4ucyggfGnkhHOWLnddxX2xf0wa4olMzMTd2VbLANuF9Szb8bc805EtuKTzyxrCgt/GByzsK27wNWQR10PsMa7TfXeyjfwFg0CdygaSDn6ADi5zKCB8VSq4rEuTQlDAgLGi5HPbDIIvT+UNORMQoUXR6IDn/3ME2DcsMtfZlAWDQJ3KBpIOSxWonF3FK3DgddvbdX6MFbUXfYiX6zhRSORD7oAyhb755eJe5a/PXlM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw9/SH/kfW8Kmvfe9BUWVacDcc7WB6YSrzgCLmfIM/UTQLuZWZvb5BOW7GNtU97kTE1HZ9WYTKq9U6ODkWV7yhQiIGR/z632+sOlaqHQ6HYhZTNc+Ti7rrdc99O/uKD1+pNCI7WaAKu7dJSmz4/fohxpqUwHTMG+qxQUtlKIpmwMxF4JAwcpRs2w1ZmiKIU3ioevUCBeDMp+9ViCACHbNjEqs6bgY2Nlcm3i4XgOVDPh/08MDQF/7jEYzasixnaPUTISW9VF0VD+7x3MlbIhFGnUEjboyxTc6guwT8X/oXxNlWKlDeM0NhdLnRpRErudjt6Pa8hQIu2MdliCACHbNjEqs6bgY2Nlcm114MgsNq16RoJ6HzkK0z2ePsEepaclp1zWJYkQfLASlaw9aDoVJ6fI6m3ZnKEGKjz8BVvBnRzJscLg4TLFSlMPsUJYN6b3gXtij/6YhOIJtm+0363IHGe1bHw/TgDTHhmx5cebPGCxzEDhRVcgwpvj7GNtU97kTE1HZ9WYTKq9Ux3MlbIhFGnUTeY85nAP6AgkUVqGJt3PInHO1gemEq84Ai5nyDP1E0AH0c/sN122PuxjbVPe5ExNR2fVmEyqvVMdzJWyIRRp1E3mPOZwD+gIAtjXpwrEp0GPaJ1wSxBbGlMzMTd2VbLAOkoH8fk64rYvBxFRCj5i39DHspvqm9uL5mT2hz2VUTde8gHhuo5/I1TM/LO5RPzdCa1xN53e85ZtRd9iJfrOFFwX1VcRZhYfBdCW24yIRfZXwYV/YJp8kEIUGh1sl2hPdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDy+e20YBwTMxQMh0h/c9gEFkP0muh7dxwseXHmzxgscwWiW/fZWFdbOxjbVPe5ExN4UHRF2FP0mw455NQelIqO7wLWxJRj1vLV0pGt5hZIZ3/EnNF8wz1b6Ic/j4NtRsPsNMwfWlh5XL8ernI8tWt7mbo3TeQ57vp3g86caSD1DYNs+RMmCND0sb2a3wBSeOcYo/+mITiCbZvtN+tyBxntWx8P04A0x4ZlM7FV/qoydkji9MrIcEZzw91bZfIhUf8VFYclhD8d4dBboDWT8dzIy8HEVEKPmLf0Meym+qb24t6wH+C2xtIBA1jOungVNZtwgpAf3FqkpYUiOnUM637J8lSdRHSbQuyx3Ki6aiOBv2gBtrqkXN7BDA7z0L52nuKIIvT+UNORMRBboDWT8dzIy8HEVEKPmLf0Meym+qb24vmZPaHPZVRNyAvZetnnrzMUzMxN3ZVssAr5MLZhS3k9gZNgkwu7nTyvxFUNS/UPOT4zpNPO5YgWbio0GtoX/Btzc2icvd1bNG+XEJO7hU6yxxHLifkb0sGhVUg9RSnF7QJvTdg2CjOa8dyoumojgb9/W4v/XdWrrFf7zJnV0piQDlmsLGCk0KdWIIAIds2MSryTKIkUcCMHe7RX6e0WZRBf/j/uyHCLVWb+orvOP9ecF7SWiKSZw/o1ZmiKIU3ioevUCBeDMp+9ViCACHbNjEq8kyiJFHAjB3u0V+ntFmUQdJNkmtHVLFwxHh3M/7l8Fmvh48WgeAe+K0edPGUxp3REpgAIGjw+8XhwyaAxLfQPQoNPNjpfmM0WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNw301UyWjFl91ZbuY+n6jy10mll5AvlasuR0cZVb9tSLCgt/GByzsKOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHKZVhEt1a4dxGkmZKZxGELEhDLwVhRFmb3R8WdJFTO+nSY2/TYeUf1yaSZkpnEYQsRiHW7aO5vxU6/78KYYJzZNaDHA85r5sJlgPHSgvyImSlqk89/pi6AIv9281ooBjDYfILcYi00x4h991K5Rjd5QAgRr7UzjYUyoNfGWRcbK3xxd+IAGZeat6QoGFUtdHnuoNfGWRcbK3/RcTsJJ8QYw5o94szA1qLuzxO7EBtu+KPzk0seZwX46GUMQ26CV9ZyoNfGWRcbK39zHLiU0HIspy041qprKfGy/3bzWigGMNsT2P1AbHH2oU8ChHu9j2s8i+PxZxyAsv2Y8kpni2j7KnUyy6YcmI8RLTpAqdXgC+VTszs8iePtfihqTq5TohFfIgh23HomE7LUffbA2vmQPM1z5OLuut1z307+4oPX6k0IjtZoAq7t0lKbPj9+iHGkIQxJWNPcBHe6gnuh/ZnB50ESaE7bHR/HrLdk6xCRreJ7JkW377qQR1Kqe/h8ErS/Qx7Kb6pvbi+Zk9oc9lVE34QIrqGEqX6zVmaIohTeKh5un7lHWnxT4TeY85nAP6AivvrsKqjSAqiBlpncqvXb2wnTnW/vJGXE+MMucS0eT2JvG0WizjqoT4jey/TkwTw2xQlg3pveBewRxMkPH3rMdoqDp5/6OfnmepmnNDYHvQh3MlbIhFGnUEjboyxTc6gvsmSO3WiJ9KGDUy0bAGUzIHcyVsiEUadQ3iGnW7Zak29+R+U+mkAaqjXKO4yh+XN+L0+ewznAFam0teJyG8k3w2ui9m17lwjeoNfGWRcbK33XgyCw2rXpGx3Ki6aiOBv3noVSnIQatPa36XsVf8dJBDJRo7zJdbmg94PgCmNLgmckQpThCFeIsg1YFRsRCSxYU+ZOe7mk+Se2Nhkx7Il6t4UhL0KhpJ38bcNzpKwLX1AyUaO8yXW5oPeD4ApjS4JmkH9NYKFxnQag18ZZFxsrfdeDILDatekbHcqLpqI4G/akIn4nmGBpITiBBA/fC90J14MgsNq16Rsdyoumojgb9HS2X739wjpEULPS1lugrtqg18ZZFxsrfdeDILDatekbHcqLpqI4G/akIn4nmGBpICR3Kc/rCFUB14MgsNq16Rsdyoumojgb9HS2X739wjpHFEm8S+fTTaKg18ZZFxsrfdeDILDatekbHcqLpqI4G/fxoyKKxJMhHiVblzfGmBcJ14MgsNq16Rsdyoumojgb9HS2X739wjpGGtqRii5E3AKg18ZZFxsrfdeDILDatekbHcqLpqI4G/fxoyKKxJMhHcHvbVgXuI+F14MgsNq16Rsdyoumojgb9HS2X739wjpGb6I8P/0Lpa6g18ZZFxsrfdeDILDatekbHcqLpqI4G/aAG2uqRc3sEm74Izq1+Jp2qU3zeZD4TfeD3oLb/XEQKaAbKeHAIb90GPUiUezMBVAyUaO8yXW5oPeD4ApjS4JlOfHBU1oPAvhMj/SBH0KPLTeY85nAP6AivvrsKqjSAqjcgfXEg9tLEXBfVVxFmFh+qU3zeZD4TfeD3oLb/XEQKQUzIUYkn2ybztvsrnUGVHL8RVDUv1Dzk+M6TTzuWIFlQiFKdx+yNPWDUy0bAGUzIHcyVsiEUadSE1w9p75u9Z0v7BcKJm44OEyP9IEfQo8uE1w9p75u9ZwwIOVo+saRwZjySmeLaPsovBxFRCj5i3ypCuc76fiTIx+eOQ8PDT3hnAwBH26HYtMbNprK4LYgbrh9/sx4J4Zfy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOFJZfy2x9508vnttGAcEzMvxFUNS/UPORkDlE+6f2frvyClNc+FMtjMVC7VNuCUoUU+ZOe7mk+Se2Nhkx7Il6tLvf5l/HvL+PszYnLau54RmKP/piE4gm2b7TfrcgcZ7UMCSj+ZiZ5RS8HEVEKPmLf0Meym+qb24slw0GaAd5zqnJ3oG7RzGOQf/j/uyHCLVWb+orvOP9ecLednca2bpdJ+hVxEg4lpoYF0JbbjIhF9lfBhX9gmnyQWpoJfdxr4eYvBxFRCj5i3ypCuc76fiTIEr+2qBBPvXMxULtU24JShYvT57DOcAVqk2kPZutRC5sbodo5ViUGwpdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmP58q1NiVv8c4vgTtOK5VSRleRIfiaIYRsOQP0eQmhULV/ZDDSjCStsmeCRzsMz1a8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTIGEjBijipE0SUcRnmdZ5Sr8lnN6ToyxXE1GyEI8J76Ug8QQ46zmxgkWGz5Pqa8LcGnkhHOWLndfkJGrPv+AUqh9TFW4JdLljfY+SK17iu0YpD1cpko4vTY1VxarjbYSyYVxXqkpAiBi/EVQ1L9Q85PjOk087liBZWxF3Y/ii2q5AhoDL61JMcTfs2T3tv7quaLqzJmflsPSXt14nAyWWX0NaRZr5dtq7lcwbKRQEQlmWnABkhfYwG9iuoTHUj00c9RtFt/kJVCzmJ3jtfpYQHM6pQZIsT/k4vCDbezovTlKzxO7EBtu+KHzCuCEWjwuex3Ki6aiOBv3noVSnIQatPSZnEJezfXs9y5PpLEgYovQYa77f8vmAHaEdVcCihkLlPeD4ApjS4JlHLZ/lRM5hy7twcZyZxxott1OLXHeZwhiQ0Q8ygJvXejYkeoCQpLdmFPmTnu5pPkntjYZMeyJerY0fJhxugN4fkV9gUsiqwrNxCvea/bRFrP9VOEEPlSHPvxFUNS/UPOT4zpNPO5YgWaCeQxK1Q7FeVMz8s7lE/N0vBxFRCj5i39DHspvqm9uL5mT2hz2VUTezpuBjY2VybfcaLydpsQM0LwcRUQo+Yt/Qx7Kb6pvbixMP5hb5t5DaETuc2nyyzNzmIqollrQmagWTiPQ0N7bd7Y2GTHsiXq1YicvCQgrerJ7Rh4kaLURo7Y2GTHsiXq1YicvCQgrerGV42WujtM9gvasFSgZCszDjdhVjvvgpIWFmjN23bm9wM1ILnQKCFfPmjKghd4lsW+un3f3QvH4/K6EhIz/oZ7nhT/oGmF1lXzokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyA2f5OWNrScEU+ZOe7mk+Se2Nhkx7Il6tWInLwkIK3qye0YeJGi1EaO2Nhkx7Il6tpBpOzomdoGcMihLJdAxE+aIc/j4NtRsPsNMwfWlh5XJmqNNMdXpyChSVTkv8zn4wH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3LQVlKofHHLJtrrWYvsHNnIzsey4CsrGdYqBAckRbuav5vX7RwU2rinlHrBC07kStu9J5gHlaVqiqr4MCPcf7rXUMUP9aNywiw3SPTlUXbzjkGwgGfgT6nEqWiSDJVsh3Z4d3j5Em1GJijk6f10lHPQFYYhl+XAKgJ1Kc+iCax6YZnynTrgorqLBsEY5rCh9x+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCxOkt2vc9ZNFnlFEOez9nWfw9MlWEq9WakLp/n2nSKsklM7FV/qoydlVr5987fmvr+erqih1M4/juhK1yHWe8Eecluno/rLjFjJakekrNK1qUt/ZazNBY4eCeBlNilgh9jJakekrNK1qAzhYZ40TFYEjbPf3JibGSxuqimyh3chz3jKlVr5PnBkjA4Ul7SfdWts7gbstDN5adU4OTYdMe3ABLmdLVRh/xFvVIAgx1sm4aDcb8kPEFtZTA+jtY2bE9m3gjXOEok0Sqf+pnFXZBCQJuaglfeAYmwicGGCIg0gkNrBKvbSWGzgfkn6GBxXQ4ClT50JpQ6IZBmmNrOWyAJ0xPrlasMDNvCvIow6cmO01ngV18WB6UPvJN5N3UJEcrdvOOWEzN8OBB+IQ17Q66D0NlONtS4gi6SMDhSXtJ91aaN+L75UVHu+CibNiHARz8SvkwtmFLeT2KWRseQJNfzi8C1sSUY9bywIOwtTcXwUBBHEyQ8fesx17MgNFn1iXUJxqJIHSnBRTtZs5Ri1VsAoxPrlasMDNvNLDI3FnuJoScsFvPBiMwXstMZHWzYyLJ6n/qZxV2QQkCbmoJX3gGJsInBhgiINIJEa3zjj0aHVEb7CKGgQd+Im7n0AJwgNkC3P5I5WTGaea99GvZaLhYDteGO/gp+2qSfWG/YX5hDGIEjboyxTc6gsy57o8DQoM2Fo+25FgObr5FIjp1DOt+ycaNFlXzF9E/5tm8h3jKpl6RRkTm9rFTNL8BVvBnRzJscLg4TLFSlMP50r/6zZg8QngL06kmsumvzWDp3sTkzViaZ+cHv+AQvXm1fRD6ARM9ysE6EgXdjLiFIjp1DOt+ydqv4JmAN7Yo8cNdJjNmzYFr2nM1TdOPxp4YUNMIn4SDFiCACHbNjEq8kyiJFHAjB1ciKBtGkJ7V3bH5RAW+rQ4APUSqEkqfEA6rVgu/t5LXjjgq5bS0R06bUXfYiX6zhRvsIoaBB34iYXBd8WHtillCONgulB3uAY6rVgu/t5LXjjgq5bS0R06bUXfYiX6zhRvsIoaBB34iYXBd8WHtillPUK39uQ74XY6rVgu/t5LXjjgq5bS0R06bUXfYiX6zhRvsIoaBB34icMfw/ustf9RW2mt/IUi6tMFwgdNOoiIzRxHLifkb0sGhVUg9RSnF7QhQsoGMdsL1sZMuMqSUt+2r2nM1TdOPxp4YUNMIn4SDFiCACHbNjEqQLw4iiueoOJvsIoaBB34iekQ1oe8LDK56Jzm+JTZIoGmYftLJ89blfwFW8GdHMmxwuDhMsVKUw/nSv/rNmDxCZ8tDrlph67IhyJu09TkcB9iYAEqiFN1Aj+H1ckGx1PGa9CKQlY8TsIr5MLZhS3k9iwjF6cd+1c7Q2+wrYI7E/NdOYpq2r5bZQAB4LgJfBif5tX0Q+gETPdUVhyWEPx3h0FugNZPx3Mjwq/E6KuC5WH3TjxpmeIoIXn6nZOGYC936ja7qAz/lfFYggAh2zYxKvJMoiRRwIwdXIigbRpCe1fwncYjNsqPX8bXe09SFZZkYmABKohTdQI/h9XJBsdTxmvQikJWPE7CK+TC2YUt5PYQ0i/VF+eUlLP96qOblb2/e3yG802Gi7sabNF7pGEbiM5tsGZyE+TH4cMmgMS30D0UiOnUM637JywkOTnN3PTBKgYxFtDBT6Bbaa38hSLq0+o2u6gM/5XxWIIAIds2MSryTKIkUcCMHVyIoG0aQntX8I1EQsuDpQbqyGODYemtaQAB4LgJfBif5tX0Q+gETPcrBOhIF3Yy4orz7xR5vZrL0KyVEYCjTvuE5B2e4Roiw4bWnDTum0T3DsMHTjZeXWOD+dw5rplWpXWS5ang/xfHuc+DrplHeHXmbDxANfJCsR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC8O+zhfXeKzlr5fZTZKviHa1+k9DaRcW1iHPN0Q9IlPlr7uCvDZS6KHnQ2vP0U0BAQ+vYtuw8VBz/zmFdEeLXeq9+phO5VgpWXS7gBu3zNPtNZRaCcRjFL55tWE/gsBuNbW7uczLhdNjrTExBvUE7t6Ux6WCFBtxH3PQhLPU/v3pnBZlDDWPRc0fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv19JhV0Bg8FAX8cYC1vw6ZInrSOdnQKWp0tGcGsxfg0omtQ797AIb1pn5zUaoL+FImERhWsm5kQkFnNNo97vtpDsuOAuWahUAp+b8/epKVm2q5gyM5K/Ntm+rPKsEBPe9BDw5nl0nob9ZJwV5YQzzoI2z39yYmxkvSgIrk3Duj8dZJwV5YQzzonSggCnu4qDywUBTkL2d8olY1tXzOO1m7Jjb9Nh5R/XIAupHEAvr/j8oAxG2oU6OZtfJjinfBJCHC/Akftdwe1zE+uVqwwM2893jaDoJOdejtG1k0bLNkma5YLeqOZKQRUxKtFKe1H5zD6ZycAbPtkYsr+xQjjpXxh2NLxFc1XinkOwfUh5x028BYLB37rmkwYbo5NtfjTJPWmH0QnDKBipTvgT5Y3Pp5449n2RHU5anAuGDhsFoG18N+zASgf4D+YOXiu5r1A9YP2rrHdb1eRrR3f3Mf0P/X7Y2GTHsiXq3Nxe0HbovEqGHW9k/xEsA/PBo4bk72mikh/wM+xCDWlH1oCKIur7f0WsAEiNoPPIvb2/T/MLAx8PszoAcSSMB5nwOmAujGGLoiTYgnaEY9ipwtqEPKcLSowR+mm+pxTPoBq8OYNNE4kdKDEt0ZXQvCabaYySE8y06sPWg6FSenyE7slFv/HsQ4SLLlIdizBEylVI5U9r6HGrT//Islk0UTlXeHI7I2QVs1epxaUq4HuDbwCp+NvTJ+AWDQJ3KBpIOfoAOLnMoIH5oOnpptJ7Ig8bsTdDFOIKDsLS6NijTT1RxHLifkb0sGc8rFJQKPIgNIsuUh2LMETELb3Tom5psazUXhaLMpmYRhfQeIFI3IYtSMm8EQGs7zQhQaHWyXaE+qkA96vqRo0RxHLifkb0sGc8rFJQKPIgON+6jE6JHeCzHcDu8XMKjbH0km0H4E0GIpim5dgZrhdGvQikJWPE7CNuF9Szb8bc9geRD7LDFinycNF6Xh9oRrcICN93vFAvaNs9a1jKePK8TZrR9MdAnrsraGiqK4eHXBH6ab6nFM+q0edPGUxp3R1D8XUnf5aNBN5jzmcA/oCNdY61XS4HJTWIIAIds2MSqzpuBjY2VybWSR3DO4+l0JvikGWcuEr9RRVIBa+SRHIclQhwwd/5HsD7DkI+4jM/Jr0IpCVjxOwh2DWy5n0Tr/HnR5XoeMh83g96C2/1xECkVOThjF2eJ8UzZu75YUdPVDgkyyDP8+zMLg4TLFSlMPKqLBu3yOMdqEqM2ibohLc25XSi3zeRFCMCAsaLkc9sMCLmfIM/UTQAfRz+w3XbY+7GNtU97kTE2foAOLnMoIH9t0NliArEXrPeD4ApjS4Jkpa8rPfcFPWKw9aDoVJ6fITuyUW/8exDjZsyA953UF6u2Nhkx7Il6tWInLwkIK3qzxuxN0MU4goDlmsLGCk0KdWIIAIds2MSoRuLG4+wILq/BwnZcmTAaA0Meym+qb24vWcrLWwUl/M+SOCFwaOINhKN+o8Y3BzwtwVH0b77Yhk2+0363IHGe1PWu08ROnR1SWBYt/A1hOvyCKiooIc76tm6HrtbffkzZiSiR2u+FIv/zmMgugc2g+kfvD/Qfi4tJTtWTJEG5oqA7wnkJqcvIWb7TfrcgcZ7XCWmZ9OnA28BxHLifkb0sGhVUg9RSnF7RdR+uEUgMpq4huYtKdSZDtTHfyjKY6dJ6cOmNUNiQp+dDHspvqm9uLnDyTxmdIM4rhwyaAxLfQPRSI6dQzrfsncmugrqLgp8ykcbJHbQgsfb2ZfnkyPxNaniv+1iNSrX9N5jzmcA/oCKEgdOTgzP7Ca9CKQlY8TsIr5MLZhS3k9gFo363P2P865tde/T0vyyBl63Nwo349CjxYyQKcLncOt/XtuqXLQQxvtN+tyBxntdTSRCRalyta4cMmgMS30D0UiOnUM637J+N+Fun2/LF8ceKYvi5QGz3Ku3bBzjLZXi13IUxTLzX+nDpjVDYkKfnQx7Kb6pvbi63pTOsxQmwu7GNtU97kTE0pwUOeZhNxAcwywBB2p8jzb7TfrcgcZ7WJMjrMeW1IpUoNKiewNIBWAa+cch8jSnhYggAh2zYxKvJMoiRRwIwdSXFnkheyCSU94PgCmNLgmSAvZetnnrzMUzMxN3ZVssAr5MLZhS3k9pDBcKEp/OLdI/M13JkvEV3gq05SGeU6HZTOxVf6qMnZI4vTKyHBGc88/86HSkKUDe2Nhkx7Il6t/CSiwSGFTOTC4OEyxUpTD+dK/+s2YPEJUxKtFKe1H5zjz21g8nqpA0PqPg72vnt7zc2icvd1bNFrNMEJkNLPxeC7noJyhgLObUXfYiX6zhSnJ6defzt03f5OdJ2k4EJN+M6TTzuWIFluVZtPPGIBbjaxjIxorNUKHEcuJ+RvSwaFVSD1FKcXtF1H64RSAymr5mT2hz2VUTeMUfrFsQAMFtI1uCBKva8tvZ0cin6BSwJ+VawGUS6tvOxjbVPe5ExNnGokgdKcFFP4MMNVGwB+imx8P04A0x4ZlM7FV/qoydkji9MrIcEZzzz/zodKQpQN7Y2GTHsiXq38JKLBIYVM5MLg4TLFSlMP50r/6zZg8QlTEq0Up7UfnK++uwqqNICqCXFf19TCX2Lbrw8/02YrL2YWUEPoesfEI/tL8RalmbxYggAh2zYxKkC8OIornqDiC8g1E4M0/TYD5eTr4S7FDvSjPdZPbMmLnDpjVDYkKfnQx7Kb6pvbi63pTOsxQmwu7GNtU97kTE2caiSB0pwUU3RQ37ViZzvFKX54BpvuYKnvfieJNHKPypi1H3hoELT1PeD4ApjS4JlB42W2Gx38R8Lg4TLFSlMP50r/6zZg8QllHo16KJwxA+TE2EslXO6M0jW4IEq9ry29nRyKfoFLAiuhk12RnH0iHEcuJ+RvSwaFVSD1FKcXtOjTGBzE51pHVhWiDUWOHsxkqNYjBwGHKTz/zodKQpQN7Y2GTHsiXq1SXuzV2VDDRmvQikJWPE7CK+TC2YUt5PYQsUqzOpOPbSoJ9VoTsZR9+SYm1G2g6p6YtR94aBC09T3g+AKY0uCZQeNlthsd/EfC4OEyxUpTD+dK/+s2YPEJpFRrV+tIZZS34X8xDSDsR9uvDz/TZisvZhZQQ+h6x8SlpzJ7lSVPqzjgq5bS0R06bUXfYiX6zhTAk8yfFtp1ednmw0WWmZaZzDIG2wgILyWcOmNUNiQp+dDHspvqm9uLrelM6zFCbC7sY21T3uRMTZxqJIHSnBRTgL5c+0ismyEpfngGm+5gqYTu0N2252e/mLUfeGgQtPU94PgCmNLgmUHjZbYbHfxHwuDhMsVKUw/nSv/rNmDxCZuyMtQ4si3HUiOA+a1tHuUYiMpUi4oPIbf17bqly0EMb7TfrcgcZ7XU0kQkWpcrWuHDJoDEt9A9FIjp1DOt+yc85qYyNC6bUm11Qv3exBQ49jJ9UGXP55c8/86HSkKUDe2Nhkx7Il6tUl7s1dlQw0Zr0IpCVjxOwivkwtmFLeT2f5PoyaZ2lL2U7j1xL+CkiWfBQ6EYMMsEPP/Oh0pClA3tjYZMeyJerVJe7NXZUMNGa9CKQlY8TsIr5MLZhS3k9n+T6MmmdpS9GXtRpcLGKjJnwUOhGDDLBDz/zodKQpQN7Y2GTHsiXq1SXuzV2VDDRmvQikJWPE7CK+TC2YUt5PbSBHSPBzUZsdV72z6hEmMOD0d6pSj9f/6eK/7WI1Ktf03mPOZwD+gI11jrVdLgclNYggAh2zYxKvJMoiRRwIwdTUPDHmnSGO8XLShb4QznFkx+kvJC4kT0268PP9NmKy9mFlBD6HrHxKWnMnuVJU+rOOCrltLRHTptRd9iJfrOFAvINRODNP02xfxF2xPWDu/ExTNIirtarpw6Y1Q2JCn50Meym+qb24ut6UzrMUJsLuxjbVPe5ExNnGokgdKcFFOUY1JmcmIsPCl+eAab7mCp7zex2TjmveyYtR94aBC09T3g+AKY0uCZQeNlthsd/EfC4OEyxUpTD+dK/+s2YPEJ9vZi+XBIz7jRDKF8K3NC1sIKQH9xapKW+ZiKT0jJRQvWU/GeOAeHmjiAxNBKTmIgSg0qJ7A0gFb8KXwtoYo3y/GoM0GWbfn9ln9JahpkI1kw0mP3skyStFRWHJYQ/HeHQW6A1k/HcyN79feNevrNapFwwOV6kcYWUuvyRTQzJ42eK/7WI1Ktf03mPOZwD+gII/p+o9rck6E44KuW0tEdOtGKG/xtD4e950r/6zZg8QlnAj4FcqgLAJ0iIW2HJOoVuFpuOk8Ny/lZvmYggtqVAuHDJoDEt9A9FIjp1DOt+ycoVD2Qz0+RwLhCSwkCGnKYrWVFDcYY55LrQSE+TTIjoWvQikJWPE7CK+TC2YUt5PZ1aQcrSvsbNGLFBj9Q1z1b7E7iAOxKA56DRwMyBDAMnexjbVPe5ExNnGokgdKcFFOvp5lIcrY8qlPChwfC3RnRhAn75rgJ22hV9lIU4e11XViCACHbNjEq8kyiJFHAjB3mzJGdnxFZA+DH+WIo91q8koejOOHQ5KOm0AkieOvdaOHDJoDEt9A9FIjp1DOt+ycoVD2Qz0+RwIJkbFKREvOui0kWLnusckLgu56CcoYCztGKG/xtD4e90kfhGIVJ+sqXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZt6/+445Yo4pKLRL53Na22LML8H3LkfDQVkHA9osP92YLPXto4VbtxOfZE9UU/BHjKaqUsONv48Y1vFPMEedBPgy4dleL5gYQgkqynyK4dCEN4Ppi1Sx9wpWnP++ZTqHJp9kT1RT8EeMzasixnaPUTI0VldX/5MjiwzdVkA/y8eO0rc6Oul9+DKkzOcC9/gJnpdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmDX/aUb2X9hZ2woXz0TKgOyZeaT/v8OS1YPDP1zxxfajkJGrPv+AUqh9TFW4JdLljl7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHNaowTzld5YjOIDE0EpOYiDvhiQO1qY9SMcNdJjNmzYFiJZ8gG/bdpTHDXSYzZs2BRa7zoMzwU8uQYrSQJBv7P7tyEloUAZhvmxHoMmoJRXKaPJhJU/mJxFxwf0uM9v696g18ZZFxsrfvtk5SKcFdH8aGmou/8QwOhOi5IghwOCq/z7svFHqk+Ujpg4yMtebifGP8129pjHbQPVHMmkNW9PsY21T3uRMTdVqmPXCNsfaPfrjP69VQDQ2FMDmFkneugRM5a3QoG6cNv1C5IcM1159+qWmlydBZquwSwszM3a5YSBlwfxDgEHDPI4Y22ZnyfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln5Ojh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2WpiLgVtcz+6yMokQ8Xzmo9ObcPamcengk16VxjrDT0MK8tz1QEMzvvrYQn+0aiyBMMRv5acdDkl6N0UV6eTY8RUjdBXjqPjgJf5A2djcky68QCYtECgVBPg7Kdb0s9rI4aphD75swo+qYtuHA1qT4jSThHACCR/41nKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTjJ/OxMxCwDDlUUIrHUaZqVCu+mR2vgpwqjmrgqPScEShYWAR161KjWdq6q+4iv7MalCoso7qGU4npv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWslfZCyA0NLGA94PgCmNLgmTXoi8p+1sklLwdkQahPEIPBPkYA06LX7SPzNdyZLxFdGkiNv4oOALK7cHGcmccaLbdTi1x3mcIYkNEPMoCb13pTEq0Up7UfnOPPbWDyeqkDMJducXsWsZZAhoDL61JMcTfs2T3tv7quVVtw4ikZM8L+TnSdpOBCTfjOk087liBZWxF3Y/ii2q5AhoDL61JMcTfs2T3tv7quG3ynRfQJ0PbtjYZMeyJerQiVEkxlqWvzldmD65voKkpAhoDL61JMceRAr9Y3JhT7GmM340wuvpHo0u8+V8CORvGED6cYfjdoNrlzvRZ41imTysGfIDZrZ5jY2T67Es+9y5PpLEgYovQbfKdF9AnQ9u2Nhkx7Il6t6TJZvc0qKnbZsyA953UF6u2Nhkx7Il6tX9/RxVkxG7TJZIJ3xSMlN2+0363IHGe12m1vAK0Tcmn2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTJXlwbgmXVaZeD3oLb/XEQKbYTaQi9UxxTL8ElX1S2Iid9yIvxc5OLJ0Meym+qb24ucv8T+ZT1F8N/EzAsb4Xos/k50naTgQk0SUcRnmdZ5Si57sf1umrHmzGRGnucXhCmgBtrqkXN7BLB5JIIdSKgV1S3+/aM4X15vtN+tyBxntVEAxF+JRliszGRGnucXhCnnoVSnIQatPTjax/h7OrMLMuayWMqNqvHnoVSnIQatPSMBSHeyBizv7Y2GTHsiXq0IlRJMZalr80NS5kH2JRrhMNJj97JMkrTKPwX8ZGi/bdt0NliArEXrPeD4ApjS4JlFmo0KuYTpQhJao7CnWxLZTeY85nAP6AivvrsKqjSAqpYAC4pvx9kr/k50naTgQk34zpNPO5YgWSl9m5P6d5QoajkcM0HTJMWiAiNHs4agN4V/WU3qpupr9c0Et+l9X/8Nxe2QllSjW9/0R5oi6Y2ycCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHoSIsomI/+g6gkLJdr3Dz9+HR6wgyZ2KDzmt2ko6MMbby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8VUplQXIBHQn8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOUuVvumBoEQRlt/8KBI/GYtAjus0rNARigkLJdr3Dz96+kdq4nChGnY6C1JXq5n6GmBGCwtpd4/hypOO84iHzgwLUWde3Bh2oQtkFbC4U27AnfutdISm/jq3yd/PALGm+gomfx5cpBl/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk9kQUBDhdQ0ETtJE+F0feJkXW78NTiYfDcBYLB37rmkwwFgsHfuuaTDAWCwd+65pMDoFVVo/YPIZlL03ZswhwxggrLEnFT8WA5ODjhOcs98irYBq+ZVKcB6hAb5FCZiaMtwJyRAwlWAnauzov06c+m0YUFZlBvjdrmk81lE3TidBfs68pZAp+Q7tGKadmRcej036/d9UylwapEHU72SpwbvT9MgH/iBDX7kKqsiGMrkXmc8UN3rYjOR5KAjcU3G/A9d5k03BA28ydjlhQ6Tow9n0g2shWVfD2HBk246PxgOcIX0fiB5F/kSUuVvumBoEQZ9SjlWG/itCLofZLPmqhrCNSkndxJgh/EU+JUjU1wy2I8qlv/sDuZ9d+faJVVJpq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTj3xHKw7Y5etwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk5Amhzf3ng0L5mT2hz2VUTdvoEC7z1edMBnWng+1mx0boWFgEdetSo1nauqvuIr+zGpQqLKO6hlOJ6b+11OiNzEAGkuTHgN5IB8gtxiLTTHixi1yExziaZRxCvea/bRFrGNQnSbq+UXfWInLwkIK3qw0nN0fx0OZ3Tkh1dWah2CZUQlm3kjqGg20C28BNr6eaRBDmFrgBPP4rwzQccgjIuj2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTL3Gi8nabEDNEu+dfYO6F+PdRYolDpH0bOmt+QzqmdAq78RQpZeJabnqDXxlkXGyt/noVSnIQatPWxnHwi4UUX4bPz/c6/JJ/2iPRAJAhOGHuuwrupyCFw2Q/i9SenvYJ+4QHkjGNhy5k3mPOZwD+gIdao27wru/NVdkINk58cbdxYIrgHFJbfVnwPfoCo/23wlAjXh6w8auSzYBVHs218nBPsvgTeYHoHtjYZMeyJerX+2TT/d4e3JD+wStopmLoLmd92JXPyKJ5x+AS9XSZa9Aali67BC4/6wFdAbRARLaBhrvt/y+YAdO9HxPyntJRzsSITjDzblWL2dHIp+gUsCo1yHmga2QjHqLEJknZBvSXMai7FEdqtBv9XuzqdyIujQx7Kb6pvbi7CtinIM1HSjqDXxlkXGyt8oD5Ox2vaw2UCTFANmNP+SarJHaLTH5gRN5jzmcA/oCFZBW481cEtUuWDl+4FOsmjMQT5ndyMiZ9mzID3ndQXq7Y2GTHsiXq0mwYphmOBmEuNTtdERx66+GGu+3/L5gB1jUJ0m6vlF38mAFdJz89hnLhg6QtYxBZVnRXa9faaECMbByddibIgds6bgY2Nlcm0WnOIbR1Um54MoNZA6HRxHwFgsHfuuaTD9bi/9d1ausXyjZbp9CZN57J9nPDNHgoo/SvJtuzsGM8pi11qMuj9p7Gfhw9lEZps2/ULkhwzXXsBYLB37rmkwrTIP0x/AMDAYa77f8vmAHW1zIw3oNll+iYsXHI05xDydBJEKRY6cDa0tOBEbY0UMyQKM93pQCgn95JsW2KW5gY9La0Y4HBprglqz+vy98s/AWCwd+65pME2WeN266KtHTeY85nAP6AivDNBxyCMi6L+5us15GAOW5iKqJZa0JmpjUJ0m6vlF3wRbnhTMYuZiDj/oLYYe9+mQ0Q8ygJvXehD0ExRs9ghbdwwqZv6zyy7HVbaI9yUfqqiElkWPOTuYYWaM3bdub3AzUgudAoIV8+aMqCF3iWxb66fd/dC8fj9HuOphjrTHNEb+jsZ+iiMUcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxH2WGmXFrr17cIJD/3/E3KGS3Ua1MeI8lgFO4KCBYYOICWy5HHtjmD+m4go2IHP5VmS1Qf3OouMY/y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8drnMYhhGMP6hnI7LwFZoySFf1lN6qbqazCBT/1Aeq2TUQckFapdvvdN5jzmcA/oCK++uwqqNICqusdtqK88M9RpTNEAUiIqBy8V8b58GG7aG1QhNxWUqndD+L1J6e9gn7hAeSMY2HLmTeY85nAP6Ah1qjbvCu781V2Qg2Tnxxt3/+DXU56Az20EW54UzGLmYu871r0UQiAQ4SSlnUTC2QjJZIJ3xSMlN2+0363IHGe12jv5Er6c5R9fWADTFbkpBE3mPOZwD+gIr767Cqo0gKoue7H9bpqx5tYubd4q3g5PwFgsHfuuaTDQx7Kb6pvbi+Zk9oc9lVE3eMMHzF9kVHuvvrsKqjSAqqyd79yEa96/AEpUG6CU5b5rHszq1lh4rsdVtoj3JR+qw1CJGvLT0E5iCjv/vpJYcEb5NXIrNUWEkhCnosRnLI5LuRgyX6MnyvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk2wB+7h+Ops6cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJP0e81vVW9ueHBGIYlBna68rTExBvUE7t6Ux6WCFBtxH/UU7oZD+AIKl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGYkjxSbwT8TYW+0363IHGe1SWkWqmH1kvcETGOhmusAcThRF75Ga1Np0Meym+qb24sFLpGvYNhwGBq0oC5+4w/QPeY46do02cY94PgCmNLgmTaMWyOJnvaYpmRSLqrDyOGC1TjSiQZSENJH4RiFSfrKQvZOoeWO9V9SZHPQQDrFWqfEb3WHMzLgUWPn5y6uxfwczSDxcOSOcrlg5fuBTrJojATQ++vsEuvQx7Kb6pvbiw3SpwqG3ZfcElvsOF4XWHDGDh/j4G18UOYiqiWWtCZqY1CdJur5Rd9Qo44irhrrWFJTuU3JkJFITOo8YE9G74yvvrsKqjSAqozzeEpU+0a6MuayWMqNqvGgBtrqkXN7BNWxV+32rY/V7Gfhw9lEZps2/ULkhwzXXsBYLB37rmkw2XXEtJhIU/GHHaJFRC7K1WfqQhGqky6vSHiRAVn+cSQbnFxjjXEudT3g+AKY0uCZKLZmRhS+HlPo0u8+V8CORhD0ExRs9ghbdwwqZv6zyy72iuplgCAem2un0oXkzpyqb7TfrcgcZ7V0HvmOxjI4bzXR6dfO/9nfk5vDWDoY7XDtjYZMeyJerT5c5iaKWu3+8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWX8BneAa15M97nZwbX/dmE3b+WL68jVja06pKGjH5A/8kmLf5cqSfGpOUrjzKLCkW+QtAfnChtyP6S/LYWaM6lQ9LT2agh0TWajyrgAj6DfckZXoljzqrYCKSf92MKceG8cDzAedhnDN8rixIvI3Gh9XAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTm4ZZr1nx3iny/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUck7SRPhdH3iZeRB+SSl6egy0CO6zSs0BGF60a68EpnDBfad1uKmdKYFO0kT4XR94meHWMJbeo2PDrPJ4C/6Rq19+zrylkCn5DuBsjv3AGrSPCsT530b4fzby/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPZEFAQ4XUNBE7SRPhdH3iZF1u/DU4mHw3AWCwd+65pMMBYLB37rmkwfad1uKmdKYFO0kT4XR94mcA8FaiksCn/pof1ZPst0KrAgRpueqiAtMUrCUjw/yUuTtJE+F0feJm70LjCSmzaNKaH9WT7LdCqwIEabnqogLTFKwlI8P8lLk7SRPhdH3iZyhUnCGw0tmus8ngL/pGrX8CBGm56qIC0xSsJSPD/JS5O0kT4XR94mR4URTY76PskrPJ4C/6Rq19+zrylkCn5DsUrCUjw/yUuTtJE+F0feJn1oQo2aNryRazyeAv+katffs68pZAp+Q7gbI79wBq0j7eGkY48Lf0+8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGYIflgfoI4z2Oun3f3QvH4/H77FF1YKRnPW4VbMTLTe84V/WU3qpupr7Z36IFzy/QUfILcYi00x4udtI/0UeRgdZFdkSnhQ3bdyErauFowuZk/kMqEp6+Cp4YUHeRv16uTmIqollrQmajdUEiFAlz/sl4BuHx+ia1c0nN0fx0OZ3Tkh1dWah2CZUQlm3kjqGg20C28BNr6eaVVbcOIpGTPCEGrPghc2Psda7FjBiYUt7faqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+gGwFmQkytbgP1ziX8hdVw2N7AhKNvBXLfCf1a1PYXmtrLsSh2Hw2xeEkpZ1EwtkInt7wAqyJilkETGOhmusAcThRF75Ga1Np0Meym+qb24sWWnhoar7wZpROKHG0m4e4QvZOoeWO9V/Qx7Kb6pvbi3rAf4LbG0gECydMKLoRPvF6n9iIdRbgqKg18ZZFxsrfcbwwikB6wzHZdcS0mEhT8YcdokVELsrVshKv3NWfVZ4NUYmPjK7iaxhrvt/y+YAdvbd/0eK55LLAWCwd+65pMDdUEiFAlz/sbMetH+lXVyH4NuuE0jGdN1rsWMGJhS3tJIvRPwe8MVPAWCwd+65pMK0yD9MfwDAwl+VJtD/uv6CWIfqIs0eBJ6g18ZZFxsrfDEHKq52jrwnm1179PS/LIB7cwCB+W0ejceKYvi5QGz0CLCps9PQdpmo5HDNB0yTFogIjR7OGoDeFf1lN6qbqa/XNBLfpfV//C+XNPBlySxSmMqc2evm4FFnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTQxLD92or0ceXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZheq+uebihxHyAHdSTe0HeZW8lRgNdMUbTBQ5Ch+AcOcCSrKfIrh0IQ3g+mLVLH3Cn+JCU+ad8W92XwjiM/gVTTDufJVvaSyZ0TNOPLQbLu3dF2MLFXGMaBZspnCMagpFPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyBhIwYo4qRNDof5RJ6fzZAg8QQ46zmxgojojbGMMRDcLxXxvnwYbtrLApOQol6t30u+dfYO6F+PdRYolDpH0bOmt+QzqmdAq78RQpZeJabnqDXxlkXGyt+XEYhV5OZR+Ya31l+4dBcL8agzQZZt+f2Wf0lqGmQjWbhLmDiLqTUvGGu+3/L5gB3kd+NSJQdfWdl6MBcfTccuNp/C+/jHUhfcABiEC3Cb4LCCehpaHt7ETE5SsWIahHzeDL6dNoD/r76uAJDCpPpBBQLNz0lER0TEAdm/7hcVLA4np+Fuk9fRXrWEYoRRpjjWp/5pn5zLqkB8uoZqwNyn6NLvPlfAjkYrNkUdqsgVVphzLVkrcvDftNd3+Ny1F6x/VxQ2viUoEdl1xLSYSFPxwKrX53Q9TAaq/1Je712ZK5DRDzKAm9d6+D/oW6NM1wFEyxyfFy2sCTFQu1TbglKFEGrPghc2Psda7FjBiYUt7WNGRgWqGd3NnCQEQbCmj+umYURHNrLDk16KmzmB8rstNsserZTdptzkd+NSJQdfWYu0rJ5GizcCGMwJHpKxslioNfGWRcbK34x5jSsPHYitRMscnxctrAkK3tBvBB1c93DJ8ZXI557yStTdK/qWRYymYURHNrLDk16JN6CzdglfXriVNXski/jHDXSYzZs2BRjS5F2cgeLfZiohxoSGxljdKhmPOWS04UzBmFHAOwS0DcITCqE4bbFS5Fhn4vBKCWKi9NUPhDRQwFgsHfuuaTC4EQXmPpeno8wvwfcuR8NBRai/hw89L1cYa77f8vmAHbCkbeAj8ssBIgXZZSR0jLlshP7KPeFQFKITy/e2KwCk8cV8W39jWMBNOcPqVvJryiVFTR4bmwnQr5JQpIAdF8biRElPR3NRSud3wtZJUJN8lxV6QatEYR9Ct0yeerDdRjBImKUFCEXuYcBFZ42sF+lT4EQUuyU2Z6394hjSIavC37cEVTJFRrSC9TX5sAYwGuCOueztBkGp+bY1nBIQ1LI1LZdt0TTB8JDRDzKAm9d64MvUaj21Sl5XnNmeKozYWuuRDpYJOjph3thCIxGtwVmC9TX5sAYwGpIXu9Fr24Bvgp8yzhk87I6BxxdBe9PiXMpi11qMuj9pX4CHGxF1gxPJw4Nr43cAi9qnSd+PxqOn69X5XEwE68kCgedoCuA+3byJFBV/LwZjhRsBEP+9W/MCGEfdpdFYcTMh4mDQjfoC9QCLXoO8JB7gofqfTM1QiqhdqE7lTFOPNS2XbdE0wfAzmdlYvBT9lMBYLB37rmkwLkSjkYzaph9yWDO1b+iPhyJhx+c7I9vp/3lfsRDvNEXXMoHOiCAj/f9yMxJYmuerDfZ/L94i3SDXMoHOiCAj/ZDRDzKAm9d6WGtfBT+QcumhTlob0CDHW60yD9MfwDAwm7Cl/JGm4dRMzOo1oB5ATV/RxpMENFILl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkzn2Cf6wkDYmUcMsw4JWTAbElEauj3VXm9qNWZ+SFyc++HeaDf62ttVcoWr7neF1uvwynX2c8/G+2yHxffVSi5kfsNQFrMbl67wHpAnIjSLH3gKDWYvH7RgktnsSGOYYNATYtOoT7nIVR54boltAh86EJKXf3iCoXIM40BRQKurwBe+B5GNr6KkWoX6eEfn2Ug9Au7GZ1uJpOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHLMi/Z9y6rv88EINEXysZB6hX9ZTeqm6mvtnfogXPL9BR8gtxiLTTHi520j/RR5GB1kV2RKeFDdt3IStq4WjC5mT+QyoSnr4KnhhQd5G/Xq5OYiqiWWtCZqkngGnGfhgZo0nN0fx0OZ3Tkh1dWah2CZUQlm3kjqGg20C28BNr6eaZ7WNoaMRI3Ytp7kMdSI+R+7cHGcmccaLau89FjbHlF3E9c1gpRGLR+OL9z0IaBXzAwrjVQlO79KZcxmz9AAC0ynxG91hzMy4FFj5+cursX8ETuc2nyyzNzmIqollrQmaukkKpWfySGq8kVan6uHiAGYtR94aBC09T3g+AKY0uCZgAj7l/iVZXWoNfGWRcbK3y3c9dka9WadxNmtH0x0CevtoXtuk72geykJuMch/Os1uWDl+4FOsmi7DCpmgfhZV8GO7LwMPI7EHlbhmQhfdoMXEGMWfEHdKlA6mBBxzyj/FzIuTzuQM1bAWCwd+65pMAOiVc1Q0DVa2mDXuHxzGRU6VHcnaTQTmwOiVc1Q0DVaR6KnrgY/JqXAWCwd+65pMKl8+09yWfa4wFgsHfuuaTDalGjUNcuOE0Sn9vmOMxGYbPz/c6/JJ/2iPRAJAhOGHsBYLB37rmkw76mp6Ah4PjtfG33d7c5AOFEJZt5I6hoN5iRnMMMFpPvAWCwd+65pMK0yD9MfwDAwl+VJtD/uv6CWIfqIs0eBJx+pBQUd/IzhvoiGCRllu1SRftjjGWJHTTrwQPJBxam4FEiZ5C1cWVf/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk1vBvlGgaYRlOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHLbIfF99VKLme6Vbqd1dOK6R0ztKm6j0PFhi4xl6ZktLVm6NWMJS8uDKG4dxRtWCYFkEu0bW5bZUvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyBhIwYo4qRNqdRtUO++o5V6Hu9O0DpjbPxScREvltrsHDZMRgFfe1OrGISi5pGmy/7rFS/YCcMms4LkgELa378aTiTc6HMjoAfxaBjrX27puDMwYXLoEPiIhdTrbbAMB1RWHJYQ/HeHJ3ow1ybKT4w8cdVdGEDSz1nX8J/7J+1ONYOnexOTNWL0PJ+X2fy9z4HGXTL4rBS7bUXfYiX6zhTSR+EYhUn6yngsHxKdieRYm6EfCirzLRNjn0y093vawblg5fuBTrJoOuIYo/f2D8DYMoTYU5HxijSc3R/HQ5ndOSHV1ZqHYJlRCWbeSOoaDbQLbwE2vp5pEelJFGUuidkAAzdkf+JEEUBxARvQm1MnJV9ui98xHoOIeAXRfAiNJWS/vNeMNayWrJD8Sy/vIH1hzmCobOs//DPPxyTJWJp78erlt9uTitJs/P9zr8kn/SVfbovfMR6DCZrVxtmjyhmQ0Q8ygJvXemcCPgVyqAsAKSDojujB2Tk0OvP90zT1HixfGI9/oyonbPz/c6/JJ/0zJ/bYDVRTMKnDRjqcd8g4QoNNOoenXDrx6uW325OK0mz8/3OvySf9oj0QCQIThh6zRGdrPOVnAcIf+Ax3a0gC9qoHINnqNTQT1zWClEYtH4XLjiOTjsUy9xovJ2mxAzRLvnX2Duhfj3UWKJQ6R9GzprfkM6pnQKu/EUKWXiWm56g18ZZFxsrfbJYWSVT7RZ+oEXDTEvwCQNM/IDej5ATiNiAaYT8fxOjYh1BCfOPQGUr15D2mwrLWLJ+TtsdRtZ68197s23yhybtwcZyZxxotq7z0WNseUXcT1zWClEYtH44v3PQhoFfMUAbSjVcAROkaTiTc6HMjoIrMhDJ8h7hkJV9ui98xHoOIeAXRfAiNJWS/vNeMNayWrJD8Sy/vIH0GY0NzhgYSbFnX8J/7J+1OtNo6E8jNFVK9nRyKfoFLAiuhk12RnH0iHEcuJ+RvSwYEbVgC2qNq51vdoW/0sn1LUAbSjVcAROkaTiTc6HMjoLGlyNlJK9HrZhZQQ+h6x8SlpzJ7lSVPqzjgq5bS0R06hLTvtFBaWuA0+3dHKmEX2qg18ZZFxsrfWyY3gKarmfzzy9/ocWiuDsdvv+2BTmcjRYAR5glqdZXP2IWIk85JlsBYLB37rmkwLJ+TtsdRtZ4b26QCci5mEax3W73WWWwNjT7YRXs13sfKXoCJJkzFhLHJKXFkkppYuBLNYgSP2e+sWjoPqEC7Ui/m/LUJQgEyK7mC5X5SWTCzpuBjY2VybWHOYKhs6z/8gF07HWFlZ8BEyxyfFy2sCfIfFKmnxE42Wdfwn/sn7U65BCN3vs0znJBK1+Ij3uqfGv7VJ/STSYI/AaikY3kVDj8TjtH703KJFKbZMim8lWqDKkvY++ZbwXH06B2eQclnnwDziWeYZMxFAl2kc/PTz5mP5+TWtcwA6SQqlZ/JIap2LWt9YGv/5uC8J9pII1u3kbt3wfQLWjMAAzdkf+JEEZ2dztqlDtBrUk3hgaBzAWEAAzdkf+JEETivdrk6lKQddYobP4gyVh64YragtYXl5bKoTVgs61uDiGXIKjq8HYwj8Yi2s3f/YZG7d8H0C1ozAAM3ZH/iRBGWUfBfW6m7plJN4YGgcwFhAAM3ZH/iRBHJh+RMU61RM3WKGz+IMlYeuGK2oLWF5eWAXTsdYWVnwCNAR7eDv0atI/GItrN3/2EASlQboJTlvhLubMjDCne3RN7coAtNOaQj3godUGkEVag18ZZFxsrfLJ+TtsdRtZ5ZLLXks2tPasMER6L/UoxtYsUGP1DXPVuvJr7TUPUQSdPFnlTm89XDNqNUk/03fnBGKMGcxfKDwXPKxSUCjyID8FPB8WT8BcdP6wUL1mayzi2DKeo4lUXhNqNUk/03fnB+HftKVLPq9lB9wchIIhkn4O3bPEuSu2C6mAJ6OQzVt+LkxM8KWrfovasFSgZCszC+cTnAo1owFGIKO/++klhwkFS45SEGu1OzLzf7kXdlezokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyMj1EomkBOXDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8Y5nH7tHlcp0q18fGnEjbL5ZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkxLIL9TF1yaItfNaX9JCLjgltvwaKfnW3SDxBDjrObGCRYbPk+prwtwaeSEc5Yud1+Qkas+/4BSqH1MVbgl0uWN9j5IrXuK7RikPVymSji9NjVXFquNthLJg1MtGwBlMyLZZzmiwPIDzqfGpLh8RcwNAhoDL61JMcTfs2T3tv7quYNTLRsAZTMi2Wc5osDyA8x+uHWPs/vISQIaAy+tSTHE37Nk97b+6rmi6syZn5bD0l7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHKDJFSWdxsGBqsOoW0atmaESNujLFNzqC/0WqMgNUJzn5iOYf8n1yOKoNfGWRcbK380nLhPTehIoyTMWzs4hE/uujeYOu9Pds6cLcQrv4Vv8xtd7T1IVlmTGDUrUHXao0R3MlbIhFGnUhNcPae+bvWdJ97MyAr7tlzKLBMAY28JyNV9NkJ3IgcyVhqsillAnUn7zkdl5xa5VbPz/c6/JJ/2iPRAJAhOGHjF9B9IdWyuosR10XrjdKUSnC3EK7+Fb/MbXe09SFZZk7+i5nuKN2JviuZN+oLRoUeDH+WIo91q8IwLgaoSjBJkPvdZNxVnlCxhrvt/y+YAdjfuoxOiR3gsee83d/nVokXXaKtbgW/t42sDjs+wTFF+mkNSNuTw+Vvor0BFbSohZLVkUaUEPea4ASlQboJTlvmsezOrWWHiuajkcM0HTJMWiAiNHs4agN4V/WU3qpupr41nPGV3Y6TXw9GCLAz0CcP+o6hWtmGM88v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk6AOksM/8I1x8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTbAH7uH46mzpwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkzXJ0x7MafQ411wcvqAkiUBEmm3xCd8NkwSYd5GkkAmBGf4YnEaS9txs2lJ26ewe1vL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZpMgNlQbpC1BX2SE7VNdvUKz2YvovkAtYrOBnT9RdRgfB7eb1JQyS/0yObog6RQ0v473IRwcQ1EcBqWLrsELj/rfsD+cs1GJqAali67BC4/5rJsnfKlvHrWa6DRuzrj8afguSor3iZH4tQK9hADT0fyy0L+xyfY2XLxXxvnwYbtoAFjRhzGDuIjMwNFIJnmJW/uWnbOerDpE0OvP90zT1Hglga+5SqahCu0ekMY82N2FfmFNVaT4O43/ltmg1QS2VNJzdH8dDmd37zv2mpBufb6W6IOb4qfh6+VLK8seYNEcoM6yNJL0tWnqZ401uSJ4NJV9ui98xHoP6VU10G8wPdELn3320Md3Svtk5SKcFdH+1GeF4Si6Wd/aqByDZ6jU0k/tNCZ/aJVWzpuBjY2VybWxHRwpZ1wMlRdXRhrhNplWBRUaVK6H+WlEJZt5I6hoNbUXfYiX6zhRTYudYE/V+fljPkr0erOkoepnjTW5Ing0lX26L3zEeg/pVTXQbzA90QufffbQx3dJuYDDnBCDalnXtMOX+a8Osu3BxnJnHGi080P9Cl/ZvZAAWNGHMYO4iY/jKogrB5sT+5ads56sOkTQ68/3TNPUeCWBr7lKpqEJxIurGghkjiWL6OwOWFQ/LgTBG9KOf57W9nRyKfoFLAiuhk12RnH0i4Lwn2kgjW7fJ1sawggAx/TMwNFIJnmJWb09PynwLIq6BMnUsLXnpay9DQhuHiJm+2pRo1DXLjhPo0u8+V8CORkoQjcQ0YgtNXsXTUZz5XV3d5Maz1rRTm8JtgoS4weo0mOKfowoW+ahzuGqjhemxi5DRDzKAm9d6MqNzV3NT3KmPkfSV8TSHu29PT8p8CyKugTJ1LC156WsvQ0Ibh4iZvnv19416+s1qP0rybbs7BjPYkKoSzvZCqULn3320Md3Svtk5SKcFdH+1GeF4Si6Wd3jDB8xfZFR7y/BJV9UtiIksRSJshh+sXv8+7LxR6pPlgO8SRjlp6mXJ1sawggAx/X4igDS2/7NN6ihOEYXlsHH6UWWojamjFFJTuU3JkJFITIOnSECLhxqA7xJGOWnqZcnWxrCCADH9/3lfsRDvNEXqKE4RheWwcfpRZaiNqaMUUlO5TcmQkUiMrAeylkdSiIDvEkY5aeplydbGsIIAMf1PuFDQfNhSNG9PT8p8CyKugTJ1LC156WsvQ0Ibh4iZvvZ1ix81CJrq6NLvPlfAjkZl/lsUehay7kZf/QH7nSII3eTGs9a0U5vCbYKEuMHqNE54tjlDdovFBuuhctBCF18ETOWt0KBunJYh+oizR4EnM1ILnQKCFfP35BbVn6rNwf+41YaofDYGfm9BEi96ay8cbi0ijlgSm/03qOIzJ5d08v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTjq/W/DnY7h/q3YFFR2s4AFQEo83cZQQWl/ux5LaKvyLSu5NX3VJkLh+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC4kq3srN7+p8SDYYEZZ2nr5tri1hIYa7vqDpZWXNzWXSk5Ok5wGBoKhccAKiMeC1ZbF3uU2H/DCyQO8ZxWsk4lK1bfk3tLW1g39e2VsGp8X0crH0S+o222lQulnY1n4OaArbEW9wUUhXAMq5V9IKK+rTc1BAUKC0PB+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwty09P8htiA7a5WfCD8gy7r/pfcYVzcVjdk+/6CBSpoQ+9c4Zcw0m9czc2icvd1bNFLnqqfezW6ZZj0EJIIrJfLWBa/jGXMVR2l9JlDWvKVW+0bWTRss2SZnlFEOez9nWfwPApFPJfc0sL8CR+13B7XRrMkkuIJQ4G18mOKd8EkIcL8CR+13B7XLlk89pyoh1QKcIdUpPLmJTRs7EO/weafO0+iUPoaTRHN/jys/Hw1bLBQFOQvZ3yiVjW1fM47WbtJi8mo3u4XzqNUbehcOlfX6pOtkR5QI7rnkyOhxNuHYvuKiazyQ07CygDEbahTo5m18mOKd8EkIcL8CR+13B7XMT65WrDAzbz/Pwx6skM0PyNs9/cmJsZL7wr+i+5ntM2iFnIMegDHVIcqqiDGcCkSZ+CulQJw8O09JiKzD8Imx+Hqxs2JxBciLlaEv1OfgYXAWCwd+65pMFwo8iTPXgTza6sMkM+revcAvUSs1lj6hRJXmGt6H2IFVK+VCqi2ieWYCNJDPeQzSGIGWLcbAeNGLwL0gn1Absu9nRyKfoFLAgZ5rjNF7xI7DPbkBzQdmF5ozpLjZcXpTgBuhDVR39T5E6RAzhAj/jcrWK08TVYnH5CIcvGdXEvF5MB2D6eLykhTApSq93f73Vh5E0gkpomTYDx0oL8iJkpmAmFR3LKaecIKQH9xapKWm5wIy7VEbo3tIPi8/JGwoF4JAwcpRs2wpWqh0Oh2IWWWGOmg9F0eMyi8nY8DaDPkAvSQSN0gihcdg1suZ9E6/4+SAElTCEGyNm1NPq7LqJTBH6ab6nFM+gGrw5g00TiREtRfj9IyqtXeEjXO9/j/Nx3bcYOqDhgjKJnyGPmNyWbhwyaAxLfQPadxdvymQ2UtQkP1FgSCfe//N2MTaHVG9xFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybekbiNfBS06ImACD1HOvDAa0//yLJZNFE6cLcQrv4Vv8e66BPmKRG8X3yLFENI5ayaw9aDoVJ6fITuyUW/8exDiN+6jE6JHeCzQ7e1k80QpnH0km0H4E0GIpim5dgZrhdGvQikJWPE7COkoH8fk64rYMHZNkdaymPSsoshgLutmaNWYnM+lVTIQoJyPBu6KPyFRWHJYQ/HeHIHo30Cu57AfeHD/Xt+YMt1KmP/44N2Ur00RGcH1v3HWPaJ1wSxBbGs3NonL3dWzRF/O8s64DUvK6maR0RWksW21F32Il+s4UJGTiO4QTk9YF/eDlOHv3ONSqnv4fBK0vUMVJnXwC3aifAo4nHH+TJzAgLGi5HPbDIIvT+UNORMR6KJwYfaUHKD4wy5xLR5PYm8bRaLOOqhPiN7L9OTBPDcFOlKqDpMwoMT65WrDAzbwJXZAhY8A6KydQKgT5HtzBAWDQJ3KBpIOSxWonF3FK3DgddvbdX6MFbUXfYiX6zhTBTpSqg6TMKNTVqIMPVmlu7It+N8s5jtvO1wO9faAMx8EfppvqcUz6rR508ZTGndESmAAgaPD7xeHDJoDEt9A9m5wIy7VEbo3+TnSdpOBCTWQOUT7p/Z+uQpenfM2t/MWeuCv8EL5+zg91bZfIhUf8VFYclhD8d4fmoETK2hidRk3mPOZwD+gIsraGiqK4eHXBH6ab6nFM+q0edPGUxp3RruSmgqSTU9Jr0IpCVjxOwh2DWy5n0Tr/HnR5XoeMh83g96C2/1xECuS3dzsckfdslM7FV/qoydnBYUSx7a+c9tUt/v2jOF9eb7TfrcgcZ7Xx+2VROkD97wYIH6B0tKspr5EQVKqlJmfsY21T3uRMTZ+gA4ucyggfHcyVsiEUadSE1w9p75u9Z6A9PRfdxrzkHdtxg6oOGCMomfIY+Y3JZuHDJoDEt9A9m5wIy7VEbo2L0+ewznAFapNpD2brUQubxFu4E03+Cv5UzPyzuUT83Tjgq5bS0R067N9ax/BvGXN+TFSQ0YK9gN2PgnOG3gnzWXbbTKHNIjStmTbdvekH8lQEo83cZQQWgpvZrikp48q8C1sSUY9byx8pWXSZSj1OTc+2J5/NvU9sdRRleC9UaDQ8NUcz0oJwmo59SWkrRX43h97F8QR2vxuofeqqBDYthdcP5rXzimWfsrlKyYgDb3sDzbt9n/3hIJBpxOyBDyXET/gv9cMW9Qwr+bgpFBz+KkK5zvp+JMhffZCb6FM75pqOfUlpK0V+4bCC/vGL6oHSTZJrR1SxcFKYnU1vXRMSUJGs/haPEoTksfIdYTmdZPJ6/nou/PGxHA8aowldih1IwM4TVqUcszawSr20lhs4Ct8SvCt1vNrDAsjo9oSIbdEJJhArXtOpzHuyememPFJHXemX/sBPK2N7nopOgvSGR+2F/tKtrZbP34Hlu/oQqJ64K/wQvn7OiIXU622wDAdUVhyWEPx3h0FugNZPx3MjVFQf51dFuydByPWgy+P8E4NxIMYhzmp74cMmgMS30D0UiOnUM637J33X0A/a/canHAISymnVJt9UzPyzuUT83fwKGpys6MCqVFYclhD8d4dBboDWT8dzI/kE66qo6GUKuJtF/EYKv84xk8wvrRXYtexjbVPe5ExNnGokgdKcFFOQAX8ZQKQb5lHiC0UNN4IyMDvPQvnae4ogi9P5Q05ExEFugNZPx3MjYSBlwfxDgEE3xUva11WZWPSJ52KAGWjkgiTgKVADo8A/AaikY3kVDo8akDvDFsQrWIIAIds2MSryTKIkUcCMHWlAqlLKErBpiKx9BSOhCks1g6d7E5M1YmOvvVYKodJr+lsWumkQKDoJbxjfsvZQ028+re2pHp494cMmgMS30D0UiOnUM637J7KxeGQcqauwMHiwATbD+KiXv44E5MyRAM3NonL3dWzR2rxXc96ZmxfNXPFu6k6ved+qVChex818q+H8f8FSTy/C4OEyxUpTD+dK/+s2YPEJSATDtgUv1yQ2sEq9tJYbOPzmMgugc2g+JRLCGPqyGfgcDxqjCV2KHUjAzhNWpRyz4JW1MwKc75n/QiY+QmZbGq2LiTlmATyVv3T+/Q7PTTlwrlUyUpbX0v2CsIMYRyvGPwGopGN5FQ41Hkx1gZXsVyvkwtmFLeT2tJF+uavjAu4iQpHci9AjyDVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3h0FugNZPx3MjlTUrDTQILBI9LaGidc4WLxFrKC0Tmdo5WIIAIds2MSryTKIkUcCMHUlxZ5IXsgklf/BMyL01X6N/rmlOCs+pkSjSrOYz7E2R7GNtU97kTE2caiSB0pwUUw96uxB8fpVr9048aZniKCFjuqaY4wcJjimKbl2BmuF0a9CKQlY8TsIr5MLZhS3k9k7rPVFPrbfv7QnN/bBZVR2LSRYue6xyQoHGXTL4rBS7bUXfYiX6zhTbA8chY5Tt3PvuBv+mkgT5Y7qmmOMHCY7qfUNT01XmRmvQikJWPE7CK+TC2YUt5PYztvDHYsTTMYXQY7khYfYai0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+InZrtBfc+pw72O6ppjjBwmOD7DkI+4jM/Jr0IpCVjxOwivkwtmFLeT2T5+wWP+EdwWdf6nBsXgvDuJMAqrxFw2na9CKQlY8TsIr5MLZhS3k9k+fsFj/hHcFo6Fxp5dO7pXiTAKq8RcNp2vQikJWPE7CK+TC2YUt5PZPn7BY/4R3BQXLDiN0wNsZ4kwCqvEXDadr0IpCVjxOwivkwtmFLeT2T5+wWP+EdwW3ab7bgqPU2OJMAqrxFw2na9CKQlY8TsIr5MLZhS3k9kbDk5mdUyTuDles2xfXwOmfoVOgPrJwDliCACHbNjEq8kyiJFHAjB1wC4ndpowqb6YMr33hCFL5KX6FkM9GFm44HXb23V+jBW1F32Il+s4UncaLrFKUm4cJ6tqYqc21hg5XrNsX18DpOIzwpEsi3BFYggAh2zYxKvJMoiRRwIwdwljjrqUrWVetifjYzngz52O6ppjjBwmOHCmANQf1H19r0IpCVjxOwivkwtmFLeT2ziQ4naM5jK5XqIj6MJT+q8IIPxBr+NBQ1hAIlb2xXDLC4OEyxUpTD+dK/+s2YPEJgRmzYoq7PH2mDK994QhS+Sl+hZDPRhZuAYCZgsLQ7uZtRd9iJfrOFKcnp15/O3Tds/3qo5uVvb80O3tZPNEKZ6P33I5QEiCsZHXZPv29g4ZtRd9iJfrOFKcnp15/O3Tds/3qo5uVvb8x3A7vFzCo26P33I5QEiCsZHXZPv29g4ZtRd9iJfrOFG+wihoEHfiJ2yooR3rR3bFjBfVosytm4ymKbl2BmuF0a9CKQlY8TsIr5MLZhS3k9v2s1D2kyMWnMdwO7xcwqNuLSRYue6xyQgmtcTed3vOWbUXfYiX6zhRvsIoaBB34ibwLWxJRj1vL3T3qOLnPAV0wO89C+dp7igIuZ8gz9RNAHChBkRHlDB5r0IpCVjxOwivkwtmFLeT2JmzTkaATZsi8C1sSUY9by9096ji5zwFdMDvPQvnae4oCLmfIM/UTQBwoQZER5Qwea9CKQlY8TsIr5MLZhS3k9sav0b7CzNyrB+CZbzfAuFIBYNAncoGkg29zv0N7Jz4/pIRh8L25QCUumDR3Gts2lAa7pznMtw3ROjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2R+JOhZGjs2qfBzt+PhrTzkgFxsc7HdT9fL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk6xambyK5ZxNCQ3bmdTTHwSU9XczSMtPKB0nUY3H7fwi3/5iZdU5+2h40l1lb1OXtEisFUyYgp+4QZMeFQwgW5KeuCv8EL5+znckWoY56cgvX/VuTF7etTeuD2pzivrOKu6gnuh/ZnB5q0SLj91Ue6/VmaIohTeKhzh9A8064LSKe1TYiCbn8biUzsVX+qjJ2SOL0yshwRnPQnjH9mQ9QSGuH3+zHgnhl/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4Ull/LbH3nTg/ncOa6ZVqVl3/JOXLbMggimqlb30GztUQlm3kjqGg3pxNuRzzOsSMTZrR9MdAnr7whiIHij6dZQOwMiM8LK2CMDhSXtJ91aJOBXqtLt38tsm124DgR058TZrR9MdAnrRpQvZGe7I5DWxBg7V9yl67wLWxJRj1vL3T3qOLnPAV2scQE1hVaQ5/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx3NytrwMXzq39GHaSvEAEy1D/pkSL3Ck8oJw1b4i9AlPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPdYOKzBbKsR7Zlh55SO90ReF/if0p7KnTZJCN37lemMsy5NmanRy8FgfzBNpXKiyOgnDVviL0CU9yZ5m3LYOxnSW7iwRLiwVVPkJK4xKvxsAYGsMjn6WTZgrEB2sHJXujlLtWFFFLAuAePxLG2o3WY6dZEDtKimZy3Z2eIQiWHAGkjwuV23KD8Ld0RaCT/cJAD45zU2m2Hr1Fj5+cursX8PU31359fs/CoNfGWRcbK35ciTUmVl2NykxGQ5DlU5Nw63KRBzNiNf7PE7sQG274owx88GWye2AtpqE8auG9/XtUHj58x068MqDXxlkXGyt/BSZctyWYz9nZJiru1KFI0iuBZrA0FO1azxO7EBtu+KD8BqKRjeRUOfvr28kEsfd9sR6DJqCUVys++rW9+bixxqDXxlkXGyt8VBFNCDVDPUGyr7gXK2UTWPwGopGN5FQ5TPAJSXOY2s5V3hyOyNkFbPVHhZqWGaMyGQ9GMRcfna7GGk90gjqWqRN7coAtNOaQnHJK7K5aHezzRsi96Gpp88hJqX57rjKdhfQeIFI3IYjxStOXLI6x84BfQhOSDF/P0sPfoNAGcc7/5cgVXFR2tYX0HiBSNyGJCwH/1ob0ps5gWzBccA5VUHXrULF91ybyoNfGWRcbK3/4ndrcguBFsbgaw7SvbuK23zksPIxe5DMTd5fHu6/15l2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkzn2Cf6wkDYml/EDOfVfo6o/nPGhn6hGYoQkpd/eIKhcgUQpVDhBElXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMzRXvCR3DN0G+0363IHGe1K7v8TeBT4K3cskGuRzF0Lqj3wGdt6if2gyXBNg5UGkNz6RQbUJEjH6nCVTc3M8USqDXxlkXGyt/jWBp/Wq2ELzTvD6BOH7n/T5CSuMSr8bCYtR94aBC09T3g+AKY0uCZlvEqUDwhQIVmFlBD6HrHxOkbkEPW4zzky0YT4BhZbefQq6vvWj9+6Kg18ZZFxsrfWLfuNP5FCVhn+djsM4CPbbPE7sQG274oGnkhHOWLndfXqX1BcT19fpeVSw8eeK1BRN7coAtNOaQriyPp1ahjhotDm2SkoC7m+fu3S3MoLDAS1F+P0jKq1cMd2hdfixOdFsHnHAppJ7VR4gtFDTeCMr/dvNaKAYw2bEegyaglFcrr+tKYXNgMSB161Cxfdcm8qDXxlkXGyt/pG4jXwUtOiJgAg9RzrwwGtP/8iyWTRRM1X02QnciBzNsqKEd60d2xTUoy/TGCk6x/8EzIvTVfo1M8AlJc5jazpwtxCu/hW/xMVz5kVthoXzWcGAPK0V46wh/4DHdrSAK/3bzWigGMNnTSnCmLL8pXMW1IP+hPk/wG3SJPCawg3py20QfQAbjTSzfvRkyAUokJXZAhY8A6K/MxOyzyBlmzu2EpzdE/7SZl3/JOXLbMglq4EdcFYjuQ5qBEytoYnUZ/+P+7IcItVZv6iu84/15wkxGQ5DlU5Nxs3Qp6R0IR63PeoGGTEiybRNdit7e3UtYqosG7fI4x2oSozaJuiEtz56FUpyEGrT0a1ENvqr53g/5OdJ2k4EJNZA5RPun9n662HHNbW9CXUOagRMraGJ1GTeY85nAP6AjPCEqjHSZRAtUt/v2jOF9eb7TfrcgcZ7WIk/350jaeX8FOlKqDpMwo0Meym+qb24sTD+YW+beQ2k7gS1r63R5D0Meym+qb24tIDrLKTtzWVLPE7sQG274o23Q2WICsRes94PgCmNLgmU58cFTWg8C+2bMgPed1BertjYZMeyJerR1fzzHTTChP/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNbwb5RoGmEZTokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRy8OhdHeSatRpXvxEyKrRaoWJcflCBAP5NFgDLnvCTtyK3gxOHXjh0z9IIlUsHIlfpipL/2CO4stc6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUckXQE/WWLPjpiKx9BSOhCks2jFsjiZ72mKZkUi6qw8jhtrLqfBnyQDMNBQUlLIPgxdTj4HLci4iSZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYwZO9Yy3tQ3ehKlCAG3SxEiA3IsFghRLd9Gu11ZTq/jTAWgaVGAwawWxHoMmoJRXKC15MEywTNkCSoGtWHrMQoIisfQUjoQpLPErZMKxxufumABk2dOpUihUEU0INUM9QuKPqxC7RtK/FkHJ1/mvrNXENawMGez8Ukkgl9/s3LB0fXVUrveNjQvGTg7NduaAadnJ9malVwu48NHhaUBQbNU/rBQvWZrLOYGxxPxltFAHrmtzLenEkep9mQ4Wktpgjs6bgY2Nlcm2tMg/TH8AwMJuwpfyRpuHUTMzqNaAeQE0/AaikY3kVDqtJq3Ejr16sl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkzn2Cf6wkDYmedXCV/38kOdJL/KburqFcgjeZ9ZJ8cmR228aV8mHTkvAlCJBb+anty3CGF5nDx2yiZjvtPUD3cQ6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUckXQE/WWLPjpiKx9BSOhCkuti4k5ZgE8leaMqCF3iWxbsDbvaSa+SnqXIk1JlZdjcg3Fg828WMI6IKLVRP+gR5C0Tn30WE92R1UX+GZmgzz/ytYQDdKpC4RIYQ4pQCMNLfpbFrppECg6CW8Y37L2UNM0g3l8ZIe6XMnwQn5HMaOUpssqxz22YnL+6xUv2AnDJtOzjAXFxvcUFTGB6w7KoFvGPbG4bYuGlkXn8EctYzTULXGgDy3/zrryFchVcU6H8A8+rMr90dyqBXbcYW79+rQYkw79JL0RLG8KaPHf++t9DQUFJSyD4MVNhDOo5YPnV/ML3EO/WvzNjhwIGUocy7GoNfGWRcbK364UwxpT64E0bgHGiKZwURSGWPttRvxKNzct4uUjQIxzDY1iAzS0/iLW6GR/nSUEpDB4sAE2w/ioldmD65voKkpAhoDL61JMcTfs2T3tv7quaLqzJmflsPRZvMPH8q+ASWN7AhKNvBXLfCf1a1PYXmsvaMWHyZ3xknEK95r9tEWsQvZOoeWO9V/2iFgisxvhsWPX+/DM2Fc07akzeH9Wt1Gh+pQtBcKOBtiuoTHUj00ch4hSVNwEjRjHr9xBLHM1uZFDTb0YSVoWb5lhdorn5WioNfGWRcbK35N5A/ogEMdEE7pC89/+gBNvPguC5mNDfs6Y0n7XqYAlEPQTFGz2CFt3DCpm/rPLLv/T1vKOzVz/Z+/Svll0ePMNGqnTTkK9GaZhREc2ssOTdrLr7XHPBx71viLCyT7lmPaIWCKzG+GxHa0KJuCFwkf/ORp12Hykb9bEGDtX3KXrUDIdIf3PYBDhFKCN6NmkhbPE7sQG274o/hp0j/T3vlOu7pE3AQPuKc1c8W7qTq9536pUKF7HzXwFZY3SpS4oxMBYLB37rmkwrhTDGlPrgTRwOfDfS97jg9lAi4NgHX0dzVzxbupOr3nfqlQoXsfNfLy95nBhp5Cq1i5t3ireDk/AWCwd+65pMK4UwxpT64E0cDnw30ve44OVF7bvv+7oUQBKVBuglOW+yaF0zM9PAM6hKlCAG3SxEvrulmFJfXtIIC1mSktdDCCSSCX3+zcsHbxiooMp8WxajMLLxsQny9w1epxaUq4HuHbNeEqJ2HthB/0N7qXtgUuCFfgvXHzSERcjFoDC4x78wx3aF1+LE50ETOWt0KBunDb9QuSHDNdeffqlppcnQWarsEsLMzN2uWEgZcH8Q4BBM5V7vxl6SJb/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyPXyMGM0AOBdKU1eiC1V3IonbrQyp6yo+z+rSyRgpHm2ORIAnEKnqt/5/InIEaeQ1J8mHG3rjn3X0tk1hU4H4JjfVtWtGMN6sIf+Ax3a0gCOpohsAwkhiKTT9nj/iUo9ZzXgZ2p0Z11lTUrDTQILBIXgCM814Ju2YT4X36zRhgVx2NGG0h3rs5JFqDMGrNoZGt2IWtDebHnOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHK7V2ObpTkM5gQx+/QQpBHCvd/P1Ff7hG2sfx89aGbWJTQbPr9FivoV/N7n82cN5/tlpcHtu7xS9d7RLHkYpbTg8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTIGEjBijipE2+ifnZ4SKPdrUda/Df4hrj5oyoIXeJbFssqisAKpLZ9Cem/tdTojcxABpLkx4DeSDf2Gv1VRyY95CsWg2rHz6bYv0GcUwNsoLENeksuzUqtNiuoTHUj00ceiicGH2lByiyPilougH/hSv3EGN2Uc6Y4r2TfVzeBQ90pTV6ILVXcq/KKj79mo3iFaC6+bC2tC6oNfGWRcbK37m+Q914Yne8O7ynueTP0rbBD5tH9ZtoSdmu0F9z6nDvTKVS+fDCQUIcP6m2H10prSsdqq64ZQeSZ3cPvv/yKnPNJ+YYRCcWoxeAIzzXgm7Zg3D9ypd69YhGT/oQ8kyzcVRGMsxgLxhBDIAPNh59rU4yDMJnGS3tOag18ZZFxsrfvX6wOe1vxRKCsw5l+Vg+cvlCm7f0w4BO+I9lCC0nhdcqwwIr3m3FxCY4H+AJFAaTOWqR6YvN8kJv6qUwOF2sJIPdwd9zyGAfk0vOqY+3Vq3jq5Hw4anVxJzKnuejMauXvasFSgZCszC+cTnAo1owFGIKO/++klhwNwlulwgnidvAFDSYFL4Js0St62alONtI8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCThSWX8tsfedMrVwrc300F7xhwSrMeIlNela/HrVedTdhtLXichvJN8BkNGj54zAwZ1fjaJT/ij14J6tqYqc21hlksteSza09qa5pyonMfqRtXzt8WiAJU+juBUYL9KuNxrYn42M54M+e7rUQwr5O4qWb182whRLcE3W3lShrJOaQ6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZchfmhCxn1pnx5n+2CwYtJ1O+FoYYQh23l2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGahejh7pY1JT+yLfjfLOY7bJTl8/fTcwAgg8QQ46zmxgkWGz5Pqa8LcGnkhHOWLndfkJGrPv+AUqh9TFW4JdLljfY+SK17iu0YpD1cpko4vTY1VxarjbYSy6My141/1x+nkNRJQg2YhY6nxqS4fEXMDQIaAy+tSTHE37Nk97b+6rujMteNf9cfp5DUSUINmIWMfrh1j7P7yEkCGgMvrUkxxN+zZPe2/uq5ourMmZ+Ww9Je3XicDJZZfQ1pFmvl22ruVzBspFARCWZacAGSF9jAb2K6hMdSPTRyct66d0DJZamSR3DO4+l0JgnofOQrTPZ4+wR6lpyWnXMwStDVzf86kHmWvyhCceuiacRksE/8TIGhU56WSokhn4kRJT0dzUUrkNRJQg2YhY7MacMvqox5wbplQI+OUr2v2cFPsPBLzDO8hoGSxBhpUe3hqEB2OSd/AWCwd+65pMAlwZq6GWDZ8neP0N/uBkPNmDmarMzI9a/fiWhaYfnp3p2QUyLF9II1d1JF4gmT8DR5lr8oQnHrohGnVc56yB9loVOelkqJIZ+JESU9Hc1FK5DUSUINmIWOzGnDL6qMecODnDvG6Gh33nfwQPIkiYeCTSjpatecfuicjgeVVuCXb4kRJT0dzUUrkNRJQg2YhYyHbx7iNNVS+4OcO8boaHfed/BA8iSJh4J3/JI9BHpnSJyOB5VW4JdukBz+FUA62mJcRaHwDcIfmaFTnpZKiSGfiRElPR3NRSuQ1ElCDZiFjWSy15LNrT2oJ6tqYqc21hheAIzzXgm7ZwFgsHfuuaTAJcGauhlg2fJ3j9Df7gZDzy+j4OUQtrnjQxjvZI/ggvwBKVBuglOW+XtMm5Dtaery9qwVKBkKzML5xOcCjWjAUYgo7/76SWHAa5uKIY/O4dFuzFkAKLG9pEipV0iWaBZ46JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcjI9RKJpATlw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwt2nglrGm/E9WPtaBNmxroM40BRQKurwWcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMSyC/UxdcmiLXzWl/SQi44Jbb8Gin51t0g8QQ46zmxgkWGz5Pqa8LcGnkhHOWLndfkJGrPv+AUqh9TFW4JdLljfY+SK17iu0YpD1cpko4vTY1VxarjbYSyVVtw4ikZM8Kz/eqjm5W9v5CGwyPdZ4tcu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6U/ODLJ/5ShxMVz5kVthoXzSc3R/HQ5ndZL+814w1rJYvxMuc4I56TiIQWBwpLzSMkIbDI91ni1y7cHGcmccaLbdTi1x3mcIYkNEPMoCb13ouxPUN2+8SQh+uHWPs/vISQIaAy+tSTHE37Nk97b+6rmDUy0bAGUzItlnOaLA8gPPDKs7TWGVK9XaoYn9Prc449xikmyUKNrP3gRvClmu+NJCsWg2rHz6bYv0GcUwNsoIpCbjHIfzrNblg5fuBTrJo+1KC2JQX44Utul1WCB0BCyxRMGNmpkmPhpwBPpy08Yi3vWY9SllqwBP+4XuuaQmQoRt+3LBo7m62Wc5osDyA8y55r8llU0/ZrPQ+NCK9aHLwN83ru1m6GeDLWBziTG2LxmaTqZuuAWyoNfGWRcbK35ZPS1/oJxSYKCCmunWnM5QZIBxpTeGKdMWY6ModpxG/p2QUyLF9II1UfalmxjPZqqLPvKheOBdNAAytXkAZIRP67pZhSX17SBjw3rHtyzD6j5IASVMIQbIKd+5bHLOu759/H8nlmqDAKQm4xyH86zW5YOX7gU6yaDGc3nODWG+mF5TvcqXOBv2KOoV32B9NRHWrM16ZTDZB2yooR3rR3bE2lc2U2lpm6Rhrvt/y+YAdLsT1DdvvEkIh28e4jTVUvgMJfh4Q4NFolk9LX+gnFJhEjG8SumzCXw4IgyW8+QWOZjySmeLaPsoMHZNkdaymPUdN/wHf7/99FpYxxog+HqYxfQfSHVsrqLEddF643SlEIhBYHCkvNIyQhsMj3WeLXLtwcZyZxxott1OLXHeZwhiQ0Q8ygJvXeiIQWBwpLzSMHnvN3f51aJG7cHGcmccaLbdTi1x3mcIYkNEPMoCb13qnC3EK7+Fb/HuugT5ikRvF3O7dk5YeTiJ6c9O0Bg63Vmo5HDNB0yTFBEzlrdCgbpw2/ULkhwzXXn36paaXJ0Fmq7BLCzMzdrnaLBLsYs+9qZ2eoXVhTTpfOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHJanN3RpC24j9sqKEd60d2xo9Sz2ROrnOLCxkfGYxEhttDnumNqBSSRHNYQoPY+k1ez8hPZk9AeGbReBOnbSegyOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2Scckrsrlod7htsEJq8gOaX2qFdVP8L/mHkDSvrx2tRcC9/atjq3bzHy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8V+zhAWVmL5N+OkmS/0g18es9mL6L5ALWNhnSUVsTvDFvAtbElGPW8ujHXuTgWAjAGgKKyLBBcfgpH+iYXN2p5bZc0hgaXrT7MCUIkFv5qe3PHrYr99U5d+ZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjOyGzJ84JlP4hMY7OSSvyJ22N71FU5195jjbP1PE3yMXysR4oKvE8eWcTxE7hd+vD4JDYB2RmqX0HB8UTeMQO7rZlBIjvxIe9Wwo9mk8m5UvDi8sDixjycgKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTyNOGBYR8d3lP/QA2hnD6g7LT9KQ3pbn9Gu2EpzdE/7SY0DDZRAYBhdCrBIK2a2rrVLEXGmfgOzLMpGPVwIBlRWRW+d+8qtxiYsOf19bmX7AAnenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvroSb6BlUFCI0YMP94Bmjpk3vYq/yHVGJ72xmBfkJZtCUwOnAhonrC5b48tYcnBx2ygqZVyAs0jFkVLDpjziJ0oF/6AsqgYPVWQiO7VtkSldPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuv4Rn9g03rmWQ7/GCLlfEsaQ0qZVTtRlgTVl9AgiCXh12jfX96yewauUWAEeYJanWVt/XtuqXLQQxvtN+tyBxntXpD9uGXz4gcGrSgLn7jD9CL4CnVhh/Zh7wLWxJRj1vLox17k4FgIwAfBactKxaMDwkNgHZGapfQcHxRN4xA7usuQMf/mEHfwCCc0IDM3C7ITYP2BaKjE7bRp6MwmT5LXCM4c/S7Mace5jf3mVivngs+3wUp4AHlaZpBVhazntdDmUWeMkXenwAVAW4LwKrLdlF3o7IHwq++s6bgY2Nlcm3jbP1PE3yMXysR4oKvE8eW/dbflPc4IAx1nQvWtGCDoixFxpn4DsyzKRj1cCAZUVnsDEDhnJsiFEQ0g9fitX04rP9dKfjvo7xwd5/XVcjawpSzvf+Ei06Nh/OtHz0A/7/4aIi/A+pRzn7e4xvVnKJT+VLK8seYNEcoM6yNJL0tWt8sZ8UtQYXMpbog5vip+Hq7n0AJwgNkC7FbctI76sneikkDt4Xdxb1zFq6NmjTDgmXmK7xcbFXjNgG8aKR6EU73G5mVe/CLYAActdTOjqUY54NARHvgdqpb8lZHdGhSIgRaKkigQKicmWM7sg7m9pItp3y7fmTZdWEIpEEohUVnow4N0lW1I5ZRd6OyB8KvvrOm4GNjZXJt42z9TxN8jF8rEeKCrxPHlv3W35T3OCAM8tRgADsBQNMsRcaZ+A7MsykY9XAgGVFZ2yrNEMZFKpoAHLXUzo6lGOeDQER74HaqW/JWR3RoUiIEWipIoEConJljO7IO5vaSLad8u35k2XVPQes58MXDlAGLmLc6c3vQ3yxnxS1BhcyluiDm+Kn4erufQAnCA2QLsVty0jvqyd6KSQO3hd3FvV5gMk3W1mKcZeYrvFxsVeM2AbxopHoRTixdgfHvkmEzb+PGmbCCNZbng0BEe+B2qlvyVkd0aFIiBFoqSKBAqJyZYzuyDub2ki2nfLt+ZNl1YQikQSiFRWf2ZrvKUqlVl1F3o7IHwq++s6bgY2Nlcm3jbP1PE3yMXysR4oKvE8eW/dbflPc4IAwJyuFRLt//vCxFxpn4DsyzKRj1cCAZUVmlMJ3BzZDoj2/jxpmwgjWW54NARHvgdqpb8lZHdGhSIgRaKkigQKicmWM7sg7m9pItp3y7fmTZdU9B6znwxcOURl/9AfudIgjfLGfFLUGFzKW6IOb4qfh6u59ACcIDZAuxW3LSO+rJ3opJA7eF3cW9NpT7TnEJf7xl5iu8XGxV4zYBvGikehFOGgAW8cjr1u0EWitRPGZDlsqzt/VKiRlfMb1+qwA4chQEWtzfF9J0tqPA8XIE0tuMKaIn7NYNLGKAaS6fqqpcMZuHa7Es8geLI/ja5RlEu+u7R6QxjzY3YQRxMkPH3rMdJ6y6pZzR8W2aTStjH6x7uz7JxAwuEmQkpH+iYXN2p5bZc0hgaXrT7O+pqegIeD47TYP2BaKjE7bRp6MwmT5LXCM4c/S7Mace5jf3mVivngs+3wUp4AHlaZpBVhazntdD4C9OpJrLpr8wF9adUZkNPtZJYDDz/BQ0jl5YD7ZmhyYIMEmt5aG1PeAwa8Ni+6HHd5xAZmZC80i7n0AJwgNkC7FbctI76sne8wMcs0KZN2UJDYB2RmqX0HB8UTeMQO7rRz5DCifoymXa2KQlAIYf9qJGCPTekGzXmWM7sg7m9pItp3y7fmTZdcVSVVRNYpozvzIhHbIESW/a2KQlAIYf9hiU/p0DOgMLY6FG8xkcuRojA4Ul7SfdWuooThGF5bBx0Qk33mkBR8akf6Jhc3anltlzSGBpetPsdl8pqchiP0ei31hILaS1AEGZftECsE+Iq4j0S+aVfp5Lek8xFmzmIlJTuU3JkJFIbgnd/TfQURx/RVlmrd5Dp7T9KQ3pbn9Gu2EpzdE/7SY0DDZRAYBhdJ/PdKQSi7mFsOW9w8BUFblrS1TXObGJTkQ4daPsguOMZAQZ7dlaAviH860fPQD/v/hoiL8D6lHOMZaJukqSckHL8ElX1S2Iidn4NnqHjnv7U3OeAaB0Udi4ugDXg6fOPzE+uVqwwM28w3jAwnCbrr9iLumdgI34KSxFxpn4DsyzKRj1cCAZUVnUA23qltv4rqLfWEgtpLUAQZl+0QKwT4iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUg8usmgs1Mv/UUjTNUrsZdT2GdJRWxO8MW8C1sSUY9by6Mde5OBYCMAV06xwO9FNXRl5iu8XGxV4zYBvGikehFOz1lCvexYxk14XgLSZRtKdQ/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg8EmZGuEoHlf2yooR3rR3bHY3vUVTnX3mONs/U8TfIxfKxHigq8Tx5b2wMLV/TWN3lvjy1hycHHbKCplXICzSMXKNqKpH6TgK5WGqyKWUCdScqS0oJ9iCfI+3wUp4AHlaZpBVhazntdDFXX9LD/Bi695zs5PRIUJlqwbTrb/HNEQEpqvazg/7vIsuz6XhOjIDoTkHZ7hGiLD8tbuCI8byk7y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPGxkGe0pm8RZxz38vshk4xKN+o8Y3BzwtEVRlw+CYWvdcB9u/qWYJQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LuByd/PverQFaqS53zBtL8hnLXdIfXO1vNpQQWf5HvYU+eoa6rFNJu/QSH2YZFW3xFeE6ZypoaFfbWmxzHlS9XPhY+xAPB4d3kggVfaYiee1xj+Tqgb1vVOY/1kk5C7FasHhv35Z6JyYj+JZkAow9qRygSbqelUaTXPKeD36xX4xW9EiFfraz+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/SOUqXqc4IdsI6Op4SZut/nDzHsULEgQUFnNNo97vtp0uXiEffkxxqc/Jhw+MxWm+0bWTRss2SZ7boMQ9kCHfmtp4PKx0pUXc3+PKz8fDVsdU4OTYdMe3CMw98LvuzZj4G3eXrLjNqthYgNYxe7wxTTREZwfW/cdcBYLB37rmkwwFgsHfuuaTB2Gzbvha9BMobvWnk0VbzsRgZsYqWWnjZu6Sd61SUWtDjCgNQSVdmTE+lrgtFc1crdHQ5BG+ZDmZLFsfdigeEoe6zI6+pUlAzAWCwd+65pMKvvciyv21W/bYiDHSwIOawInIRsqE7jQmbQFTYqvlIwTc+2J5/NvU+pkEbAltJTXcLCIxa0aOLzWotQEC/VFa/AWCwd+65pMFwNT4Su+gmAv3T+/Q7PTTnZ0pn6axGRmhYZ/vTCkqXK+3UCQ6/Os9obqH3qqgQ2LeEwJz0lgV1+BsHXHqEjaVfRVKRms1ftdMBYLB37rmkwSmIo5j8yCJGJWbp1N0EuioBxG/arAspjag9o9V03daeMw98LvuzZj4G3eXrLjNqthYgNYxe7wxSruDnuKlgiycBYLB37rmkwwFgsHfuuaTB2Gzbvha9BMobvWnk0VbzspGlNYMKGK5f6AkhmLx3jR9r9NS/2J1eOxB0dI1EaCdwuxinGJGN23y+3qZdYvE57i+CAxW59BpMJj1sdy5O8AQbB1x6hI2lXyRscHKFYmPPjwZx15J6L+Yjn7Uiajytw4wW4eWngNMCuWh8UlluuUmHW9k/xEsA/z1R7kBiKD29YggAh2zYxKhKar2s4P+7ywsIjFrRo4vOlbOdzqU7cM+PBnHXknov5iOftSJqPK3AM23Pn5bqBCP/7r49FSN7PaBkzWVro+7j3MVxRVqxruhy73ZaAmNJsCY9bHcuTvAEGwdceoSNpV5QMhwBBDOJLM2166FXwotZFffRzpT6CYrDl1Bw7HnEHYdb2T/ESwD8cH2ZPWsfkLBxHLifkb0sGtrE4T8eKGtRVVHZWTNJI9IeGrVsTrhltx6Mxajn3SOQP7cmuv6OeJrSCXgofxdjQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Ltx5v2R/2i7QW6cR3ugt84yOSikUR84Jm6vt7lh6NPTEyIl9tcDvIrKwQFMBrptmFt2FocRTvBr2+YkbIMZ8A+du/y3mwoDlqvnujeI7UaGwAyrlX0gor6voinbaxZqbTkV25AI4Ixd6a2bDCOSH9j1GVkb0YUfE/iwbBGOawofcfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsTpLdr3PWTRZ5RRDns/Z1n8PTJVhKvVmpC6f59p0irJJTOxVf6qMnZVa+ffO35r680bOxDv8Hmn1DDYZLKoha/iQAQOxef0k61YdP0BXT70DGQv3X6heHUWyemHUYw8wDnkyOhxNuHYqEwGrWml3M+x6Mxajn3SOQjbPf3JibGS+8K/ovuZ7TN02kadUJHIbAymT6ykczkCWC+J75ggO3xrRGSu5IrBBIdg1suZ9E6/wTJWSiPyNhKrD1oOhUnp8hO7JRb/x7EOB8gtxiLTTHiGvuCZChpPFyUzsVX+qjJ2cFhRLHtr5z2HF34gAZl5q3pCgYVS10eex2DWy5n0Tr/RU5OGMXZ4nysPWg6FSenyE7slFv/HsQ4Y/3FFXKQO95mAmFR3LKaecIKQH9xapKWixdRZESkTMKO5K8dh3pLdaw9aDoVJ6fI6m3ZnKEGKjwoco184hoJLMLg4TLFSlMPyvZhKluyThlNbFwOWiv+X8EfppvqcUz6rR508ZTGndGpcg1sRIlPCWvQikJWPE7COkoH8fk64rbZdQdps8ZOyWKlDeM0NhdLnRpRErudjt6lr9eQQZ3jNxxHLifkb0sGc8rFJQKPIgN1TGReX5j+UI9onXBLEFsaUzMxN3ZVssA24X1LNvxtz1ninZk5BIlNO6CkLF8CmfSXqvcJKNs5fpmrRWrRZOUy7qCe6H9mcHlxX2xf0wa4os3NonL3dWzRF/O8s64DUvK6maR0RWksW21F32Il+s4UpIAH3GDGpAcM23Pn5bqBCAMf5L1RVeMOlM7FV/qoydkji9MrIcEZzzgLIkEoIHZdVFYclhD8d4eZq0Vq0WTlMshkEnLnkXkHGL5BUOX+1xgwICxouRz2wwIuZ8gz9RNAs6riPrEhekRr0IpCVjxOwjbhfUs2/G3P+eN/hBVIbTMnDRel4faEa3CAjfd7xQL2dWTJ1KHwjnoxJT+Am07gFzJS9tMv+/wwoq9ojlmavqCUzsVX+qjJ2SOL0yshwRnPOAsiQSggdl1UVhyWEPx3hwY9SJR7MwFUD1pWD0DZnyXSj47rm8Yq3tgsZshfLtydrD1oOhUnp8hO7JRb/x7EOEKFPp+74f6IE35JoD5HJZdZ36WaPk0oGyXoPohMQjK5rR508ZTGndGpcg1sRIlPCWvQikJWPE7COkoH8fk64rY9D6YhvSdkvKu4Oe4qWCLJQhQaHWyXaE8BYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3hwY9SJR7MwFUD1pWD0DZnyU7XVmVJn3woCBkf8+t9vrDry+gfaMV2Br63I2TU/dOm6CeZ0nsT+2C9Hf01UlyyqrAC8/lj5kKjVrgSNBvfq0OZf11sV/DEVTqlhapxtMHHY6C/Exo+RCSaMSTESCu1grAk8yfFtp1eSgaRNLNiI+VNz3gAPE1y+XnSv/rNmDxCR+lFIzyhXH2NcLAKWIy4N3VmaIohTeKhyUGtg9pP9WQ7GNtU97kTE2caiSB0pwUU4Ke3RH6KbgnPB33uCU9gsmdGlESu52O3qWv15BBneM3HEcuJ+RvSwaFVSD1FKcXtBMFz68YcXSzNGERh5UHqB+laqHQ6HYhZedK/+s2YPEJC4aCMXedht5TMzE3dlWywCvkwtmFLeT2MLHXl0A1q5CUzsVX+qjJ2ToUI3EUh971pyenXn87dN0xJT+Am07gFzJS9tMv+/wwNcLAKWIy4N3VmaIohTeKh8+Vbs8zyvfK7GNtU97kTE2caiSB0pwUU8nghxtgSf/dwsIjFrRo4vMkQjeavmdzPzXCwCliMuDdpWqh0Oh2IWXnSv/rNmDxCa3uRShdZDwvMriQusSU8tU9zQjfrwajONWZoiiFN4qHr1AgXgzKfvVYggAh2zYxKvJMoiRRwIwd7tFfp7RZlEEPWlYPQNmfJakVFNTeICNOlM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCa3uRShdZDwvf666Tkuiwn81wsApYjLg3aVqodDodiFl5v3z4BoloQNZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWXsHhv35Z6JyZ0/zvTlgbGk1nKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTwUZ0OCl52YgxWDHBfoP5+RAuXF+x4SDo3LJBrkcxdC65BAP/YCJG9mUmo93yjcAY2tWZ4ublbysOjshum56CyS+595hQ5cfijMsvaH75WwlZTKAgnBK099N+9hMV9g88T+QyoSnr4KkzBv3q1rE56vP050jzw4zuaPuY0ytJXcx0ipyWLszxhiuQjVJvX3zI27wNWQR10PtUfxXF83AvLrYcc1tb0JdQPbEZ6naIcP7vLq5wEfd55MuhlKJ/OiHPX9jyCjXAW/euhhtPcIagUS5HanjcYjPwvKpMsm2TwyYx8+fSCxlRIMT2P1AbHH2ovouOyzR2lpcrldI+4X6yN4Wxy4iwpZ8+LacqIrCCWniyImF4gLRZAX6l+UWRND8K6QoGFUtdHnuoNfGWRcbK35jo3NMZR7zraAbKeHAIb90YjDI2ctzIMG+gZaWqKFW9ZjySmeLaPsp76s3YnyjNbQ5/Vu3HKKHWv9281ooBjDZhH99VyTSp3ouQMlSkoQRfl5RhnkA+4iOXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZiMvbJ5KuI8YITb9aoC7ldGG79eKMzZ6uVTM/LO5RPzdDn9W7ccoodbftwRVMkVGtJdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmeWqSY/V8J8gDp6JqC8S5aHRsqR31kDb8szHT3smYOULy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8caBAzOFbh3Ctin84MpLvtsmf0g7T8uikTmdjCz+epvdf0N2LXKhc5/X88nixuUVIMk0flCMwg9o1dZ0prWwPdDsynjmpITlE1eYB5ioJUYgkcehumNwmTX9v20Po1mDRqmm1dNs4x8F9qoHINnqNTQT1zWClEYtH4XLjiOTjsUysUJYN6b3gXv9v20Po1mDRqmm1dNs4x8FNeiLyn7WySUvB2RBqE8Qg/VoTfJXkX+sE35JoD5HJZep8akuHxFzA0CGgMvrUkxxN+zZPe2/uq5VW3DiKRkzwjElP4CbTuAXIrFPH/HX6kE0nN0fx0OZ3WS/vNeMNayWL8TLnOCOek4GPUiUezMBVA9aVg9A2Z8lRcLpVFUzJoMvZwDlzKIgxAwrjVQlO79KZcxmz9AAC0ynxG91hzMy4FFj5+cursX8ETuc2nyyzNzmIqollrQmakKFPp+74f6IE35JoD5HJZc16IvKftbJJS8HZEGoTxCDBj1IlHszAVQPWlYPQNmfJdKPjuubxirellYfXr/5N5h6c9O0Bg63Vn5o5KD4eBcYKQm4xyH86zW5YOX7gU6yaC7qGu31ag43ayk2vHGtIuqoNfGWRcbK33mI+vqzK689qZBGwJbSU13CwiMWtGji80lhkicgI27dSMGkaYCErkSC9TX5sAYwGjElP4CbTuAXMlL20y/7/DA7q7UYMY19q9RRVJDpaF2+wsIjFrRo4vMOE64xrnjCO6g18ZZFxsrfZjySmeLaPso9D6YhvSdkvAzbc+fluoEIuABHWkUrJawWljHGiD4epsBYLB37rmkw35uVDSA9htO7v5CueOv1izK4kLrElPLVS1+9WeDzVnTAWCwd+65pMGOekVfcBzwjBsHXHqEjaVfukZUgm5l+T2CljEGCQ2OFD1pWD0DZnyXlS2V743wsV8BYLB37rmkw/1g4hWW9x0mFiA1jF7vDFKu4Oe4qWCLJaFTnpZKiSGfAWCwd+65pMK3uRShdZDwvKhBzSnCQ4Zvne5heOPpqZtRRVJDpaF2+wsIjFrRo4vMNhglDt1esTcBYLB37rmkwQoU+n7vh/ogTfkmgPkcllzXoi8p+1sklcPeNm59NMYEeZa/KEJx66PbAFiPCP9Aa7N/b5JbcqHzAWCwd+65pMN2JTYjsYtAYqDXxlkXGyt+fIwYpG+dc1S2YloElx8fqEPQTFGz2CFt3DCpm/rPLLq0yD9MfwDAwm7Cl/JGm4dRMzOo1oB5ATQsteX/pLtfRUr4s0iddEK3y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPFpbEnY3Ckt1nKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTcN9NVMloxZeweG/flnonJg+cMn9BgdFKao3NSLHGzcOXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZvXFOhOCzn7oG78uzJtzcoQg8QQ46zmxgkWGz5Pqa8LcGnkhHOWLndfkJGrPv+AUqh9TFW4JdLljfY+SK17iu0YpD1cpko4vTY1VxarjbYSyYNTLRsAZTMjC1gLXUG6EtTSc3R/HQ5ndZL+814w1rJYvxMuc4I56TvGED6cYfjdoNrlzvRZ41imTysGfIDZrZ5jY2T67Es+9y5PpLEgYovRg1MtGwBlMyMLWAtdQboS1NJzdH8dDmd1kv7zXjDWslsqXWf7HESECwNSgROhYtQu+6dBkYMzRxIm81zCsbjdDJGt93FLnFxYRO5zafLLM3OYiqiWWtCZqnLeundAyWWpvbEeOIXIN/Bhrvt/y+YAdeDspfEuZJsr344wggLikq54k+1u6yqrnawtzpqCyYSHAWCwd+65pMI2aUZ9CPIbWOVvkfSuBliursF+kKdIWSFMfE/cwJiXawFgsHfuuaTDfm5UNID2G07u/kK546/WLyGQScueReQcnn/eRhT9Sxag18ZZFxsrfOvzm46oTw3GUUHQYVZ+36Pa2WsouxPRPksWx92KB4Sh+DbmFakobSg9aVg9A2Z8lKfaITWj4BHx+UXDQdGONeFrL2xd/GFnka2fhra+8NHrdHQ5BG+ZDmamm1dNs4x8FaFTnpZKiSGfAWCwd+65pMNgyf6f+E6976gFp5T294R0M23Pn5bqBCHqZI07S4q+pD1pWD0DZnyVnQsqeq1f2T6g18ZZFxsrfeYj6+rMrrz2pkEbAltJTXcLCIxa0aOLzvOwD/61naXAYa77f8vmAHYNWBUbEQksWqZezZPkxilXCwiMWtGji85Pju3Rqjz0E/b9tD6NZg0ZWsM3QiHD0pRhrvt/y+YAdeDspfEuZJsr344wggLikqxN+SaA+RyWX5uMv12qGDYjAWCwd+65pMH9If+R9bwqawwx1Y9Kiz4ATfkmgPkcll19YANMVuSkED1pWD0DZnyVFehOJaeEBhMBYLB37rmkwhdPZ5y/hF35RCWbeSOoaDag18ZZFxsrfL34jfyAKTSye3/v8nWoHdABKVBuglOW+XtMm5DtaeryDKkvY++Zbwb6IhgkZZbtUEPQTFGz2CFss0q2Qk0aD5bgSQbjEJG3ML/44EZn9q5SF0bY309F5+5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm7M2Jy2rueEb9v20Po1mDRqmm1dNs4x8F/FIPAS8qijfCwiMWtGji83Y/toYFNVE2cnegbtHMY5APWlYPQNmfJYnhaT+BVij2re5FKF1kPC8yuJC6xJTy1QsX4lP0nDbaPQ+mIb0nZLyruDnuKlgiyfxSDwEvKoo3wsIjFrRo4vM+0pd7O1Y9+UdLiAHUHL0Svt0W25erGITJibuQ934z3OZsPEA18kKxH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8Lw77OF9d4rOWvl9lNkq+IdrX6T0NpFxbWIc83RD0iU+Wvu4K8NlLooedDa8/RTQEBD69i27DxUHP/OYV0R4td6r36mE7lWClZdLuAG7fM0+01lFoJxGMUvmTlFV1SR22TwURxqfShO1MDW6tcf0NOEx1gX59vE719/3qMvpJ11Z9W9EiFfraz+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC/SOUqXqc4IdsI6Op4SZut/nDzHsULEgQUFnNNo97vtp0uXiEffkxxqc/Jhw+MxWm4J4GU2KWCH2o7IgfUbYao66E0Ypsh6pbTKbtlqu6/gxhqfiesrmPWgl9BK0MsVDTVY1tXzOO1m70Wn0KhqZOKmwUBTkL2d8olY1tXzOO1m763z+s8h6wpuOgvxMaPkQkgpwh1Sk8uYlrnrDy9x642jW/oELsAX0EgFcsWN4jUhLwFfzu/pgaLrRdlEeUweax6Prf0CC1QVulmAsj5iny4sIGh6GIRYdrTCX/pV9xny3q+9yLK/bVb8fum945sPLeWnflm2GWPztaDHA85r5sJm5fcLCHADv2jAgLGi5HPbDIIvT+UNORMQ73kiJl9dwNPl0uiV+r/FjwR+mm+pxTPoBq8OYNNE4kUj57B3LdGdrhoQvMVl4vr5AdXnF4vjGJyQgN42ztupWMCAsaLkc9sMgi9P5Q05ExD2xGep2iHD+sie8IHhclNMBYNAncoGkg5+gA4ucyggfrYuJOWYBPJUwICxouRz2wwIuZ8gz9RNAHChBkRHlDB5r0IpCVjxOwh2DWy5n0Tr/4VQLknJoeu9eCQMHKUbNsNWZoiiFN4qHr1AgXgzKfvVYggAh2zYxKrOm4GNjZXJtSPZCjBZnXw1CFBodbJdoTwFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHihqTq5TohFcb6fWz5DNEYJTOxVf6qMnZwWFEse2vnPYBjsOiGyB4sluyWR/fbfv31eHKnnBEGeeUgj9hxhl6454k+1u6yqrnYm7S8NbLioiUzsVX+qjJ2SOL0yshwRnPTkGSJu/s69jC4OEyxUpTD4eiwO9xP+5his56PQm0umWY3JjE6+3cOPWqEdoGn7o3cCu8ryHrFY7tIsPYmpLgc5hcRIPQMbYrIGR/z632+sOlaqHQ6HYhZf8TfVvBgTEMBsHXHqEjaVeAmefhmnKSoPSJ52KAGWjkniv+1iNSrX8PWlYPQNmfJajntpcAlJr+a9CKQlY8TsI6Sgfx+TritsLCIxa0aOLznZsRGrnGEqzKjsB1J/ogsduvDz/TZisvjtjuLVBB+XpzUsA4WQFmBliCACHbNjEqEbixuPsCC6vwcJ2XJkwGgK2ng8rHSlRdV0pGt5hZIZ3/EnNF8wz1b6Ic/j4NtRsPsNMwfWlh5XL4yL8WosqVv/R39NVJcsqqQVlWo4auvX0F7pVL7p7RG+7RX6e0WZRBD1pWD0DZnyXSj47rm8Yq3g1jOungVNZtwgpAf3FqkpYUiOnUM637JzEugNrPMCslBsHXHqEjaVcNYzrp4FTWbcIKQH9xapKWFIjp1DOt+ycxLoDazzArJQbB1x6hI2lXhauMtfc3NEsBYNAncoGkg5LFaicXcUrcupmkdEVpLFttRd9iJfrOFJ3Gi6xSlJuHE35JoD5HJZeti4k5ZgE8lVM2bu+WFHT1NobcwiHYDNXC4OEyxUpTD+dK/+s2YPEJre5FKF1kPC8yuJC6xJTy1T3NCN+vBqM41ZmiKIU3ioevUCBeDMp+9ViCACHbNjEq8kyiJFHAjB3u0V+ntFmUQQ9aVg9A2Z8lqRUU1N4gI06UzsVX+qjJ2SOL0yshwRnPTkGSJu/s69jC4OEyxUpTD+dK/+s2YPEJvyBp6CCyHuYp9ohNaPgEfL++fVVIhOx6tACV4q1xv5bsY21T3uRMTfrzcrVPrhZXcrpLydPnYbDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJM59gn+sJA2JpfxAzn1X6OquP9Sg89xHJKnaWEOBQNVw+kKBhVLXR57WcqT4xF2Vxjy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJP7FnK3UwEB9DKZPrKRzOQJo2DDkVTO+A0/G8MS9PnKJGOJKd5hF3+U9Hf01UlyyqpiHW7aO5vxU6/78KYYJzZNaDHA85r5sJlgPHSgvyImSlqk89/pi6AIv9281ooBjDYfILcYi00x4h991K5Rjd5QAgRr7UzjYUyoNfGWRcbK3xxd+IAGZeat6QoGFUtdHnuoNfGWRcbK3/RcTsJJ8QYw5o94szA1qLuzxO7EBtu+KPzk0seZwX46GUMQ26CV9ZyoNfGWRcbK39zHLiU0HIspy041qprKfGy/3bzWigGMNsT2P1AbHH2oU8ChHu9j2s8i+PxZxyAsv2Y8kpni2j7KnUyy6YcmI8RLTpAqdXgC+VTszs8iePtfihqTq5TohFfIgh23HomE7LUffbA2vmQPM1z5OLuut1z307+4oPX6k0IjtZoAq7t0lKbPj9+iHGmZq0Vq0WTlMu6gnuh/ZnB51GL2IZWXr8qb0dcNAokWN57JkW377qQRpIAH3GDGpAcM23Pn5bqBCI37iPb5nUVizc2icvd1bNG4+HOgwKwt7hN+SaA+RyWXu0a1A3VjyGWzxO7EBtu+KA9aVg9A2Z8lKfaITWj4BHwjiSU2rxMiSp0aURK7nY7eFgXYlvHGlvAGwdceoSNpV5pBVhazntdDqDXxlkXGyt/i4XgOVDPh/08MDQF/7jEYzasixnaPUTJ8gPwsN5c8KkKFPp+74f6IE35JoD5HJZdOfHBU1oPAvq3uRShdZDwv/WczRISouxnASdLvMqoB3bFCWDem94F7/b9tD6NZg0apptXTbOMfBXTF9b0wdUvcMSU/gJtO4BcyUvbTL/v8MOQQRns8txCxg1YFRsRCSxYxJT+Am07gFxB+VaJBV3EILaEkrSAVqcATfkmgPkcll1By0nrdhs43sUJYN6b3gXv9v20Po1mDRpWStaC/+Ito9BYedILm4ZUGwdceoSNpV/BdPgDYCdLDBj1IlHszAVQPWlYPQNmfJR06TI+L8vmjre5FKF1kPC9/rrpOS6LCf41HDMcBDxHL8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWX6iOMcDwrlMsu1h6RFkM0nWYKlakzehx7DCWlZXCPhBuIwpTVG4MzpPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4Jaxpvx4A1xBXqnXN5VA5KvKHmUxyDxBDjrObGCRYbPk+prwtwaeSEc5Yud1+Qkas+/4BSqH1MVbgl0uWN9j5IrXuK7RikPVymSji9NjVXFquNthLKX5Um0P+6/oBN+SaA+RyWXRy2f5UTOYcu7cHGcmccaLbdTi1x3mcIYkNEPMoCb13q3hSg4mUlTlRB+VaJBV3EINJzdH8dDmd05IdXVmodgmVEJZt5I6hoNtAtvATa+nmlg1MtGwBlMyA9aVg9A2Z8ltV3JxQSIfM27cHGcmccaLau89FjbHlF3E9c1gpRGLR+OL9z0IaBXzGWVgzT9cOAbE35JoD5HJZcoviA8nPFl62Q6arWa36ObaLqzJmflsPSXt14nAyWWX0NaRZr5dtq7lcwbKRQEQlkpCbjHIfzrNblg5fuBTrJoF6r655uKHEetMTEG9QTu3hV5mShiH+JTBt0iTwmsIN4ctas+oPi1vKaMgaeoROMWwsIjFrRo4vMkQjeavmdzPwpjzpCsXKdk4SSlnUTC2QgbeHu3NebJjwbB1x6hI2lXNy3i5SNAjHOeuCv8EL5+zm7oSYKhGe9x/WczRISouxnHRIkZMDEnfTF9B9IdWyuoFFPMs7ICBMITfkmgPkcll9M9uxQ07dhRV5gHmKglRiDAWCwd+65pMEmuIp1ug90YMlL20y/7/DAKBKI3H/vNGQh60+nnb8N/TTG0uAJhe/PYrqEx1I9NHOxn4cPZRGabE35JoD5HJZdHLZ/lRM5hy7twcZyZxxott1OLXHeZwhiQ0Q8ygJvXepvhQT+f1furGGu+3/L5gB3tqB/XZXJTgTJS9tMv+/wwRLlur4NsaI/9ZzNEhKi7GTq/b+Rd+GciqDXxlkXGyt9qORwzQdMkxZDRDzKAm9d6YWaM3bdub3Dj5RcgwgjQhReq+uebihxHrTExBvUE7t4G3SJPCawg3py20QfQAbjT3PPK93m2DfNs1MLIczSl/G/nZ8vIefdvSc+YnhH5GrR/W1GecHngSTElP4CbTuAX8zRofA2lBo4pCbjHIfzrNblg5fuBTrJo/xN9W8GBMQwGwdceoSNpV+B39dwXU/8+IzTVVgkBqzgGwdceoSNpV7RpfTwkqql3tNd3+Ny1F6xu6EmCoRnvcTK4kLrElPLV4vTbZ33JAvhllYM0/XDgGxN+SaA+RyWXNSspm+Ofd8jPv/1si5pHVhN+SaA+RyWX5qiLi71Bj9fwCST4xkKSPFUgETDDv25WBsHXHqEjaVeYG1py1sf2zsxBPmd3IyJnvyBp6CCyHuZOVCkWvMetfj77vTzzbraPwsIjFrRo4vMCWoIflgdmdeYiqiWWtCZqZZWDNP1w4BsTfkmgPkcllyi+IDyc8WXrBrunOcy3DdEYa77f8vmAHWFmjN23bm9wqDXxlkXGyt+tMg/TH8AwMIM+aEC2mLhmax7M6tZYeK72iuplgCAem3v/O9MAL9tNrxaqwvYfP/v/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyPXyMGM0AOBwsIjFrRo4vMcFYaXr9ZqJSxNqNqoDz23VMz8s7lE/N1xYL5f0eHOqK8WqsL2Hz/7FpRWcIMbKOeSxbH3YoHhKEGj0wPc42WeVnPSnmzzGo7q3YFFR2s4AFQEo83cZQQWl/ux5LaKvyLSu5NX3VJkLh+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC4kq3srN7+p8SDYYEZZ2nr5tri1hIYa7vqDpZWXNzWXSk5Ok5wGBoKhccAKiMeC1ZbF3uU2H/DCyQO8ZxWsk4lK1bfk3tLW1g39e2VsGp8X0lWEJ6KfY0nLzFn1/kYFYVi0bluF31BjZe+ToSZEujRSpP+Wem6+qbcSdxR8LiiPb2bSy/ssm1qcfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu84Qta0VhokDGQv3X6heHUAAcouGPgvdGNanhf98S2FY2x2rG/JzSm++E74jtv3CjXqdpuCbaDKLCOjqeEmbrfNg0ZOIlCNdkv94TlSlGhCUZ6CCfYNpaWND5/1YD7AQ8v94TlSlGhCWL0YIzvLQ8VIqrp3xKIxtDtG1k0bLNkme26DEPZAh35raeDysdKVF2XLoi95JK1wOxJbku+DGjGivPvFHm9msvQrJURgKNO+4TkHZ7hGiLDNnr+NhM2pvBNz7Ynn829T+smzz5674GmmoaPu15mwu8InBhgiINIJDawSr20lhs4emyoaVsNeoEpU+dCaUOiGQZpjazlsgCdraeDysdKVF28KYGKV1qjLsndCD0/RgZs0trTxM/mtAyylsmzXHZzx14Y7+Cn7apJTKW8qsIVrLzYvZ7+qnnvuk+NDMtblj/lwTQuk7lnHyznSv/rNmDxCcii33v/fBqayAM8T53RmMqN6/v2LlbCwvMWfX+RgVhWt/F5lUyR5ghBboDWT8dzI+quOeptdosl8C/MhI5SRFL30a9louFgO14Y7+Cn7apJTKW8qsIVrLzYvZ7+qnnvuk+NDMtblj/lwTQuk7lnHyznSv/rNmDxCcii33v/fBqaRXlV6pv9awckQU3a48Xf2gfiENe0Oug94v/KUh2YV6UBXLFjeI1ISzLnujwNCgzYWj7bkWA5uvmK8+8Ueb2ay9CslRGAo077hOQdnuEaIsOG1pw07ptE9w7DB042Xl1j+iKdtrFmptP/Pwx6skM0Pw/tya6/o54mtIJeCh/F2NAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu3Hm/ZH/aLtBbpxHe6C3zjI5KKRRHzgmbq+3uWHo09MTIiX21wO8isrBAUwGum2YW3YWhxFO8Gvb5iRsgxnwD527/LebCgOWq+e6N4jtRobADKuVfSCivq8dauuWrPHf/87xs4Igtz+ft/5Fw87SHagCvMDmp2o5MfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvGsVqECQ9P1fMK16swBak6aDrV0SaupysaHlTmKsmfKgFg0CdygaSDdwS7MS5Y9KzSgIrk3Duj8Y+YStKhYVkrvWyKpZe+sEzXqdpuCbaDKLCOjqeEmbrfNg0ZOIlCNdkv94TlSlGhCUZ6CCfYNpaWND5/1YD7AQ8v94TlSlGhCXjazt+6rrfB+Ko8VlHmIOiCeBlNilgh9jJakekrNK1qQkb41xZ0+zJ532mKjRs8AuQ9zsKk8AIidXQoFv1vZWCiB9WB76XcZLBQFOQvZ3yiVjW1fM47WbuugXT7eLWvflucMDlUgErFND5/1YD7AQ8v94TlSlGhCTvxtcK6gyzu/z8MerJDND8jbPf3JibGS+8K/ovuZ7TN02kadUJHIbDBNXEhzns0vNJCZTW10xy+0kpBS5r4LY4+/8gGLek9mi+nta1340811ph9EJwygYqU74E+WNz6eX+OoqL6yzGhylkAVKjW7xxPVhhC7z2gtK3NoBUN/erA20ZgPF2W9Z4aKd3IU1VzAeAXWmedi1yI07ZvP/PYbvGmXHkMIxSa1yH/Az7EINaU+Mi/FqLKlb/1rkCRBNBMQOviItnNbTHvWHkTSCSmiZNgPHSgvyImSmYCYVHcspp5wgpAf3FqkpabnAjLtURuje0g+Lz8kbCgXgkDBylGzbClaqHQ6HYhZRzIjmkRPghqXMZyHBq//8zBXmRQxKUEuD8BqKRjeRUO6mycOFNXsoMwICxouRz2wyCL0/lDTkTElXeHI7I2QVtAUjqf8aFBxclQhwwd/5HsKYpuXYGa4XRr0IpCVjxOwh2DWy5n0Tr/0BiPpbsi2bpyfFt1tmECVqqQD3q+pGjRHEcuJ+RvSwZzysUlAo8iA0kAGDAq7+VAcuTCtH6/xJL49dKirrGTNojEpQP5hfCVjtQiGLJgL5txztYHphKvOCCL0/lDTkTEpwtxCu/hW/zG13tPUhWWZEwiL+7bR3NuEWsoLROZ2jlYggAh2zYxKrOm4GNjZXJt/id2tyC4EWzuoTejPGnBubkOsWPaq9s5KJnyGPmNyWbhwyaAxLfQPWpGPxRfAM1oJuXBVwKnjiL/E31bwYExDJvR1w0CiRY3j7GeEBde/DuUzsVX+qjJ2SOL0yshwRnPTkGSJu/s69jC4OEyxUpTD+0hvUBC+7PRO+8giOLw1uEtYAA5kqse/gbB1x6hI2lXvXolK5pzHUZeCQMHKUbNsKVqodDodiFlLWAAOZKrHv4GwdceoSNpV1KUnG7T12N59KM91k9syYucOmNUNiQp+QWYHEHuOOgu7GNtU97kTE2foAOLnMoIHw9aVg9A2Z8lqRUU1N4gI0460qRV9sVQrNuvDz/TZisvlRgTnlgd4ig44KuW0tEdOuzfWsfwbxlzfkxUkNGCvYBpmUPUVMhtGandfhFa3l8R5I4IXBo4g2Eo36jxjcHPC1HKay3IZ/ge5j/WSTkLsVqaMs1s/8Z3eBuofeqqBDYtRytZtfKGYoI2sEq9tJYbOM55pewN4e8yXiu5UQV8FEMIeHeJyIgr0xNdnFsInRFoVMz8s7lE/N2Bxl0y+KwUu21F32Il+s4U2vT/xxzABuHuxsvB00awOFM2bu+WFHT1/jJ9evvwc5rC4OEyxUpTD+dK/+s2YPEJvyBp6CCyHuaORbBg3WAZBPSjPdZPbMmLnDpjVDYkKfkFmBxB7jjoLuxjbVPe5ExNnGokgdKcFFNa4DKPbOmTfau4Oe4qWCLJDWSX1+HDlqTbrw8/02YrL5UYE55YHeIoOOCrltLRHTptRd9iJfrOFG+wihoEHfiJ/RR3NYigAxyym6TZ+4ZAL8TFM0iKu1quNKw7lJGkWWWVGBOeWB3iKJjiCQ0HNKypVFYclhD8d4dBboDWT8dzI9AYj6W7Itm61Rax6caHSJl7td2RznPfJAfI63n40WDTUIhTjrAFHFrOG+f7BdZNEcLg4TLFSlMP50r/6zZg8QnAlCJBb+ant6tKDDDIltpJ+QTvuMLqRE6dGlESu52O3o3MCALtK1/SUIhTjrAFHFoOmvV3gZiMhVRWHJYQ/HeHQW6A1k/HcyPygFi2Xk65vUaC32k5ERpLjiFu246anN2Ns4NBVtFnV0HjZbYbHfxHwuDhMsVKUw/nSv/rNmDxCQtR5JnFhgjIy4kEYPmGHzuG25WMDLJL+htoVsRktZ6NRWQfiSrBvSvhwyaAxLfQPRSI6dQzrfsnS5IF/DrN16sowpG0bJjuO4CXl3h8nhtKhGkiShnkr5Kb9BwLc9xme2vQikJWPE7CK+TC2YUt5PZKxi/QrsF3O551Frg5x1/ccOmUg5H4/5ScOmNUNiQp+QWYHEHuOOgu7GNtU97kTE2caiSB0pwUUx5PreZaz39V/2Pl6xLAifC4Wm46Tw3L+Z4r/tYjUq1/hNtI11oVuVFYggAh2zYxKvJMoiRRwIwdBnT/fzTooEvlOobQYJQDia1lRQ3GGOeS0jW4IEq9ry1vev70hjoafxxHLifkb0sGhVUg9RSnF7QB/atx6Gb2s+8/aVQzBSScO22mXiN3cm3brw8/02YrL5UYE55YHeIoOOCrltLRHTptRd9iJfrOFNVVQjB0a0gQAqp7yWmw8cCu2GeVxrSCsLeAcpCiywfCUIhTjrAFHFow0mP3skyStFRWHJYQ/HeHQW6A1k/HcyN8ZPiNFLrDyxKBBq97ivdIjiFu246anN2Ns4NBVtFnV0HjZbYbHfxHwuDhMsVKUw8r5MLZhS3k9rc/abVWqH62QeUPnyAo29Fw6ZSDkfj/lJw6Y1Q2JCn5BZgcQe446C7sY21T3uRMTZxqJIHSnBRTc23KWnbOQ/RKYgmd853BOrhabjpPDcv5niv+1iNSrX+E20jXWhW5UViCACHbNjEq8kyiJFHAjB18cOoLIX1tFNO7wRUiU/9VrWVFDcYY55LSNbggSr2vLW96/vSGOhp/HEcuJ+RvSwaFVSD1FKcXtLVuaovWGxGbBvuRh4ZTJ6w7baZeI3dybduvDz/TZisvlRgTnlgd4ig44KuW0tEdOm1F32Il+s4UC8g1E4M0/TawLJfHz6qRkWTWU1Lsp7f7t4BykKLLB8JQiFOOsAUcWjDSY/eyTJK0VFYclhD8d4dBboDWT8dzIwzdOH/XAMU1YYHQ2XVJnVKOIW7bjpqc3Y2zg0FW0WdXQeNlthsd/EfC4OEyxUpTD+dK/+s2YPEJl8FmqpKYCRGw5GxFcqdKGCt9JQ0lrBJ7G2hWxGS1no1FZB+JKsG9K+HDJoDEt9A9FIjp1DOt+ycA2kfmSyZvGq7uyUnV3Pl9SvNQx6fDevGEaSJKGeSvkpv0HAtz3GZ7a9CKQlY8TsIr5MLZhS3k9klEdxqOirYno3R/tSRh50vQSVDkiTbSp5w6Y1Q2JCn5BZgcQe446C7sY21T3uRMTZxqJIHSnBRTY1cNecz3//czqUP2CcH12Mct/N01i7ZXw6Dttv2iywdQiFOOsAUcWjDSY/eyTJK0VFYclhD8d4dBboDWT8dzIyKg+vl56cpkBZ/YVsPsMWHQSVDkiTbSp5w6Y1Q2JCn5BZgcQe446C7sY21T3uRMTZxqJIHSnBRTY1cNecz3//caQyfpAiC+3cct/N01i7ZXw6Dttv2iywdQiFOOsAUcWjDSY/eyTJK0VFYclhD8d4dBboDWT8dzI66d/k78+swjUiOA+a1tHuUrfSUNJawSextoVsRktZ6NRWQfiSrBvSvhwyaAxLfQPRSI6dQzrfsnRpVc1B/in/QMMAxMLFAlw9BJUOSJNtKnnDpjVDYkKfkFmBxB7jjoLuxjbVPe5ExNnGokgdKcFFMFTZEF+DDDKZjB68ztlxeS0kIcb1K/xltBN5++Ce9cppw6Y1Q2JCn5BZgcQe446C7sY21T3uRMTZxqJIHSnBRTBU2RBfgwwymYwevM7ZcXkgwwDEwsUCXDQTefvgnvXKacOmNUNiQp+QWYHEHuOOgu7GNtU97kTE2caiSB0pwUU6+nmUhytjyqm5s8z1DwV71AQ31CyYTADtI1uCBKva8tb3r+9IY6Gn8cRy4n5G9LBoVVIPUUpxe0pWGb78OwoqKcbndff9XWWwhH02k8SOOhw6Dttv2iywdQiFOOsAUcWjDSY/eyTJK0VFYclhD8d4dBboDWT8dzIwwdk2R1rKY9f65pTgrPqZExk8wvrRXYtexjbVPe5ExNnGokgdKcFFMEqBWW0JLx7oB2QMhvPCeJNWYnM+lVTIQovhtOCX0ZQCsE6EgXdjLiivPvFHm9msvQrJURgKNO+4TkHZ7hGiLDNnr+NhM2pvBNz7Ynn829T7VRbMaU9R3EbPAzUDuqMnQXWgy0b6ZB3ZELeDiO4EYROvCthHYYtLAeZszbmnxUrk65bNWSRgdXfBIDRqGKAPqogwm4UoeHsqExlKxSUW3tOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2R+JOhZGjs2qfBzt+PhrTzkgFxsc7HdT9fL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk6xambyK5ZxNCQ3bmdTTHwSU9XczSMtPKOojpHBDUBIMjpys13y/ZAh40l1lb1OXtEisFUyYgp+4QZMeFQwgW5KeuCv8EL5+znckWoY56cgvX/VuTF7etTcRfx/sKVZT8+6gnuh/ZnB5q0SLj91Ue6/VmaIohTeKhzh9A8064LSKe1TYiCbn8biUzsVX+qjJ2SOL0yshwRnPQnjH9mQ9QSGuH3+zHgnhl/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4Ull/LbH3nTl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGazHE0TLcm3h76KBVUhxEgorTExBvUE7t4dUmLyHTtKMnAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTR2QLyaRZrsOvFqrC9h8/+zaMWyOJnvaYpmRSLqrDyOGA61zq5LyRKADNFTHDXYzPUaXl6z3PdmQf2/k5reashCyJl+6w7q+Bi0kWLnusckK6maR0RWksW3+YnvcDjB1JE0b2mIA/m0PJKftaojQLOUr6PyH2nimcDQUFJSyD4MVNhDOo5YPnV/ML3EO/WvzNjhwIGUocy7GoNfGWRcbK35cRiFXk5lH5hrfWX7h0FwtQiFOOsAUcWrhLmDiLqTUvGGu+3/L5gB0MvHoJrtpKj4RpIkoZ5K+Sy4k/HDus2etxCvea/bRFrMBYLB37rmkwvyBp6CCyHubTK/m8BpEC8yVvJ6a0QeUXzzxKVqaHvijAWCwd+65pMKl8+09yWfa4wFgsHfuuaTDCwiMWtGji85PeydIoIHrQNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpOAEpUG6CU5b5rHszq1lh4rr2rBUoGQrMwopCZHa9+O/FyjaZc3+cyiyoQc0pwkOGbfvOR2XnFrlVs/P9zr8kn/SVfbovfMR6DCZrVxtmjyhkETOWt0KBunJJ3ezUKUQNvZs35wr6U5PW4XQ4ypfxM+3BFUL5mbOGYcQr3mv20RaxC9k6h5Y71X+SbmEZbeoxyvTkbkiw8QdgyBX2aIP47pXEK95r9tEWs7Gfhw9lEZpsTfkmgPkcll1G5mylj9mW/D1pWD0DZnyWZqkZGIEsWzsBYLB37rmkwwsIjFrRo4vNXKYJnDCCQGeSbmEZbeoxymRrgjnwrJbqX5Um0P+6/oDb9QuSHDNdevasFSgZCszC+cTnAo1owFGIKO/++klhwBZ1hnzatIOdtIjyaD7uHRlnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTQxLD92or0ceXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZt6/+445Yo4p+CDoKHjQUubML8H3LkfDQVnKk+MRdlcY8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTmDQ7hHxSyV568NVAsXZ40TaMWyOJnvaYpmRSLqrDyOGA61zq5LyRKADNFTHDXYzP5v3z4BoloQOwb5BE4LPl1hp5IRzli53XmFInidWHoGXYrqEx1I9NHDfqZVk0CUssUIH2xnbSDJLx6uW325OK0mz8/3OvySf9JV9ui98xHoMJmtXG2aPKGZDRDzKAm9d6wJQiQW/mp7cQasdgistmEzSc3R/HQ5ndOSHV1ZqHYJlRCWbeSOoaDbQLbwE2vp5pYVxXqkpAiBgFSl7jwbxSJ70/byzNr6MK9qoHINnqNTQT1zWClEYtH4XLjiOTjsUy9xovJ2mxAzRLvnX2Duhfj3UWKJQ6R9GzprfkM6pnQKu/EUKWXiWm56g18ZZFxsrfJtNkV8Glhre2OivC5aHEE0zDBcOZL/WDkqBrVh6zEKA9Aaus/LRVh1fQsuy7XWp2/RR3NYigAxy0rCGMeKg5mXOj+a8t9l483KjZPqsRiGA2n6KkkWCc7x/s+IeSLTJoFQRTQg1Qz1AXgCM814Ju2TGc3nODWG+mK7icYRi0cpDoHBUH6cekqNzUcTNyiZjljMLLxsQny9wjuQen7Od6z0NS5kH2JRrhMNJj97JMkrTKPwX8ZGi/bT8BqKRjeRUOsjXH8JsuUqE36mVZNAlLLLxiooMp8WxayLp3vGdAsWuPkgBJUwhBsgp37lscs67v04RImX88lRYweLABNsP4qENS5kH2JRrhMNJj97JMkrTKPwX8ZGi/bT8BqKRjeRUOS8m86eC3M/O9qwVKBkKzML5xOcCjWjAUYgo7/76SWHAP2cqmlErUmhL35b5RcOz5cCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJOTm0c0jNHELPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxH5yPtMKXTpSoOzonD0/SHt5dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm4Fel1NOPPfyKjlw6QYeYkZbawVdxIXDxoWFgEdetSo1OgFKyacnuL9JH4RiFSfrKeCwfEp2J5FinGTQoBpT15m4JQmX6vUqjr52FJW9ZFldXmAeYqCVGIETe3KALTTmk1G10OVJSLFb6BlnsWKpjH3yA/Cw3lzwq6SQqlZ/JIaryRVqfq4eIAY2zg0FW0WdXgAj7l/iVZXWoNfGWRcbK31CTkalDCbMy44uvLco0E0BNTDL00vCUkAv5vYgaZr/dPUVcsgFwY5tghCbCqX0xiVIXgI7OMDNM+EHZ2JSAnxZy+5nx1JzUfCqV5UkVMW+VWuHzQuAYPLwER7mZEvaajbOm4GNjZXJtUheAjs4wM0z1VzFZ6LgbWnL7mfHUnNR8KpXlSRUxb5XzcKm9J13JTwRHuZkS9pqNs6bgY2Nlcm1SF4COzjAzTNQH/61hfQNtcvuZ8dSc1HwwX8+RloSREzU/ySJhxWxQOpohsAwkhiKoNfGWRcbK39Ft5GvSMzX5t5XV1u1e6Svkz8hwVK7P7xN+SaA+RyWXxSbvrIeNnsjXEzoiAC0FgCv3EGN2Uc6YfmCwuaSzqdcCGEfdpdFYcWExJ0bC9VdMA3vtrwnv1wHH+5AvWAbiH6g18ZZFxsrf0W3ka9IzNfkaWbG2uetPTim5jLl4xkZQ/RR3NYigAxwGyVNHKesLncf7kC9YBuIf4+UXIMII0IVSF4COzjAzTDYp/b1hEdqBcvuZ8dSc1HwwX8+RloSRE9Mr+bwGkQLzOpohsAwkhiLAWCwd+65pMHxk+I0UusPL5Tvoo04A5/RADntIZNywiSoQc0pwkOGbVGWVBfeXYOezpuBjY2VybVIXgI7OMDNMuov6qqwCFlFy+5nx1JzUfCqV5UkVMW+V83CpvSddyU8ER7mZEvaajUC8OIornqDi37jP9zzxZSCR0dku4b/Z9wOSjMOQAQEYAIb4/DEp4BOgh2qck/cJTwCG+PwxKeATOzlk7+mTce++rgCQwqT6QaoR01lDfqdjQIEwp/DfklXygFi2Xk65vQMZVBQu5Ab3qDXxlkXGyt8e8sS6TROxebeV1dbtXukrUZNLB5L+NNVR74NcCBMrWb8VSTBiNrBxDsAxsh0cWyCQ0Q8ygJvXeqiGe7owBpmNM9vQHkvRFKCr0acoB63Nn7i8Y/80DGthQLw4iiueoOLfuM/3PPFlIPWXugkUq3sOA5KMw5ABARgCqnvJabDxwPRD73Gd61Q3Aqp7yWmw8cA7OWTv6ZNx776uAJDCpPpBsCyXx8+qkZFAgTCn8N+SVXxk+I0UusPLAxlUFC7kBveoNfGWRcbK32e7aJbN79NjJpYVH2VbcbqiKbH5TiQCO/pXm+r6LNZIGrWZydbEiIOIBKbPEuhB8Rhrvt/y+YAdl8FmqpKYCRGxDtvPCXxPoRq1mcnWxIiDG7b5A3vRSJ/ER8brwJGbki597ReeT1g+wFgsHfuuaTCJ0PtkjsScopbjLYnwuhkJDN04f9cAxTUJIBrjfifl2bAsl8fPqpGRmPp/TLnx3D8Ya77f8vmAHVPE/sgT7J/p7iKtejvHhOU09co58RJEr+4irXo7x4TlkNEPMoCb13qK68E6rjNXlPLbKD1YJhvOh7mVcKMrAwzy2yg9WCYbzspi11qMuj9pX4CHGxF1gxOJ0PtkjsScopbjLYnwuhkJidD7ZI7EnKJC/cFnQv6kmxhrvt/y+YAdjKtE+AXxtGL0SG7yS6s6OyCcTrsttXGEeZ3kOXwHn8Lijvf0oUVql4nQ+2SOxJyiSre7TODSvTC8Q1K0g7GUgsPoaoWnBFreoxbIYYYZI5dTxP7IE+yf6e4irXo7x4TlG0valbzf4elPywZPUINYcHlVD42AbwkBvENStIOxlIIUSeGdgMd4fohD5dBIbxNZeMMHzF9kVHvqgopDLxrXy4hD5dBIbxNZ2rsyQafNQLeQ0Q8ygJvXelmSE0u/6TxyAQnACWcsxlFIfnKTZ32I/R5W4ZkIX3aDuPf+jsa7B00lfLMwmuiGvFoCDaeA0Ze2AEpUG6CU5b4S7mzIwwp3t72rBUoGQrMwvnE5wKNaMBRiCjv/vpJYcAWdYZ82rSDnP54Yox7mb40tanye4MTGmfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln5Ojh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2TrXNW+ggo9Ojqwd0RDmC6Z/vIBUSmMmCPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxAIGDl8WsiCr+HlE24QQ/EaFhYBHXrUqNZ2rqr7iK/sxqUKiyjuoZThuYozLwMEAyqNXzXd6GrG0sn5O2x1G1nt4SNc73+P83QTefvgnvXKZz0+sjVL57EuHDJoDEt9A9G5ijMvAwQDKo1fNd3oasbSyfk7bHUbWez4F3rcbGH0VBN5++Ce9cpnPT6yNUvnsS4cMmgMS30D0npv7XU6I3MQAaS5MeA3kgHyC3GItNMeLGLXITHOJplHEK95r9tEWss0RnazzlZwFMNkpqivOHwvaqByDZ6jU0w5PI0uBw12RAhoDL61JMcar8T3pkicx+qDXxlkXGyt9XAcLtp0uZbZXZg+ub6CpKQIaAy+tSTHHkQK/WNyYU+xpjN+NMLr6R6NLvPlfAjkYiEFgcKS80jJCGwyPdZ4tcu3BxnJnHGi23U4tcd5nCGJDRDzKAm9d6LsT1DdvvEkIfrh1j7P7yEkCGgMvrUkxxN+zZPe2/uq5ourMmZ+Ww9Je3XicDJZZfQ1pFmvl22ruVzBspFARCWZacAGSF9jAb2K6hMdSPTRwiTSnRezj4j7vlGl4H81DacvuZ8dSc1Hwx0pzH+p88U8PoaoWnBFreHcAc9YZ5tawnvS/Z5hBNum2EID8oFSgFds0VMhNr6nty+5nx1JzUfDHSnMf6nzxTw+hqhacEWt4eItKDf9WQQSe9L9nmEE26jI8rTYbbMrLxA8zvcGctU5tCl+2cZzGX4QtF+AwRQjxdkINk58cbd2HOYKhs6z/8WuHzQuAYPLweKcJItM3sIfnPPzGgVQWsz9u1oAOJUf3sD+/eSZpfzEw2SmqK84fC36hCCnKzlPLAWCwd+65pMFcBwu2nS5ltFzV5r4XGGSmI9xhdTL1o/K6d/k78+swjVeuzTB9VsNpJnytpMzu7YsbByddibIgds6bgY2Nlcm3HVbaI9yUfqqiElkWPOTuY6SuWUm1yrhymjxIrfCv56AgqreyUP7sxIhBYHCkvNIyQhsMj3WeLXG15chBRdA8sfqQKOTtxEvXX0r37z3x1n1CIU46wBRxa2e/hUrgjH2aQ0Q8ygJvXei7E9Q3b7xJCIdvHuI01VL4DCX4eEODRaFcBwu2nS5ltp+sz7olPhbVvev70hjoaf2HO5FuHl9qGgz5oQLaYuGZrHszq1lh4rvaK6mWAIB6bRxpcJCe/G10OtJxI+62IgXAjKOUl6ter8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTRlvRND2F/BQMHZNkdaymPUdN/wHf7/99wJQiQW/mp7erSgwwyJbaSYbd/hhOo6IVvGKigynxbFrcqNk+qxGIYIPnDTuEvw4ztlnOaLA8gPOtr1oAQUPw4NsqKEd60d2xCxfiU/ScNtoMHZNkdaymPUmpY1EOJIl0HNYQoPY+k1escQE1hVaQ5/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxVBRdCi75HEeRC8GLgq8kmnEbw+JV8LJzvB90DR3bIdNIBIIea8EweJdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44ZxmAS5nS1UYf8Rb1SAIMdbJuGg3G/JDxBbWwagjrIeiun15e0i0T/oG7qtxQ9HiOYFLuaZr2+J8tcosRcaZ+A7Ms+TfsxQgIklwqa6oy30WRYxafV9lbSLkie14PRYIbJCSHncx7ZFvizdYOIDpsmIDv/hoiL8D6lHOMZaJukqSckHL8ElX1S2IiXxpZJSDjlAnCoMDdDSaWK64ugDXg6fOP62ng8rHSlRdox17k4FgIwB4A9eqSnfw53ARTTIGopTtl+WnXdqlS4fSJD/qZn2kQVN82YRSaoyBwWq1AVMfsL3gS7psfl3kYg/IYWiIqjyhXlB9PcWZIklyA8lDag+GgwKqZTd3FRM1PwGopGN5FQ6DWZ0WK4xoJoKg6GIELG2UlProfl+x2nli+jsDlhUPy4EwRvSjn+e1b3r+9IY6Gn+PoZw8slvU/l2rNxDzmV8neXtItE/6Bu6rcUPR4jmBS8WmCYmoB4NxZljrmRmb9lwoKmVcgLNIxVz++vnM3GKUzrogeifzvRR8jRLnCqHAbn3lLFHUx/YW3jix45vLzXfWmH0QnDKBijzdrqjwcFWlYw1QmDWJm2lYOIDpsmIDv/hoiL8D6lHOMZaJukqSckHL8ElX1S2IiQWqRR4fYaH3j6LhGyOOUhro0u8+V8CORsii33v/fBqayTRSk7lf1Zp3lfjsi0/7VDZIZW8GYvQXpH+iYXN2p5YcbQH8dG2aqwh8gkp9XXDmoi1Hn//j9/BbLLsNkDbgVuK3HGdv0j3RlIyGaEtDN/foXtjLQPXKgLU+dvifs+5ux8ukv8/2FIA+3wUp4AHlaZpBVhazntdDFXX9LD/Bi68e3DdqPZeU3vNwqb0nXclPr9CS0QsBhNGtEIFQyXhkUnPumg84OM9+dZ0wkesP4yG0/SkN6W5/RiOY3ivuHiY0w3jAwnCbrr8Enc4+cT19OGXmK7xcbFXjWbh/xwwWuVqK4G6uKl+FgqEM6PsRQw3r8DhOAb9OTiAvuopUtWZLu1g4gOmyYgO/+GiIvwPqUc4xlom6SpJyQcvwSVfVLYiJ2+rEPYCrNpNBrkJgewmeTu4VPjsGFB+p8xZ9f5GBWFbqKE4RheWwcV0q0LFEsSKlcBFNMgailO2X5add2qVLh9IkP+pmfaRBU3zZhFJqjIE6O+s7hQ1C0j/pKbRms9PqJ3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb4MHZNkdaymPYNZnRYrjGgmVPGqq10AvUNvse8LNKlEp+prxooDEabJIBcbHOx3U/Xy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPWsQ/0g/i8LaIc/j4NtRsPsNMwfWlh5XKIg4iknzwWu9cB9u/qWYJQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LuByd/PverQFaqS53zBtL8hnLXdIfXO1vNpQQWf5HvYU+eoa6rFNJu/QSH2YZFW3xFeE6ZypoaFfbWmxzHlS9XPhY+xAPB4d3kggVfaYiee3pVCSq8Baa3p/djRfyYKks99O/uKD1+pOawKYBavthoH2q801yQRY6YZnynTrgorqLBsEY5rCh9x+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCxOkt2vc9ZNFnlFEOez9nWfw9MlWEq9WakLp/n2nSKsklM7FV/qoydlVr5987fmvr0iU5SiHsM8OR5LFPC5jWsZu9niu5LqvH1TuwfQ5FlmVm+Cgk0cbG7E4woDUElXZkxPpa4LRXNXK6O7ph0Z4zqtTyOu6KxnYkMBYLB37rmkwwFgsHfuuaTCr73Isr9tVv22Igx0sCDmsNlGkDIAjeMFm0BU2Kr5SME3Ptiefzb1PqZBGwJbSU11xejSEavCb8GF+sW5GOPZ3wFgsHfuuaTBcDU+ErvoJgL90/v0Oz005vc5czTCXMWEWGf70wpKlyvt1AkOvzrPaG6h96qoENi2aTdjp1eIBwHTuv32Ju54cngOyi4JI5yTAWCwd+65pMEpiKOY/MgiRiVm6dTdBLorSFyKnSseqEWoPaPVdN3WnjMPfC77s2Y+Bt3l6y4zarUk0rA2POTQSliUd8H/OpnPUe4+pr40+z8BYLB37rmkwdhs274WvQTKG71p5NFW87CcMgqcQs+oW+gJIZi8d40c4woDUElXZkxPpa4LRXNXKWUKlCzwqQGonBGffsI2SR1cjp01RZXdDwFgsHfuuaTCr73Isr9tVv22Igx0sCDmsihzaWPLX/sjCX3TpPARXBdr9NS/2J1eOxB0dI1EaCdwuxinGJGN23xsFyxykc4vTGQci5RHCjtMHcvNDY7HcGnTuv32Ju54cTNFMUEGQGYHjwZx15J6L+dODWbmTzBAJOljepNphMcwFvjT6P0kEKXNPZYRDAtjxKL4bTgl9GUC5wC+2cLJEZM8XBDZ+gPOCWW/4dBdYxiKUEq4a+D7CS9RipjlsWqci4yHtrrI+VMFzRSQ0BCKfZkodg7Lws3CNS+NUGOoRoh/JeV/VJ1seV6vNMbwb34KrRvIdFJb4qjCaRp1c+dcyzqPzmJ8jav8gKx9DkkqvyjcAyrlX0gor6h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC5phREvPgpvHBpIYeA2rj5kBghSAkob+RtcYPplyneb5FgMEVi6IXblsFshSxqvZfeXR15LUBDW8Q9t/s4jiy19tVJMf5fqF0qOH/tgCkP0SSPXFdmWcYdvPFwQ2foDzgtYn+f/5OFuxA1urXH9DThOE/XzYSfYdP1b0SIV+trP6H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8L9I5Spepzgh2wjo6nhJm63+cPMexQsSBBQWc02j3u+2nS5eIR9+THGpz8mHD4zFabgngZTYpYIfajsiB9RthqjroTRimyHqltMpu2Wq7r+DGGp+J6yuY9aCX0ErQyxUNNVjW1fM47WbtHvc4YtZTD9jSCYyn8060xI2z39yYmxkvvCv6L7me0zZ3CBB9uJcsOo/OYnyNq/yAoYSWBy9stOqwcV0A9sL6eH4XBOP/gst8ISggg8rXMzpTOxVf6qMnZwWFEse2vnPaXIk1JlZdjcrInvCB4XJTTAWDQJ3KBpIMINkwj4mslX6OUB6hiZZNBpycy7UvdI8TqPUuJwIaTpUKXp3zNrfzFlM7FV/qoydnBYUSx7a+c9m8j3ZcTuY4tXgkDBylGzbClaqHQ6HYhZV/Y8go1wFv3Ax/kvVFV4w6UzsVX+qjJ2SOL0yshwRnPPu3zCk60TctUVhyWEPx3h9krICdrjHPCsRCyHo/0ifysPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPXVkydSh8I569gwBvbypc18gZH/Prfb6w9WZoiiFN4qHr1AgXgzKfvVYggAh2zYxKrOm4GNjZXJt3t81s5c/A11ipQ3jNDYXS8IKQH9xapKWakY/FF8AzWiweG/flnonJiN7/mLRrQX53hw/17fmDLeHoKHYA8AQ1NNERnB9b9x1ZgJhUdyymnmdGlESu52O3qWv15BBneM3HEcuJ+RvSwZzysUlAo8iA7dhRYqKr0THMW1IP+hPk/wG3SJPCawg3py20QfQAbjTPEj4qDeU1h907r99ibueHFnfpZo+TSgbJeg+iExCMrmtHnTxlMad0alyDWxEiU8Ja9CKQlY8TsI6Sgfx+TritlNOTXGzDJIU3Ce5aNdQQFCTiCByiFkIq5TOxVf6qMnZI4vTKyHBGc9OQZIm7+zr2MLg4TLFSlMPsUJYN6b3gXtzNp9Gswa/oX7PBDO6c/cLG+n1s+QzRGCUzsVX+qjJ2SOL0yshwRnPTkGSJu/s69jC4OEyxUpTD7FCWDem94F7czafRrMGv6EnBGffsI2SR5OIIHKIWQirlM7FV/qoydkji9MrIcEZz05Bkibv7OvYcdmIiNk4jAj63I2TU/dOm2PCuyL7hfJvC14sTL9rLUAscRRyaZLrh77dFtuXqxiEA/bXJzI/US4vbtZeeNd9T3NihUB6r+9pBe6VS+6e0RuC0f3wSX6TaTxTddWHwtmuqmA+PLbqdMrzqsUZ4hmxNuFqBOaMPNFKr4ePFoHgHvitHnTxlMad0UGWRiIb9KWh4cMmgMS30D0UiOnUM637J8I5Q3PYnxzLMDvPQvnae4oCLmfIM/UTQLuZWZvb5BOW7GNtU97kTE2caiSB0pwUU7QPAHasXVOgr4ePFoHgHvgBq8OYNNE4kejjhCoiburJNcLAKWIy4N2laqHQ6HYhZedK/+s2YPEJMwLZdSkMVVdTMzE3dlWywF4ruVEFfBRD7tFfp7RZlEFrrA7/ukzA6rOD2xl/IUBxrD1oOhUnp8jqbdmcoQYqPHPT6yNUvnsS4cMmgMS30D0UiOnUM637J00RpSB76oCzdO6/fYm7nhyF4i/YCvRBac3NonL3dWzRF/O8s64DUvK6maR0RWksW21F32Il+s4UpyenXn87dN2BY4w7hPMia1lv+HQXWMYiACbLWmUmE5+dGlESu52O3qWv15BBneM3HEcuJ+RvSwaFVSD1FKcXtMb2a3wBSeOcczafRrMGv6EnBGffsI2SR+2FMdHeDB4p1ZmiKIU3ioevUCBeDMp+9ViCACHbNjEqHggFQc16mFUFFHdQTzdYEvL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk91g4rMFsqxHTUfvZh6UJ3TNoWEV0YMbJgX94OU4e/c48v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEeGMqnYXNKpFwU8V7r9+cLd4kBOEElYdWw7T6JQ+hpNEZSM52hi903UThPClLMenoCv+/CmGCc2TWgxwPOa+bCZYDx0oL8iJkpapPPf6YugCL/dvNaKAYw2HyC3GItNMeIffdSuUY3eUAIEa+1M42FMqDXxlkXGyt8cXfiABmXmrekKBhVLXR57qDXxlkXGyt/0XE7CSfEGMOaPeLMwNai7s8TuxAbbvij85NLHmcF+OhlDENuglfWcqDXxlkXGyt/cxy4lNByLKctONaqaynxsv9281ooBjDbE9j9QGxx9qFPAoR7vY9rPIvj8WccgLL9mPJKZ4to+ymyu7djU1miZtqS4qdM4as2fAPOJZ5hkzBPjM7imPWpkEQOeBBUHdoorkI1Sb198yAm2XbSg4746V5tUtr/hz9Bg1MtGwBlMyMKpcqZiKlAmnsmRbfvupBFDZUxayoTvBfamYnzeoPQGLkdqeNxiM/Cu52PMC060hDHz59ILGVEgbGy3n645ZmL/qOoVrZhjPPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyPXyMGM0AOBNy3i5SNAjHO7ZNdaujmE8qBJP3vZnYqhR/0hgS820S0GBwE/B/lTHjo4dhv1qMaw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTAWnuxfXvy9lZ4p2ZOQSJTRPU5gyyFywJ/n/Odelz6zdwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyTrfYZxqBDKZavSrhn+PkAmXmk/7/DktWDwz9c8cX2oM3yHCRp5cv16eTMFa3S0m9JH4RiFSfrKeCwfEp2J5FiboR8KKvMtE2OfTLT3e9rBuWDl+4FOsmiukHNY9tc2/3Tuv32Ju54cqfGpLh8RcwNAhoDL61JMcTfs2T3tv7quVVtw4ikZM8IKUqKC1zajjbHm7A2lmZMT9qoHINnqNTQT1zWClEYtH4XLjiOTjsUyIfsv+SkPX9ysVA9Ijc/4YZBJZEZTuySB902+yXyUDt0uuKDMeEVk5nXACPzLjgRX8eXoQ8pE015+dvg3wN0oOjQ68/3TNPUeGmM340wuvpGzpuBjY2VybfOoYXf/L/aGpxk0KAaU9eZuCUJl+r1Ko6+dhSVvWRZXV5gHmKglRiDMQT5ndyMiZ8xkVW9vDPYGV5gHmKglRiDAWCwd+65pMGUmuIEf6izZHylZdJlKPU7AWCwd+65pMP9YOIVlvcdJSTSsDY85NBLKz0FvcL9nm0tfvVng81Z0wFgsHfuuaTCukHNY9tc2/3Tuv32Ju54cUbmbKWP2Zb9z1NE963/61CsS51jmg+x8tYWf/sEnVBjAWCwd+65pMEXzqeoqfDChmk3Y6dXiAcB07r99ibueHObjL9dqhg2IwFgsHfuuaTAh+y/5KQ9f3HF6NIRq8JvwJHslKXcBbujE9j9QGxx9qM/meoqjCqMoICYkcuhdGXCoNfGWRcbK33mI+vqzK689qZBGwJbSU12sVA9Ijc/4YZBJZEZTuySBS/wy2EPapNzAWCwd+65pMFNOTXGzDJIUliUd8H/OpnNRuZspY/Zlv3PU0T3rf/rUYoyrka4GD1yw4/AtNrVSMMBYLB37rmkw35uVDSA9htOF8tXaC7/x4DK4kLrElPLVoo68GSZW/J4Ya77f8vmAHRJao7CnWxLZXqGdW1doInyT+I/p7L2FsgDld8Ik6dHLLJIUpBXMDhPx5ehDykTTXrOm4GNjZXJtWsvbF38YWeSLQtQkmkitdcqJ+k5q9hXVwFgsHfuuaTD1iuTbXoZIwRhrvt/y+YAdw2Ym95CQ9HlRAMRfiUZYrGo5HDNB0yTFBEzlrdCgbpw2/ULkhwzXXn36paaXJ0Fmq7BLCzMzdrn9x/2wXHAq7K53VJAQUklV8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTbAH7uH46mzpwIyjlJerXq/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkyOYkaacOUfl99O/uKD1+pNh2Z7BgEuR7niUD75bNfNc8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEdu5GsWQ+CTZnqlEqoF4fNNJn9IO0/LopE5nYws/nqb3X9Ddi1yoXOf1/PJ4sblFSDJNH5QjMIPaNXWdKa1sD3Q7Mp45qSE5RNXmAeYqCVGIGY8kpni2j7K3OXkGArzLsM0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm3zqGF3/y/2hqcZNCgGlPXmbglCZfq9SqOvnYUlb1kWV1eYB5ioJUYgZjySmeLaPsrc5eQYCvMuwzQ68/3TNPUeGmM340wuvpHZlfh9SR/8Rw7oPk7qlpF/67gLJ+CTSRWoNfGWRcbK34/Nsz5O1DUPvxFCll4lpueoNfGWRcbK3ymqdgzo4ZHd/u3btpaMr8DAWCwd+65pMEXzqeoqfDChmk3Y6dXiAcBss32bt1w+qggJLz91HB5JwFgsHfuuaTB72cywEGpcnNOKCkPqOrXqidtz5nHprm4cTbRDnel3zcBYLB37rmkw/1g4hWW9x0lJNKwNjzk0EsrPQW9wv2ebS1+9WeDzVnTAWCwd+65pMHvZzLAQalyc8QkPL392NnKft4ug7bhBZPxSDwEvKoo3cXo0hGrwm/D7T5gwZSGzxsBYLB37rmkwRfOp6ip8MKGaTdjp1eIBwHTuv32Ju54c5uMv12qGDYjAWCwd+65pMH9If+R9bwqaLJIUpBXMDhP18/HUNm88hQcA+b2PnsTy42AmQ2DxbUDWicDCQk8Fiag18ZZFxsrfeYj6+rMrrz2pkEbAltJTXaxUD0iNz/hhkElkRlO7JIFL/DLYQ9qk3MBYLB37rmkwSPZCjBZnXw1I4AvLdsMvpYVYP8izPwbjy85Ms2/YvzkyuJC6xJTy1TYAfN5hr4QEwFgsHfuuaTDfm5UNID2G04Xy1doLv/HgMriQusSU8tWijrwZJlb8nhhrvt/y+YAdg1YFRsRCSxapl7Nk+TGKVaxUD0iNz/hhk+O7dGqPPQRzNp9Gswa/oScEZ9+wjZJHTKVS+fDCQUJay9sXfxhZ5ItC1CSaSK11yon6Tmr2FdXAWCwd+65pMPWK5NtehkjBGGu+3/L5gB3DZib3kJD0eVEAxF+JRlisajkcM0HTJMUETOWt0KBunDb9QuSHDNdeffqlppcnQWarsEsLMzN2uaOQKYsC2AmQ/6jqFa2YYzzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMj18jBjNADgTxI+Kg3lNYfdO6/fYm7nhwuea/JZVNP2QpSooLXNqONuLbu13agDlMZhKx9mlr7aQpSooLXNqONsebsDaWZkxP8Ug8BLyqKN3F6NIRq8JvwNVK9vGqRpzpcF9VXEWYWH6xUD0iNz/hhkElkRlO7JIH7Em/LVhMXt/Hl6EPKRNNesCUt9y2505hyd6Bu0cxjkF6hnVtXaCJ8k/iP6ey9hbL8Ug8BLyqKN6xUD0iNz/hh79AultxgZkCuX4NqRgbVYXZsepsqC2cUcyP8LAktKTFCh9UaQDXif1DHPHgFJjKgH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LAMq5V9IKK+rVSrYO2jw6FQdwchiv1QTp4it2tMizOZkUEA5tPhcluXAq0axs+DeKxT8E4X+MTvd+SnBV1xlcDSxTeuC4B+QjAMq5V9IKK+oR3YktULj5Iftv7hef05vdHxIjz5gCL21n1jfmKJE433YPa4lVG1jXnBZlDDWPRc0fpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv19JhV0Bg8FAX8cYC1vw6ZInrSOdnQKWp0tGcGsxfg0omtQ797AIb1pn5zUaoL+FImERhWsm5kQkFnNNo97vtpDsuOAuWahUAp+b8/epKVmw1fLXh+RnpyY8K7IvuF8m8LXixMv2stQO1r32W9EobICqD4nUayamL3FBVXLnrdhYLkAzBtEkvpXgkDBylGzbClaqHQ6HYhZSqiwbt8jjHaOLU5nnUugAcwICxouRz2wyCL0/lDTkTEGB6jBl007Ic8OcUvtKIUaMtTNNKBXsMOsfEoSEIM7uVeCQMHKUbNsKVqodDodiFlyvZhKluyThkfcsHapQOQ0JTOxVf6qMnZwWFEse2vnPZYXgyXk/raPV4JAwcpRs2w1ZmiKIU3ioclBrYPaT/VkOxjbVPe5ExNn6ADi5zKCB+lqmFVgZ1MPmYCYVHcspp5nRpRErudjt6lr9eQQZ3jNxxHLifkb0sGc8rFJQKPIgPYMn+n/hOve2aUWvu4AhcMlM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw9Vm/O3LQvkUuPqFpjzn2ScrD1oOhUnp8hO7JRb/x7EOE1H72YelCd04d25Ov43oRL9fWYL+PrUhR2DWy5n0Tr/idtz5nHprm65Dxmmqoeuzaw9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9akY/FF8AzWjk7vOH1LLGLR72ncro64s3bFg2Or5Tn2CxQlg3pveBe+NgJkNg8W1Ax0ozqF4iw/RMIi/u20dzbhFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybTxI+Kg3lNYfdO6/fYm7nhz3IEJC81H1gTGFM4H4efwuTkGSJu/s69jC4OEyxUpTD7FCWDem94F7czafRrMGv6F+zwQzunP3Cxvp9bPkM0Rgi0kWLnusckK6maR0RWksW21F32Il+s4UXBfVVxFmFh+sVA9Ijc/4YTJU5QDL+3syTCIv7ttHc24RaygtE5naOViCACHbNjEqEbixuPsCC6vwcJ2XJkwGgInbc+Zx6a5uWrVxQXYuSnmGH/n/2B7cK1rgSNBvfq0OZf11sV/DEVQzICZGXrCzkjSCYyn8060xoSF3Q0r6i7Yr5MLZhS3k9r3lVbkVtXI59fPx1DZvPIXe1qNZioQyIAFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHQW6A1k/HcyNTTk1xswySFNwnuWjXUEBQ7YUx0d4MHinVmaIohTeKh69QIF4Myn71WIIAIds2MSryTKIkUcCMHe7RX6e0WZRBXqGdW1doInysLYGoygqbpjA7z0L52nuKAi5nyDP1E0C7mVmb2+QTluxjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3axUD0iNz/hhMlTlAMv7ezKvh48WgeAe+K0edPGUxp3RqXINbESJTwlr0IpCVjxOwqExlKxSUW3tOjh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2epCRbrACC7PJtq8dKn8FhDlTlogd91ZDKcnMu1L3SPEcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPMV77l3sTy2gteLEy/ay1AZewjlq6V2B7cskGuRzF0Lh1nNtWiC93BkTDJhlfKOdcK3OJbrgocAiPwbd6jtD0Ks8TuxAbbvijjo7C3kNP3INLkH4dC4si1L7n3mFDlx+KboR8KKvMtE6xlrn6QXuemiccdViuS2KCRjGUlDW9J9MjKJEPF85qP0fI81agyzrE9FnxwYF5MXUBuEIh57UHU7Ili+TO6kwDK9mEqW7JOGfoRoal+XLywDVC61irCVcHuvtGY2j5/QW91zfi78Dw6bcW54N9/A+QvufeYUOXH4pVVC/ajRiRXJ5b2RqYp4khU7M7PInj7X42aUZ9CPIbWCv9ED+Y/TDG2Zoxwzadgwag18ZZFxsrfzVWgefLB9+0ntQyxMoEi6r/dvNaKAYw2TUfvZh6UJ3Th3bk6/jehEv19Zgv4+tSFqDXxlkXGyt9eTWhK4xsxKXx1o143bV27l9Ky46TX1wh6VrVJn4zOc58A84lnmGTMay79/pMxdRsf3i5JiFZy84LQ04Y/0qyIqDXxlkXGyt88SPioN5TWH3Tuv32Ju54cYs2s9iLj3jEKUqKC1zajjbi27td2oA5Tv9281ooBjDagjm3Nb4yARPXz8dQ2bzyFcHvbVgXuI+FTTk1xswySFNwnuWjXUEBQQtCGF+QhAnpcF9VXEWYWH6xUD0iNz/hhkElkRlO7JIFzSukR8JKCBvHl6EPKRNNe+PDTXCmJZ91g1MtGwBlMyMGLilyNiLjCMriQusSU8tWqfAtLY6eGvVNOTXGzDJIUliUd8H/OpnN8GGkjC/nuIpdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm7M2Jy2rueEbjYCZDYPFtQMdKM6heIsP08Akk+MZCkjyNrCWlmF07znTuv32Ju54c3wUXdvcyv0Kgjm3Nb4yARPXz8dQ2bzyFneP0N/uBkPMxULtU24JShQpSooLXNqONsebsDaWZkxNamgl93Gvh5lNOTXGzDJIUliUd8H/OpnOzGnDL6qMecNZdNsyqy9LIczafRrMGv6F+zwQzunP3C21dIJZcC7GwwYuKXI2IuMIyuJC6xJTy1XEOz+xggGuJMVC7VNuCUoWBY4w7hPMia1lv+HQXWMYisiqXjDkth61qbuITBtwgaw18//UIG53xSobEgpG71M9wukwNlc6T+h+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC3eCMgS2aQYlSf8lVN2ZZgfoxCFMy3ABQrty9SLWj9MahDVHhRSEtqXSdRsYz5JZBMnmvXHN8NcKUL5H3JR+gnQZvxh72Y6FA+VPnyoAOCdrJtrrWYvsHNmJ23Pmcemubi0bluF31BjZe+ToSZEujRSpP+Wem6+qbcSdxR8LiiPb2bSy/ssm1qcfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu84Qta0VhokDGQv3X6heHUAAcouGPgvdGNanhf98S2FY2x2rG/JzSm++E74jtv3CjXqdpuCbaDKLCOjqeEmbrfNg0ZOIlCNdkv94TlSlGhCUZ6CCfYNpaWND5/1YD7AQ8v94TlSlGhCWL0YIzvLQ8VIqrp3xKIxtDtG1k0bLNkme26DEPZAh35idtz5nHprm7bO4G7LQzeWnVODk2HTHtwAS5nS1UYf8Rb1SAIMdbJuGg3G/JDxBbWUwPo7WNmxPZt4I1zhKJNEvi54OaoeF/Z4SQKv0LJm42cxC+6eqjMUMY9sbhti4aW1a6g6wwTrBXnSv/rNmDxCTx1jO3+HDIZ0pjFGq+1smHtMEoEICHI//FoG5ZSuGPqqe/scAU9oL725uy1f6d1U61B847iMrHmRYhohQbvuYDHuhOXTeaFEQQTKhkCMCgM0RRoVXO6yLJG8h0UlviqMJpGnVz51zLOE3MZ/3HsQPDKAMRtqFOjmWao00x1enIKFJVOS/zOfjAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctBWUqh8ccsm2utZi+wc2cjOx7LgKysZ1ioEByRFu5q/m9ftHBTauKeUesELTuRK270nmAeVpWqKqvgwI9x/utdQxQ/1o3LCLDdI9OVRdvOOQbCAZ+BPqTxhZryFbn9nXWyv+HBl9+2E/XzYSfYdP1b0SIV+trP6H6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8L9I5Spepzgh2wjo6nhJm63+cPMexQsSBBQWc02j3u+2nS5eIR9+THGpz8mHD4zFabgngZTYpYIfajsiB9RthqjroTRimyHqltMpu2Wq7r+DGGp+J6yuY9aCX0ErQyxUNNVjW1fM47WbvRafQqGpk4qbBQFOQvZ3yiVjW1fM47WbtNB4xZLhbP1C7BdOXRkn+wND5/1YD7AQ8v94TlSlGhCUZ6CCfYNpaWND5/1YD7AQ8v94TlSlGhCaCqNBkpBYoKCnCHVKTy5iU0bOxDv8HmnztPolD6Gk0Ry+ka9ka/GLwjbPf3JibGS9KAiuTcO6Px1knBXlhDPOjbO4G7LQzeWrBQFOQvZ3yiVjW1fM47WbtHvc4YtZTD9vbm7LV/p3VTy2MMpwoe9ECuesPL3HrjaJMmDNgWDJggzl7Jo0CTCDkKoPidRrJqYvcUFVcuet2FguQDMG0SS+leCQMHKUbNsKVqodDodiFlKqLBu3yOMdo4tTmedS6ABzAgLGi5HPbDIIvT+UNORMQrojOorBNgIgL0kEjdIIoXHYNbLmfROv+PkgBJUwhBsjZtTT6uy6iUwR+mm+pxTPoBq8OYNNE4kRLUX4/SMqrV3hI1zvf4/zcd23GDqg4YIyiZ8hj5jclm4cMmgMS30D2ncXb8pkNlLUJD9RYEgn3v/zdjE2h1RvcRaygtE5naOViCACHbNjEqs6bgY2Nlcm1UFF0KLvkcR81F4WizKZmEYX0HiBSNyGI8UrTlyyOsfI3SSFu17+KWJeg+iExCMrkBq8OYNNE4kdz0JJUew4U+9bI4ROdRjGsHCIkzAlfR/DGTzC+tFdi17GNtU97kTE1HZ9WYTKq9U7ZZzmiwPIDz9yBCQvNR9YExhTOB+Hn8Lk5Bkibv7OvYwuDhMsVKUw+CxfZwGW1tTJeq9wko2zl+FMinNZ60OfPuoJ7of2ZweUIUGh1sl2hPAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4d6KJwYfaUHKD4wy5xLR5PYqiSqI1Y4a0DiN7L9OTBPDcFOlKqDpMwocXo0hGrwm/CH+OQE6RbVHR3bcYOqDhgjKJnyGPmNyWbhwyaAxLfQPZucCMu1RG6NClKigtc2o42x5uwNpZmTE/83YxNodUb3EWsoLROZ2jlYggAh2zYxKrOm4GNjZXJt9cYajgjHtiuZ5Vyg3Slq7EzRx7e39Um0Hdtxg6oOGCMomfIY+Y3JZuHDJoDEt9A9m5wIy7VEbo2BY4w7hPMia1lv+HQXWMYic4SNAPWFs2eLSRYue6xyQrqZpHRFaSxb7N9ax/BvGXN+TFSQ0YK9gOi344puLZ6TiH0OH0ZEmseuBmteAD/0kHMj/CwJLSkxu7QNatxTR0YeEyzQ8WsjrozD3wu+7NmPKaC9KZYGkVTuxsvB00awOMY9sbhti4aWS+otvOAZIEkr5MLZhS3k9qduh6Ccax3+aGYQK30rOQh+huMKSsoteliCACHbNjEq8kyiJFHAjB2ECyWlhTEG2yHeVQdh63s4VMz8s7lE/N2Bxl0y+KwUu9GKG/xtD4e950r/6zZg8QnAlCJBb+ant0zRx7e39Um0i0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+In9FHc1iKADHD0toaJ1zhYvEWsoLROZ2jlYggAh2zYxKvJMoiRRwIwd7tFfp7RZlEFeoZ1bV2gifKwtgajKCpumkoejOOHQ5KMomfIY+Y3JZuHDJoDEt9A9FIjp1DOt+ydNEaUge+qAs5nlXKDdKWrsWoDLYLSKRSOLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhTVVUIwdGtIENwXYbDRREPZNWYnM+lVTIRhw4ye9aQIFVRWHJYQ/HeHQW6A1k/HcyMPxzTSIVscY8IIPxBr+NBQ/JM0QwbobnXC4OEyxUpTD+dK/+s2YPEJ73cZ3DCZFxwOV6zbF9fA6YnQe5Uf6V63WIIAIds2MSryTKIkUcCMHcVNzNk/5DKQD8c00iFbHGPCCD8Qa/jQUPyTNEMG6G51wuDhMsVKUw/nSv/rNmDxCcvOTLNv2L85SQnhjGX6DAh/rmlOCs+pkTGTzC+tFdi17GNtU97kTE2caiSB0pwUU8nghxtgSf/dcXo0hGrwm/D9mg+vlZNWiItJFi57rHJCupmkdEVpLFttRd9iJfrOFG+wihoEHfiJQkP1FgSCfe+ym6TZ+4ZAL/SjPdZPbMmLdiMl3CC5FgANu9GXfU3btedK/+s2YPEJ5FD3qZeR9ZD555utOKn6IzBszIs4p133HEcuJ+RvSwaFVSD1FKcXtHIM07ImKul/E6NGL3neb/djuqaY4wcJjgnmMKtBe4c3a9CKQlY8TsIr5MLZhS3k9vUr25bkj0n67QnN/bBZVR2LSRYue6xyQgJxrYyvr9AVbUXfYiX6zhTVVUIwdGtIEEd84T3o1lkkY7qmmOMHCY4J5jCrQXuHN2vQikJWPE7CK+TC2YUt5Pb9rNQ9pMjFpzQ7e1k80Qpni0kWLnusckK6maR0RWksW21F32Il+s4Ub7CKGgQd+ImVhqsillAnUmO6ppjjBwmOD7DkI+4jM/Jr0IpCVjxOwivkwtmFLeT2h/+1DVOfI068YqKDKfFsWsuftvLrSGNFlM7FV/qoydkji9MrIcEZzzgLIkEoIHZdVht/0VhHvqQRgZf3KU7i+TokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyV1G0Y6W/jsODuBCGVCiAh9tBJuddKMmnOiRo9jXnvUPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTckrJJsGiVHIBwEEid0Xk4SIAQQY9C2veCkg+do3OI16JRUq48mlZrCDgZNW7YsKRYb45kLdWsJDInirKBcADewvvfBO/7LF6msAgkAG5f2dTJlOAccGZARcyLk87kDNWHxQr17pO3GwJDduZ1NMfBKw9aDoVJ6fI6m3ZnKEGKjxoHqLkvghI+FyL+851qizMnRpRErudjt6cepaextTSItJjQ+7kSrnPcCMo5SXq16vy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNyukvJ0+dhsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkzn2Cf6wkDYmDtqL784shMEtWoZ7GLFEjzokaPY1571D8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3JKySbBolRyhpW7cPg9EnFfcgXPscSDtiZeaT/v8OS1YPDP1zxxfajkJGrPv+AUqh9TFW4JdLljl7deJwMlll9DWkWa+Xbau5XMGykUBEJZlpwAZIX2MBvYrqEx1I9NHDfqZVk0CUss09Dv8uQU09N88Ge1xrOKSS3CepOro0C7YVxXqkpAiBj9FHc1iKADHCdRbueM7dJ7PwGopGN5FQ6fmmS/7b21AHXACPzLjgRX8eXoQ8pE016L36PK5wBCxx8Y8QTsDBkOrFQPSI3P+GF4Wx2Di67ldqg18ZZFxsrfU05NcbMMkhSWJR3wf86mcydRbueM7dJ7wYuKXI2IuMIyuJC6xJTy1bVUshcnsQ+unwDziWeYZMwWvtshoJm9jaVybwa0KtEH+OSEWtOk2Hl+aWXsl30uMWBscT8ZbRQBuLVLYsaYmwvLzkyzb9i/OTK4kLrElPLVNgB83mGvhAQ5w1mjPaNT8KV28Afnmg+YExjs5JK/InZeYc0TbKcVyoFjjDuE8yJrWW/4dBdYxiKyNcfwmy5SoYGtcUQFzb4Xt0xFngyo3EClSZ0z7Bld8JDRDzKAm9d673cZ3DCZFxzC4DX0AO4H1635MnS5THCRgz5oQLaYuGZrHszq1lh4rvaK6mWAIB6bxtzYw1dwYMtatr9VNODlif+o6hWtmGM88v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTW8G+UaBphGU6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUchdUowDY5SJp1EQq+XMXAFiocrqxY4Ln6PL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxZJjMs+JZh85ZWoH4A8ZKXuaMqCF3iWxbsDbvaSa+SnqXIk1JlZdjci2qYd2EgdKtDQUFJSyD4MVNhDOo5YPnV/ML3EO/WvzNjhwIGUocy7GoNfGWRcbK31NOTXGzDJIUys9Bb3C/Z5vx6uW325OK0mz8/3OvySf9oj0QCQIThh4SWqOwp1sS2WusDv+6TMDq/v4bE3mH3DU0OvP90zT1HhpjN+NMLr6Rs6bgY2Nlcm3W6GR/nSUEpImu+pg8kxLl9qoHINnqNTTDk8jS4HDXZECGgMvrUkxxqvxPemSJzH6oNfGWRcbK377+9m6sTA25qfGpLh8RcwNAhoDL61JMcTfs2T3tv7quVVtw4ikZM8Liilibd7xVDL5zxI7TXmNiUQlm3kjqGg3mJGcwwwWk+yv3EGN2Uc6YbZWbwjzgDjT2qgcg2eo1NBPXNYKURi0fhcuOI5OOxTKDcP3Kl3r1iAZbYNk/Mh4kNDrz/dM09R4aYzfjTC6+kbOm4GNjZXJtYK3CE4cXXxcIm+/CbkyXViVfbovfMR6DMMIMVCYg7BmoNfGWRcbK3wwdk2R1rKY9vnPEjtNeY2JRCWbeSOoaDeYkZzDDBaT7oSpQgBt0sRL67pZhSX17SCAtZkpLXQwgNJzdH8dDmd1kv7zXjDWsli/Ey5zgjnpO8YQPpxh+N2g2uXO9FnjWKZPKwZ8gNmtnmNjZPrsSz73Lk+ksSBii9FVbcOIpGTPCClKigtc2o424tu7XdqAOU0/MTsEX+1QQ42AmQ2DxbUD2/isXJoBuaag18ZZFxsrfU05NcbMMkhTcJ7lo11BAUHtZWtuiP4GaClKigtc2o42x5uwNpZmTEwKB52gK4D7dWuuEnttgnLZ+aWXsl30uMRkgHGlN4Yp0bP0QjGEtPjJucdNMECAza18xgZ1e9SeEkNEPMoCb13rkUPepl5H1kKV28Afnmg+YFWLngtvuKDrkyA/eCe0YuQGvSEvl65pFp9BGrMNZhlumYURHNrLDk1tgTPaPY4NfLnmvyWVTT9niilibd7xVDJ+aZL/tvbUACm3/7xmbcxrM30VW848PY+RQ96mXkfWQat4brw5j6CZCQ/UWBIJ9714exXekNcaRAoHnaArgPt0iEFgcKS80jJCGwyPdZ4tcddoq1uBb+3jCHPSQmbkgPkJTWrvHfodyU05NcbMMkhTKz0FvcL9nm5k2TXcn8hluYVxXqkpAiBiVhqsillAnUulu5XUa7NdTSRqvrav/w8JHfOE96NZZJNBVSvLqOS4UcXo0hGrwm/D8qmKK6MLbPdtbv+xeLKxwkqBrVh6zEKAjuQen7Od6z1fQsuy7XWp2QkP1FgSCfe+0rCGMeKg5mdzUcTNyiZjl3KjZPqsRiGA2n6KkkWCc76kKusz0wYsiFQRTQg1Qz1C4o+rELtG0rzGc3nODWG+mwx3aF1+LE51SQiTI9fxSysCUIkFv5qe3q0oMMMiW2kmG3f4YTqOiFbxiooMp8Wxa3KjZPqsRiGA2n6KkkWCc76kKusz0wYsiFQRTQg1Qz1D4Fbsq/pafJ4M+aEC2mLhmax7M6tZYeK72iuplgCAem1JGsz31sskthA/1K8xJSFRccVcmfH49K/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk4Ull/LbH3nTjfuoxOiR3gsP/9hTuIR62bPyE9mT0B4Zwx3aF1+LE51iPPbx3cBazFZM9fmLyJU+2yooR3rR3bGj1LPZE6uc4sLGR8ZjESG20Oe6Y2oFJJEc1hCg9j6TV7PyE9mT0B4ZtF4E6dtJ6DI6OHYb9ajGsPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQkwFp7sX178vZJxySuyuWh3uG2wQmryA5pfaoV1U/wv+YeQNK+vHa1FwL39q2OrdvMfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk8Ldp4JaxpvxTrls1ZJGB1d8EgNGoYoA+k86/2QZrtGwSweZ3UVRh51GqhBrmBznHjrhvS3E7tUlpH+iYXN2p5aB6lEntCuL28CUIkFv5qe3e9DNL0JiEfk+3wUp4AHlaZpBVhazntdDFXX9LD/Bi6+Y0lrrlWmnAAY3NfbQXckUwxUdIyEIHcTIiNakPA7/yWX1RNWP+Q+5ZeYrvFxsVeNij+EL4Jb83mwSQQp3vHfYvaodYXuo5QCjwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+yerg4Gueif9EJD9RYEgn3vC9UxHq3ksiZGePBVStwkpeHExRpRAhr9LEXGmfgOzLMJj2LXsH8WEtjZbKruFW/susYanHoofj0PyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoPBJmRrhKB5X9sqKEd60d2x2N71FU5195jH1yKtFNcUngVg8qsA7GjjsOW9w8BUFblrS1TXObGJTqZC0iaX6mJKGC1UJbFNTrYnenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvgwdk2R1rKY9g1mdFiuMaCY8dYzt/hwyGSth/xoxHItyXh44Eru+G2/DFdE/EjAVqFsM7Bn8/nJSa6wO/7pMwOoAiS9cHv8PeSd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+9cYajgjHtit07r99ibueHBiU/p0DOgML1b9VfrL9uF6dYzRILyXK7wAIENq7GEAzcHxRN4xA7uu2sBF7DcfTs+NgJkNg8W1AIiFUSb5Bm9fLyclcgJ/T+KuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSJX37UfHsVfx9fPx1DZvPIWcJARBsKaP68l4XyPlR7lWNVZGb6vNC+YoSLm/Hcy9hygqZVyAs0jFf5hX1cNB9hyBY4w7hPMia1lv+HQXWMYie9DNL0JiEfk+3wUp4AHlaZpBVhazntdDFXX9LD/Bi69969UIqW36JHM2n0azBr+hfs8EM7pz9wvY3vUVTnX3mMfXIq0U1xSeWCKf/pFB1z+w5b3DwFQVuWtLVNc5sYlOsxbsDvRZdZKsVA9Ijc/4YWwQvjzMDdHky8nJXICf0/iriPRL5pV+nkt6TzEWbOYiUlO5TcmQkUiV9+1Hx7FX8fHl6EPKRNNeU5H9GC0Wk3cSmq9rOD/u8tXyXX2KMXIhDJ9LeExL72R/x+iCgxSc9pdgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxmam7iEwbcIGsNfP/1CBud8a6AK0y7DOlC5mw8QDXyQrEfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwvDvs4X13is5a+X2U2Sr4h2tfpPQ2kXFtYhzzdEPSJT5a+7grw2Uuih50Nrz9FNAQEPr2LbsPFQc/85hXRHi13qvfqYTuVYKVl0u4Abt8zT7TWUWgnEYxS+p6Bxh5dCP3ueUPML9TIc5yYo5On9dJRz0BWGIZflwCoCdSnPogmsemGZ8p064KK6iwbBGOawofcfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsTpLdr3PWTRZ5RRDns/Z1n8PTJVhKvVmpC6f59p0irJJTOxVf6qMnZVa+ffO35r6/nq6oodTOP47oStch1nvBHnJbp6P6y4xYyWpHpKzStagM4WGeNExWBI2z39yYmxksbqopsod3Ic94ypVa+T5wZPWSA7yLFqU0a2PDz7v9VBOUN5Pq3V+oLAW4EXs3c+9NcIJECOL9wK2g3G/JDxBbWOrNdZEEJcukhQsoGMdsL1msfbEm4KgCU0R2biQCYPlxVxXZny2UoGUg9iON0OTU69CAeWVvvRXVRpjNvcV01fPgH6mKA8iOZqIMJuFKHh7Lss5dabj+Yg94ypVa+T5wZPWSA7yLFqU0a2PDz7v9VBA/tya6/o54mtIJeCh/F2NAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwu3Hm/ZH/aLtBbpxHe6C3zjI5KKRRHzgmbq+3uWHo09MTIiX21wO8isrBAUwGum2YW3YWhxFO8Gvb5iRsgxnwD527/LebCgOWq+e6N4jtRobADKuVfSCivqYrwr8Zr4As/LN7EBYOe22mj/7jB7SARWtDPLtgm1BiPaObPiUIfhsR+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCy9lfO8WMOT8TyMKatMDfgQK55YaiicrcZj0EJIIrJfLWJ2KnGVS4jRLfeFRTmgh0QRYfj4vCt1JjWp4X/fEthVl3pEEo0zoSKn0kHG8CNQXnAz/tY0NP4e3cejq3/OveSygZpjnuuyyO0+iUPoaTRGiNFH2NtD6fjRs7EO/weafO0+iUPoaTREV+wVeeATG83nfaYqNGzwC5D3OwqTwAiJ1dCgW/W9lYKIH1YHvpdxksFAU5C9nfKJWNbV8zjtZu66BdPt4ta9+W5wwOVSASsU0Pn/VgPsBDy/3hOVKUaEJfnnYXugKDA1qOuOvdVDCHsoAxG2oU6OZ16nabgm2gygUDq8zao+Gqrr8J8oS8aJb5qJWUQRvcWSLK/sUI46V8YdjS8RXNV4pGindyFNVcwHCwiMWtGji87fCS7R4NrAvmo59SWkrRX7W5eVBSW67U1QpZ+tnWt5YJqWbEMG9PrJxX2xf0wa4olMzMTd2VbLAHYNbLmfROv+boR8KKvMtE2YCYVHcspp5wgpAf3FqkpYIPrN5gXWc15kLg62wnfIElf087lBdQfkwICxouRz2wyCL0/lDTkTE0eLVINCmTFZ5s63yiIExvXLkwrR+v8SSp3F2/KZDZS0FSl7jwbxSJ1xLzhnLPbnBrD1oOhUnp8hO7JRb/x7EOGxHoMmoJRXKqQ9E78HC2+We89mzNgf3y05Bkibv7OvYwuDhMsVKUw8B/WwMvpibSmVsn5R87rmOi32YOSX61agxk8wvrRXYtexjbVPe5ExNCDZMI+JrJV9nQA9Bc3p4/Scckrsrlod7I8v8JpqqcQbc9CSVHsOFPiKcIW0S4ke4j7GeEBde/DuUzsVX+qjJ2cFhRLHtr5z2/id2tyC4EWx0t5l/KSVXDLkOsWPaq9s5KJnyGPmNyWbhwyaAxLfQPfj10qKusZM2lYarIpZQJ1KTiCByiFkIq4tJFi57rHJCupmkdEVpLFttRd9iJfrOFLzR89UNRM5NlKbPj9+iHGnkcnkKrnpDwxS2UoimbAzEYqUN4zQ2F0udGlESu52O3qWv15BBneM3HEcuJ+RvSwZzysUlAo8iA7eFKDiZSVOVFLZSiKZsDMRipQ3jNDYXS50aURK7nY7epa/XkEGd4zccRy4n5G9LBnPKxSUCjyIDN3ncyBj5kQIUtlKIpmwMxGKlDeM0NhdLnRpRErudjt6lr9eQQZ3jNxxHLifkb0sGc8rFJQKPIgPQVQhCSehFqhS2UoimbAzEYqUN4zQ2F0udGlESu52O3qWv15BBneM3HEcuJ+RvSwZzysUlAo8iA4CAxv9na6VITGnZ8m8TbE7Dhxg6ak1chprJYspl083tCJ7LlVGvUlq0WVUtAOZfnvfIsUQ0jlrJrD1oOhUnp8hO7JRb/x7EOO64dCfBbeDVIkKR3IvQI8gHCIkzAlfR/DGTzC+tFdi17GNtU97kTE1HZ9WYTKq9U6He0LYURydZK0PhJuLRlye5DrFj2qvbOSiZ8hj5jclm4cMmgMS30D1qRj8UXwDNaAuxizP2bUcBp3F2/KZDZS28C1sSUY9by9096ji5zwFdcV9sX9MGuKJTMzE3dlWywDbhfUs2/G3PYHkQ+ywxYp8nDRel4faEa3CAjfd7xQL2m5wIy7VEbo3uqzrUUL6jA1kP0muh7dxwHdtxg6oOGCO5mKZPaRBfYMLg4TLFSlMPKqLBu3yOMdoEcTJDx96zHaKg6ef+jn55ZTHmGcAOxiysPWg6FSenyOpt2ZyhBio8KHKNfOIaCSzC4OEyxUpTDyqiwbt8jjHaUuneTJL9hFy9zIVVBTd7poDz7x/K4WMMXgkDBylGzbDVmaIohTeKh9cmIYqSm9q57GNtU97kTE2foAOLnMoIHx3MlbIhFGnUTeY85nAP6AivDNBxyCMi6BBcYyRrjy2Po/fcjlASIKwcRy4n5G9LBnPKxSUCjyID1sQYO1fcpeu/EVQ1L9Q85HT1OMxyaa4kXgkDBylGzbDVmaIohTeKhzIRSWTDxSHxWIIAIds2MSqzpuBjY2VybWSR3DO4+l0Jx3Ki6aiOBv2gBtrqkXN7BHFfbF/TBriiUzMxN3ZVssAdg1suZ9E6/y8HEVEKPmLf0Meym+qb24vmZPaHPZVRNxBcYyRrjy2PNrGMjGis1QocRy4n5G9LBnPKxSUCjyID1sQYO1fcpesHhDgYvs7CIO8AC8tnYUSJi32YOSX61agxk8wvrRXYtexjbVPe5ExNn6ADi5zKCB8dzJWyIRRp1MnwQn5HMaOUuDPJL5MM2pZTNm7vlhR09eBQM0cBZ0KcwuDhMsVKUw8tYAA5kqse/gbB1x6hI2lXvXolK5pzHUZeCQMHKUbNsKVqodDodiFlLWAAOZKrHv4GwdceoSNpV1KUnG7T12N59KM91k9syYucOmNUNiQp+cLCIxa0aOLzS9JKC+EaKPzhwyaAxLfQPZSCP2HGGXrjE35JoD5HJZfO2tIEHj2/xPSJ52KAGWjkniv+1iNSrX8PWlYPQNmfJajntpcAlJr+a9CKQlY8TsIdg1suZ9E6/1NOTXGzDJIUys9Bb3C/Z5snUCoE+R7cwXVgpvDe2lFKHEcuJ+RvSwZzysUlAo8iA3LQrjN2ZRXu9fPx1DZvPIX/ibx74/aph57z2bM2B/fLTkGSJu/s69jC4OEyxUpTDyqiwbt8jjHaczafRrMGv6F+zwQzunP3CydQKgT5HtzBdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDctCuM3ZlFe7x5ehDykTTXowe45iwHqh3yVCHDB3/kewPsOQj7iMz8q6E6k0oCYu0+EluFqiHje8QmDD1ZmbxHz1kgO8ixalNlQw9Z6/6lQFa4EjQb36tDmX9dbFfwxFUJPHaThUAXmIFid0AHkg1uAXulUvuntEb9g85bOuv9pvgx/liKPdavJKHozjh0OSjKJnyGPmNyWbhwyaAxLfQPRSI6dQzrfsn/0VFJniP9y2CZGxSkRLzrotJFi57rHJCupmkdEVpLFttRd9iJfrOFG+wihoEHfiJj44EHcmWcLvqbJw4U1eyg5TOxVf6qMnZnRPJTL8CXosaVwlQ67rnaODH+WIo91q8koejOOHQ5KPveW98boqideHDJoDEt9A9FIjp1DOt+yfXAE5hDbOljoJkbFKREvOui0kWLnusckIJrXE3nd7zlm1F32Il+s4UncaLrFKUm4dYj89OQCzh2OpsnDhTV7KDlM7FV/qoydmdE8lMvwJeiwA/UJGcuuQV4Mf5Yij3WrySh6M44dDkoyiZ8hj5jclm4cMmgMS30D0UiOnUM637J1O1hzaDNeLxgmRsUpES866LSRYue6xyQrqZpHRFaSxbbUXfYiX6zhTISQALWFAgvFSW1B46GEvM6mycOFNXsoOUzsVX+qjJ2Z0TyUy/Al6L3Ue+sVPao9Pgx/liKPdavJKHozjh0OSjKJnyGPmNyWbhwyaAxLfQPRSI6dQzrfsnjEUeOBs8HnqCZGxSkRLzrotJFi57rHJCupmkdEVpLFuNdQh89Yc9medK/+s2YPEJg/ncOa6ZVqVl3/JOXLbMgqGNz6f6pw+jnRpRErudjt6Pa8hQIu2MdliCACHbNjEqIvyDxlgqBzbbA8chY5Tt3Gk68EBfYWYYxNmtH0x0Cetf4nFInuvbJQFg0CdygaSDksVqJxdxStw4HXb23V+jBW1F32Il+s4UXv9yBR+/ijDTgI+gsDxqVTA7z0L52nuKAh7GJdVdRXcRgZf3KU7i+Xe5+Pg0gAw6gkXTrB5PTrHmnWkGLugJ85dgPw53gZIl8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk+FRkIk44Zxm2wHhkpjJuW7ItzCLx/anPpIDt4/x8hndl2A/DneBkiXy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT4VGQiTjhnGZTLX+5CB5ul/WHb5n7CD8xOaruDmZXmMLiQE4QSVh1bMJIBjvr8UD0jA+OnBq18uJvaTYvfvLB7LLNfbZhUPHlJ9iYlPGJoeX+Zfjrga4Apz7/yAYt6T2aJeha2uICFNfLRhPgGFlt59Crq+9aP37oqDXxlkXGyt9Yt+40/kUJWGf52OwzgI9ts8TuxAbbvigaeSEc5Yud19epfUFxPX1+l5VLDx54rUEvufeYUOXH4ln6Cb21JXNZxPNyWnEsWwaUytPcZGSb9eY4yvlTLgmQv9281ooBjDY7LFBnXdjbx3M6vb13oGie9FkT/f+3TGxOXXxxNZK6ipGMZSUNb0n0i0ObZKSgLuZWYuTZOUuk8CzlFL6DMU+kbkp0z2Z7gpWoNfGWRcbK3xUEU0INUM9QbKvuBcrZRNY/AaikY3kVDlM8AlJc5jazlXeHI7I2QVs9UeFmpYZozIZD0YxFx+drsYaT3SCOpapE3tygC005pCcckrsrlod7I8v8JpqqcQZhfQeIFI3IYtSMm8EQGs7zwb31UJ2GHyjY5EgCcQqeq6g18ZZFxsrf/id2tyC4EWxwe9tWBe4j4UH3SRcPn5N+fBhpIwv57iKXYD8Od4GSJfL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPhUZCJOOGcZnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiZDQIny+n+4gtIl9iCT0SzUnUSdnSVmnNnVguiwp5cHh/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk6MOrxET/cLaYUE3gRWQ3UwSNujLFNzqCzR7x7YVGOZYjnCw3frpxtUC7YKbRCnvybHkJ+pYPBZSKNIsS9eN4Cct3RFoJP9wkAPjnNTabYevUWPn5y6uxfw9TfXfn1+z8Kg18ZZFxsrflyJNSZWXY3KTEZDkOVTk3DrcpEHM2I1/nwDziWeYZMwgg5X3i7JF+CPL/CaaqnEGAf1sDL6Ym0pxu3YnQvJHIaXwDXiHKmaLwx88GWye2AtXmM/1PwQfAag18ZZFxsrfFQRTQg1Qz1Bsq+4FytlE1j8BqKRjeRUOUzwCUlzmNrOVd4cjsjZBWz1R4WalhmjMhkPRjEXH52uxhpPdII6lqkTe3KALTTmkJxySuyuWh3sjy/wmmqpxBmF9B4gUjchiPFK05csjrHyS+y3WIrgMxqHe0LYURydZfok7hsiyXpuoNfGWRcbK3/4ndrcguBFsiVblzfGmBcI9Imyz4w6NGEp+eaQ/bo0WZjySmeLaPsoMHZNkdaymPX8edvUP4ccEa+j9RwRAM83/HNN5W3do94LF9nAZbW1Ml6r3CSjbOX4+FuXQiofxf4i3VUeawOTkrE4hkseJlr1lvFFOl+mP7PaHZPSlN8aT7SG9QEL7s9E77yCI4vDW4S+595hQ5cfi/8Qp1S2I2UBEmi7s8XjtDE7gS1r63R5DAu2Cm0Qp78nKv0zCfTayifL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk92f7CJyEln5Ojh2G/WoxrDy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJMBae7F9e/L2YP53DmumVal3z1d3inx7vzy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPC3aeCWsab8TE+uVqwwM28ayVSuQ4vRAPR8WdJFTO+nSY2/TYeUf1ykgO3j/HyGd1z6RQbUJEjH6nCVTc3M8USqDXxlkXGyt/jWBp/Wq2EL3j0HmvhRi0+JOezvosXp2L7nDoPIfO6cvp3I5i7aEg4w9vTzlT0czHlLtWFFFLAuPGoM0GWbfn9ln9JahpkI1nj6V7oaPPsU1ujWqee8sUAb7TfrcgcZ7XAhgFepJXW0ZrgHTNiKjwkRtVIfZAaxOImpZsQwb0+srpYUQZ2Hk/seGPF6pWKLSvSgxLdGV0LwtA075UKDQ6lGnkhHOWLnde/3bzWigGMNkiy5SHYswRMpVSOVPa+hxq0//yLJZNFE09Z2VwlPbyNBUpe48G8Uif+LZg0n7IakNOAj6CwPGpVv9281ooBjDZsR6DJqCUVypwc2UXDo+z9QfdJFw+fk35QctJ63YbONwH9bAy+mJtKZWyflHzuuY5BirwsO+3oug0Xf4rZOEuMnwDziWeYZMxnQA9Bc3p4/Scckrsrlod7I8v8JpqqcQZhfQeIFI3IYjxStOXLI6x8Qo5We0LU/XuPjgQdyZZwu4Hgowb2FukwZjySmeLaPsoMHZNkdaymPYUpKESyg+vQddjWUPwzqneIk/350jaeX9z0JJUew4U+uiQpG6ujY5s5AM09dgSnXnPis7cGEN7FRN7coAtNOaTV4cqecEQZ52DUy0bAGUzItuoKi9MTT9iEh99ZOx+TGIV4+QItDQMg3q9tvrw6O29E3tygC005pGgLnMoJSJnyqDXxlkXGyt9N10wk9JOFq6Kg6ef+jn554mOv8wBomL67YSnN0T/tJmXf8k5ctsyCWrgR1wViO5B6KJwYfaUHKD4wy5xLR5PYm8bRaLOOqhPiN7L9OTBPDSqiwbt8jjHaBHEyQ8fesx2ioOnn/o5+eeJjr/MAaJi+HcyVsiEUadQSNujLFNzqC+yZI7daIn0os8TuxAbbvigdzJWyIRRp1DeIadbtlqTb35H5T6aQBqpHVLs+GwZ//YvT57DOcAVqbS14nIbyTfDa6L2bXuXCN6g18ZZFxsrf1S3+/aM4X15vtN+tyBxntRA6j8HaVmif1sQYO1fcpeu/EVQ1L9Q85GQOUT7p/Z+uthxzW1vQl1DmoETK2hidRk3mPOZwD+gIzwhKox0mUQJkkdwzuPpdCcdyoumojgb9DUBF9QCbWRsvufeYUOXH4h50eV6HjIfN4Pegtv9cRAp6SFhGbR23UC8HEVEKPmLf0Meym+qb24tIDrLKTtzWVLPE7sQG274o23Q2WICsRes94PgCmNLgmU58cFTWg8C+1sQYO1fcpeu/EVQ1L9Q85PjOk087liBZwEnS7zKqAd0qosG7fI4x2t2zvhdmk0B6V8tzyRa4W0QmQGT0Wk5p9C8HEVEKPmLfJIRI5vx5XOI1Os+qASClLdN+9hMV9g88i9PnsM5wBWqTaQ9m61ELm7S70PPs/Ll2i9PnsM5wBWqTaQ9m61ELm5JfeLpM/lYD8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTxaWxJ2NwpLdZypPjEXZXGPL/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk3DfTVTJaMWX6iOMcDwrlMvVguiwp5cHh/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk7ZzqBBzETjaAVyxY3iNSEs0e8e2FRjmWI5wsN366cbVraeDysdKVF2kab8tyNYGPyfYmJTxiaHl/mX464GuAKc+/8gGLek9mkt3qWvzTXgqSWXO1VYueuO8X+mIO/UwK9qJJfozAccGT1YYQu89oLTau0999S+iSxop3chTVXMBZ8GRu+sv6Z9xYL5f0eHOqK8WqsL2Hz/7aSPC5XbcoPwt3RFoJP9wkAPjnNTabYevUWPn5y6uxfw9TfXfn1+z8Kg18ZZFxsrflyJNSZWXY3KTEZDkOVTk3DrcpEHM2I1/nwDziWeYZMwgg5X3i7JF+CPL/CaaqnEGAf1sDL6Ym0r67pZhSX17SHgypQCv3vHyIyhBMhl8JNp3JjemjG0NjE9Z2VwlPbyN/RR3NYigAxx8wTOlwT5BINjkSAJxCp6rqDXxlkXGyt8VBFNCDVDPUP0M+UGvyt0Zj44EHcmWcLvwXT4A2AnSw+krllJtcq4cibWHIFPZElCKPVGY51VV1o37qMTokd4LD//YU7iEetkqmPBnHCNKcrRZVS0A5l+eYk+ciHfVdO6nC3EK7+Fb/MbXe09SFZZkXXFL/tGDKxD89FXxiUvhUmDUy0bAGUzItlnOaLA8gPMi0xnBqhv/UFiPz05ALOHY8F0+ANgJ0sMgejfQK7nsB94cP9e35gy3/xN9W8GBMQyb0dcNAokWN34RaLTzCg1VniT7W7rKqudiT5yId9V07vLDnoQtds5MMWoMMEapAuY++RUutOnuTxN+SaA+RyWXKL4gPJzxZesd6FVy/VZuS+0iw9iakuBzbSKp3ktAkWAvufeYUOXH4sLCIxa0aOLzg4rppOdra6zkm5hGW3qMcm9EOYGlmaMJs8TuxAbbvigPWlYPQNmfJTVSL35l37IkAlvd8DrMGZusUdwpYNO+f/+o6hWtmGM88v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTW8G+UaBphGU6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcgdy80NjsdwaM/Rtmhlh9QI6JGj2Nee9Q/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJNySskmwaJUcqm5ISuvYuJUJjM5EW9x6s8/G8MS9PnKJPwDt87oUwnhfvpCk4VcQLMSNWNrcAyGzv5l+OuBrgCnDwbn6gg9H1g0io35VsxJ9WD1sf0QqXLIO95IiZfXcDRf7GSoCDOSwZciTUmVl2NyqVPvVDE1+0Nklm0yLGFEkHLkwrR+v8SSs8TuxAbbvig/AaikY3kVDn769vJBLH3fjcaRRWWlkpR+iTuGyLJem6g18ZZFxsrfFQRTQg1Qz1A+Mh/JVUGIbViPz05ALOHYUzwCUlzmNrOVd4cjsjZBWz1R4WalhmjMLB/wUPYIRh5z4rO3BhDexUTe3KALTTmkJxySuyuWh3sjy/wmmqpxBmF9B4gUjchiPFK05csjrHyA6BCNA34JfVSW1B46GEvMgeCjBvYW6TBmPJKZ4to+ygwdk2R1rKY9rcDdB8fMKCuWXSeXODUEVoiT/fnSNp5f3PQklR7DhT66JCkbq6NjmyJQ7s7ixE1Dc+KztwYQ3sVE3tygC005pNXhyp5wRBnnYNTLRsAZTMhGqhBrmBznHoSH31k7H5MYHxQr17pO3Gzer22+vDo7b0Te3KALTTmkYHkQ+ywxYp8Tm0pPe/4M6nCAjfd7xQL2s8TuxAbbvijBi4pcjYi4wkkJ4Yxl+gwIKm0doPtSltdTTk1xswySFMrPQW9wv2ebiJP9+dI2nl/BTpSqg6TMKHF6NIRq8JvwM6LBEk0NA+ly0K4zdmUV7vXz8dQ2bzyFDV5fLgsPbb7TfvYTFfYPPIFjjDuE8yJrWW/4dBdYxiIqbR2g+1KW11NOTXGzDJIUliUd8H/OpnNQctJ63YbONyqiwbt8jjHaczafRrMGv6EnBGffsI2SR+G/UqP5ZSRagWOMO4TzImtZb/h0F1jGIpgbWnLWx/bO8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3Z/sInISWfnORTQOSZQ9af/B8PknsyJvAvSQSN0gihfQ57pjagUkkTxStOXLI6x8oyWa2Iw8GMxUltQeOhhLzEvJvOngtzPz3PQklR7DhT4XlO9ypc4G/TqqyfQhfd5RfAfBCy+Ha6Xc9CSVHsOFPiggprp1pzOUOqrJ9CF93lHKozpNDeqVLnK6S8nT52Gw8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCTOfYJ/rCQNiZEfwOqUUUJloUkXSGwKudVVE8Ebn6RXJynRi6WSalTmzMlfuRRpczm8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT3WDiswWyrEe/q5DVtD5XU/mD7dVSTCwEo/ooX7TTzaae3f/94nn6mGsfbEm4KgCUSRL6TBLGB8CxG8gTR1hwNigqZVyAs0jF/n0xr1ojJqTnKegXN/1nkPVHwEGHekIjwFgsHfuuaTAnenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvqrDqFtGrZmhPwGopGN5FQ7+xVfWHEepO7Y1/USzen0gu98wr8b9aEQHVKsG75GdKkLtKRtVRiqeiW3QJarOahjMxCQBz9dzu8WLAnrKFIAKmZD76Wf40+ZAG/EfEl/qkEGZftECsE+Iq4j0S+aVfp5Lek8xFmzmIlJTuU3JkJFIfwGtZARwlNkVBFNCDVDPUIbulSkxHOO0IvyDxlgqBzbjbP1PE3yMXz3L9eNYRTOMMQyxxx8ClY2kf6Jhc3anltlzSGBpetPsi6RLPDkLTF+N51rtCk3uP6JojZ50H8S0WDiA6bJiA7/4aIi/A+pRzn7e4xvVnKJTmOQCVyLExfkO5kh72uncVwCrOM60P1E43cvZs/pdu99RgprYb7ScV9NbG1bkVCvcsOW9w8BUFblrS1TXObGJTgmIFG0SQTghG3y9fwy8xpW+qsQgC2kTKzI6FHp5AgQVo8DxcgTS24wpoifs1g0sYtjX8CS6wl+wqORYhzctgv5VOR7IaAU8nJ7d//3iefqYax9sSbgqAJRvxOJpxKvc/1vjy1hycHHbKCplXICzSMX+fTGvWiMmpOcp6Bc3/WeQ4R07VhoSEEv6hlhPJZpcHCd6ekNIuEEQdyBsTm1jDkXOi4moCnkAQC9DQhuHiJm+YyuDuKHW/mTDdRsRfG1bWhRjVvRan2GsYlUgMXwVHfhYcruwXrqAcAkNgHZGapfQcHxRN4xA7utplZGKAkcBMRa4jI48uxgko1FMVEi/wYbN0mkgwGM+1Q/IYWiIqjyhXlB9PcWZIklyA8lDag+Gg2XQozfpEWWQfVu30zj8EX3nRtsmIhkLd+8XFxMTF5ftuvwnyhLxolu9Bz92p984IV4eOBK7vhtvwxXRPxIwFailDUjT2Ykae3CBv8M7nxhzCU8rf8mdmO+yp8vU4+WvrZljO7IO5vaSLad8u35k2XXFUlVUTWKaM+QScWujNYFnddjWUPwzqneclqFbMFRCimOhRvMZHLkaPWSA7yLFqU3yVgdEyxOfvixFxpn4DsyzKRj1cCAZUVknFfRZAXkKu8T8DcAotGDshYqEwCBQ3Koky15w/MTbiz7fBSngAeVpmkFWFrOe10MVdf0sP8GLr5eDyIelXCim0+MWElIggdoi/IPGWCoHNuNs/U8TfIxfPcv141hFM4yWNTWi08yegqR/omFzdqeW2XNIYGl60+yLpEs8OQtMXyjtcPPVw7bUZE03TzDMaqRYOIDpsmIDv/hoiL8D6lHOMZaJukqSckHL8ElX1S2IiU1KwQL72mw8U3OeAaB0Udie3f/94nn6mGsfbEm4KgCUvx5mmeBW9IRb48tYcnBx2ygqZVyAs0jF/n0xr1ojJqTnKegXN/1nkDC/ekOWoPEwGYXUxK3UkN0nenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvpyeRijwt/wt50bbJiIZC3fvFxcTExeX7br8J8oS8aJbvslryu//ChJeHjgSu74bb8MV0T8SMBWopQ1I09mJGnuL8R+SGuh6Lv6QJzD/XShLsqfL1OPlr62ZYzuyDub2ki2nfLt+ZNl1xVJVVE1imjMjmBZWthnmsJZdJ5c4NQRWnJahWzBUQopjoUbzGRy5Gj1kgO8ixalNvfc2exSR+1YsRcaZ+A7MsykY9XAgGVFZJxX0WQF5CrusgSyqxjZj+4WKhMAgUNyqJMtecPzE24s+3wUp4AHlaZpBVhazntdDFXX9LD/Bi69+iy7Nc6mXuNPjFhJSIIHaIvyDxlgqBzbjbP1PE3yMXz3L9eNYRTOMewr1t39QQ/6kf6Jhc3anltlzSGBpetPsi6RLPDkLTF/kNgsJPS9kLI16M+ScCbWLWDiA6bJiA7/4aIi/A+pRzjGWibpKknJBy/BJV9UtiInfciL8XOTiydWYYYKPNgs1E/ZeNlEoL6/WUtto+kmW+d3L2bP6XbvfUYKa2G+0nFcC1Vz0HtXCrLDlvcPAVBW5a0tU1zmxiU4JiBRtEkE4IbuqlcoKdghmEWjR2ks/Qu5zy9ZY4pGLVqPA8XIE0tuMKaIn7NYNLGIL5ZgXVjx77GtnWDGfJZnXGaSFRmu4bnh+lEs+bXF73BGJDVIolLY2nt3//eJ5+phrH2xJuCoAlJ0JoNzlideh4JqNUH0ax5QoKmVcgLNIxf59Ma9aIyak5ynoFzf9Z5BJKkXIC1vaib6G+J+T6yR9J3p6Q0i4QRB3IGxObWMORc6LiagKeQBAL0NCG4eImb7Q9Iz6BwHdItD6SFeltyPgmzfyKTkjxb66j/DkQn3raTe9ir/IdUYnQgfeht6B/8juQVtFoE/6hGXmK7xcbFXjNgG8aKR6EU7ynfyowpB3fWW2UnZi5pcc656fPX95n6U4vLA4sY8nIClRennIJyfmdIMKBdj+g1C7ZNdaujmE8vVeRl6QOREF5c53VVWpRXBblxhN7uaZ/GjuX+MdfH2dFGNW9FqfYaxiVSAxfBUd+MYDvtmSv6JyAAgQ2rsYQDNwfFE3jEDu62mVkYoCRwEx7a5p0CvexHGIXFDrlna7nlAE1hMdrIRLD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDAqplN3cVEzWI8Fr57XLiYi8jKhI7hEwpOvnqAzq55s66j/DkQn3raTe9ir/IdUYnQgfeht6B/8gyT482ArlQ0GXmK7xcbFXjNgG8aKR6EU7ynfyowpB3fWW2UnZi5pccCzwbr5ouFEM4vLA4sY8nIClRennIJyfmdIMKBdj+g1C7ZNdaujmE8vVeRl6QOREF5c53VVWpRXBblxhN7uaZ/OVsM5W+dxjTFGNW9FqfYaxiVSAxfBUd+GgxvOX2bQ3BAAgQ2rsYQDNwfFE3jEDu62mVkYoCRwEx7a5p0CvexHFwOToL2navpf5h0Aqb1inbD8hhaIiqPKFeUH09xZkiSXIDyUNqD4aDAqplN3cVEzWI8Fr57XLiYj8BqKRjeRUOMcbuefjHIy2e3f/94nn6mGsfbEm4KgCUnQmg3OWJ16FVcVFIG5VOrygqZVyAs0jF/n0xr1ojJqTnKegXN/1nkC+4TwZHXtxf74I9e3WKMIknenpDSLhBEHcgbE5tYw5FzouJqAp5AEAvQ0Ibh4iZvtD0jPoHAd0iqORYhzctgv6snuJ8cdyYPCL8g8ZYKgc242z9TxN8jF89y/XjWEUzjJwGMn9cA5BxpH+iYXN2p5bZc0hgaXrT7IukSzw5C0xftvUWbRQzGpTFytmgscVIeofzrR89AP+/+GiIvwPqUc4xlom6SpJyQcvwSVfVLYiJy+RZzUu5Uqpn5CTe8uxjXLORbtp68Tr3A9dE52dTkJZZU5NGj2O4tGOhRvMZHLkaPWSA7yLFqU2P+zQZFzTvOyxFxpn4DsyzKRj1cCAZUVknFfRZAXkKu1si0cTxM1v6XBiDcCxLj9qk0l8wp5aSyD7fBSngAeVpmkFWFrOe10MVdf0sP8GLr0W1/kraY6inwSAbVKu+WLTXnf1lW33QV6eWBGo/tZLb+HHWkys7uwgWNo0Wigo337qP8ORCfetpN72Kv8h1RidCB96G3oH/yFNGVH40JWF2ZeYrvFxsVeM2AbxopHoRTvKd/KjCkHd9515rbKRGMXiqfSiSNkUrNmxy+MXltnCpKVF6ecgnJ+Z0gwoF2P6DULtk11q6OYTyskWDAfl5Q0j31b1qz7eRCCtLfyNBEnlG94APv36K8aazJxUy2AnSkd3L2bP6XbvfUYKa2G+0nFcX/jJPpRiAObDlvcPAVBW5a0tU1zmxiU4JiBRtEkE4IVXM/XnFL3XnFTITrSFGIO8zhYFPBfwvZqPA8XIE0tuMKaIn7NYNLGIL5ZgXVjx77JeHLXwK7n9Vggz7lcQ+wKLfYMfb0t7NpSxNFldc1k8y6dsVEcbCcQmSQOM6YKUvFllTk0aPY7i0Y6FG8xkcuRo9ZIDvIsWpTQilUt9/eo6MLEXGmfgOzLMpGPVwIBlRWScV9FkBeQq7MFhDBms4zUyZFMcuPokF9ISwiggU7lMmPt8FKeAB5WmaQVYWs57XQxV1/Sw/wYuvUqRL9JIgy+8QyQZBwQXoHSkFb2NrxNkooPq8dYvXBDgwtWBYl0SQyO8XFxMTF5ftuvwnyhLxolvQR6L1lwZ2U14eOBK7vhtvwxXRPxIwFailDUjT2Ykae/QrsB8XXwX8kOD3u1GlSyKKeSPmhfDv0ZljO7IO5vaSLad8u35k2XXFUlVUTWKaMwhF2ceu/1WGUH1QSdhfNqSnG/y4VKCNj2zchFs+323y5Tmu6uudbGW/nRZXo0nfqez2j1/VWjKf3cvZs/pdu99RgprYb7ScVxeFU7OinkijsOW9w8BUFblrS1TXObGJTgmIFG0SQTgh7PTCLShGAhUvvfYSdCeicTI6FHp5AgQVo8DxcgTS24wpoifs1g0sYh+w9KTakyfBFEB+jvEgReFWpWmLDQU+wp7d//3iefqYax9sSbgqAJR2A5SrKOmP4e67v/WYzPlPKCplXICzSMX+fTGvWiMmpOcp6Bc3/WeQ8wqA+6pYlEICnc/whay4hCd6ekNIuEEQdyBsTm1jDkUSm8uJmjX3PBM3fs/sBgyj0BiPpbsi2bqoaUDFpgVI9je9ir/IdUYnQgfeht6B/8goSDTPO1n0+WXmK7xcbFXjNgG8aKR6EU7ynfyowpB3fYFuYkPkhESn2obei4ROJO44vLA4sY8nIClRennIJyfmdIMKBdj+g1Dm6n85lBOtfwwdk2R1rKY9QZ5MnWTLhsnvFxcTExeX7br8J8oS8aJbOaqRM6VImoteHjgSu74bb8MV0T8SMBWopQ1I09mJGnuW8WjX274zJ+ukG3oKaduJNQn3c57EXW6ZYzuyDub2ki2nfLt+ZNl18ssgR/LIf8SIJ+VFi0eGOlbwMDv6LuM+tjX9RLN6fSC73zCvxv1oRAdUqwbvkZ0qs54kCpWz2iFwEU0yBqKU7czEJAHP13O7xYsCesoUgApE3Q7nAG7fs6ip8R4HKNTsQZl+0QKwT4iriPRL5pV+nrg+8x841apwxDOnbRINvwNxguPqG4CKq1BBajxn9izjY6FG8xkcuRo9ZIDvIsWpTWAdDXfkegtSLEXGmfgOzLMpGPVwIBlRWScV9FkBeQq74OUyJKvpxCljQd0O6TeIr8fLpL/P9hSAPt8FKeAB5WmaQVYWs57XQxY0ENmV2aTGtlnOaLA8gPPJnVgyMW1c0xRjVvRan2GsYlUgMXwVHfga8UvkI7qTcAAIENq7GEAzcHxRN4xA7utplZGKAkcBMeEGffWUumAmxb8HhiKV17iR8queASAYvA/IYWiIqjyhXlB9PcWZIkm2/EZjdJpceuTjfgXGuW/L2yooR3rR3bEU6QX0zYZX/ze9ir/IdUYnQgfeht6B/8jsXWFYD79hYWXmK7xcbFXjNgG8aKR6EU7ynfyowpB3fVd3K4lvEFUdI3WNEChNgWE4vLA4sY8nIClRennIJyfmdIMKBdj+g1DjMCCJDBx2Wyj9qJndmR6S/KmTZPpfbagUY1b0Wp9hrGJVIDF8FR34Xepgnw8ATKMACBDauxhAM3B8UTeMQO7raZWRigJHATEWuIyOPLsYJOrWiJ61vLihtrsZJ1ubFZ0PyGFoiKo8oV5QfT3FmSJJcgPJQ2oPhoNl0KM36RFlkP5p6pw8ruA06bFxQGIZ89G2Nf1Es3p9ILvfMK/G/WhEB1SrBu+RnSoqzlliDJYXunARTTIGopTtzMQkAc/Xc7vFiwJ6yhSACodGXQrtK92Te9fiGoVgtUfLyclcgJ/T+KuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSKicFLtRGYDoNw+lzy19SQq6j/DkQn3raTe9ir/IdUYnQgfeht6B/8ghXvyWOD/0eGXmK7xcbFXjNgG8aKR6EU7ynfyowpB3fduigANTI3CtqKnxHgco1Oy+AvgBoStECylRennIJyfmdIMKBdj+g1C7ZNdaujmE8ljW0R6SfOtn/CYBED0ltRFZU5NGj2O4tGOhRvMZHLkaPWSA7yLFqU0jovkm4yKW5SxFxpn4DsyzKRj1cCAZUVknFfRZAXkKu1A1JrtMy9IOhYqEwCBQ3Koky15w/MTbiz7fBSngAeVpmkFWFrOe10MVdf0sP8GLr7+EEKKVMADIoKwvSUtJnWbWUtto+kmW+d3L2bP6XbvfUYKa2G+0nFeZjNF+49nkJLDlvcPAVBW5a0tU1zmxiU4JiBRtEkE4IT0p3Gw+Zu9AEATw4DETZKur2j1pVYmbZKPA8XIE0tuMKaIn7NYNLGIL5ZgXVjx77JeHLXwK7n9Vggz7lcQ+wKIgqM2eF+wkgpkLg62wnfIEoXgjHbV5iEO2Nf1Es3p9ILvfMK/G/WhEB1SrBu+RnSr7InfBnEI+WXARTTIGopTtzMQkAc/Xc7vFiwJ6yhSACryvD7K5JQ1TwFgsHfuuaTBBmX7RArBPiKuI9EvmlX6eS3pPMRZs5iJSU7lNyZCRSKembJ8RnIRAfVB9pA0HQXs7LFBnXdjbxxJXXuZsCxiU2kTBR+ETmI7dy9mz+l2731GCmthvtJxXXNYeT1bckhaw5b3DwFQVuWtLVNc5sYlOCYgUbRJBOCE9KdxsPmbvQBWRrqI2WlRFq9o9aVWJm2SjwPFyBNLbjCmiJ+zWDSxiC+WYF1Y8e+yXhy18Cu5/VYIM+5XEPsCiIKjNnhfsJIKZC4OtsJ3yBN2R+vkuI8RREpqvazg/7vIsuz6XhOjIDoTkHZ7hGiLD8tbuCI8byk7y/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPy/9mX4ssQk/L/2ZfiyxCT8v/Zl+LLEJPGxkGe0pm8RZxz38vshk4xKN+o8Y3BzwtEVRlw+CYWvdcB9u/qWYJQH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LuByd/PverQFaqS53zBtL8hnLXdIfXO1vNpQQWf5HvYU+eoa6rFNJu/QSH2YZFW3xFeE6ZypoaFfbWmxzHlS9XPhY+xAPB4d3kggVfaYiee279akWKpg6U/OZcmWYYs/E/c7CircjkIvSx1r+VLCLlIT9fNhJ9h0/VvRIhX62s/ofpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwv0jlKl6nOCHbCOjqeEmbrf5w8x7FCxIEFBZzTaPe77adLl4hH35McanPyYcPjMVpuCeBlNilgh9qOyIH1G2GqOuhNGKbIeqW0ym7Zaruv4MSqMOvQjEZxU8Y7e1CufhUAynnyV3bs0mq6lw5RRYKNd3Jnmbctg7GekjEo6w0GvcWtES93EBEy0E35JoD5HJZeuOTBnkKfyaJ4txg4dyQbFSBAjOODOs0uDEjmNBHtvdqkKd4lwG18cjurekoIcRxhp35Zthlj87WgxwPOa+bCZxW8Oc8L0MvfAWCwd+65pMMBYLB37rmkwyr55SjUCQwqUzsVX+qjJ2cFhRLHtr5z2OGdD8dBHJYT6nY9cDso9N8BYLB37rmkwyr55SjUCQwqUzsVX+qjJ2cFhRLHtr5z2lyJNSZWXY3KkGqMpcrzT6MBYLB37rmkwyr55SjUCQwqUzsVX+qjJ2cFhRLHtr5z2lyJNSZWXY3IyB2pThxVbcsBYLB37rmkwyr55SjUCQwqUzsVX+qjJ2cFhRLHtr5z2lMrT3GRkm/XmOMr5Uy4JkMBYLB37rmkwyr55SjUCQwqUzsVX+qjJ2cFhRLHtr5z26RuI18FLTojxGTNAT9OPCCPL/CaaqnEGEtRfj9IyqtXDHdoXX4sTncBYLB37rmkwnbRqRLVzwSvBH6ab6nFM+gGrw5g00TiREtRfj9IyqtVbvUphMl/AaMBYLB37rmkwnbRqRLVzwSue89mzNgf3y05Bkibv7OvYwuDhMsVKUw8B/WwMvpibSmVsn5R87rmOwFgsHfuuaTBhujk21+NMk8lQhwwd/5HsD7DkI+4jM/Jr0IpCVjxOwjbhfUs2/G3PK4sj6dWoY4ZRx8k0NEWRjFCCcmaBVJKejfuoxOiR3gsP/9hTuIR62cBYLB37rmkwdQbDXgsLRtkl6D6ITEIyuQGrw5g00TiR3PQklR7DhT7/wrOkJ1lLo8BYLB37rmkwWOQXn4xhYDq5DrFj2qvbOSiZ8hj5jclm4cMmgMS30D349dKirrGTNpWGqyKWUCdSVyOnTVFld0PAWCwd+65pMEwiL+7bR3NuEWsoLROZ2jlYggAh2zYxKrOm4GNjZXJtBbapp/JRLtKLtOqSsYaxGf/B8PknsyJvFhCPWhSUC5nuuHQnwW3g1UaaNVc4GpZaHOti4yAQJxl1BsNeCwtG2SXoPohMQjK5AavDmDTROJEInsuVUa9SWnENawMGez8UwFgsHfuuaTBY5BefjGFgOrkOsWPaq9s5KJnyGPmNyWbhwyaAxLfQPeNmm5Lr1p2pYhJ8WOeA6efPPNjzPIH+K8BYLB37rmkwTCIv7ttHc24RaygtE5naOViCACHbNjEqs6bgY2Nlcm2gOdmIOZ5ujGV+ciC9trJaTddMJPSThauioOnn/o5+eWst6CpWA+sFyr55SjUCQwqUzsVX+qjJ2cFhRLHtr5z2HF34gAZl5q3pCgYVS10eex2DWy5n0Tr//GAxA/UaCRbAWCwd+65pMMBYLB37rmkwcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/yW20jIkTGnjAWCwd+65pMMBYLB37rmkwcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr//AuEAaXgkojAWCwd+65pMMBYLB37rmkwcV9sX9MGuKLNzaJy93Vs0f4EvhrV3uedHEcuJ+RvSwZzysUlAo8iA8T2P1AbHH2oTr25ZjJjJtDAWCwd+65pMO8sFERkGzIprD1oOhUnp8jqbdmcoQYqPHPT6yNUvnsS4cMmgMS30D11ZMnUofCOetRgt+Jt54RjwFgsHfuuaTDAWCwd+65pMI9onXBLEFsazc2icvd1bNEX87yzrgNS8rqZpHRFaSxbbUXfYiX6zhQrldI+4X6yN8BYLB37rmkwwFgsHfuuaTBY5BefjGFgOnHO1gemEq8464RU5Vx7mf/DUgxQnnMPO3ta4ysjEri7TXGGAda61w4uc92gsVwEKrCOjqeEmbrfNg0ZOIlCNdkv94TlSlGhCUZ6CCfYNpaWND5/1YD7AQ8v94TlSlGhCaCqNBkpBYoKCnCHVKTy5iWvK9NWInNX9lrgSNBvfq0OZf11sV/DEVQk8dpOFQBeYk1xhgHWutcO5V4HH/RrsN/5mIpPSMlFC7rQ6zrLR5iG8IuW/pqHZ5TNzaJy93Vs0dq8V3PemZsXb/HBCwSJLTgGJVGYi5tDsYF7kKGW2QSaS8uHYtzf8Vz2aEsqrG9ztDC7LZ9mNvu1aSZkpnEYQsSN7SdIsYVmbZnQHPSEFy5P50r/6zZg8QnWE0GVhbVM/V7SWiKSZw/opWqh0Oh2IWXnSv/rNmDxCdmvG2ivsk7ANcLAKWIy4N3VmaIohTeKhyUGtg9pP9WQ7GNtU97kTE2caiSB0pwUU7rQ6zrLR5iG4VQLknJoeu+sPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPRSI6dQzrfsnM0oR3xn/Tt39dttIfq43CQFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHQW6A1k/HcyMpulwKMYH5DTA7z0L52nuKIIvT+UNORMRBboDWT8dzI+lwCf/Z0pA7PB33uCU9gsmdGlESu52O3qWv15BBneM3HEcuJ+RvSwaFVSD1FKcXtAm9N2DYKM5rYhx5Xg+Lo7UwO89C+dp7igIuZ8gz9RNAu5lZm9vkE5bsY21T3uRMTZxqJIHSnBRTWuAyj2zpk33ZdQdps8ZOyaw9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9FIjp1DOt+yehog3BwCaDFP1220h+rjcJAWDQJ3KBpIOSxWonF3FK3Ci+G04JfRlAVFYclhD8d4dBboDWT8dzI8Ytn2qOlhtCMDvPQvnae4ogi9P5Q05ExEFugNZPx3MjPl7b1kKTcjcwO89C+dp7iiCL0/lDTkTEQW6A1k/HcyOrwnWqSnx4BTA7z0L52nuKIIvT+UNORMRBboDWT8dzI249uZkj+imSMDvPQvnae4qf1Ly4rVHjsBSI6dQzrfsn5zknYQn7uwxhQTeBFZDdTJKHozjh0OSjuZimT2kQX2DC4OEyxUpTD+dK/+s2YPEJEyP9IEfQo8sSNujLFNzqC7BPxf+hfE2VrD1oOhUnp8jqbdmcoQYqPChyjXziGgkswuDhMsVKUw/nSv/rNmDxCRMj/SBH0KPLN4hp1u2WpNvfkflPppAGqv3+YEl8JkNJ1ZmiKIU3iofXJiGKkpvauexjbVPe5ExNnGokgdKcFFPJ4IcbYEn/3apTfN5kPhN94Pegtv9cRAqKBrJedLKNZ6P33I5QEiCsHEcuJ+RvSwaFVSD1FKcXtMb2a3wBSeOcYo/+mITiCbZvtN+tyBxntT3NCN+vBqM41ZmiKIU3iocyEUlkw8Uh8ViCACHbNjEq8kyiJFHAjB3u0V+ntFmUQQyUaO8yXW5oPeD4ApjS4JkgL2XrZ568zFMzMTd2VbLAK+TC2YUt5PYGTYJMLu508r8RVDUv1Dzk+M6TTzuWIFluVZtPPGIBbjaxjIxorNUKHEcuJ+RvSwaFVSD1FKcXtMb2a3wBSeOc3bO+F2aTQHpXy3PJFrhbRPnbJj3hpKE7MZPML60V2LXsY21T3uRMTZxqJIHSnBRTyeCHG2BJ/91K7b3LNGkdrPjHhtwRYHNqUzZu75YUdPXgUDNHAWdCnMLg4TLFSlMP50r/6zZg8Qm/IGnoILIe5l3nN8rZ3/VpPc0I368GozilaqHQ6HYhZedK/+s2YPEJvyBp6CCyHuaORbBg3WAZBPSjPdZPbMmLnDpjVDYkKfnCwiMWtGji80vSSgvhGij84cMmgMS30D0UiOnUM637J2YR3kJe1z5ocX0eIVKkqev0iedigBlo5J4r/tYjUq1/D1pWD0DZnyWo57aXAJSa/mvQikJWPE7CK+TC2YUt5Pa95VW5FbVyOfXz8dQ2bzyF3tajWYqEMiB1YKbw3tpRShxHLifkb0sGhVUg9RSnF7TG9mt8AUnjnONgJkNg8W1AsxT3i2+x4ivCCD8Qa/jQUE5Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCcvOTLNv2L85MriQusSU8tUyInjWJvR8WnVgpvDe2lFKHEcuJ+RvSwaFVSD1FKcXtMb2a3wBSeOcczafRrMGv6EnBGffsI2SR2O6ppjjBwmOD7DkI+4jM/Jr0IpCVjxOwivkwtmFLeT2NXETs1GlA+QUtlKIpmwMxKw9aDoVJ6fI6m3ZnKEGKjxz0+sjVL57EuHDJoDEt9A9FIjp1DOt+ycZBl+11sOVHM/fgeW7+hColM7FV/qoydkji9MrIcEZz05Bkibv7OvYwuDhMsVKUw/nSv/rNmDxCXiaDcSXtR/IO0m6H650vKIBYNAncoGkg5LFaicXcUrcKL4bTgl9GUBUVhyWEPx3h0FugNZPx3MjZbxRTpfpj+zVeA9o7RaLis3NonL3dWzRF/O8s64DUvK6maR0RWksW7aJ8/lTY3NynAnqRY0tzpnoaY6yLWGnPBPCZumaDXGV4kBOEElYdWzXZxhq9dA2Fz1kgO8ixalNmXhVc80BBXOj639AgtUFbo/ive0PzKRfycFbLWpFUOKO2O4tUEH5eooB1PBzyS/ma0RL3cQETLQTfkmgPkcllwLpRAauV7n+r/vwphgnNk1oMcDzmvmwmWA8dKC/IiZKWqTz3+mLoAi/3bzWigGMNh8gtxiLTTHiH33UrlGN3lACBGvtTONhTKg18ZZFxsrflMrT3GRkm/XmOMr5Uy4JkL5IhN3EmD7rOuzshnXKlCFrteGTdCZOu5GMZSUNb0n0PLXN2EDq885cxnIcGr//zIo9UZjnVVXWbEegyaglFcrS+DkO8fYpMRbMZAwlNQRlNXqcWlKuB7ieyZFt++6kERLUX4/SMqrVUERbWOXMtNdsR6DJqCUVyjleJwmkc0wsT1nZXCU9vI1CQ/UWBIJ97yY9EvBAEIvmouLZ+ATHA0CoNfGWRcbK3+kbiNfBS06ImACD1HOvDAa0//yLJZNFEzVfTZCdyIHMiMSlA/mF8JUFPGYARHVhHP4ndrcguBFspa8DwFyFzLyoNfGWRcbK3/4ndrcguBFsiVblzfGmBcL+J3a3ILgRbDY1jvGMqZMANV9NkJ3IgcyVhqsillAnUr/X0fW1H4DylYarIpZQJ1JC0IYX5CECerzR89UNRM5NlKbPj9+iHGnRy4dND93dh+6gnuh/ZnB5fMEzpcE+QSDl7BTXTEk6g6g18ZZFxsrflRwUrVf0HBF8daNeN21duyKwoR3vfaj6/W0Z7tf4gNyR+HmBRsGWpW72eK7kuq8fskNM1WyjJWFss32bt1w+qp7JkW377qQRCJ7LlVGvUlrTREZwfW/cdfEG3XqCiYSYela1SZ+MznOfAPOJZ5hkzNF5I7Y8f/OnlynNs5RRMG6FtNohxU2WZAnGrfRVZV1uCJ7LlVGvUlq0WVUtAOZfnqxOIZLHiZa9a+j9RwRAM839aW9Cy7WhxWDUy0bAGUzIod7QthRHJ1n1yFn65YULtj0ibLPjDo0YSn55pD9ujRZmPJKZ4to+ymvo/UcEQDPNQCinyBBLvjuh3tC2FEcnWUSbAtwNeaZdkYxlJQ1vSfQLsYsz9m1HAbPE7sQG274ou2EpzdE/7SZl3/JOXLbMghHUDJLAZU35MT65WrDAzbwJXZAhY8A6K4iT/fnSNp5fAKtuCg390GLjES9EfGyAKJis8nXcgBlZsrgO018QId/moETK2hidRm/xwQsEiS04oUyD8zKG9dvuqzrUUL6jA/keQdkGX1zJL7n3mFDlx+IvBxFRCj5i31DFSZ18At2ob7wggUCVjBkTI/0gR9CjyxI26MsU3OoL7Jkjt1oifSizxO7EBtu+KB3MlbIhFGnUN4hp1u2WpNvfkflPppAGqj01XPCuGRyBQS23IkbDemdbsxZACixvadcsbK8fM8aBL7n3mFDlx+IvBxFRCj5i39DHspvqm9uLJVc6h4vwlzPztvsrnUGVHL8RVDUv1DzkZA5RPun9n662HHNbW9CXUOagRMraGJ1GDJRo7zJdbmg94PgCmNLgmZu+CM6tfiadqlN83mQ+E30UdtogReyh8ag18ZZFxsrfZJHcM7j6XQnHcqLpqI4G/aAG2uqRc3sEm74Izq1+Jp2qU3zeZD4TfeD3oLb/XEQKaAbKeHAIb93moETK2hidRgyUaO8yXW5oPeD4ApjS4JlOfHBU1oPAvhMj/SBH0KPLTeY85nAP6AivvrsKqjSAqjcgfXEg9tLEwU6UqoOkzCgF0JbbjIhF9lfBhX9gmnyQm74Izq1+Jp0F0JbbjIhF9lfBhX9gmnyQv9281ooBjDbWxBg7V9yl61AyHSH9z2AQB59eXk9x5vETI/0gR9Cjy8nwQn5HMaOUAGx7KqFmVDEtYAA5kqse/gbB1x6hI2lXIBJMN1Es1hoM/zPhlXVnyb05G5IsPEHYGWmw/Pq6wg+Zq0Vq0WTlMjK4kLrElPLVxWnU73DnOiwyuJC6xJTy1YiT/fnSNp5fpIAH3GDGpAeruDnuKlgiySqY8GccI0pyq7g57ipYIsm/3bzWigGMNnLQrjN2ZRXu9fPx1DZvPIWJVuXN8aYFwlNOTXGzDJIUys9Bb3C/Z5uIk/350jaeX8FOlKqDpMwocXo0hGrwm/AzosESTQ0D6cvOTLNv2L85SQnhjGX6DAjwXT4A2AnSw+agRMraGJ1GXqGdW1doInysLYGoygqbppu+CM6tfiadrFQPSI3P+GENL87u5+sZIag18ZZFxsrf9cYajgjHtiuZ5Vyg3Slq7HX8vRGTDnO4y85Ms2/YvzkyuJC6xJTy1TotoNbS4PggqeSYoivzWC0MdPmA7qIZ8DGu6anjPS6G2SQjd+5XpjKTRBNl1SEPd8WpcfJ6DDBE3uSqnP5e2hl3/s2S3/AcnNtFH8awFvWeaDHA85r5sJlYLbd5Jmn5klAP5royjNU0zz5bVmpaSFW7YSnN0T/tJmoX7D9ZCBeyedqtiy+m99lDgidxJvFYSadTNlDuVSuBUA/mujKM1TTPPltWalpIVW/xwQsEiS04BiVRmIubQ7GBe5ChltkEmkvLh2Lc3/FcWQ6MbX8gbuSv+/CmGCc2TWgxwPOa+bCZkbmwnoS8qa0mQGT0Wk5p9NrlVRlgRSW/qDXxlkXGyt8D9bKlyQKyzQafdJWfhyeIYPWx/RCpcsg73kiJl9dwNJLm9l/kv09VrGWufpBe56ZOUV0x4upUH7/dvNaKAYw2HyC3GItNMeLyrqj8yZgXOTMG/erWsTnq8/TnSPPDjO5QDx4rh3D1S9uyBK2DNHi0sKC38YHLOwovufeYUOXH4gQE9l397Yn0VH8VxfNwLy62HHNbW9CXULlTaR50VJkMtq4pcoVZfcYCapzjWGoI3KlT71QxNftD1/WkQFWySPXhgPie2HHU4ctONaqaynxsv9281ooBjDaUyMpMFu/g+6WqYVWBnUw+mBdAEbtIgEAUcHXO09MXFMmgRuZRQteWzFBE4Cthej654wTl0gKsu2gtTHbsyiD7YNTLRsAZTMggQLozWXkxVfxQFvkEtyk6aep3wUVLBkpE3tygC005pNgq7mZpXNDCzlHt9oQ4rx6xHXReuN0pRGETpzZc2/VMAmATUzco9W+FyJUZ8qdEG7/dvNaKAYw2YROnNlzb9UzC1lf1PnuJKYLa8L52mtZQwQS/n0cCeEV3f9ioyitj+tWBWu08fNX706OvW+YNEoAuR2p43GIz8IHm83qUyivsTTib+DQieAqT2QQbTYkLPrloCWNwO1TiVOzOzyJ4+1+5U2kedFSZDGkVvHFMW6mVmCMBStr7MMxv26g2/OX//L/dvNaKAYw2EmMk3iVz5AqrkLpT0TNcFovPSv/c01Xm8CY83mAYs6T4XopKX4c+BSfQD2F7fPktahfsP1kIF7Jl+Rc4A54IbuJAThBJWHVslGl9q0T8UWhhQTeBFZDdTBI26MsU3OoLwFfzu/pgaLr0BJRgEJ4OGy3dEWgk/3CQA+Oc1Npth69RY+fnLq7F/D1N9d+fX7PwqDXxlkXGyt+XIk1JlZdjcpMRkOQ5VOTcOtykQczYjX+fAPOJZ5hkzKOUB6hiZZNBpycy7UvdI8SzxO7EBtu+KLqqcKWCb+S94QHDuhuSDzBP2AwfIhAnSifQD2F7fPktahfsP1kIF7J52q2LL6b32Zdg1818K3MVyvZhKluyThlUSO5DZHH5Riwt+ugE7hVKs8TuxAbbvihOfHBU1oPAvtmvG2ivsk7ANyB9cSD20sRSORD7oAyhb5gjAUra+zDMrUkC7LYDZCO/3bzWigGMNtgyf6f+E697xcRKDPmkby22Zoxwzadgwag18ZZFxsrfzVWgefLB9+2WAimIQhaQoC2nKiKwglp4FOhwqLeiYvCGnGZm0K9VJVpf1m+gl7py+GpcnNosxo6z8IMycnmZ5NNERnB9b9x18QbdeoKJhJh6VrVJn4zOc58A84lnmGTMay79/pMxdRsf3i5JiFZy84LQ04Y/0qyIqDXxlkXGyt+MmBmoI4SmBWFBN4EVkN1Mm74Izq1+Jp0C7YKbRCnvydEvw+OmFkBzosnzqGkBrSyx9+KGCXaa2Xc6dlD9mz9P2SQjd+5XpjICKvBmcLSfELwLWxJRj1vLV0pGt5hZIZ1Fqr4J81dRsprgHTNiKjwkRtVIfZAaxOImpZsQwb0+srpYUQZ2Hk/seGPF6pWKLSvSgxLdGV0LwtA075UKDQ6lGnkhHOWLnde/3bzWigGMNiua7IPsybiHzlHt9oQ4rx6xHXReuN0pRMdAsIJP9jW2yD440lMU6uaDRQpi9SD45Gbo3TeQ57vpgD3lzUPAEKxkMMWH4Pmee7PE7sQG274o/OTSx5nBfjrWE0GVhbVM/alT71QxNftDDy0I+VfMnMbTo69b5g0SgC5HanjcYjPwvKpMsm2TwyYx8+fSCxlRIA7l7Ruj8iMyFHB1ztPTFxR/SH/kfW8KmpPZBBtNiQs+z3a8Y6iNyHlU7M7PInj7X4oak6uU6IRX+PlPLE2KlMZp6nfBRUsGSkTe3KALTTmkWeKdmTkEiU07oKQsXwKZ9Jeq9wko2zl+T1nZXCU9vI18fWqIKGwXjHgypQCv3vHy6y3ZOsQka3ieyZFt++6kEeUXWaUTU3wN4xEvRHxsgCiYrPJ13IAZWbK4DtNfECHfBj1IlHszAVS7YSnN0T/tJmXf8k5ctsyCOWkn1mupLPsEcTJDx96zHaKg6ef+jn55NRjP9Z260P2xQlg3pveBe1Lp3kyS/YRcvcyFVQU3e6bLB19/I/LGWlyJgvIexFuBgnofOQrTPZ4+wR6lpyWnXPI/RvSbSQrZBj1IlHszAVQMlGjvMl1uaD3g+AKY0uCZuqpwpYJv5L0vBxFRCj5i39DHspvqm9uL7H2ZIUpil7WoNfGWRcbK33XgyCw2rXpGx3Ki6aiOBv3ZBLCz24cOrxMj/SBH0KPLTeY85nAP6Ag/vtvpFCnj3YNWBUbEQksWFPmTnu5pPkntjYZMeyJerdlre+IE2a1fEyP9IEfQo8tN5jzmcA/oCDAV1IQBH7KfqDXxlkXGyt914MgsNq16Rsdyoumojgb9/W4v/XdWrrHKm8UuA/SnKGKP/piE4gm2b7TfrcgcZ7Uyh4ydZdqI1WDUy0bAGUzIHcyVsiEUadSE1w9p75u9Z0v7BcKJm44OEyP9IEfQo8uE1w9p75u9ZwwIOVo+saRwZjySmeLaPsovBxFRCj5i3ypCuc76fiTIx+eOQ8PDT3hnAwBH26HYtMbNprK4LYgbQLw4iiueoOKtp4PKx0pUXVdKRreYWSGdC31lxCh4My0/G8MS9PnKJGOJKd5hF3+U9Hf01UlyyqrEE/vBiMQ/rXf+zZLf8Byc20UfxrAW9Z5oMcDzmvmwmRop3chTVXMBwsIjFrRo4vMoK39j8wc+abucsNsJ2uoUeeqtTp4HFk4K3OJbrgocAiPwbd6jtD0Ks8TuxAbbvijjo7C3kNP3INLkH4dC4si1L7n3mFDlx+KboR8KKvMtE6xlrn6QXuemiccdViuS2KCRjGUlDW9J9MjKJEPF85qP0fI81agyzrE9FnxwYF5MXeEdgCe+xNqSW/VisDTKv1qtp4PKx0pUXSey/ZCypF6BAIY3o68Oed8r6UhuhHB4P0z4vQS8JRtc06OvW+YNEoANULrWKsJVwe6+0ZjaPn9BVnQl2Y7WQOp+7yZOIOnN+Kg18ZZFxsrfbnn+2wcSbtLTo69b5g0SgJpb1tIBC0VVYNTLRsAZTMjC1gLXUG6EtUbwuwJZevVnw1rgTYtyBHxmPJKZ4to+ymyu7djU1miZq8J1qkp8eAW/3bzWigGMNk1H72YelCd04d25Ov43oRL9fWYL+PrUhag18ZZFxsrfvCI8np9xX/h8daNeN21duyKwoR3vfaj6/W0Z7tf4gNyRjGUlDW9J9OTu84fUssYtHvadyujrizdsWDY6vlOfYGY8kpni2j7KwsIjFrRo4vMELUAbq3Qw6SqY8GccI0pybNTCyHM0pfxd9zK8MJxCc2WVgzT9cOAbE35JoD5HJZc+Mh/JVUGIbRN+SaA+RyWXUHLSet2Gzjf/E31bwYExDAbB1x6hI2lX6GceRn/xG+oGwdceoSNpV7Iql4w5LYet8KJqa0NkkKBkZtQlldKqY3S2Kwp+Pvo48HCdlyZMBoD+WJMejt+5AKPzmJ8jav8gxBP7wYjEP60K3OJbrgocAiPwbd6jtD0Ks8TuxAbbvijjo7C3kNP3INLkH4dC4si1L7n3mFDlx+KboR8KKvMtE6xlrn6QXuemiccdViuS2KCRjGUlDW9J9MjKJEPF85qP0fI81agyzrE9FnxwYF5MXeEdgCe+xNqSW/VisDTKv1qJ23PmcemubjWLkJ9nQ4JLgv+r2BwWYHa/3bzWigGMNmP9xRVykDverx6WIJXkULjLoZSifzohz1/Y8go1wFv3uwcRay4Oudl0qq/ZPM64f7PE7sQG274opaphVYGdTD6vHpYgleRQuCL4/FnHICy/ZjySmeLaPsqdTLLphyYjxCz4lDkL7KOyNk/hRZZ21vQ1X02QnciBzA7DdhbnCZp3pOeZUI3kkFSoNfGWRcbK3wGOw6IbIHiyW7JZH99t+/fV4cqecEQZ57PE7sQG274oRqoQa5gc5x6Eh99ZOx+TGInbc+Zx6a5u9odk9KU3xpOHosDvcT/uYYrOej0JtLplmNyYxOvt3Dj1qhHaBp+6N4NWBUbEQksWClKigtc2o424tu7XdqAOU5u+CM6tfiadcXo0hGrwm/BjLr/hJ4BKIGY8kpni2j7KU05NcbMMkhTcJ7lo11BAUM35uz5odFtAa6wO/7pMwOpNZEMKSrudw2DUy0bAGUzIwYuKXI2IuMIyuJC6xJTy1XyvZtfJfx7FU05NcbMMkhSWJR3wf86mc1By0nrdhs43sUJYN6b3gXtzNp9Gswa/oScEZ9+wjZJHzfm7Pmh0W0BeoZ1bV2gifJP4j+nsvYWyQLw4iiueoOJUyzdbVM/TrW7omRQM+vi1FfxY8Sp+iJqEOcKpDvFtToRC/UeD9xII3hREv4iEjWv5MNVETavMkJA//4qmhneIV5CuVDAMcDq31PHUpBdxSJD9xRvzxkLcM5NKrNJrCAaWZoioH5pKq45uuMWLS5cA4VTO4xSW6/28dRUBtXEZKgyKEsl0DET5ohz+Pg21Gw+w0zB9aWHlcmao00x1enIKFJVOS/zOfjAfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LctBWUqh8ccsm2utZi+wc2cjOx7LgKysZ1ioEByRFu5q/m9ftHBTauKeUesELTuRK270nmAeVpWqKqvgwI9x/utdQxQ/1o3LCLDdI9OVRdvOOQbCAZ+BPqUbuRIJm2GvPhkdhTY1r6yGjT10NNlst5kj0ev7uhfA7+3/kXDztIdqAK8wOanajkx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PCx+mA30VTw8LH6YDfRVPDwsfpgN9FU8PC8axWoQJD0/V8wrXqzAFqTpoOtXRJq6nKxoeVOYqyZ8qAWDQJ3KBpIN3BLsxLlj0rNKAiuTcO6Pxj5hK0qFhWSu9bIqll76wTNep2m4JtoMoFA6vM2qPhqpBMzQimTdiBuaiVlEEb3Fkiyv7FCOOlfGHY0vEVzVeKfPxUuxmn4rWta6m0McaVwfrngkB1+IcwSDzcsAxjJBkS7V5fZC1CesIx4RleAtOAZBoBOmfxQ+rz5xpXs71TMPR03DvDUKeAZPc4efDTTzUhnDq8RgF5MWimZzjQEhc7Vwo8iTPXgTz1KnEtfKCz5Uh/wM+xCDWlMgrHOieNU1dQlaX9H3PCuDD8WwGiTOKV1QEo83cZQQWRvd4IpKK8l8I6iv2LelJtHwfMSIeSJj06Z5+NEcaAVkM9uQHNB2YXirPy6PIIrxXthgUfk6efO2jDDW0uDLVVyS1ZZwkYnkNW4aJtCdFqoAmQqZuTxy3jcBsxjJO0HzVnh05PBA/u5KU8bAXtrXJQtaYfRCcMoGKVUggGYQH9/4ARSuw1bMwk8KQowZpmIDFAe8hcqMYE+wubuGKVBN2duQvv76PZGY9tSdyoY6N4JKKH4/yj+If+ViI0yhOYoEBIPNywDGMkGQMHQwXOl2lGNHz0brRV14uvIhTf0r0kntd73vksJ/7u4MQLhpxmxu6L288j+CeMMDXbt5G5rFPBWDHTBgTqXIz3sjlPbKKDcLixS0fZB1znzdEspXdWi8xgt08FGkSxVbR03DvDUKeAZkQelFZ/eLjI94KHVBpBFUI6iv2LelJtOhSWVWm+TdEsNo+4wfcbnYM9uQHNB2YXirPy6PIIrxXs/44G2kt1zGjDDW0uDLVVyS1ZZwkYnkNW4aJtCdFqoAmQqZuTxy3jUQ/3xdLebc3VMu/+92bZBwk5BAT+rKygdaYfRCcMoGKmx1t7HnTjv06MWLd6UpJ7MKQowZpmIDFAe8hcqMYE+wubuGKVBN2duQvv76PZGY9clwL3R+wizaVzEWP7b63NBOltzDxZk5RIPNywDGMkGQjWwlcGOESrhgAsWbnkLLWvIhTf0r0kntd73vksJ/7u4MQLhpxmxu6L288j+CeMMCptWn9VuGbznBHgQfi3ncpMJ95Mz24b3HixS0fZB1znw66jFvtkhwp7071zLPJz7TR03DvDUKeAZkQelFZ/eLjI94KHVBpBFUI6iv2LelJtLucsNsJ2uoU1DEPau+MSXk2sEq9tJYbOFeCTK/H4ULSs/44G2kt1zFZERUgID87kL7Yq4sorIMnrTExBvUE7t4KoPidRrJqYvcUFVcuet2FguQDMG0SS+leCQMHKUbNsKVqodDodiFlDwbn6gg9H1i2jreTA/DukTAgLGi5HPbDIIvT+UNORMQ73kiJl9dwNPl0uiV+r/FjwR+mm+pxTPoBq8OYNNE4kdKDEt0ZXQvCoqKhoANAWexmAmFR3LKaecIKQH9xapKWCD6zeYF1nNeZC4OtsJ3yBJX9PO5QXUH5MCAsaLkc9sMgi9P5Q05ExKXZ7WLKC+D7u3JcPYzt4rszoeYB/Je6qqw9aDoVJ6fITuyUW/8exDg7LFBnXdjbxxJXXuZsCxiUuE89Q78DJLEBYNAncoGkg5+gA4ucyggfwx88GWye2AtKydNv6CTNi3FfbF/TBriiUzMxN3ZVssAdg1suZ9E6/1n6Cb21JXNZBjqhfL5iLWpmAmFR3LKaecIKQH9xapKWakY/FF8AzWg8tc3YQOrzzlzGchwav//MwV5kUMSlBLg/AaikY3kVDl2ntTTj/8rdnvPZszYH98tOQZIm7+zr2MLg4TLFSlMPAf1sDL6Ym0oI5S79pPi0dHJ8W3W2YQJWdWCm8N7aUUocRy4n5G9LBnPKxSUCjyIDbEegyaglFcp+4t6rXZc88slQhwwd/5HsD7DkI+4jM/Jr0IpCVjxOwh2DWy5n0Tr/SqIV4oOEBmTO2tIEHj2/xDVmJzPpVUyEKL4bTgl9GUBUVhyWEPx3h5V3hyOyNkFbd/SRbAOsi23/N2MTaHVG9xFrKC0Tmdo5WIIAIds2MSqzpuBjY2VybRUEU0INUM9Q7nxhi9heT94d23GDqg4YIyiZ8hj5jclm4cMmgMS30D2ncXb8pkNlLU7a+m9o2eVLUpScbtPXY3mLSRYue6xyQrqZpHRFaSxbbUXfYiX6zhQS1F+P0jKq1eGAd2x1OiLxi32YOSX61agxk8wvrRXYtexjbVPe5ExNCDZMI+JrJV9nQA9Bc3p4/Scckrsrlod7I8v8JpqqcQbc9CSVHsOFPvWyOETnUYxrBwiJMwJX0fwxk8wvrRXYtexjbVPe5ExNR2fVmEyqvVO2Wc5osDyA8/cgQkLzUfWBMYUzgfh5/C5OQZIm7+zr2MLg4TLFSlMPgsX2cBltbUyXqvcJKNs5flnlgC6aLpiMQSzqy9UUwd/yGyyc3dV6AZbyZVpsQEqZJeg+iExCMrmtHnTxlMad0UGWRiIb9KWh4cMmgMS30D1qRj8UXwDNaAuxizP2bUcBH4XBOP/gst/O1vv0WSUjnN096ji5zwFdcV9sX9MGuKJTMzE3dlWywB2DWy5n0Tr/hr/7NekDA/riROEB4O4qE3FfbF/TBriiUzMxN3ZVssAdg1suZ9E6/zE+uVqwwM28CV2QIWPAOisnUCoE+R7cwQFg0CdygaSDCDZMI+JrJV+jlAeoYmWTQacnMu1L3SPE6j1LicCGk6VCl6d8za38xZTOxVf6qMnZwWFEse2vnPZvI92XE7mOLV4JAwcpRs2wpWqh0Oh2IWVf2PIKNcBb9wMf5L1RVeMOlM7FV/qoydkji9MrIcEZz5lVBEjCxWaEVFYclhD8d4fZKyAna4xzwrEQsh6P9In8rD1oOhUnp8jqbdmcoQYqPHPT6yNUvnsS4cMmgMS30D11ZMnUofCOevYMAb28qXNfIGR/z632+sPVmaIohTeKh69QIF4Myn71WIIAIds2MSqzpuBjY2Vybd7fNbOXPwNdYqUN4zQ2F0vQzGX31fjqc8ReZFtDC5/JfYlKVrrtuCtCB96G3oH/yFif3L+FiXhivt0W25erGIQD9tcnMj9RLnEaxK8U960+k0aTKe+Wl6FhEABmpbOO11h/TEZfw21wDB2TZHWspj1/rmlOCs+pkY+ECzyoDEkO7GNtU97kTE2caiSB0pwUU1h/TEZfw21wDB2TZHWspj390Cr4XAixz4+ECzyoDEkO7GNtU97kTE2caiSB0pwUU5bxIJEMlI4bDB2TZHWspj1/rmlOCs+pkTGTzC+tFdi17GNtU97kTE2caiSB0pwUU5bxIJEMlI4bDB2TZHWspj390Cr4XAixzzGTzC+tFdi17GNtU97kTE2caiSB0pwUU1h/TEZfw21w2XUHabPGTsmsPWg6FSenyOpt2ZyhBio8c9PrI1S+exLhwyaAxLfQPRSI6dQzrfsn83sskUR7aCn9dttIfq43CQFg0CdygaSDksVqJxdxStwovhtOCX0ZQFRWHJYQ/HeHQW6A1k/HcyPPdrxjqI3IeTwd97glPYLJnRpRErudjt6lr9eQQZ3jNxxHLifkb0sGhVUg9RSnF7QnCfb4od+M6tv/OPjQwid7rD1oOhUnp8h3gCAXaX5vscf/QTe4OAnKl9WcS3HRv6SsPWg6FSenyHeAIBdpfm+xCb03YNgozmva5bIjtEyZNKw9aDoVJ6fId4AgF2l+b7GISx6ocjkhJy6YNHca2zaUr4ePFoHgHvhGDO5jrD3WTZwJ6kWNLc6Zpewtr2lM+p0yNyaN+ibVXOIv8vZq+ewAgOhy8YLAPDirbZZrywUVSpNuqJ+R/2A20fFnSRUzvp1e/K2OqFt23j3L9eNYRTOMK/3TS4xfaGQOoV5ciNV9Q4/ive0PzKRfRbI5MTZTA1yEF0TvcY0ReHJyfR9zMs9YDwbn6gg9H1h2jxBP15tzLkhPieK3qr606qm3XMv4wdY73kiJl9dwNF/sZKgIM5LBlyJNSZWXY3KpU+9UMTX7Q9KDEt0ZXQvCoqKhoANAWeysZa5+kF7npk5RXTHi6lQfv9281ooBjDY7LFBnXdjbxxJXXuZsCxiU2ykrhcsaIu6ZC4OtsJ3yBGDkDuspKpjAL7n3mFDlx+JZ+gm9tSVzWSa6WbzyOHvUK6xTjPn6TjyxeSmMOxMQec7HaWlsiLNgpdntYsoL4Pu7clw9jO3iu3tZfZheOnjtwx88GWye2Avyk9RXJBZObqg18ZZFxsrflMrT3GRkm/Uudhg6xCrch39AuaRQ1fBsmQuDrbCd8gSN/el7M3CuVLPE7sQG274owx88GWye2AsQqXirCFbXlb5IhN3EmD7rOuzshnXKlCFC/imLXpqQd0Te3KALTTmkK4sj6dWoY4aLQ5tkpKAu5vn7t0tzKCwwEtRfj9IyqtX+hmqpirqtsxbMZAwlNQRl7ejU3k1c0ra/3bzWigGMNmxHoMmoJRXKEJgZiWPfTEGGQ9GMRcfna4lVYToGJFJOqDXxlkXGyt8VBFNCDVDPUHn0gyjCmkiYbEegyaglFcrgsPFoE5DRmLPE7sQG274oPwGopGN5FQ50MwoMQQIOaBUEU0INUM9Qz5BUckJrI7ovufeYUOXH4qvV8ZIoYFr4bKvuBcrZRNY/AaikY3kVDmyl7wnC8iPwT1nZXCU9vI2Ww1RP2jllshSt7apcRCOKq9XxkihgWvj/HNN5W3do9wH9bAy+mJtKcrmFvgaAcBX0OvMHvDYg/E7a+m9o2eVLUzwCUlzmNrOVd4cjsjZBWzUb5x+EX7UBJj0S8EAQi+ZB1eW/EwchxULQhhfkIQJ66vwdSZBVz3uFtNohxU2WZHLkwrR+v8SSYNTLRsAZTMi2Wc5osDyA89pvXPIilMnChGLZSTTAd+Zq1l/GsS89hmY8kpni2j7KDB2TZHWspj0sSfV2DQd4B0fzCHzVovFBDV5fLgsPbb6RjGUlDW9J9MjKJEPF85qP0fI81agyzrE9FnxwYF5MXUBuEIh57UHU7Ili+TO6kwDK9mEqW7JOGfoRoal+XLywDVC61irCVcHuvtGY2j5/QW91zfi78Dw6bcW54N9/A+QvufeYUOXH4pVVC/ajRiRXJ5b2RqYp4khU7M7PInj7X42aUZ9CPIbW/NQlqESvKGZ+D6x/KQk/0b6Ljss0dpaXK5XSPuF+sjf7IRyw9tabr9W2+xhmgf38kZTvEB0ucXvR768ZeCgbj2X5FzgDnghu4kBOEElYdWzyP5RBVXdjddHvrxl4KBuPK/3TS4xfaGRz6RQbUJEjH6nCVTc3M8USqDXxlkXGyt/DkZ7J29H4sNtyqkh7VNEbjxRlahtDi8HB19WHuPejwtjPPaA3Qcd2qDXxlkXGyt+gpI+oj25gFOvrPHWItcTvfI9sR+RpffGZzEU9ofVWWmWRAxiszVICT5CSuMSr8bCVzEWP7b63NFX4D5pKHLZBHvOxFd+Zu5I3V8WVOYGSZ9IHp2DEvi+HqDXxlkXGyt/Xbt5G5rFPBWDHTBgTqXIzrKgi6qQ2/Od8HzEiHkiY9BclTTAQGT81v9281ooBjDbq6av9CaIXlspFAKM9WD4wrJMSGyvUWg6VzEWP7b63NFX4D5pKHLZBicBM2G+IVyG1J3Khjo3gkoofj/KP4h/5Ixfr0G8YMMDXbt5G5rFPBWDHTBgTqXIz2UllyUlXgbR1MO+W8n0Wo9ztx7v42bgQApdfdT16waoRKro5GXzlN3wfMSIeSJj0a5FlNQw8LRlyXAvdH7CLNpXMRY/tvrc0IHGhtRlFLAOptWn9VuGbznVOxSw+bqJRv9281ooBjDYRKro5GXzlN3wfMSIeSJj06FTocgxR6VgtZyDB6R0ucRr/0QQUDIF5qDXxlkXGyt+ptWn9VuGbznBHgQfi3ncpfI9sR+RpffHoUllVpvk3RGzzURLLajm2CtziW64KHAIj8G3eo7Q9CrPE7sQG274o46Owt5DT9yDS5B+HQuLItS+595hQ5cfiiELh5CtS3k1apPPf6YugCOjtB9vfRxkX0372ExX2DzxP5DKhKevgqTMG/erWsTnq8/TnSPPDjO4qosG7fI4x2oMeYwbJbELEkxGQ5DlU5Nx6nDPYWVBQKwezedDC0hir0eLVINCmTFZ5s63yiIExvXLkwrR+v8SSs8TuxAbbvig/AaikY3kVDn769vJBLH3fOyxQZ13Y28cSV17mbAsYlInATNhviFchEtRfj9IyqtVQRFtY5cy01504Yox6N4gW0oPW/uFoIpqoNfGWRcbK3xUEU0INUM9Q/Qz5Qa/K3RmEYtlJNMB35oeocJ8U7bIORN7coAtNOaQriyPp1ahjhlHHyTQ0RZGMUIJyZoFUkp6nC3EK7+Fb/HuugT5ikRvFcD9qmszl86TBBL+fRwJ4RacLcQrv4Vv8xtd7T1IVlmTQz5AjeYpyZ9sqKEd60d2xiJP9+dI2nl/c9CSVHsOFProkKRuro2ObhchILHYmhXMc1hCg9j6TV7/dvNaKAYw2bW5ec5Qv+Jr4alyc2izGjnD3DMUc/da/NV5eLQMVlL61S4MS/PZkgnTmtsRAhcTlTnsJf44REAeLyNilbh+0cc32gqqToy/0nwDziWeYZMyXZ1kdq40uGFGGS3zKBooEMpcev8pQg+zE2a0fTHQJ688ISqMdJlECDCIWhhTCDVaioOnn/o5+eTUYz/WdutD9KnNj3pkyIuT04SclxQUmldFkk4qMsZDxsz9joM+yYRxdGYFcVyWNtQb7fS/8zs0kkYxlJQ1vSfTIyiRDxfOaj9HyPNWoMs6xPRZ8cGBeTF1AbhCIee1B1OyJYvkzupMAyvZhKluyThn6EaGpfly8sA1QutYqwlXB7r7RmNo+f0Fvdc34u/A8Om3FueDffwPkL7n3mFDlx+KVVQv2o0YkVyeW9kamKeJIVOzOzyJ4+1+NmlGfQjyG1jlewXUoPBy8jdEGTG6A+1q+i47LNHaWlyuV0j7hfrI3Jm3LgZz5FuXVtvsYZoH9/NqB6K+5pKC5PWSA7yLFqU25skJQ29v+3zR7x7YVGOZYjnCw3frpxtW6/CfKEvGiWxGO5gMMvo/AiVJqEyAe7Vsn2JiU8Ymh5f5l+OuBrgCnLwL0gn1AbssIetPp52/Df8WP3DiKPlZ1cWC+X9HhzqivFqrC9h8/+2kjwuV23KD8Ld0RaCT/cJAD45zU2m2Hr1Fj5+cursX8PU31359fs/CoNfGWRcbK3zhnQ/HQRyWE6Pf0JKm26TvgUSTw8uMa/LPE7sQG274oGnkhHOWLndfXqX1BcT19fpeVSw8eeK1BL7n3mFDlx+KR2oL8nuFWz/idPcnRWI2moQpAMATGjcohbxV3AF2ZFo+JumCeYkcomQuDrbCd8gTuTotTi6DcnjssUGdd2NvHElde5mwLGJSJwEzYb4hXIer8HUmQVc97wQ+vUjvBdjzNReFosymZhC+595hQ5cfij5IASVMIQbIFPGYARHVhHEt6ximsPJZn4rM4TttidQcS1F+P0jKq1VBEW1jlzLTXZax0spYeFH3Sg9b+4Wgimqg18ZZFxsrfFQRTQg1Qz1DX6ALqQqn8dogn5UWLR4Y6h6hwnxTtsg5E3tygC005pCuLI+nVqGOGUcfJNDRFkYxQgnJmgVSSnqcLcQrv4Vv8e66BPmKRG8VwP2qazOXzpMEEv59HAnhFpwtxCu/hW/zG13tPUhWWZCtqyXD/qKKY0oPW/uFoIpqoNfGWRcbK3/4ndrcguBFscHvbVgXuI+H+J3a3ILgRbA1eXy4LD22+kYxlJQ1vSfQLsYsz9m1HAbPE7sQG274ou2EpzdE/7SZl3/JOXLbMghHUDJLAZU35MT65WrDAzbwJXZAhY8A6K4iT/fnSNp5fSPnsHct0Z2uGhC8xWXi+vkB1ecXi+MYnMVN4UCyUmVY2z8hmOe+/PL/dvNaKAYw2Y/3FFXKQO94CapzjWGoI3KlT71QxNftDDy0I+VfMnMaLyld6BlNZOQI3SdDE0ozW2SsgJ2uMc8IVpnuM8FXowjDIRANadAGjqDXxlkXGyt9I9kKMFmdfDXzBM6XBPkEgaC1MduzKIPtg1MtGwBlMyD1Okt2cq3elRD3r/lTasadLzGYdxnJGeosCLRNrMsuPzVnJqBaH/N/OUe32hDivHikG6JBDwo7s3OXkGArzLsO4zmBdi/5v8vkw1URNq8yQUA1QEL+Z9g8ligUqx4fvHWIceV4Pi6O1Vkz1+YvIlT5SnJHd7EB6d8oZsJ9DfUfMXRju5BytK8Qzk0qs0msIBn3OJF94egtdDIoSyXQMRPmiHP4+DbUbD7DTMH1pYeVykNEPMoCb13o=
%%% protect end_protected
