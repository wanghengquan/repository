// Library - io, Cell - PDUW08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 17:52:32 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module PDUW08DGZ ( C, PAD, I, OEN, REN );
output  C;

inout  PAD;

input  I, OEN, REN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - nvcm_cell_334x232, View - schematic
// LAST TIME SAVED: Jun 26 10:51:17 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module nvcm_cell_334x232 ( bl, bl_dummyl, bl_dummyr, bl_test, wp,
     wp_dummyb, wp_dummyt, wr, wr_dummyb, wr_dummyt );


inout [335:0]  bl;
inout [1:0]  bl_test;
inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;

input [1:0]  wp_dummyb;
input [1:0]  wp_dummyt;
input [227:0]  wp;
input [1:0]  wr_dummyt;
input [227:0]  wr;
input [1:0]  wr_dummyb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_336x8_8f Invcm_cell_336x8_26_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[221:214]),
     .wp(wp[221:214]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_25_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[213:206]),
     .wp(wp[213:206]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_24_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[205:198]),
     .wp(wp[205:198]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_23_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[197:190]),
     .wp(wp[197:190]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_22_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[189:182]),
     .wp(wp[189:182]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_21_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[181:174]),
     .wp(wp[181:174]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_20_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[173:166]),
     .wp(wp[173:166]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_19_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[165:158]),
     .wp(wp[165:158]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_18_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[157:150]),
     .wp(wp[157:150]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_17_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[149:142]),
     .wp(wp[149:142]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_16_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[141:134]),
     .wp(wp[141:134]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_15_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[133:126]),
     .wp(wp[133:126]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_14_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[125:118]),
     .wp(wp[125:118]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_13_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[117:110]),
     .wp(wp[117:110]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_12_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[109:102]),
     .wp(wp[109:102]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_11_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[101:94]),
     .wp(wp[101:94]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_10_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[93:86]),
     .wp(wp[93:86]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_9_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[85:78]),
     .wp(wp[85:78]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_8_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[77:70]),
     .wp(wp[77:70]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_7_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[69:62]),
     .wp(wp[69:62]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_6_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[61:54]),
     .wp(wp[61:54]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_5_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[53:46]),
     .wp(wp[53:46]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_4_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[45:38]),
     .wp(wp[45:38]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_3_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[37:30]),
     .wp(wp[37:30]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_2_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[29:22]),
     .wp(wp[29:22]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_1_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[21:14]),
     .wp(wp[21:14]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_0_ ( .bl({bl_test[1:0],
     bl[335:0]}), .bl_dummyr(bl_dummyr[1:0]), .wr(wr[13:6]),
     .wp(wp[13:6]), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_t ( .bl({bl_test[1:0], bl[335:0]}),
     .bl_dummyr(bl_dummyr[1:0]), .wr({wr[5:0], wr_dummyt[1:0]}),
     .wp({wp[5:0], wp_dummyt[1:0]}), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_336x8_8f Invcm_cell_336x8_b ( .bl({bl_test[1:0], bl[335:0]}),
     .bl_dummyr(bl_dummyr[1:0]), .wr({wr_dummyb[1:0], wr[227:222]}),
     .wp({wp_dummyb[1:0], wp[227:222]}), .bl_dummyl(bl_dummyl[1:0]));

endmodule
// Library - NVCM, Cell - ml_testdec_columnsx336, View - schematic
// LAST TIME SAVED: Jun 26 10:47:22 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_testdec_columnsx336 ( bl, bl_dummyl, bl_dummyr, bl_test,
     dec_det_even_25, dec_det_odd_25 );

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl_dummyl;
inout [335:0]  bl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_testdec_columns Itestdec_columns_dml (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyl[1:0]));
ml_testdec_columns Itestdec_columns_167_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[335:334]));
ml_testdec_columns Itestdec_columns_166_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[333:332]));
ml_testdec_columns Itestdec_columns_165_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[331:330]));
ml_testdec_columns Itestdec_columns_164_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[329:328]));
ml_testdec_columns Itestdec_columns_163_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[327:326]));
ml_testdec_columns Itestdec_columns_162_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[325:324]));
ml_testdec_columns Itestdec_columns_161_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[323:322]));
ml_testdec_columns Itestdec_columns_160_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[321:320]));
ml_testdec_columns Itestdec_columns_159_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[319:318]));
ml_testdec_columns Itestdec_columns_158_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[317:316]));
ml_testdec_columns Itestdec_columns_157_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[315:314]));
ml_testdec_columns Itestdec_columns_156_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[313:312]));
ml_testdec_columns Itestdec_columns_155_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[311:310]));
ml_testdec_columns Itestdec_columns_154_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[309:308]));
ml_testdec_columns Itestdec_columns_153_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[307:306]));
ml_testdec_columns Itestdec_columns_152_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[305:304]));
ml_testdec_columns Itestdec_columns_151_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[303:302]));
ml_testdec_columns Itestdec_columns_150_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[301:300]));
ml_testdec_columns Itestdec_columns_149_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[299:298]));
ml_testdec_columns Itestdec_columns_148_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[297:296]));
ml_testdec_columns Itestdec_columns_147_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[295:294]));
ml_testdec_columns Itestdec_columns_146_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[293:292]));
ml_testdec_columns Itestdec_columns_145_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[291:290]));
ml_testdec_columns Itestdec_columns_144_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[289:288]));
ml_testdec_columns Itestdec_columns_143_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[287:286]));
ml_testdec_columns Itestdec_columns_142_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[285:284]));
ml_testdec_columns Itestdec_columns_141_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[283:282]));
ml_testdec_columns Itestdec_columns_140_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[281:280]));
ml_testdec_columns Itestdec_columns_139_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[279:278]));
ml_testdec_columns Itestdec_columns_138_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[277:276]));
ml_testdec_columns Itestdec_columns_137_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[275:274]));
ml_testdec_columns Itestdec_columns_136_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[273:272]));
ml_testdec_columns Itestdec_columns_135_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[271:270]));
ml_testdec_columns Itestdec_columns_134_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[269:268]));
ml_testdec_columns Itestdec_columns_133_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[267:266]));
ml_testdec_columns Itestdec_columns_132_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[265:264]));
ml_testdec_columns Itestdec_columns_131_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[263:262]));
ml_testdec_columns Itestdec_columns_130_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[261:260]));
ml_testdec_columns Itestdec_columns_129_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[259:258]));
ml_testdec_columns Itestdec_columns_128_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[257:256]));
ml_testdec_columns Itestdec_columns_127_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[255:254]));
ml_testdec_columns Itestdec_columns_126_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[253:252]));
ml_testdec_columns Itestdec_columns_125_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[251:250]));
ml_testdec_columns Itestdec_columns_124_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[249:248]));
ml_testdec_columns Itestdec_columns_123_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[247:246]));
ml_testdec_columns Itestdec_columns_122_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[245:244]));
ml_testdec_columns Itestdec_columns_121_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[243:242]));
ml_testdec_columns Itestdec_columns_120_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[241:240]));
ml_testdec_columns Itestdec_columns_119_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[239:238]));
ml_testdec_columns Itestdec_columns_118_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[237:236]));
ml_testdec_columns Itestdec_columns_117_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[235:234]));
ml_testdec_columns Itestdec_columns_116_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[233:232]));
ml_testdec_columns Itestdec_columns_115_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[231:230]));
ml_testdec_columns Itestdec_columns_114_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[229:228]));
ml_testdec_columns Itestdec_columns_113_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[227:226]));
ml_testdec_columns Itestdec_columns_112_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[225:224]));
ml_testdec_columns Itestdec_columns_111_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[223:222]));
ml_testdec_columns Itestdec_columns_110_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[221:220]));
ml_testdec_columns Itestdec_columns_109_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[219:218]));
ml_testdec_columns Itestdec_columns_108_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[217:216]));
ml_testdec_columns Itestdec_columns_107_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[215:214]));
ml_testdec_columns Itestdec_columns_106_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[213:212]));
ml_testdec_columns Itestdec_columns_105_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[211:210]));
ml_testdec_columns Itestdec_columns_104_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[209:208]));
ml_testdec_columns Itestdec_columns_103_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[207:206]));
ml_testdec_columns Itestdec_columns_102_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[205:204]));
ml_testdec_columns Itestdec_columns_101_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[203:202]));
ml_testdec_columns Itestdec_columns_100_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[201:200]));
ml_testdec_columns Itestdec_columns_99_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[199:198]));
ml_testdec_columns Itestdec_columns_98_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[197:196]));
ml_testdec_columns Itestdec_columns_97_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[195:194]));
ml_testdec_columns Itestdec_columns_96_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[193:192]));
ml_testdec_columns Itestdec_columns_95_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[191:190]));
ml_testdec_columns Itestdec_columns_94_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[189:188]));
ml_testdec_columns Itestdec_columns_93_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[187:186]));
ml_testdec_columns Itestdec_columns_92_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[185:184]));
ml_testdec_columns Itestdec_columns_91_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[183:182]));
ml_testdec_columns Itestdec_columns_90_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[181:180]));
ml_testdec_columns Itestdec_columns_89_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[179:178]));
ml_testdec_columns Itestdec_columns_88_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[177:176]));
ml_testdec_columns Itestdec_columns_87_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[175:174]));
ml_testdec_columns Itestdec_columns_86_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[173:172]));
ml_testdec_columns Itestdec_columns_85_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[171:170]));
ml_testdec_columns Itestdec_columns_84_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[169:168]));
ml_testdec_columns Itestdec_columns_83_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[167:166]));
ml_testdec_columns Itestdec_columns_82_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[165:164]));
ml_testdec_columns Itestdec_columns_81_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[163:162]));
ml_testdec_columns Itestdec_columns_80_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[161:160]));
ml_testdec_columns Itestdec_columns_79_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[159:158]));
ml_testdec_columns Itestdec_columns_78_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[157:156]));
ml_testdec_columns Itestdec_columns_77_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[155:154]));
ml_testdec_columns Itestdec_columns_76_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[153:152]));
ml_testdec_columns Itestdec_columns_75_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[151:150]));
ml_testdec_columns Itestdec_columns_74_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[149:148]));
ml_testdec_columns Itestdec_columns_73_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[147:146]));
ml_testdec_columns Itestdec_columns_72_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[145:144]));
ml_testdec_columns Itestdec_columns_71_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[143:142]));
ml_testdec_columns Itestdec_columns_70_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[141:140]));
ml_testdec_columns Itestdec_columns_69_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[139:138]));
ml_testdec_columns Itestdec_columns_68_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[137:136]));
ml_testdec_columns Itestdec_columns_67_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[135:134]));
ml_testdec_columns Itestdec_columns_66_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[133:132]));
ml_testdec_columns Itestdec_columns_65_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[131:130]));
ml_testdec_columns Itestdec_columns_64_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[129:128]));
ml_testdec_columns Itestdec_columns_63_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[127:126]));
ml_testdec_columns Itestdec_columns_62_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[125:124]));
ml_testdec_columns Itestdec_columns_61_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[123:122]));
ml_testdec_columns Itestdec_columns_60_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[121:120]));
ml_testdec_columns Itestdec_columns_59_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[119:118]));
ml_testdec_columns Itestdec_columns_58_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[117:116]));
ml_testdec_columns Itestdec_columns_57_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[115:114]));
ml_testdec_columns Itestdec_columns_56_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[113:112]));
ml_testdec_columns Itestdec_columns_55_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[111:110]));
ml_testdec_columns Itestdec_columns_54_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[109:108]));
ml_testdec_columns Itestdec_columns_53_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[107:106]));
ml_testdec_columns Itestdec_columns_52_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[105:104]));
ml_testdec_columns Itestdec_columns_51_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[103:102]));
ml_testdec_columns Itestdec_columns_50_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[101:100]));
ml_testdec_columns Itestdec_columns_49_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[99:98]));
ml_testdec_columns Itestdec_columns_48_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[97:96]));
ml_testdec_columns Itestdec_columns_47_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[95:94]));
ml_testdec_columns Itestdec_columns_46_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[93:92]));
ml_testdec_columns Itestdec_columns_45_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[91:90]));
ml_testdec_columns Itestdec_columns_44_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[89:88]));
ml_testdec_columns Itestdec_columns_43_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[87:86]));
ml_testdec_columns Itestdec_columns_42_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[85:84]));
ml_testdec_columns Itestdec_columns_41_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[83:82]));
ml_testdec_columns Itestdec_columns_40_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[81:80]));
ml_testdec_columns Itestdec_columns_39_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[79:78]));
ml_testdec_columns Itestdec_columns_38_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[77:76]));
ml_testdec_columns Itestdec_columns_37_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[75:74]));
ml_testdec_columns Itestdec_columns_36_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[73:72]));
ml_testdec_columns Itestdec_columns_35_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[71:70]));
ml_testdec_columns Itestdec_columns_34_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[69:68]));
ml_testdec_columns Itestdec_columns_33_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[67:66]));
ml_testdec_columns Itestdec_columns_32_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[65:64]));
ml_testdec_columns Itestdec_columns_31_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[63:62]));
ml_testdec_columns Itestdec_columns_30_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[61:60]));
ml_testdec_columns Itestdec_columns_29_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[59:58]));
ml_testdec_columns Itestdec_columns_28_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[57:56]));
ml_testdec_columns Itestdec_columns_27_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[55:54]));
ml_testdec_columns Itestdec_columns_26_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[53:52]));
ml_testdec_columns Itestdec_columns_25_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[51:50]));
ml_testdec_columns Itestdec_columns_24_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[49:48]));
ml_testdec_columns Itestdec_columns_23_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[47:46]));
ml_testdec_columns Itestdec_columns_22_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[45:44]));
ml_testdec_columns Itestdec_columns_21_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[43:42]));
ml_testdec_columns Itestdec_columns_20_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[41:40]));
ml_testdec_columns Itestdec_columns_19_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[39:38]));
ml_testdec_columns Itestdec_columns_18_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[37:36]));
ml_testdec_columns Itestdec_columns_17_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[35:34]));
ml_testdec_columns Itestdec_columns_16_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[33:32]));
ml_testdec_columns Itestdec_columns_15_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[31:30]));
ml_testdec_columns Itestdec_columns_14_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[29:28]));
ml_testdec_columns Itestdec_columns_13_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[27:26]));
ml_testdec_columns Itestdec_columns_12_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[25:24]));
ml_testdec_columns Itestdec_columns_11_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[23:22]));
ml_testdec_columns Itestdec_columns_10_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[21:20]));
ml_testdec_columns Itestdec_columns_9_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[19:18]));
ml_testdec_columns Itestdec_columns_8_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[17:16]));
ml_testdec_columns Itestdec_columns_7_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[15:14]));
ml_testdec_columns Itestdec_columns_6_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[13:12]));
ml_testdec_columns Itestdec_columns_5_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[11:10]));
ml_testdec_columns Itestdec_columns_4_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[9:8]));
ml_testdec_columns Itestdec_columns_3_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[7:6]));
ml_testdec_columns Itestdec_columns_2_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[5:4]));
ml_testdec_columns Itestdec_columns_1_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[3:2]));
ml_testdec_columns Itestdec_columns_0_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[1:0]));
ml_testdec_columns Itestdec_columns_dmr (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyr[1:0]));
ml_testdec_columns Itestdec_columns_tst (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_test[1:0]));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x16, View - schematic
// LAST TIME SAVED: Jun 26 10:50:42 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_x16 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp2, yp2_b_25, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [15:0]  bl;

input [7:0]  yp3_25;
input [7:0]  yp3_b_25;
input [1:0]  yp2;
input [1:0]  yp2_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M0 ( .D(net49), .B(GND_), .G(yp2[1]), .S(bl_out));
nch_hvt  M2 ( .D(net53), .B(GND_), .G(yp2[0]), .S(bl_out));
nch_25  M11 ( .D(net49), .B(GND_), .G(yp2_b_25[1]), .S(vblinhi_rdo));
nch_25  M20 ( .D(net53), .B(GND_), .G(yp2_b_25[0]), .S(vblinhi_rde));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]), .bl_out(net53),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_1 ( .bl(bl[15:8]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .vdd_tieh(vdd_tieh), .bl_out(net49), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x336, View - schematic
// LAST TIME SAVED: Jun 26 10:50:57 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_x336 ( bl, bl_dummyl, bl_dummyr, bl_out, bl_test,
     vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh,
     pgminhi_dmmy_b_25, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25,
     yp_test, yp_test_25, yp_test_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25;

inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;
inout [1:0]  bl_test;
inout [335:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp2;
input [7:0]  yp2_b_25;
input [10:5]  yp1_b_25;
input [7:0]  yp3_25;
input [1:0]  yp_test_25;
input [10:5]  yp1;
input [1:0]  yp_test;
input [1:0]  yp_test_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:10]  blx8_out;

wire  [5:9]  blx64_out;



ml_ymux_bls_x16 Iml_ymux_bls_x16 ( .bl(bl[335:320]),
     .yp2_b_25(yp2_b_25[1:0]), .yp2(yp2[1:0]), .bl_out(blx8_out[10]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_r ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyr[1:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_l ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyl[1:0]));
pch_25  M7 ( .D(bl_test[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M8 ( .D(bl_test[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
ml_ymux_bls_x64 Iml_ymux_bls_x64_0 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[5]), .bl(bl[63:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_2 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[7]), .bl(bl[191:128]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_4 ( .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]), .bl(bl[319:256]),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .bl_out(blx64_out[9]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo));
ml_ymux_bls_x64 Iml_ymux_bls_x64_1 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[6]), .bl(bl[127:64]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_3 ( .yp2(yp2[7:0]), .bl_out(blx64_out[8]),
     .bl(bl[255:192]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .yp2_b_25(yp2_b_25[7:0]), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));
nch_hvt  M21 ( .D(net224), .B(GND_), .G(yp_test[1]), .S(bl_out));
nch_hvt  M19 ( .D(net228), .B(GND_), .G(yp_test[1]), .S(net224));
nch_hvt  M23 ( .D(net232), .B(GND_), .G(yp_test[0]), .S(bl_out));
nch_hvt  M28 ( .D(net236), .B(GND_), .G(yp1[10]), .S(bl_out));
nch_hvt  M0 ( .D(blx64_out[7]), .B(GND_), .G(yp1[7]), .S(bl_out));
nch_hvt  M22 ( .D(net244), .B(GND_), .G(yp_test[0]), .S(net232));
nch_hvt  M24 ( .D(blx64_out[5]), .B(GND_), .G(yp1[5]), .S(bl_out));
nch_hvt  M30 ( .D(blx8_out[10]), .B(GND_), .G(yp1[10]), .S(net236));
nch_hvt  M3 ( .D(blx64_out[9]), .B(GND_), .G(yp1[9]), .S(bl_out));
nch_hvt  M4 ( .D(blx64_out[8]), .B(GND_), .G(yp1[8]), .S(bl_out));
nch_hvt  M2 ( .D(blx64_out[6]), .B(GND_), .G(yp1[6]), .S(bl_out));
nch_25  M27 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[5]),
     .S(blx64_out[5]));
nch_25  M26 ( .D(vblinhi_rdo), .B(GND_), .G(yp_test_b_25[1]),
     .S(bl_test[1]));
nch_25  M25 ( .D(bl_test[1]), .B(GND_), .G(yp_test_25[1]), .S(net228));
nch_25  M18 ( .D(vblinhi_rde), .B(GND_), .G(yp_test_b_25[0]),
     .S(bl_test[0]));
nch_25  M29 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[10]),
     .S(blx8_out[10]));
nch_25  M17 ( .D(bl_test[0]), .B(GND_), .G(yp_test_25[0]), .S(net244));
nch_25  M1 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[7]),
     .S(blx64_out[7]));
nch_25  M20 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[6]),
     .S(blx64_out[6]));
nch_25  M5 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[9]),
     .S(blx64_out[9]));
nch_25  M6 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[8]),
     .S(blx64_out[8]));

endmodule
// Library - NVCM, Cell - ml_core_336x232, View - schematic
// LAST TIME SAVED: Jun 26 10:53:25 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_core_336x232 ( dec_ok_25, bl_out, vblinhi_pgm_25,
     vblinhi_rde, vblinhi_rdo, vdd_tieh, pgminhi_dmmy_b_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp, wr, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25,
     yp3_b_25, yp_test, yp_test_25, yp_test_b_25 );
output  dec_ok_25;

inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25, testdec_en_b_25, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b_25;

input [7:0]  yp3_b_25;
input [1:0]  yp_test_b_25;
input [1:0]  yp_test;
input [10:5]  yp1;
input [227:0]  wp;
input [7:0]  yp3_25;
input [10:5]  yp1_b_25;
input [7:0]  yp2_b_25;
input [227:0]  wr;
input [7:0]  yp2;
input [1:0]  yp_test_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  bl_dummyr;

wire  [1:0]  bl_test;

wire  [1:0]  bl_dummyl;

wire  [335:0]  bl;



nvcm_cell_334x232 Invcm_cell_334x232 ( .bl(bl[335:0]),
     .bl_dummyr(bl_dummyr[1:0]), .wr_dummyt({net100, net100}),
     .wr_dummyb({net100, net100}), .wr(wr[227:0]), .wp_dummyt({net100,
     net100}), .wp_dummyb({net100, net100}), .wp(wp[227:0]),
     .bl_test(bl_test[1:0]), .bl_dummyl(bl_dummyl[1:0]));
ml_testdec_columnsx336 Itestdec_columnsx336 ( .bl(bl[335:0]),
     .bl_dummyr(bl_dummyr[1:0]), .bl_dummyl(bl_dummyl[1:0]),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl_test(bl_test[1:0]));
ml_ymux_bls_x336 Iml_ymux_bls_x336 ( .bl(bl[335:0]), .yp1(yp1[10:5]),
     .yp1_b_25(yp1_b_25[10:5]), .yp2_b_25(yp2_b_25[7:0]),
     .yp2(yp2[7:0]), .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .bl_dummyl(bl_dummyl[1:0]),
     .bl_dummyr(bl_dummyr[1:0]), .bl_test(bl_test[1:0]),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_25(yp_test_25[1:0]),
     .yp_test(yp_test[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3_25[7:0]), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_out(bl_out));
vdd_tielow I47 ( .gnd_tiel(net100));
ml_testdec_bgen Itestdec_bgen ( .dec_ok_25(dec_ok_25),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25), .dec_det_25(dec_det_25),
     .dec_bias_25(dec_bias));
ml_testdec_rowsx228 Itestdec_rowsx228 ( .dec_bias_25(dec_bias),
     .dec_det_25(dec_det_25), .wr(wr[227:0]), .wp(wp[227:0]),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp_x4, View - schematic
// LAST TIME SAVED: Jan 23 10:17:05 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x4 ( wp, gwl_b_sup_25, ngate_25, gwl_b_25,
     gwl_b_gnden_25, gwp_hv, s_b_25, s_b_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_25, gwl_b_gnden_25, gwp_hv;

output [3:0]  wp;

input [3:0]  s_b_25;
input [3:0]  s_b_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwl_b_25(gwl_b_25), .gwl_gnd_25(gwl_gnd_25));
ml_rock_lwldrv_wp Iml_lwldrv_1 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[1]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[1]), .wp(wp[1]));
ml_rock_lwldrv_wp Iml_lwldrv_2 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[2]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[2]), .wp(wp[2]));
ml_rock_lwldrv_wp Iml_lwldrv_3 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[3]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[3]), .wp(wp[3]));
ml_rock_lwldrv_wp Iml_lwldrv_0 ( .gwl_gnd_25(gwl_gnd_25),
     .s_b_hv(s_b_hv[0]), .gwp_hv(gwp_hv), .gwl_b_25(gwl_b_25),
     .ngate_25(ngate_25), .s_b_25(s_b_25[0]), .wp(wp[0]));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp_x228, View - schematic
// LAST TIME SAVED: Mar 28 09:57:53 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp_x228 ( wp, gwl_b_sup_25, ngate_25, s_b_25,
     s_b_hv, gwl_b_25, gwl_b_gnden_25, gwp_hv );

inout  gwl_b_sup_25, ngate_25;

input  gwl_b_gnden_25;

output [227:0]  wp;

inout [3:0]  s_b_25;
inout [3:0]  s_b_hv;

input [56:0]  gwl_b_25;
input [56:0]  gwp_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_56_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[56]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[227:224]), .gwl_b_25(gwl_b_25[56]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_55_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[55]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[223:220]), .gwl_b_25(gwl_b_25[55]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_54_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[54]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[219:216]), .gwl_b_25(gwl_b_25[54]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_53_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[53]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[215:212]), .gwl_b_25(gwl_b_25[53]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_52_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[52]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[211:208]), .gwl_b_25(gwl_b_25[52]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_51_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[51]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[207:204]), .gwl_b_25(gwl_b_25[51]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_50_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[50]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[203:200]), .gwl_b_25(gwl_b_25[50]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_49_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[49]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[199:196]), .gwl_b_25(gwl_b_25[49]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_48_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[48]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[195:192]), .gwl_b_25(gwl_b_25[48]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_47_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[47]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[191:188]), .gwl_b_25(gwl_b_25[47]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_46_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[46]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[187:184]), .gwl_b_25(gwl_b_25[46]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_45_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[45]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[183:180]), .gwl_b_25(gwl_b_25[45]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_44_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[44]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[179:176]), .gwl_b_25(gwl_b_25[44]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_43_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[43]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[175:172]), .gwl_b_25(gwl_b_25[43]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_42_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[42]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[171:168]), .gwl_b_25(gwl_b_25[42]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_41_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[41]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[167:164]), .gwl_b_25(gwl_b_25[41]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_40_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[40]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[163:160]), .gwl_b_25(gwl_b_25[40]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_39_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[39]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[159:156]), .gwl_b_25(gwl_b_25[39]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_38_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[38]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[155:152]), .gwl_b_25(gwl_b_25[38]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_37_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[37]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[151:148]), .gwl_b_25(gwl_b_25[37]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_36_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[36]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[147:144]), .gwl_b_25(gwl_b_25[36]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_35_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[35]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[143:140]), .gwl_b_25(gwl_b_25[35]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_34_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[34]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[139:136]), .gwl_b_25(gwl_b_25[34]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_33_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[33]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[135:132]), .gwl_b_25(gwl_b_25[33]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_32_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[32]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[131:128]), .gwl_b_25(gwl_b_25[32]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_31_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[31]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[127:124]), .gwl_b_25(gwl_b_25[31]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_30_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[30]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[123:120]), .gwl_b_25(gwl_b_25[30]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_29_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[29]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[119:116]), .gwl_b_25(gwl_b_25[29]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_28_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[28]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[115:112]), .gwl_b_25(gwl_b_25[28]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_27_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[27]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[111:108]), .gwl_b_25(gwl_b_25[27]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_26_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[26]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[107:104]), .gwl_b_25(gwl_b_25[26]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_25_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[25]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[103:100]), .gwl_b_25(gwl_b_25[25]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_24_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[24]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[99:96]), .gwl_b_25(gwl_b_25[24]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_23_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[23]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[95:92]), .gwl_b_25(gwl_b_25[23]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_22_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[22]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[91:88]), .gwl_b_25(gwl_b_25[22]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_21_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[21]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[87:84]), .gwl_b_25(gwl_b_25[21]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_20_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[20]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[83:80]), .gwl_b_25(gwl_b_25[20]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_19_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[19]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[79:76]), .gwl_b_25(gwl_b_25[19]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_18_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[18]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[75:72]), .gwl_b_25(gwl_b_25[18]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_17_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[17]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[71:68]), .gwl_b_25(gwl_b_25[17]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_16_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[16]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[67:64]), .gwl_b_25(gwl_b_25[16]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_15_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[15]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[63:60]), .gwl_b_25(gwl_b_25[15]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_14_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[14]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[59:56]), .gwl_b_25(gwl_b_25[14]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_13_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[13]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[55:52]), .gwl_b_25(gwl_b_25[13]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_12_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[12]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[51:48]), .gwl_b_25(gwl_b_25[12]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_11_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[11]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[47:44]), .gwl_b_25(gwl_b_25[11]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_10_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[10]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[43:40]), .gwl_b_25(gwl_b_25[10]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_9_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[9]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[39:36]), .gwl_b_25(gwl_b_25[9]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_8_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[8]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[35:32]), .gwl_b_25(gwl_b_25[8]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_7_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[7]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[31:28]), .gwl_b_25(gwl_b_25[7]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_6_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[6]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[27:24]), .gwl_b_25(gwl_b_25[6]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_5_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[5]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[23:20]), .gwl_b_25(gwl_b_25[5]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_4_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[4]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[19:16]), .gwl_b_25(gwl_b_25[4]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_3_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[3]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[15:12]), .gwl_b_25(gwl_b_25[3]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_2_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[2]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[11:8]), .gwl_b_25(gwl_b_25[2]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_1_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[1]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[7:4]), .gwl_b_25(gwl_b_25[1]), .s_b_hv(s_b_hv[3:0]));
ml_rock_lwldrv_wp_x4 Iml_rock_lwldrv_wp_x4_0_ (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[0]), .ngate_25(ngate_25), .s_b_25(s_b_25[3:0]),
     .wp(wp[3:0]), .gwl_b_25(gwl_b_25[0]), .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - NVCM, Cell - ml_core_654x232_top, View - schematic
// LAST TIME SAVED: Sep 23 11:13:28 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_core_654x232_top ( nv_dataout, bl_pgm_glb, gwl_b_sup_25,
     ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpxa,
     ysup_25, fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, gwl_b_25, gwp_hv, pgminhi_dmmy_b_25,
     sa_ngate_25, sa_pgate_vpxa, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, wr );
output  nv_dataout;

inout  bl_pgm_glb, gwl_b_sup_25, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi_rde, vblinhi_rdo, vpxa, ysup_25;

input  fsm_gwlbdis_b_25, fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     pgminhi_dmmy_b_25, saen_25, saen_b_vpxa, testdec_en_b_25,
     testdec_even_b_25, testdec_odd_b_25, testdec_prec_b_25,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr;

input [1:0]  fsm_rowadd;
input [9:0]  fsm_coladd;
input [4:1]  sa_ngate_25;
input [227:0]  wr;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefrd;
input [56:0]  gwp_hv;
input [56:0]  gwl_b_25;
input [2:0]  fsm_trim_rrefpgm;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  yp_test_b_25;

wire  [1:0]  yp_test_25;

wire  [1:0]  yp_test;

wire  [7:0]  yp3_b_25;

wire  [7:0]  yp3;

wire  [7:0]  yp2;

wire  [7:0]  yp2_b_25;

wire  [227:0]  wp;

wire  [3:0]  s_b_hv;

wire  [3:0]  s_b_25;

wire  [10:0]  yp1;

wire  [10:0]  yp1_b_25;



ml_core_ctrl_spare_right Iml_core_ctrl_spare_right ( );
ml_core_ctrl_spare_left Iml_core_ctrl_spare_left ( );
ml_core_ctrl_top_8f Icore_ctrl_top ( .tm_allbank_sel(tm_allbank_sel),
     .fsm_coladd(fsm_coladd[9:0]), .dec_ok_25_r(dec_ok_25_r),
     .dec_ok_25_l(dec_ok_25_l), .yp1(yp1[10:0]),
     .yp1_b_25(yp1_b_25[10:0]), .yp2_b_25(yp2_b_25[7:0]),
     .yp2(yp2[7:0]), .fsm_tm_trow(fsm_tm_trow), .tm_dma(tm_dma),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .gwl_b_gnden_25(gwl_b_gnden_25),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .bl_pgm_glb(bl_pgm_glb),
     .vdd_tieh(vdd_tieh), .tm_testdec_wr(tm_testdec_wr),
     .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .tm_allbl_l(tm_allbl_l),
     .tm_allbl_h(tm_allbl_h), .testdec_en_b_25(testdec_en_b_25),
     .saen_b_vpxa(saen_b_vpxa), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_ymuxdis(fsm_ymuxdis),
     .fsm_wpen(fsm_wpen), .fsm_vpxaset(fsm_vpxaset),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_blkadd(fsm_blkadd[3:0]), .yp_test_b_25(yp_test_b_25[1:0]),
     .yp_test_25(yp_test_25[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .nv_dataout(nv_dataout_in), .ysup_25(ysup_25),
     .vpxa(vpxa), .vblinhi_pgm_25(vblinhi_pgm_25),
     .sbhvsup_hv(sbhvsup_hv), .sb25sup_25(sb25sup_25),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .bl_out(bl_out),
     .yp_test(yp_test[1:0]));
ml_core_320x232 Iml_core_320x232 ( .dec_ok_25(dec_ok_25_l),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .wp(wp[227:0]),
     .wr(wr[227:0]), .vdd_tieh(vdd_tieh), .bl_out(bl_out),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .yp3_25(yp3[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25), .yp1(yp1[4:0]),
     .yp1_b_25(yp1_b_25[4:0]));
ml_core_336x232 Iml_core_336x232 ( .dec_ok_25(dec_ok_25_r),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_25(yp_test_25[1:0]),
     .yp_test(yp_test[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3[7:0]), .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]),
     .yp1_b_25(yp1_b_25[10:5]), .yp1(yp1[10:5]), .wr(wr[227:0]),
     .wp(wp[227:0]), .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vdd_tieh(vdd_tieh),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_rde(vblinhi_rde),
     .vblinhi_pgm_25(vblinhi_pgm_25), .bl_out(bl_out));
inv_hvt I131 ( .A(nv_dataout_in), .Y(net232));
inv_hvt I45 ( .A(net232), .Y(nv_dataout));
ml_rock_lwldrv_wp_x228 Iml_rock_lwldrv_wp_x228 (
     .gwl_b_gnden_25(gwl_b_gnden_25), .gwl_b_sup_25(gwl_b_sup_25),
     .gwp_hv(gwp_hv[56:0]), .gwl_b_25(gwl_b_25[56:0]), .wp(wp[227:0]),
     .s_b_hv(s_b_hv[3:0]), .s_b_25(s_b_25[3:0]), .ngate_25(ngate_25));

endmodule
// Library - NVCM, Cell - ml_hv_invx3_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:19:36 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hv_invx3_enhance ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh
     );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_switch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 14:46:53 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_lshv_6v_switch_enhance ( out_b_hv, out_hv, in_hv, sel_25,
     sel_b_25, vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M11 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));

endmodule
// Library - misc, Cell - vpp_clamp, View - schematic
// LAST TIME SAVED: Jun  5 16:48:52 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module vpp_clamp ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vpp_clamp_finger I3 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I1 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I2 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I5 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I6 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I7 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I8 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I9 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I0 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));
vpp_clamp_finger I4 ( .VSS(VSS), .VDDIO(VDDIO), .VPP(VPP));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv_hotsw_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:16:13 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw_enhance ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3_enhance Ihv_invx3 ( .vddp_tieh(vddp_tieh),
     .out_b_hv(out_b_hv), .sel_25(sel_25), .in_hv(in_hv),
     .sel_hv(sel_hv));
ml_lshv_6v_switch_enhance Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM, Cell - ml_hv_hotswitch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:15:29 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hv_hotswitch_enhance ( hv_in_hv, hv_out_hv, selhv_25,
     vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw_enhance Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M7 ( .D(net12), .B(GND_), .G(selhv_25), .S(net15));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
pch_25  M0 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_hotswitch_enhance, View - schematic
// LAST TIME SAVED: Apr 30 11:28:27 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch_enhance ( hvin_a_hv, hvin_b_hv, out_hv,
     sel_hv_a_25, sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch_enhance Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_logic, View - schematic
// LAST TIME SAVED: May  9 14:35:36 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_logic ( gnv, gred, gwl_misc, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, s, sa_trim, saen, testdec_en_b, testdec_even_b,
     testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen,
     wrsup_2vdd, fsm_coladd, fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv,
     fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_tm_allbl_h, fsm_tm_allbl_l,
     fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_trow, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_dma, tm_testdec, tm_testdec_wr );
output  gwl_misc, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, saen, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [1:0]  gred;
output [3:0]  s;
output [2:0]  sa_trim;
output [5:0]  gnv;

input [2:0]  fsm_trim_rrefpgm;
input [0:0]  fsm_coladd;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_b;

wire  [5:0]  gnv_b;

wire  [1:0]  xadd_b;

wire  [1:0]  gred_b;

wire  [1:0]  xadd;

wire  [0:2]  net390;

wire  [2:0]  sa_trim_b;

wire  [0:1]  net386;



vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
anor21_hvt I109_1_ ( .A(net386[0]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I109_0_ ( .A(net386[1]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
oai22x2_hvt I93 ( .A1(fsm_rd), .Y(net196), .A0(fsm_pgmvfy),
     .B0(gnd_tiel), .B1(gnd_tiel));
ml_pump_a_clkdly I230 ( .in(net0231), .out(net0232));
ml_pump_a_clkdly I208 ( .in(net200), .out(net201));
ml_pump_a_clkdly I202 ( .in(net202), .out(net203));
ml_pump_a_clkdly I198 ( .in(net204), .out(net205));
ml_pump_a_clkdly I207 ( .in(net206), .out(net207));
nor4_hvt I175 ( .D(fsm_tm_allwl_h), .B(fsm_pgmvfy), .Y(net211),
     .A(fsm_pgmvfy), .C(fsm_rd));
nor4_hvt I176 ( .D(testdec_wp), .B(fsm_nvcmen_b), .Y(net216),
     .A(fsm_wren_b), .C(net331));
nor4_hvt I218 ( .D(net282), .B(fsm_tm_allbl_l), .Y(net0258),
     .A(fsm_tm_allbl_l), .C(fsm_nvcmen_b));
nor4_hvt I191 ( .B(pgm_hvpulse), .Y(wrsup_2vdd_int), .D(fsm_nvcmen_b),
     .A(pgm_hvpulse), .C(testdec_wr));
nor4_hvt I171 ( .D(fsm_wpen_b), .B(fsm_nvcmen_b), .Y(net226),
     .A(testdec_wr), .C(fsm_tm_allwl_l));
nor2_hvt I233 ( .A(fsm_pgm), .B(fsm_pgmvfy), .Y(net0176));
nor2_hvt I228 ( .A(fsm_pgmdisc), .B(fsm_pgmhv), .Y(net0231));
nor2_hvt I231 ( .A(net0258), .B(tm_testdec), .Y(pgminhi_dmmy_b));
nor2_hvt I165 ( .B(fsm_nv_sisi_ui), .Y(x1_desel_b),
     .A(fsm_nv_rri_trim));
nor2_hvt I186 ( .A(fsm_pgmvfy), .B(fsm_pgm_b), .Y(stress2));
nor2_hvt I216 ( .A(fsm_nvcmen_b), .B(tm_dma), .Y(saen));
nor2_hvt I203 ( .A(net203), .B(net351), .Y(gwlbsup_vpxa));
nor2_hvt I209 ( .A(net207), .B(net246), .Y(gwphv_vppint));
nor2_hvt I214 ( .A(net0232), .B(fsm_nvcmen_b), .Y(net246));
nor2_hvt I210 ( .A(net359), .B(net201), .Y(gwphv_vddp));
nor2_hvt I226 ( .A(net0288), .B(net0390), .Y(gwlb_en));
nor2_hvt I201 ( .A(net196), .B(net205), .Y(gwlbsup_vddp));
nor3_hvt I182 ( .B(fsm_tm_allwl_l), .Y(net330), .A(fsm_tm_allwl_l),
     .C(fsm_tm_allwl_l));
nor3_hvt I105 ( .B(fsm_tm_allwl_h), .Y(net0288), .A(fsm_tm_allwl_h),
     .C(fsm_tm_allwl_h));
nor3_hvt I162 ( .Y(net0274), .B(fsm_tm_trow), .C(fsm_nv_sisi_ui),
     .A(fsm_nv_rri_trim));
anor31_hvt I121_3_ ( .A(net365), .D(net345), .B(xadd[1]), .Y(s_b[3]),
     .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net365), .D(net345), .B(xadd[1]), .Y(s_b[2]),
     .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net365), .D(net345), .B(xadd_b[1]), .Y(s_b[1]),
     .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net365), .D(net345), .B(xadd_b[1]), .Y(s_b[0]),
     .C(xadd_b[0]));
nand3_hvt I167 ( .B(fsm_nvcmen), .Y(gwlb_dis), .A(net0332),
     .C(testwr_wpgnd_b));
nand3_hvt I184 ( .Y(net274), .B(fsm_tm_allwl_h), .C(fsm_tm_allwl_h),
     .A(stress2));
nand3_hvt I125 ( .C(fsm_ymuxdis), .A(tm_testdec), .Y(testdec_prec_b),
     .B(fsm_rd));
nand3_hvt I195 ( .Y(net282), .B(net341), .C(fsm_lshven), .A(fsm_pgm));
nand3_hvt I154 ( .Y(net286), .B(fsm_pgm), .C(fsm_tm_allwl_h),
     .A(fsm_wren));
nand3_hvt I122 ( .A(fsm_nvcmen), .C(net307), .Y(net292),
     .B(tm_allwl_l_b));
nand2_hvt I170 ( .A(tm_testdec_wr), .Y(testwr_wpgnd_b),
     .B(tm_testdec));
nand2_hvt I188 ( .A(testdec_en), .Y(testdec_odd_b), .B(fsm_coladd[0]));
nand2_hvt I189 ( .A(net355), .Y(testdec_even_b), .B(testdec_en));
nand2_hvt I155 ( .A(net377), .Y(net307), .B(tm_testdec));
nand2_hvt I89 ( .A(fsm_rd), .Y(testdec_en_b), .B(tm_testdec));
inv_hvt I232 ( .A(net0176), .Y(net0365));
inv_hvt I174 ( .A(net211), .Y(wp_frcen));
inv_hvt I163 ( .A(net0274), .Y(gwl_misc));
inv_hvt I187 ( .A(fsm_pgm), .Y(fsm_pgm_b));
inv_hvt I131 ( .A(testdec_en_b), .Y(testdec_en));
inv_hvt I178 ( .A(net307), .Y(testdec_wp));
inv_hvt I196 ( .A(net282), .Y(pgm_hvpulse));
inv_hvt I185 ( .A(net274), .Y(wr_frcen));
inv_hvt I206 ( .A(gwlbsup_vpxa), .Y(net204));
inv_hvt I177 ( .A(net216), .Y(wr_dis));
inv_hvt I183 ( .A(net330), .Y(net331));
inv_hvt I192 ( .A(wrsup_2vdd_int), .Y(net333));
inv_hvt I179 ( .A(fsm_wpen), .Y(fsm_wpen_b));
inv_hvt I194 ( .A(testwr_wpgnd_b), .Y(testdec_wr));
inv_hvt I212 ( .A(gwphv_vddp), .Y(net206));
inv_hvt I197 ( .A(fsm_pgmvfy), .Y(net341));
inv_hvt I205 ( .A(gwlbsup_vddp), .Y(net202));
inv_hvt I152 ( .A(net286), .Y(net345));
inv_hvt I120_5_ ( .A(gnv_b[5]), .Y(gnv[5]));
inv_hvt I120_4_ ( .A(gnv_b[4]), .Y(gnv[4]));
inv_hvt I120_3_ ( .A(gnv_b[3]), .Y(gnv[3]));
inv_hvt I120_2_ ( .A(gnv_b[2]), .Y(gnv[2]));
inv_hvt I120_1_ ( .A(gnv_b[1]), .Y(gnv[1]));
inv_hvt I120_0_ ( .A(gnv_b[0]), .Y(gnv[0]));
inv_hvt I172 ( .A(net226), .Y(wp_dis));
inv_hvt I204 ( .A(net196), .Y(net351));
inv_hvt I160_1_ ( .A(gred_b[1]), .Y(gred[1]));
inv_hvt I160_0_ ( .A(gred_b[0]), .Y(gred[0]));
inv_hvt I190 ( .A(fsm_coladd[0]), .Y(net355));
inv_hvt I150_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I150_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I215 ( .A(net246), .Y(net359));
inv_hvt I225 ( .A(pgm_hvpulse), .Y(net0390));
inv_hvt I213 ( .A(gwphv_vppint), .Y(net200));
inv_hvt I161_1_ ( .A(fsm_rowadd[3]), .Y(gred_b[1]));
inv_hvt I161_0_ ( .A(fsm_rowadd[2]), .Y(gred_b[0]));
inv_hvt I151 ( .A(net292), .Y(net365));
inv_hvt I119_5_ ( .A(fsm_rowadd[7]), .Y(gnv_b[5]));
inv_hvt I119_4_ ( .A(fsm_rowadd[6]), .Y(gnv_b[4]));
inv_hvt I119_3_ ( .A(fsm_rowadd[5]), .Y(gnv_b[3]));
inv_hvt I119_2_ ( .A(fsm_rowadd[4]), .Y(gnv_b[2]));
inv_hvt I119_1_ ( .A(fsm_rowadd[3]), .Y(gnv_b[1]));
inv_hvt I119_0_ ( .A(fsm_rowadd[2]), .Y(gnv_b[0]));
inv_hvt I157 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I153 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I193 ( .A(net333), .Y(wrsup_2vdd));
inv_hvt I181 ( .A(fsm_wren), .Y(fsm_wren_b));
inv_hvt I156 ( .A(tm_testdec_wr), .Y(net377));
inv_hvt I147_3_ ( .A(s_b[3]), .Y(s[3]));
inv_hvt I147_2_ ( .A(s_b[2]), .Y(s[2]));
inv_hvt I147_1_ ( .A(s_b[1]), .Y(s[1]));
inv_hvt I147_0_ ( .A(s_b[0]), .Y(s[0]));
inv_hvt I25_2_ ( .A(sa_trim_b[2]), .Y(sa_trim[2]));
inv_hvt I25_1_ ( .A(sa_trim_b[1]), .Y(sa_trim[1]));
inv_hvt I25_0_ ( .A(sa_trim_b[0]), .Y(sa_trim[0]));
inv_hvt I24_2_ ( .A(net390[0]), .Y(sa_trim_b[2]));
inv_hvt I24_1_ ( .A(net390[1]), .Y(sa_trim_b[1]));
inv_hvt I24_0_ ( .A(net390[2]), .Y(sa_trim_b[0]));
mux2_hvt I180_1_ ( .in1(fsm_rowadd[1]), .in0(fsm_rowadd[1]),
     .out(net386[0]), .sel(fsm_nv_rrow));
mux2_hvt I180_0_ ( .in1(fsm_rowadd[0]), .in0(fsm_rowadd[0]),
     .out(net386[1]), .sel(fsm_nv_rrow));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net390[0]), .sel(net0365));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net390[1]), .sel(net0365));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net390[2]), .sel(net0365));
mux2_hvt I221 ( .in1(fsm_wpen), .in0(fsm_wgnden), .out(net0332),
     .sel(pgm_hvpulse));

endmodule
// Library - NVCM, Cell - ml_hv_invx3, View - schematic
// LAST TIME SAVED: Jan 25 09:27:09 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hv_invx3 ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M40 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_switch, View - schematic
// LAST TIME SAVED: Feb  1 16:53:01 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_lshv_6v_switch ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M4 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(gnd_), .G(vddp_tieh), .S(net132));
nch_25  M13 ( .D(net132), .B(gnd_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net140));
nch_25  M11 ( .D(net140), .B(gnd_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hv_ls_inv_hotsw, View - schematic
// LAST TIME SAVED: Jan 24 11:18:40 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hv_ls_inv_hotsw ( in_hv, out_b_hv, sel_25, sel_b_25,
     vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_invx3 Ihv_invx3 ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));
ml_lshv_6v_switch Ishv_6v_hold ( .vddp_tieh(vddp_tieh),
     .out_b_hv(net61), .in_hv(in_hv), .sel_b_25(sel_b_25),
     .sel_25(sel_25), .out_hv(sel_hv));

endmodule
// Library - NVCM, Cell - ml_hv_hotswitch, View - schematic
// LAST TIME SAVED: Jan 25 09:27:57 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hv_hotswitch ( hv_in_hv, hv_out_hv, selhv_25, vddp_tieh );
inout  hv_in_hv, hv_out_hv;

input  selhv_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_t_b), .in_hv(hv_in_hv),
     .vddp_tieh(vddp_tieh));
ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppb ( .sel_b_25(net35),
     .sel_25(selhv_25), .out_b_hv(sbhv_b_b), .in_hv(hv_out_hv),
     .vddp_tieh(vddp_tieh));
nch_25  M7 ( .D(net12), .B(GND_), .G(selhv_25), .S(net15));
nch_25  M1 ( .D(hv_in_hv), .B(GND_), .G(vddp_tieh), .S(net12));
nch_25  M2 ( .D(net15), .B(GND_), .G(vddp_tieh), .S(hv_out_hv));
pch_25  M0 ( .D(net26), .B(hv_out_hv), .G(sbhv_b_b), .S(hv_out_hv));
pch_25  M5 ( .D(net26), .B(hv_in_hv), .G(sbhv_t_b), .S(hv_in_hv));
inv_25 I114 ( .IN(selhv_25), .OUT(net35), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_hotswitch, View - schematic
// LAST TIME SAVED: Jan 26 19:35:53 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hvmux_hotswitch ( hvin_a_hv, hvin_b_hv, out_hv, sel_hv_a_25,
     sel_hv_b_25, vddp_tieh );
inout  hvin_a_hv, hvin_b_hv, out_hv;

input  sel_hv_a_25, sel_hv_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch Ihv_hotswitch_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_b_25), .hv_in_hv(hvin_b_hv), .hv_out_hv(out_hv));
ml_hv_hotswitch Ihv_hotswitch_vddp ( .vddp_tieh(vddp_tieh),
     .selhv_25(sel_hv_a_25), .hv_in_hv(hvin_a_hv), .hv_out_hv(out_hv));

endmodule
// Library - NVCM, Cell - ml_gwlwr_bldrv, View - schematic
// LAST TIME SAVED: Apr  9 11:04:12 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr_bldrv ( bgr, bl_pgm_glb, bl_frc_gnd, fsm_din, fsm_pgm,
     fsm_pgmien, fsm_trim_ipp, tm_dma );
inout  bgr, bl_pgm_glb;

input  bl_frc_gnd, fsm_din, fsm_pgm, fsm_pgmien, tm_dma;

input [3:0]  fsm_trim_ipp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net0152;

wire  [0:3]  net0172;

wire  [0:3]  net0156;

wire  [0:7]  net0115;

wire  [0:1]  net0180;

wire  [0:1]  net0160;



nand2_hvt I71 ( .B(fsm_din), .A(fsm_pgmien), .Y(fsm_pgmien_b_buf));
nor2_hvt I121 ( .A(net086), .B(fsm_pgmien_b_buf), .Y(pgm_trim0_en));
nor2_hvt I114 ( .B(tm_dma), .Y(net0116), .A(tm_dma));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
nor4_hvt I105 ( .D(fsm_trim_ipp[0]), .B(fsm_trim_ipp[2]), .Y(net086),
     .A(fsm_trim_ipp[3]), .C(fsm_trim_ipp[1]));
nch_hvt  M36 ( .D(net0173), .B(GND_), .G(pgm_trim0_en), .S(net0107));
nch_hvt  M37 ( .D(net0107), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M31_7_ ( .D(net0115[0]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[0]));
nch_hvt  M31_6_ ( .D(net0115[1]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[1]));
nch_hvt  M31_5_ ( .D(net0115[2]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[2]));
nch_hvt  M31_4_ ( .D(net0115[3]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[3]));
nch_hvt  M31_3_ ( .D(net0115[4]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[4]));
nch_hvt  M31_2_ ( .D(net0115[5]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[5]));
nch_hvt  M31_1_ ( .D(net0115[6]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[6]));
nch_hvt  M31_0_ ( .D(net0115[7]), .B(GND_), .G(fsm_trim_ipp[3]),
     .S(net0152[7]));
nch_hvt  M19 ( .D(net0135), .B(GND_), .G(fsm_trim_ipp[0]),
     .S(net0131));
nch_hvt  M38_7_ ( .D(net0152[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_6_ ( .D(net0152[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_5_ ( .D(net0152[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_4_ ( .D(net0152[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_3_ ( .D(net0152[4]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_2_ ( .D(net0152[5]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_1_ ( .D(net0152[6]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M38_0_ ( .D(net0152[7]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_3_ ( .D(net0156[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_2_ ( .D(net0156[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_1_ ( .D(net0156[2]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M39_0_ ( .D(net0156[3]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_1_ ( .D(net0160[0]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M40_0_ ( .D(net0160[1]), .B(GND_), .G(fsm_pgmien_buf),
     .S(gnd_));
nch_hvt  M26 ( .D(net0131), .B(GND_), .G(fsm_pgmien_buf), .S(gnd_));
nch_hvt  M33 ( .D(bl_pgm_glb), .B(GND_), .G(net0187), .S(gnd_));
nch_hvt  M30_3_ ( .D(net0172[0]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[0]));
nch_hvt  M30_2_ ( .D(net0172[1]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[1]));
nch_hvt  M30_1_ ( .D(net0172[2]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[2]));
nch_hvt  M30_0_ ( .D(net0172[3]), .B(GND_), .G(fsm_trim_ipp[2]),
     .S(net0156[3]));
nch_hvt  M34 ( .D(net089), .B(GND_), .G(pgm_trim0_en), .S(gnd_));
nch_hvt  M27_1_ ( .D(net0180[0]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[0]));
nch_hvt  M27_0_ ( .D(net0180[1]), .B(GND_), .G(fsm_trim_ipp[1]),
     .S(net0160[1]));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net0114), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net0114), .PLUS(net0141), .BULK(GND_));
inv_hvt I115 ( .A(net0116), .Y(net0187));
inv_hvt I58 ( .A(pgmen_b), .Y(pgmen));
inv_hvt I131 ( .A(fsm_pgm), .Y(pgmen_b));
inv_hvt I72 ( .A(fsm_pgmien_b_buf), .Y(fsm_pgmien_buf));
ml_ls_vdd2vdd25 I56 ( .in(pgmen), .sup(vddp_),
     .out_vddio_b(pgmen_b_25), .out_vddio(pgmen_25), .in_b(pgmen_b));
nch_25  M20 ( .D(net0173), .B(GND_), .G(pgm_inhi_bias),
     .S(bl_pgm_glb));
nch_25  M21 ( .D(pgm_inhi_bias), .B(GND_), .G(pgm_inhi_bias),
     .S(gnd_));
nch_25  M12_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[0]));
nch_25  M12_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0180[1]));
nch_25  M13_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[0]));
nch_25  M13_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[1]));
nch_25  M13_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[2]));
nch_25  M13_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0172[3]));
nch_25  M6 ( .D(net0164), .B(GND_), .G(net0164), .S(gnd_));
nch_25  M3 ( .D(dec_bias_p), .B(GND_), .G(bgr), .S(net0141));
nch_25  M10 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net089));
nch_25  M18_7_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[0]));
nch_25  M18_6_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[1]));
nch_25  M18_5_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[2]));
nch_25  M18_4_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[3]));
nch_25  M18_3_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[4]));
nch_25  M18_2_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[5]));
nch_25  M18_1_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[6]));
nch_25  M18_0_ ( .D(bl_pgm_glb), .B(GND_), .G(net0164),
     .S(net0115[7]));
nch_25  M9 ( .D(bl_pgm_glb), .B(GND_), .G(net0164), .S(net0135));
nch_25  M8 ( .D(net0164), .B(GND_), .G(pgmen_b_25), .S(gnd_));
pch_25  M11 ( .D(pgm_inhi_bias), .B(vddp_), .G(vdd_tieh), .S(net0259));
pch_25  M14_1_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M14_0_ ( .D(net0259), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M5 ( .D(net0164), .B(vddp_), .G(dec_bias_p), .S(net0199));
pch_25  M7_1_ ( .D(net0199), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M7_0_ ( .D(net0199), .B(vddp_), .G(pgmen_b_25), .S(vddp_));
pch_25  M4 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p), .S(net0199));

endmodule
// Library - io, Cell - pvpp, View - schematic
// LAST TIME SAVED: Jun  6 10:27:24 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module pvpp ( vpp, vppin );
inout  vpp, vppin;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



rppolywo_m  R1 ( .MINUS(vpp), .PLUS(vppin), .BULK(gnd_));
vddp_tiehigh I60 ( .vddp_tieh(net81));
vpp_clamp I59 ( .VSS(gnd_), .VDDIO(net81), .VPP(vpp));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_wr_sup, View - schematic
// LAST TIME SAVED: Jan 24 10:11:13 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_wr_sup ( wr_sup_25, wrsup_2vdd, wrsup_2vdd_25 );
inout  wr_sup_25;

input  wrsup_2vdd, wrsup_2vdd_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I120 ( .A(net19), .Y(wrsup_vdd_in));
inv_hvt I131 ( .A(wrsup_2vdd), .Y(net19));
inv_25 I119 ( .IN(net20), .OUT(wrsup_vdd_in_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(wrsup_2vdd_25), .OUT(net20), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_2_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_1_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));
ml_ymux_vblinhi_pgm_drv Iymux_vblinhi_pgm_drv_wr_0_ ( .ysup_25(vddp_),
     .en_blinhi_pgm_b_ysup_25(wrsup_vdd_in_25),
     .vblinhi_pgm_25(wr_sup_25), .en_blinhi_pgm_b(wrsup_vdd_in));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_ls25_1b, View - schematic
// LAST TIME SAVED: Jan 23 16:20:39 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25_1b ( out_25, in );
output  out_25;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I145 ( .A(in), .Y(net45));
inv_25 I153 ( .IN(out_b_25), .OUT(out_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I112 ( .in(in), .sup(vddp_), .out_vddio_b(out_b_25),
     .out_vddio(net025), .in_b(net45));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl_ls25, View - schematic
// LAST TIME SAVED: May  1 10:33:06 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl_ls25 ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25,
     gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25, s_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wrsup_2vdd_25, fsm_gwlbdis, gnv, gred, gwl_misc, gwl_nvcm,
     gwl_red, gwlb_dis, gwlb_en, gwlbsup_vddp, gwlbsup_vpxa,
     gwphv_vddp, gwphv_vppint, pgminhi_dmmy_b, s, testdec_en_b,
     testdec_even_b, testdec_odd_b, testdec_prec_b, wp_dis, wp_frcen,
     wr_dis, wr_frcen, wrsup_2vdd );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, gwlbsup_vddp_25, gwlbsup_vpxa_25,
     gwphv_vddp_25, gwphv_vppint_25, pgminhi_dmmy_b_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wrsup_2vdd_25;

input  fsm_gwlbdis, gwl_misc, gwl_nvcm, gwl_red, gwlb_dis, gwlb_en,
     gwlbsup_vddp, gwlbsup_vpxa, gwphv_vddp, gwphv_vppint,
     pgminhi_dmmy_b, testdec_en_b, testdec_even_b, testdec_odd_b,
     testdec_prec_b, wp_dis, wp_frcen, wr_dis, wr_frcen, wrsup_2vdd;

output [5:0]  gnv_b_25;
output [3:0]  s_25;
output [1:0]  gred_25;
output [5:0]  gnv_25;
output [1:0]  gred_b_25;

input [5:0]  gnv;
input [3:0]  s;
input [1:0]  gred;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I_1_ ( .IN(gred_25[1]), .OUT(gred_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I_0_ ( .IN(gred_25[0]), .OUT(gred_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I143 ( .IN(net101), .OUT(fsm_gwlbdis_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_5_ ( .IN(gnv_25[5]), .OUT(gnv_b_25[5]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_4_ ( .IN(gnv_25[4]), .OUT(gnv_b_25[4]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_3_ ( .IN(gnv_25[3]), .OUT(gnv_b_25[3]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_2_ ( .IN(gnv_25[2]), .OUT(gnv_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_1_ ( .IN(gnv_25[1]), .OUT(gnv_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_0_ ( .IN(gnv_25[0]), .OUT(gnv_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
ml_gwlwr_ctrl_ls25_1b I133 ( .in(testdec_en_b),
     .out_25(testdec_en_b_25));
ml_gwlwr_ctrl_ls25_1b I139 ( .in(gwlb_dis), .out_25(gwlb_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_frcen ( .in(wr_frcen),
     .out_25(wr_frcen_25));
ml_gwlwr_ctrl_ls25_1b I144 ( .in(gwlb_en), .out_25(gwlb_en_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vpp ( .in(gwphv_vppint),
     .out_25(gwphv_vppint_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwlb_vddp ( .in(gwlbsup_vddp),
     .out_25(gwlbsup_vddp_25));
ml_gwlwr_ctrl_ls25_1b ls25_gwlb_vpp ( .in(gwlbsup_vpxa),
     .out_25(gwlbsup_vpxa_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_vdd ( .in(wrsup_2vdd),
     .out_25(wrsup_2vdd_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wr_dis ( .in(wr_dis), .out_25(wr_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwphv_vddp ( .in(gwphv_vddp),
     .out_25(gwphv_vddp_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_frcen ( .in(wp_frcen),
     .out_25(wp_frcen_25));
ml_gwlwr_ctrl_ls25_1b Ils25_wp_dis ( .in(wp_dis), .out_25(wp_dis_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gwl_red ( .in(gwl_red),
     .out_25(gwl_red_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_nvcm ( .in(gwl_nvcm),
     .out_25(gwl_nvcm_25));
ml_gwlwr_ctrl_ls25_1b Ils25_glw_misc ( .in(gwl_misc),
     .out_25(gwl_misc_25));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_1_ ( .in(gred[1]),
     .out_25(gred_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gred_0_ ( .in(gred[0]),
     .out_25(gred_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_5_ ( .in(gnv[5]), .out_25(gnv_25[5]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_4_ ( .in(gnv[4]), .out_25(gnv_25[4]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_3_ ( .in(gnv[3]), .out_25(gnv_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_2_ ( .in(gnv[2]), .out_25(gnv_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_1_ ( .in(gnv[1]), .out_25(gnv_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_gnv_0_ ( .in(gnv[0]), .out_25(gnv_25[0]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_3_ ( .in(s[3]), .out_25(s_25[3]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_2_ ( .in(s[2]), .out_25(s_25[2]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_1_ ( .in(s[1]), .out_25(s_25[1]));
ml_gwlwr_ctrl_ls25_1b Ils25_s_0_ ( .in(s[0]), .out_25(s_25[0]));
ml_gwlwr_ctrl_ls25_1b I134 ( .in(testdec_prec_b),
     .out_25(testdec_prec_b_25));
ml_gwlwr_ctrl_ls25_1b I136 ( .in(pgminhi_dmmy_b),
     .out_25(pgminhi_dmmy_b_25));
ml_gwlwr_ctrl_ls25_1b I140 ( .in(fsm_gwlbdis), .out_25(net101));
ml_gwlwr_ctrl_ls25_1b I137 ( .in(testdec_even_b),
     .out_25(testdec_even_b_25));
ml_gwlwr_ctrl_ls25_1b I138 ( .in(testdec_odd_b),
     .out_25(testdec_odd_b_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_npgate_gen, View - schematic
// LAST TIME SAVED: Sep 15 17:15:47 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_core_sa_npgate_gen ( dec_trim, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, vpxa, fsm_tm_testdec, saen, satrim,
     vddp_tieh );
output  saen_25, saen_b_vpxa;

inout  vpxa;

input  fsm_tm_testdec, saen, vddp_tieh;

output [4:1]  sa_ngate_25;
output [4:1]  sa_pgate_vpxa;
output [7:0]  dec_trim;

input [2:0]  satrim;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net0122;

wire  [4:1]  trim_b;

wire  [4:1]  pgate_in;

wire  [7:0]  dec_trim_b;

wire  [0:3]  net48;

wire  [0:3]  net53;

wire  [4:1]  ngate_in_25_b;

wire  [2:0]  ydec_b;

wire  [2:0]  ydec;

wire  [4:1]  trim;



nor4_hvt I102 ( .D(fsm_tm_testdec), .C(dec_trim[7]), .A(dec_trim[5]),
     .B(dec_trim[6]), .Y(net47));
ml_hv_invx3 I135 ( .sel_hv(net048), .sel_25(net048),
     .vddp_tieh(vddp_tieh), .out_b_hv(saen_b_vpxa), .in_hv(vpxa));
ml_hv_invx3 I130_4_ ( .sel_hv(pgate_in[4]), .sel_25(pgate_in[4]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[4]), .in_hv(vpxa));
ml_hv_invx3 I130_3_ ( .sel_hv(pgate_in[3]), .sel_25(pgate_in[3]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[3]), .in_hv(vpxa));
ml_hv_invx3 I130_2_ ( .sel_hv(pgate_in[2]), .sel_25(pgate_in[2]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[2]), .in_hv(vpxa));
ml_hv_invx3 I130_1_ ( .sel_hv(pgate_in[1]), .sel_25(pgate_in[1]),
     .vddp_tieh(vddp_tieh), .out_b_hv(sa_pgate_vpxa[1]), .in_hv(vpxa));
inv_25 I149 ( .IN(net052), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I153_4_ ( .IN(ngate_in_25_b[4]), .OUT(sa_ngate_25[4]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_3_ ( .IN(ngate_in_25_b[3]), .OUT(sa_ngate_25[3]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_2_ ( .IN(ngate_in_25_b[2]), .OUT(sa_ngate_25[2]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I153_1_ ( .IN(ngate_in_25_b[1]), .OUT(sa_ngate_25[1]),
     .P(vddp_), .Pb(vddp_), .G(gnd_), .Gb(gnd_));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec[2]));
nand3_hvt I37_4_ ( .Y(dec_trim_b[4]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec[2]));
nand3_hvt I37_3_ ( .Y(dec_trim_b[3]), .B(ydec[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_2_ ( .Y(dec_trim_b[2]), .B(ydec[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nand3_hvt I37_1_ ( .Y(dec_trim_b[1]), .B(ydec_b[1]), .C(ydec[0]),
     .A(ydec_b[2]));
nand3_hvt I37_0_ ( .Y(dec_trim_b[0]), .B(ydec_b[1]), .C(ydec_b[0]),
     .A(ydec_b[2]));
nor2_hvt I75_4_ ( .Y(net48[0]), .B(dec_trim[4]), .A(sa_high_res));
nor2_hvt I75_3_ ( .Y(net48[1]), .B(dec_trim[3]), .A(trim[4]));
nor2_hvt I75_2_ ( .Y(net48[2]), .B(dec_trim[2]), .A(trim[3]));
nor2_hvt I75_1_ ( .Y(net48[3]), .B(dec_trim[1]), .A(trim[2]));
inv_hvt I145 ( .A(net076), .Y(net078));
inv_hvt I143 ( .A(net078), .Y(net080));
inv_hvt I146 ( .A(saen), .Y(net076));
inv_hvt I114 ( .A(net47), .Y(sa_high_res));
inv_hvt I38_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I38_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I38_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I38_4_ ( .A(dec_trim_b[4]), .Y(dec_trim[4]));
inv_hvt I38_3_ ( .A(dec_trim_b[3]), .Y(dec_trim[3]));
inv_hvt I38_2_ ( .A(dec_trim_b[2]), .Y(dec_trim[2]));
inv_hvt I38_1_ ( .A(dec_trim_b[1]), .Y(dec_trim[1]));
inv_hvt I38_0_ ( .A(dec_trim_b[0]), .Y(dec_trim[0]));
inv_hvt I40_2_ ( .A(ydec_b[2]), .Y(ydec[2]));
inv_hvt I40_1_ ( .A(ydec_b[1]), .Y(ydec[1]));
inv_hvt I40_0_ ( .A(ydec_b[0]), .Y(ydec[0]));
inv_hvt I76_4_ ( .A(net48[0]), .Y(trim[4]));
inv_hvt I76_3_ ( .A(net48[1]), .Y(trim[3]));
inv_hvt I76_2_ ( .A(net48[2]), .Y(trim[2]));
inv_hvt I76_1_ ( .A(net48[3]), .Y(trim[1]));
inv_hvt I39_2_ ( .A(satrim[2]), .Y(ydec_b[2]));
inv_hvt I39_1_ ( .A(satrim[1]), .Y(ydec_b[1]));
inv_hvt I39_0_ ( .A(satrim[0]), .Y(ydec_b[0]));
inv_hvt I78_4_ ( .A(trim[4]), .Y(trim_b[4]));
inv_hvt I78_3_ ( .A(trim[3]), .Y(trim_b[3]));
inv_hvt I78_2_ ( .A(trim[2]), .Y(trim_b[2]));
inv_hvt I78_1_ ( .A(trim[1]), .Y(trim_b[1]));
ml_ls_vdd2vdd25 I128_4_ ( .in(ngate_in_25_b[4]), .sup(vpxa),
     .out_vddio_b(pgate_in[4]), .out_vddio(net53[0]),
     .in_b(net0122[0]));
ml_ls_vdd2vdd25 I128_3_ ( .in(ngate_in_25_b[3]), .sup(vpxa),
     .out_vddio_b(pgate_in[3]), .out_vddio(net53[1]),
     .in_b(net0122[1]));
ml_ls_vdd2vdd25 I128_2_ ( .in(ngate_in_25_b[2]), .sup(vpxa),
     .out_vddio_b(pgate_in[2]), .out_vddio(net53[2]),
     .in_b(net0122[2]));
ml_ls_vdd2vdd25 I128_1_ ( .in(ngate_in_25_b[1]), .sup(vpxa),
     .out_vddio_b(pgate_in[1]), .out_vddio(net53[3]),
     .in_b(net0122[3]));
ml_ls_vdd2vdd25 I136 ( .in(net053), .sup(vpxa), .out_vddio_b(net047),
     .out_vddio(net048), .in_b(net052));
ml_ls_vdd2vdd25 I137 ( .in(net078), .sup(vddp_), .out_vddio_b(net052),
     .out_vddio(net053), .in_b(net080));
ml_ls_vdd2vdd25 I129_4_ ( .in(trim[4]), .sup(vddp_),
     .out_vddio_b(net0122[0]), .out_vddio(ngate_in_25_b[4]),
     .in_b(trim_b[4]));
ml_ls_vdd2vdd25 I129_3_ ( .in(trim[3]), .sup(vddp_),
     .out_vddio_b(net0122[1]), .out_vddio(ngate_in_25_b[3]),
     .in_b(trim_b[3]));
ml_ls_vdd2vdd25 I129_2_ ( .in(trim[2]), .sup(vddp_),
     .out_vddio_b(net0122[2]), .out_vddio(ngate_in_25_b[2]),
     .in_b(trim_b[2]));
ml_ls_vdd2vdd25 I129_1_ ( .in(trim[1]), .sup(vddp_),
     .out_vddio_b(net0122[3]), .out_vddio(ngate_in_25_b[1]),
     .in_b(trim_b[1]));

endmodule
// Library - NVCM, Cell - ml_gwlwr_ctrl, View - schematic
// LAST TIME SAVED: May  1 11:11:08 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr_ctrl ( fsm_gwlbdis_b_25, gnv_25, gnv_b_25, gred_25,
     gred_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25,
     gwlb_en_25, pgminhi_dmmy_b_25, s_25, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b_25, wp_dis_25, wp_frcen_25,
     wr_dis_25, wr_frcen_25, bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv,
     vddp_tieh, vpp_int, vpxa, wr_sup_25, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_misc_25, gwl_nvcm_25, gwl_red_25,
     gwlb_dis_25, gwlb_en_25, pgminhi_dmmy_b_25, saen_25, saen_b_vpxa,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

inout  bgr, bl_pgm_glb, gwl_b_sup_25, gwp_sup_hv, vddp_tieh, vpp_int,
     vpxa, wr_sup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [5:0]  gnv_25;
output [5:0]  gnv_b_25;
output [1:0]  gred_25;
output [4:1]  sa_ngate_25;
output [3:0]  s_25;
output [1:0]  gred_b_25;
output [4:1]  sa_pgate_vpxa;

input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
input [0:0]  fsm_coladd;
input [3:0]  fsm_trim_ipp;
input [7:0]  fsm_rowadd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  sa_trim;

wire  [3:0]  s;

wire  [1:0]  gred;

wire  [5:0]  gnv;

wire  [7:0]  dec_trim;



ml_hvmux_hotswitch_enhance Ihvmux_gwpsup_hv ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwphv_vppint_25), .sel_hv_a_25(gwphv_vddp_25),
     .out_hv(gwp_sup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_gwlwr_ctrl_logic Igwlwr_ctrl_logic ( .fsm_pgmdisc(fsm_pgmdisc),
     .gwlb_en(gwlb_en), .tm_testdec_wr(tm_testdec_wr),
     .tm_testdec(tm_testdec), .tm_dma(tm_dma),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_trow(fsm_tm_trow), .fsm_tm_allwl_l(fsm_tm_allwl_l),
     .fsm_tm_allwl_h(fsm_tm_allwl_h), .fsm_tm_allbl_l(fsm_tm_allbl_l),
     .fsm_tm_allbl_h(fsm_tm_allbl_h), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_rd(fsm_rd), .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmhv(fsm_pgmhv),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_coladd(fsm_coladd[0]), .wrsup_2vdd(wrsup_2vdd),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .testdec_prec_b(net172),
     .testdec_odd_b(testdec_odd_b), .testdec_even_b(testdec_even_b),
     .testdec_en_b(net175), .saen(saen), .sa_trim(sa_trim[2:0]),
     .s(s[3:0]), .pgminhi_dmmy_b(net179), .gwphv_vppint(gwphv_vppint),
     .gwphv_vddp(gwphv_vddp), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vddp(gwlbsup_vddp), .gwlb_dis(gwlb_dis),
     .gwl_misc(gwl_misc), .gred(gred[1:0]), .gnv(gnv[5:0]));
ml_hvmux_hotswitch Ihvmux_gwlbsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(gwlbsup_vpxa_25), .sel_hv_a_25(gwlbsup_vddp_25),
     .out_hv(gwl_b_sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_gwlwr_bldrv Igwlwr_bldrv ( .fsm_din(fsm_din), .tm_dma(tm_dma),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_pgmien(fsm_pgmien),
     .fsm_pgm(fsm_pgm), .bl_frc_gnd(gnd_), .bgr(bgr),
     .bl_pgm_glb(bl_pgm_glb));
ml_gwlwr_ctrl_wr_sup Igwlwr_ctrl_wr_sup ( .wrsup_2vdd(wrsup_2vdd),
     .wrsup_2vdd_25(wrsup_2vdd_25), .wr_sup_25(wr_sup_25));
ml_gwlwr_ctrl_ls25 Igwlwr_ctrl_ls25 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_en(gwlb_en), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwlb_dis(gwlb_dis), .gwlbsup_vpxa(gwlbsup_vpxa),
     .gwlbsup_vpxa_25(gwlbsup_vpxa_25), .wrsup_2vdd_25(wrsup_2vdd_25),
     .wrsup_2vdd(wrsup_2vdd), .testdec_odd_b(testdec_odd_b),
     .testdec_even_b(testdec_even_b),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25), .testdec_prec_b(net172),
     .testdec_en_b(net175), .pgminhi_dmmy_b(net179),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwphv_vddp(gwphv_vddp),
     .gwlbsup_vddp(gwlbsup_vddp), .gwphv_vppint(gwphv_vppint),
     .gwlbsup_vddp_25(gwlbsup_vddp_25),
     .gwphv_vppint_25(gwphv_vppint_25), .gwphv_vddp_25(gwphv_vddp_25),
     .wr_frcen(wr_frcen), .wr_dis(wr_dis), .wp_frcen(wp_frcen),
     .wp_dis(wp_dis), .s(s[3:0]), .gwl_red(fsm_nv_rrow),
     .gwl_nvcm(fsm_nv_bstream), .gwl_misc(gwl_misc), .gred(gred[1:0]),
     .gnv(gnv[5:0]), .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]));
vddp_tiehigh Ivddp_tiehigh_15_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_14_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_13_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_12_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_11_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_10_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_9_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_8_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh Ivddp_tiehigh_0_ ( .vddp_tieh(vddp_tieh));
ml_core_sa_npgate_gen Icore_sa_npgate_gen (
     .fsm_tm_testdec(tm_testdec), .satrim(sa_trim[2:0]),
     .vddp_tieh(vddp_tieh), .saen(saen), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .dec_trim(dec_trim[7:0]),
     .vpxa(vpxa));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr, View - schematic
// LAST TIME SAVED: Feb 25 14:20:48 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr ( wr, gwl_wr_25, s_25, wr_sup_25 );
output  wr;

input  gwl_wr_25, s_25, wr_sup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_25 I59 ( .A(gwl_wr_25), .Y(net27), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(s_25));
inv_25 I38 ( .IN(net27), .OUT(wr), .P(wr_sup_25), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr_x4, View - schematic
// LAST TIME SAVED: Jan 21 18:09:38 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x4 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  gwl_wr_25, wr_sup_25;

output [3:0]  wr;

input [3:0]  s_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr Iml_lwldrv_2 ( .gwl_wr_25(gwl_wr_25), .wr(wr[2]),
     .s_25(s_25[2]), .wr_sup_25(wr_sup_25));
ml_rock_lwldrv_wr Iml_lwldrv_1 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[1]), .wr(wr[1]));
ml_rock_lwldrv_wr Iml_lwldrv_3 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[3]), .wr(wr[3]));
ml_rock_lwldrv_wr Iml_lwldrv_0 ( .gwl_wr_25(gwl_wr_25),
     .wr_sup_25(wr_sup_25), .s_25(s_25[0]), .wr(wr[0]));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wr_x228, View - schematic
// LAST TIME SAVED: Jan 23 13:37:56 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wr_x228 ( wr, gwl_wr_25, s_25, wr_sup_25 );

input  wr_sup_25;

output [227:0]  wr;

input [56:0]  gwl_wr_25;
input [3:0]  s_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_56_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[227:224]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[56]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_55_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[223:220]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[55]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_54_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[219:216]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[54]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_53_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[215:212]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[53]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_52_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[211:208]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[52]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_51_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[207:204]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[51]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_50_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[203:200]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[50]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_49_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[199:196]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[49]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_48_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[195:192]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[48]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_47_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[191:188]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[47]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_46_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[187:184]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[46]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_45_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[183:180]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[45]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_44_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[179:176]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[44]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_43_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[175:172]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[43]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_42_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[171:168]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[42]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_41_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[167:164]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[41]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_40_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[163:160]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[40]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_39_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[159:156]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[39]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_38_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[155:152]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[38]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_37_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[151:148]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[37]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_36_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[147:144]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[36]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_35_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[143:140]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[35]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_34_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[139:136]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[34]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_33_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[135:132]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[33]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_32_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[131:128]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[32]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_31_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[127:124]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[31]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_30_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[123:120]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[30]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_29_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[119:116]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[29]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_28_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[115:112]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[28]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_27_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[111:108]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[27]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_26_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[107:104]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[26]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_25_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[103:100]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[25]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_24_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[99:96]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[24]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_23_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[95:92]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[23]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_22_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[91:88]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[22]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_21_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[87:84]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[21]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_20_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[83:80]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[20]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_19_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[79:76]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[19]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_18_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[75:72]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[18]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_17_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[71:68]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[17]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_16_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[67:64]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[16]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_15_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[63:60]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[15]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_14_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[59:56]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[14]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_13_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[55:52]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[13]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_12_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[51:48]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[12]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_11_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[47:44]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[11]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_10_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[43:40]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[10]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_9_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[39:36]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[9]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_8_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[35:32]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[8]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_7_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[31:28]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[7]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_6_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[27:24]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[6]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_5_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[23:20]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[5]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_4_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[19:16]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[4]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_3_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[15:12]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[3]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_2_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[11:8]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[2]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_1_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[7:4]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[1]));
ml_rock_lwldrv_wr_x4 Ilwldrv_wr_x4_0_ ( .wr_sup_25(wr_sup_25),
     .wr(wr[3:0]), .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[0]));

endmodule
// Library - NVCM, Cell - ml_ls_vddp2vpxa, View - schematic
// LAST TIME SAVED: Dec 30 20:36:23 2007
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_ls_vddp2vpxa ( out_33, out_b_33, sup, in_25, in_b_25 );
output  out_33, out_b_33;

inout  sup;

input  in_25, in_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(out_b_33), .B(sup), .G(in_25), .S(net29));
pch_25  M13 ( .D(out_33), .B(sup), .G(in_b_25), .S(net33));
pch_25  M4 ( .D(net29), .B(sup), .G(out_33), .S(sup));
pch_25  M6 ( .D(net33), .B(sup), .G(out_b_33), .S(sup));
nch_25  M9 ( .D(out_33), .B(gnd_), .G(in_b_25), .S(gnd_));
nch_25  M15 ( .D(out_b_33), .B(gnd_), .G(in_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_gwhv, View - schematic
// LAST TIME SAVED: May 16 11:27:16 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_gwhv ( gwp_hv, gwp_sup_hv, gwl_25, gwl_25_b,
     vddp_tieh );
output  gwp_hv;

inout  gwp_sup_hv;

input  gwl_25, gwl_25_b, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M10 ( .D(net0129), .B(gnd_), .G(vddp_tieh), .S(net050));
nch_25  M12 ( .D(gwp_hv), .B(gnd_), .G(vddp_tieh), .S(net034));
nch_25  M11 ( .D(net034), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M13 ( .D(net050), .B(gnd_), .G(gwl_25_b), .S(gnd_));
nch_25  M14 ( .D(net054), .B(gnd_), .G(vddp_tieh), .S(net058));
nch_25  M15 ( .D(net058), .B(gnd_), .G(gwl_25), .S(gnd_));
pch_25  M6 ( .D(net067), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M16 ( .D(gwp_hv), .B(net067), .G(gwl_25_b), .S(net067));
pch_25  M5 ( .D(net054), .B(net087), .G(gwl_25), .S(net087));
pch_25  M8 ( .D(net087), .B(gwp_sup_hv), .G(net0129), .S(gwp_sup_hv));
pch_25  M9 ( .D(net091), .B(gwp_sup_hv), .G(net054), .S(gwp_sup_hv));
pch_25  M7 ( .D(net0129), .B(net091), .G(gwl_25_b), .S(net091));

endmodule
// Library - io, Cell - topbank_f, View - schematic
// LAST TIME SAVED: Jun  6 10:46:50 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module topbank_f ( in, pad, vpp, vppin, oen, out, ren );

inout  vpp, vppin;


output [59:0]  in;

inout [59:0]  pad;

input [59:0]  out;
input [59:0]  oen;
input [59:0]  ren;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pvpp I62 ( .vppin(vppin), .vpp(vpp));
PDUW08DGZ I45_43_ ( .PAD(pad[43]), .C(in[43]), .OEN(oen[43]),
     .I(out[43]), .REN(ren[43]));
PDUW08DGZ I45_42_ ( .PAD(pad[42]), .C(in[42]), .OEN(oen[42]),
     .I(out[42]), .REN(ren[42]));
PDUW08DGZ I45_41_ ( .PAD(pad[41]), .C(in[41]), .OEN(oen[41]),
     .I(out[41]), .REN(ren[41]));
PDUW08DGZ I45_40_ ( .PAD(pad[40]), .C(in[40]), .OEN(oen[40]),
     .I(out[40]), .REN(ren[40]));
PDUW08DGZ I45_39_ ( .PAD(pad[39]), .C(in[39]), .OEN(oen[39]),
     .I(out[39]), .REN(ren[39]));
PDUW08DGZ I45_38_ ( .PAD(pad[38]), .C(in[38]), .OEN(oen[38]),
     .I(out[38]), .REN(ren[38]));
PDUW08DGZ I45_37_ ( .PAD(pad[37]), .C(in[37]), .OEN(oen[37]),
     .I(out[37]), .REN(ren[37]));
PDUW08DGZ I45_36_ ( .PAD(pad[36]), .C(in[36]), .OEN(oen[36]),
     .I(out[36]), .REN(ren[36]));
PDUW08DGZ I45_35_ ( .PAD(pad[35]), .C(in[35]), .OEN(oen[35]),
     .I(out[35]), .REN(ren[35]));
PDUW08DGZ I45_34_ ( .PAD(pad[34]), .C(in[34]), .OEN(oen[34]),
     .I(out[34]), .REN(ren[34]));
PDUW08DGZ I46_19_ ( .PAD(pad[19]), .C(in[19]), .OEN(oen[19]),
     .I(out[19]), .REN(ren[19]));
PDUW08DGZ I46_18_ ( .PAD(pad[18]), .C(in[18]), .OEN(oen[18]),
     .I(out[18]), .REN(ren[18]));
PDUW08DGZ I46_17_ ( .PAD(pad[17]), .C(in[17]), .OEN(oen[17]),
     .I(out[17]), .REN(ren[17]));
PDUW08DGZ I46_16_ ( .PAD(pad[16]), .C(in[16]), .OEN(oen[16]),
     .I(out[16]), .REN(ren[16]));
PDUW08DGZ I46_15_ ( .PAD(pad[15]), .C(in[15]), .OEN(oen[15]),
     .I(out[15]), .REN(ren[15]));
PDUW08DGZ I46_14_ ( .PAD(pad[14]), .C(in[14]), .OEN(oen[14]),
     .I(out[14]), .REN(ren[14]));
PDUW08DGZ I46_13_ ( .PAD(pad[13]), .C(in[13]), .OEN(oen[13]),
     .I(out[13]), .REN(ren[13]));
PDUW08DGZ I46_12_ ( .PAD(pad[12]), .C(in[12]), .OEN(oen[12]),
     .I(out[12]), .REN(ren[12]));
PDUW08DGZ I46_11_ ( .PAD(pad[11]), .C(in[11]), .OEN(oen[11]),
     .I(out[11]), .REN(ren[11]));
PDUW08DGZ I47_51_ ( .PAD(pad[51]), .C(in[51]), .OEN(oen[51]),
     .I(out[51]), .REN(ren[51]));
PDUW08DGZ I47_50_ ( .PAD(pad[50]), .C(in[50]), .OEN(oen[50]),
     .I(out[50]), .REN(ren[50]));
PDUW08DGZ I47_49_ ( .PAD(pad[49]), .C(in[49]), .OEN(oen[49]),
     .I(out[49]), .REN(ren[49]));
PDUW08DGZ I47_48_ ( .PAD(pad[48]), .C(in[48]), .OEN(oen[48]),
     .I(out[48]), .REN(ren[48]));
PDUW08DGZ I47_47_ ( .PAD(pad[47]), .C(in[47]), .OEN(oen[47]),
     .I(out[47]), .REN(ren[47]));
PDUW08DGZ I47_46_ ( .PAD(pad[46]), .C(in[46]), .OEN(oen[46]),
     .I(out[46]), .REN(ren[46]));
PDUW08DGZ I47_45_ ( .PAD(pad[45]), .C(in[45]), .OEN(oen[45]),
     .I(out[45]), .REN(ren[45]));
PDUW08DGZ I47_44_ ( .PAD(pad[44]), .C(in[44]), .OEN(oen[44]),
     .I(out[44]), .REN(ren[44]));
PDUW08DGZ I50_27_ ( .PAD(pad[27]), .C(in[27]), .OEN(oen[27]),
     .I(out[27]), .REN(ren[27]));
PDUW08DGZ I50_26_ ( .PAD(pad[26]), .C(in[26]), .OEN(oen[26]),
     .I(out[26]), .REN(ren[26]));
PDUW08DGZ I50_25_ ( .PAD(pad[25]), .C(in[25]), .OEN(oen[25]),
     .I(out[25]), .REN(ren[25]));
PDUW08DGZ I50_24_ ( .PAD(pad[24]), .C(in[24]), .OEN(oen[24]),
     .I(out[24]), .REN(ren[24]));
PDUW08DGZ I48_23_ ( .PAD(pad[23]), .C(in[23]), .OEN(oen[23]),
     .I(out[23]), .REN(ren[23]));
PDUW08DGZ I48_22_ ( .PAD(pad[22]), .C(in[22]), .OEN(oen[22]),
     .I(out[22]), .REN(ren[22]));
PDUW08DGZ I48_21_ ( .PAD(pad[21]), .C(in[21]), .OEN(oen[21]),
     .I(out[21]), .REN(ren[21]));
PDUW08DGZ I48_20_ ( .PAD(pad[20]), .C(in[20]), .OEN(oen[20]),
     .I(out[20]), .REN(ren[20]));
PDUW08DGZ I49_54_ ( .PAD(pad[54]), .C(in[54]), .OEN(oen[54]),
     .I(out[54]), .REN(ren[54]));
PDUW08DGZ I49_53_ ( .PAD(pad[53]), .C(in[53]), .OEN(oen[53]),
     .I(out[53]), .REN(ren[53]));
PDUW08DGZ I49_52_ ( .PAD(pad[52]), .C(in[52]), .OEN(oen[52]),
     .I(out[52]), .REN(ren[52]));
PDUW08DGZ I51_59_ ( .PAD(pad[59]), .C(in[59]), .OEN(oen[59]),
     .I(out[59]), .REN(ren[59]));
PDUW08DGZ I51_58_ ( .PAD(pad[58]), .C(in[58]), .OEN(oen[58]),
     .I(out[58]), .REN(ren[58]));
PDUW08DGZ I51_57_ ( .PAD(pad[57]), .C(in[57]), .OEN(oen[57]),
     .I(out[57]), .REN(ren[57]));
PDUW08DGZ I51_56_ ( .PAD(pad[56]), .C(in[56]), .OEN(oen[56]),
     .I(out[56]), .REN(ren[56]));
PDUW08DGZ I51_55_ ( .PAD(pad[55]), .C(in[55]), .OEN(oen[55]),
     .I(out[55]), .REN(ren[55]));
PDUW08DGZ I42_4_ ( .PAD(pad[4]), .C(in[4]), .OEN(oen[4]), .I(out[4]),
     .REN(ren[4]));
PDUW08DGZ I42_3_ ( .PAD(pad[3]), .C(in[3]), .OEN(oen[3]), .I(out[3]),
     .REN(ren[3]));
PDUW08DGZ I42_2_ ( .PAD(pad[2]), .C(in[2]), .OEN(oen[2]), .I(out[2]),
     .REN(ren[2]));
PDUW08DGZ I42_1_ ( .PAD(pad[1]), .C(in[1]), .OEN(oen[1]), .I(out[1]),
     .REN(ren[1]));
PDUW08DGZ I42_0_ ( .PAD(pad[0]), .C(in[0]), .OEN(oen[0]), .I(out[0]),
     .REN(ren[0]));
PDUW08DGZ I43_33_ ( .PAD(pad[33]), .C(in[33]), .OEN(oen[33]),
     .I(out[33]), .REN(ren[33]));
PDUW08DGZ I43_32_ ( .PAD(pad[32]), .C(in[32]), .OEN(oen[32]),
     .I(out[32]), .REN(ren[32]));
PDUW08DGZ I43_31_ ( .PAD(pad[31]), .C(in[31]), .OEN(oen[31]),
     .I(out[31]), .REN(ren[31]));
PDUW08DGZ I43_30_ ( .PAD(pad[30]), .C(in[30]), .OEN(oen[30]),
     .I(out[30]), .REN(ren[30]));
PDUW08DGZ I43_29_ ( .PAD(pad[29]), .C(in[29]), .OEN(oen[29]),
     .I(out[29]), .REN(ren[29]));
PDUW08DGZ I43_28_ ( .PAD(pad[28]), .C(in[28]), .OEN(oen[28]),
     .I(out[28]), .REN(ren[28]));
PDUW08DGZ I44_10_ ( .PAD(pad[10]), .C(in[10]), .OEN(oen[10]),
     .I(out[10]), .REN(ren[10]));
PDUW08DGZ I44_9_ ( .PAD(pad[9]), .C(in[9]), .OEN(oen[9]), .I(out[9]),
     .REN(ren[9]));
PDUW08DGZ I44_8_ ( .PAD(pad[8]), .C(in[8]), .OEN(oen[8]), .I(out[8]),
     .REN(ren[8]));
PDUW08DGZ I44_7_ ( .PAD(pad[7]), .C(in[7]), .OEN(oen[7]), .I(out[7]),
     .REN(ren[7]));
PDUW08DGZ I44_6_ ( .PAD(pad[6]), .C(in[6]), .OEN(oen[6]), .I(out[6]),
     .REN(ren[6]));
PDUW08DGZ I44_5_ ( .PAD(pad[5]), .C(in[5]), .OEN(oen[5]), .I(out[5]),
     .REN(ren[5]));
PVDD2POC I35 ( .VDDPST(vddio_topbank));
PVDD1DGZ I58_1_ ( .VDD(vdd_));
PVDD1DGZ I58_0_ ( .VDD(vdd_));
PVDD1DGZ I34_1_ ( .VDD(vdd_));
PVDD1DGZ I34_0_ ( .VDD(vdd_));
PVDD2DGZ I57 ( .VDDPST(vddio_topbank));
PVDD2DGZ I33_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ I33_0_ ( .VDDPST(vddio_topbank));
PVDD2DGZ I53_1_ ( .VDDPST(vddio_topbank));
PVDD2DGZ I53_0_ ( .VDDPST(vddio_topbank));
PVDD2DGZ I55 ( .VDDPST(vddio_topbank));
PVSS3DGZ I56_1_ ( .VSS(gnd_));
PVSS3DGZ I56_0_ ( .VSS(gnd_));
PVSS3DGZ I32_1_ ( .VSS(gnd_));
PVSS3DGZ I32_0_ ( .VSS(gnd_));
PVSS3DGZ I54_1_ ( .VSS(gnd_));
PVSS3DGZ I54_0_ ( .VSS(gnd_));
PVSS3DGZ I52_1_ ( .VSS(gnd_));
PVSS3DGZ I52_0_ ( .VSS(gnd_));

endmodule
// Library - NVCM, Cell - ml_gwl_drv, View - schematic
// LAST TIME SAVED: Apr 30 15:58:52 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwl_drv ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25,
     radd_1_25, radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );
output  gwl_b_25, gwl_wr_25, gwp_hv;

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwlb_dis_25, gwlb_en_25, gwlgrpsel_25, radd_0_25, radd_1_25,
     radd_2_25, radd_3_25, radd_4_25, radd_5_25, radd_6_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_ls_vddp2vpxa I99 ( .in_25(gwlb_25), .sup(gwl_b_sup_25),
     .in_b_25(gwlb_b_25), .out_33(out_33), .out_b_33(net053));
nor3_25 I76 ( .C(net84), .A(net68), .Y(dec_sel_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(net76));
nor2_25 I111 ( .A(net096), .Y(gwlb_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_dis_25));
nor2_25 I79 ( .A(wr_dis_25), .Y(gwl_wr_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(net056));
nor2_25 I117 ( .A(dec_sel_25), .Y(net096), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(gwlb_en_25));
nor2_25 I82 ( .A(dec_sel_25), .Y(net058), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_frcen_25));
nor2_25 I85 ( .A(net058), .Y(gwl_wp_25), .Gb(gnd_), .G(gnd_),
     .Pb(vddp_), .P(vddp_), .B(wp_dis_25));
nor2_25 I59 ( .B(dec_sel_25), .A(wr_frcen_25), .Y(net056), .P(vddp_),
     .Pb(vddp_), .Gb(gnd_), .G(gnd_));
ml_rock_lwldrv_gwhv Iml_rock_lwldrv_gwhv ( .gwp_sup_hv(gwp_sup_hv),
     .vddp_tieh(vddp_tieh), .gwp_hv(gwp_hv), .gwl_25(gwl_wp_25),
     .gwl_25_b(gwl_wp_b_25));
nand3_25 I44 ( .B(radd_4_25), .A(radd_5_25), .Y(net76), .C(radd_3_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I47 ( .B(radd_1_25), .A(radd_2_25), .Y(net84), .C(radd_0_25),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I104 ( .B(gwlgrpsel_25), .A(gwlgrpsel_25), .Y(net68),
     .C(radd_6_25), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
inv_25 I38 ( .IN(gwl_wp_25), .OUT(gwl_wp_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I100 ( .IN(out_33), .OUT(gwl_b_25), .P(gwl_b_sup_25),
     .Pb(gwl_b_sup_25), .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(gwlb_25), .OUT(gwlb_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_gwl_drv_x57, View - schematic
// LAST TIME SAVED: Apr 30 16:01:52 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwl_drv_x57 ( gwl_b_25, gwl_wr_25, gwp_hv, gwl_b_sup_25,
     gwp_sup_hv, gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25,
     gnv2_b_25, gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25,
     gnv5_b_25, gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1,
     gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gnv0_25, gnv0_b_25, gnv1_25, gnv1_b_25, gnv2_25, gnv2_b_25,
     gnv3_25, gnv3_b_25, gnv4_25, gnv4_b_25, gnv5_25, gnv5_b_25,
     gred_25_0, gred_25_1, gred_b_25_0, gred_b_25_1, gwl_misc_25,
     gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25, vddp_tieh,
     wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25;

output [56:0]  gwl_wr_25;
output [56:0]  gwl_b_25;
output [56:0]  gwp_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_gwl_drv Igwl_drv_51_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[55]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[55]), .gwl_wr_25(gwl_wr_25[55]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_50_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[54]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[54]), .gwl_wr_25(gwl_wr_25[54]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_49_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[53]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[53]), .gwl_wr_25(gwl_wr_25[53]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_48_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[52]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[52]), .gwl_wr_25(gwl_wr_25[52]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_47_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[51]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[51]), .gwl_wr_25(gwl_wr_25[51]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_46_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[50]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[50]), .gwl_wr_25(gwl_wr_25[50]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_45_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[49]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[49]), .gwl_wr_25(gwl_wr_25[49]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_44_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[48]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[48]), .gwl_wr_25(gwl_wr_25[48]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_43_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[47]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[47]), .gwl_wr_25(gwl_wr_25[47]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_42_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[46]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[46]), .gwl_wr_25(gwl_wr_25[46]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_41_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[45]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[45]), .gwl_wr_25(gwl_wr_25[45]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_40_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[44]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[44]), .gwl_wr_25(gwl_wr_25[44]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_39_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[43]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[43]), .gwl_wr_25(gwl_wr_25[43]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_38_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[42]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[42]), .gwl_wr_25(gwl_wr_25[42]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_37_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[41]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[41]), .gwl_wr_25(gwl_wr_25[41]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_36_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[40]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[40]), .gwl_wr_25(gwl_wr_25[40]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_25), .radd_1_25(gnv1_b_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_35_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[39]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[39]), .gwl_wr_25(gwl_wr_25[39]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_34_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[38]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[38]), .gwl_wr_25(gwl_wr_25[38]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25), .radd_1_25(gnv1_25),
     .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_33_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[37]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[37]), .gwl_wr_25(gwl_wr_25[37]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_25));
ml_gwl_drv Igwl_drv_32_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[36]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[36]), .gwl_wr_25(gwl_wr_25[36]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .radd_6_25(vddp_tieh), .radd_5_25(gnv5_25), .radd_4_25(gnv4_b_25),
     .radd_3_25(gnv3_b_25), .radd_2_25(gnv2_b_25),
     .radd_1_25(gnv1_b_25), .radd_0_25(gnv0_b_25));
ml_gwl_drv Igwl_drv_red_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[3]),
     .radd_0_25(gred_25_0), .radd_1_25(gred_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[3]), .gwl_wr_25(gwl_wr_25[3]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_red_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[2]),
     .radd_0_25(gred_b_25_0), .radd_1_25(gred_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[2]), .gwl_wr_25(gwl_wr_25[2]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_red_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[1]),
     .radd_0_25(gred_25_0), .radd_1_25(gred_b_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[1]), .gwl_wr_25(gwl_wr_25[1]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_red_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[0]),
     .radd_0_25(gred_b_25_0), .radd_1_25(gred_b_25_1),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_red_25),
     .gwp_hv(gwp_hv[0]), .gwl_wr_25(gwl_wr_25[0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_misc_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[56]),
     .radd_0_25(vddp_tieh), .radd_1_25(vddp_tieh),
     .radd_2_25(vddp_tieh), .radd_3_25(vddp_tieh),
     .radd_4_25(vddp_tieh), .radd_5_25(vddp_tieh),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_misc_25),
     .gwp_hv(gwp_hv[56]), .gwl_wr_25(gwl_wr_25[56]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_31_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[35]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[35]), .gwl_wr_25(gwl_wr_25[35]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_30_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[34]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[34]), .gwl_wr_25(gwl_wr_25[34]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_29_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[33]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[33]), .gwl_wr_25(gwl_wr_25[33]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_28_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[32]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[32]), .gwl_wr_25(gwl_wr_25[32]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_27_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[31]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[31]), .gwl_wr_25(gwl_wr_25[31]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_26_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[30]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[30]), .gwl_wr_25(gwl_wr_25[30]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_25_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[29]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[29]), .gwl_wr_25(gwl_wr_25[29]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_24_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[28]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_25), .radd_4_25(gnv4_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[28]),
     .gwl_wr_25(gwl_wr_25[28]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_23_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[27]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[27]), .gwl_wr_25(gwl_wr_25[27]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_22_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[26]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[26]), .gwl_wr_25(gwl_wr_25[26]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_21_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[25]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[25]), .gwl_wr_25(gwl_wr_25[25]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_20_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[24]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[24]), .gwl_wr_25(gwl_wr_25[24]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_19_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[23]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[23]), .gwl_wr_25(gwl_wr_25[23]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_18_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[22]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[22]), .gwl_wr_25(gwl_wr_25[22]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_17_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[21]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[21]), .gwl_wr_25(gwl_wr_25[21]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_16_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[20]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[20]),
     .gwl_wr_25(gwl_wr_25[20]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_15_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[19]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[19]), .gwl_wr_25(gwl_wr_25[19]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_14_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[18]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[18]), .gwl_wr_25(gwl_wr_25[18]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_13_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[17]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[17]), .gwl_wr_25(gwl_wr_25[17]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_12_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[16]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[16]), .gwl_wr_25(gwl_wr_25[16]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_11_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[15]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[15]), .gwl_wr_25(gwl_wr_25[15]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_10_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[14]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[14]), .gwl_wr_25(gwl_wr_25[14]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_9_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[13]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[13]), .gwl_wr_25(gwl_wr_25[13]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_8_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[12]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[12]),
     .gwl_wr_25(gwl_wr_25[12]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_7_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[11]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[11]),
     .gwl_wr_25(gwl_wr_25[11]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_6_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[10]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[10]),
     .gwl_wr_25(gwl_wr_25[10]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_5_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[9]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[9]),
     .gwl_wr_25(gwl_wr_25[9]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_4_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[8]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[8]),
     .gwl_wr_25(gwl_wr_25[8]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_3_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[7]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[7]),
     .gwl_wr_25(gwl_wr_25[7]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_2_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[6]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[6]),
     .gwl_wr_25(gwl_wr_25[6]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_1_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[5]),
     .radd_0_25(gnv0_25), .radd_1_25(gnv1_b_25), .radd_2_25(gnv2_b_25),
     .radd_3_25(gnv3_b_25), .radd_4_25(gnv4_b_25),
     .radd_5_25(gnv5_b_25), .radd_6_25(vddp_tieh),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .gwlgrpsel_25(gwl_nvcm_25), .gwp_hv(gwp_hv[5]),
     .gwl_wr_25(gwl_wr_25[5]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .vddp_tieh(vddp_tieh));
ml_gwl_drv Igwl_drv_0_ ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[4]),
     .radd_0_25(gnv0_b_25), .radd_1_25(gnv1_b_25),
     .radd_2_25(gnv2_b_25), .radd_3_25(gnv3_b_25),
     .radd_4_25(gnv4_b_25), .radd_5_25(gnv5_b_25),
     .radd_6_25(vddp_tieh), .wr_frcen_25(wr_frcen_25),
     .wr_dis_25(wr_dis_25), .wp_frcen_25(wp_frcen_25),
     .wp_dis_25(wp_dis_25), .gwlgrpsel_25(gwl_nvcm_25),
     .gwp_hv(gwp_hv[4]), .gwl_wr_25(gwl_wr_25[4]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25),
     .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM, Cell - ml_gwlwr, View - schematic
// LAST TIME SAVED: Apr 30 16:02:13 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr ( gwl_b_25, gwp_hv, wr, gwl_b_sup_25, gwp_sup_hv,
     gnv_25, gnv_b_25, gred_25, gred_b_25, gwl_misc_25, gwl_nvcm_25,
     gwl_red_25, gwlb_dis_25, gwlb_en_25, s_25, vddp_tieh, wp_dis_25,
     wp_frcen_25, wr_dis_25, wr_frcen_25, wr_sup_25 );

inout  gwl_b_sup_25, gwp_sup_hv;

input  gwl_misc_25, gwl_nvcm_25, gwl_red_25, gwlb_dis_25, gwlb_en_25,
     vddp_tieh, wp_dis_25, wp_frcen_25, wr_dis_25, wr_frcen_25,
     wr_sup_25;

output [227:0]  wr;
output [56:0]  gwp_hv;
output [56:0]  gwl_b_25;

input [3:0]  s_25;
input [1:0]  gred_25;
input [5:0]  gnv_b_25;
input [5:0]  gnv_25;
input [1:0]  gred_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [56:0]  gwl_wr_25;



ml_rock_lwldrv_wr_x228 Ilwldrv_wr_x228 ( .wr_sup_25(wr_sup_25),
     .s_25(s_25[3:0]), .gwl_wr_25(gwl_wr_25[56:0]), .wr(wr[227:0]));
ml_gwl_drv_x57 Igwl_drv_x57 ( .gwlb_en_25(gwlb_en_25),
     .gwlb_dis_25(gwlb_dis_25), .gwl_b_25(gwl_b_25[56:0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25_1(gred_b_25[1]), .gred_b_25_0(gred_b_25[0]),
     .gred_25_1(gred_25[1]), .gred_25_0(gred_25[0]),
     .gnv5_b_25(gnv_b_25[5]), .gnv5_25(gnv_25[5]),
     .gnv4_b_25(gnv_b_25[4]), .gnv4_25(gnv_25[4]),
     .gnv3_b_25(gnv_b_25[3]), .gnv3_25(gnv_25[3]),
     .gnv2_b_25(gnv_b_25[2]), .gnv2_25(gnv_25[2]),
     .gnv1_b_25(gnv_b_25[1]), .gnv1_25(gnv_25[1]),
     .gnv0_b_25(gnv_b_25[0]), .gnv0_25(gnv_25[0]),
     .gwp_hv(gwp_hv[56:0]), .gwl_wr_25(gwl_wr_25[56:0]),
     .gwp_sup_hv(gwp_sup_hv), .gwl_b_sup_25(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_gwlwr_top, View - schematic
// LAST TIME SAVED: May  1 11:11:13 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_gwlwr_top ( fsm_gwlbdis_b_25, gwl_b_25, gwl_b_sup_25, gwp_hv,
     pgminhi_dmmy_b_25, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wr, bgr, bl_pgm_glb, vpp_int, vpxa, fsm_coladd,
     fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma, tm_testdec,
     tm_testdec_wr );
output  fsm_gwlbdis_b_25, gwl_b_sup_25, pgminhi_dmmy_b_25, saen_25,
     saen_b_vpxa, testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25;

inout  bgr, bl_pgm_glb, vpp_int, vpxa;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_trow, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_dma,
     tm_testdec, tm_testdec_wr;

output [227:0]  wr;
output [4:1]  sa_ngate_25;
output [56:0]  gwp_hv;
output [4:1]  sa_pgate_vpxa;
output [56:0]  gwl_b_25;

input [3:0]  fsm_trim_ipp;
input [0:0]  fsm_coladd;
input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [2:0]  fsm_trim_rrefpgm;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  s_25;

wire  [1:0]  gred_25;

wire  [1:0]  gred_b_25;

wire  [5:0]  gnv_b_25;

wire  [5:0]  gnv_25;



ml_gwlwr_ctrl Igwlwr_ctrl ( .fsm_pgmdisc(fsm_pgmdisc),
     .gwlb_en_25(gwlb_en_25), .fsm_din(fsm_din),
     .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .tm_testdec_wr(tm_testdec_wr), .tm_testdec(tm_testdec),
     .tm_dma(tm_dma), .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_allwl_l(fsm_tm_allwl_l), .fsm_tm_allwl_h(fsm_tm_allwl_h),
     .fsm_tm_allbl_l(fsm_tm_allbl_l), .fsm_tm_allbl_h(fsm_tm_allbl_h),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_lshven(fsm_lshven),
     .fsm_gwlbdis(fsm_gwlbdis), .fsm_coladd(fsm_coladd[0]),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .s_25(s_25[3:0]),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_red_25(gwl_red_25), .gwl_nvcm_25(gwl_nvcm_25),
     .gwl_misc_25(gwl_misc_25), .gred_b_25(gred_b_25[1:0]),
     .gred_25(gred_25[1:0]), .gnv_b_25(gnv_b_25[5:0]),
     .gnv_25(gnv_25[5:0]), .wr_sup_25(wr_sup_25), .vpxa(vpxa),
     .vpp_int(vpp_int), .vddp_tieh(vddp_tieh), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25), .bl_pgm_glb(bl_pgm_glb), .bgr(bgr));
ml_gwlwr Igwlwr ( .gwlb_en_25(gwlb_en_25), .gwlb_dis_25(gwlb_dis_25),
     .gwl_b_25(gwl_b_25[56:0]), .wr_sup_25(wr_sup_25),
     .wr_frcen_25(wr_frcen_25), .wr_dis_25(wr_dis_25),
     .wp_frcen_25(wp_frcen_25), .wp_dis_25(wp_dis_25),
     .vddp_tieh(vddp_tieh), .s_25(s_25[3:0]), .gwl_red_25(gwl_red_25),
     .gwl_nvcm_25(gwl_nvcm_25), .gwl_misc_25(gwl_misc_25),
     .gred_b_25(gred_b_25[1:0]), .gred_25(gred_25[1:0]),
     .gnv_b_25(gnv_b_25[5:0]), .gnv_25(gnv_25[5:0]), .wr(wr[227:0]),
     .gwp_hv(gwp_hv[56:0]), .gwp_sup_hv(gwp_sup_hv),
     .gwl_b_sup_25(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_core_bank_1_8f, View - schematic
// LAST TIME SAVED: Jul 14 11:49:47 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_core_bank_1_8f ( nv_dataout, bgr, ngate_25, sb25sup_25,
     sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpp_int, vpxa, ysup_25,
     fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din, fsm_gwlbdis,
     fsm_lshven, fsm_multibl_read, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b,
     fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo,
     vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [8:4]  nv_dataout;

input [2:0]  fsm_trim_rrefpgm;
input [7:0]  fsm_rowadd;
input [3:0]  fsm_trim_ipp;
input [3:0]  fsm_blkadd_b;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefrd;
input [9:0]  fsm_coladd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:1]  sa_ngate_25;

wire  [56:0]  gwl_b_25;

wire  [227:0]  wr;

wire  [4:1]  sa_pgate_vpxa;

wire  [56:0]  gwp_hv;



ml_core_654x232_top Iblk_4 ( .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .wr(wr[227:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd[2], fsm_blkadd_b[1],
     fsm_blkadd_b[0]}), .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[4]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_654x232_top Iblk_7 ( .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .wr(wr[227:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd[2], fsm_blkadd[1],
     fsm_blkadd[0]}), .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[7]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_654x232_top blk_6 ( .tm_allbank_sel(tm_allbank_sel),
     .nv_dataout(nv_dataout[6]), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nvcmen(fsm_nvcmen), .fsm_pgm(fsm_pgm),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_rd(fsm_rd), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rowadd(fsm_rowadd[1:0]), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rst_b(fsm_rst_b), .fsm_sample(fsm_sample),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .ngate_25(ngate_25),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .gwl_b_25(gwl_b_25[56:0]), .gwp_hv(gwp_hv[56:0]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]), .saen_25(saen_25),
     .vblinhi_rdo(vblinhi_rdo), .saen_b_vpxa(saen_b_vpxa),
     .testdec_en_b_25(testdec_en_b_25),
     .testdec_even_b_25(testdec_even_b_25), .vpxa(vpxa),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_prec_b_25(testdec_prec_b_25), .tm_allbl_h(tm_allbl_h),
     .tm_allbl_l(tm_allbl_l), .ysup_25(ysup_25),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd[2],
     fsm_blkadd[1], fsm_blkadd_b[0]}), .tm_testdec_wr(tm_testdec_wr),
     .wr(wr[227:0]), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_654x232_top Iblk_5 ( .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .wr(wr[227:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd[2], fsm_blkadd_b[1],
     fsm_blkadd[0]}), .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[5]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_654x232_top Iblk_8 ( .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .wr(wr[227:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd({fsm_blkadd[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd_b[0]}), .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[8]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_gwlwr_top Igwlwr_top_0 ( .tm_testdec_wr(tm_testdec_wr),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_tm_allbl_h(tm_allbl_h),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_wren(fsm_wren), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_coladd(fsm_coladd[0]), .wr(wr[227:0]),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .vpxa(vpxa), .vpp_int(vpp_int), .bl_pgm_glb(bl_pgm_glb),
     .bgr(bgr), .gwl_b_25(gwl_b_25[56:0]), .gwl_b_sup_25(gwl_b_sup_25),
     .tm_testdec(fsm_tm_testdec), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_wpen(fsm_wpen), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_tm_allwl_l(tm_allwl_l), .fsm_tm_allbl_l(tm_allbl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .fsm_din(fsm_din), .tm_dma(tm_dma));

endmodule
// Library - NVCM, Cell - ml_core_bank_0_8f, View - schematic
// LAST TIME SAVED: Jul 14 11:49:52 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_core_bank_0_8f ( nv_dataout, bgr, ngate_25, sb25sup_25,
     sbhvsup_hv, vblinhi_rde, vblinhi_rdo, vpp_int, vpxa, ysup_25,
     fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din, fsm_gwlbdis,
     fsm_lshven, fsm_multibl_read, fsm_nv_bstream, fsm_nv_rri_trim,
     fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd, fsm_rst_b,
     fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis, tm_allbank_sel,
     tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol,
     tm_testdec_wr );

inout  bgr, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi_rde, vblinhi_rdo,
     vpp_int, vpxa, ysup_25;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  nv_dataout;

input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_trim_rrefrd;
input [7:0]  fsm_rowadd;
input [9:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [3:0]  fsm_blkadd_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [4:1]  sa_pgate_vpxa;

wire  [227:0]  wr;

wire  [56:0]  gwl_b_25;

wire  [4:1]  sa_ngate_25;

wire  [56:0]  gwp_hv;



ml_core_654x232_top Iblk_2 ( .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .wr(wr[227:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd[1],
     fsm_blkadd_b[0]}), .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[2]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_654x232_top blk_1 ( .tm_allbank_sel(tm_allbank_sel),
     .nv_dataout(nv_dataout[1]), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_nvcmen(fsm_nvcmen), .fsm_pgm(fsm_pgm),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_rd(fsm_rd), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rowadd(fsm_rowadd[1:0]), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rst_b(fsm_rst_b), .fsm_sample(fsm_sample),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .ngate_25(ngate_25),
     .fsm_tm_testdec(fsm_tm_testdec),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]), .sb25sup_25(sb25sup_25),
     .fsm_vpxaset(fsm_vpxaset), .fsm_wpen(fsm_wpen),
     .fsm_ymuxdis(fsm_ymuxdis), .sbhvsup_hv(sbhvsup_hv),
     .gwl_b_25(gwl_b_25[56:0]), .gwp_hv(gwp_hv[56:0]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .vblinhi_rde(vblinhi_rde),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]), .saen_25(saen_25),
     .vblinhi_rdo(vblinhi_rdo), .saen_b_vpxa(saen_b_vpxa),
     .testdec_en_b_25(testdec_en_b_25),
     .testdec_even_b_25(testdec_even_b_25), .vpxa(vpxa),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_prec_b_25(testdec_prec_b_25), .tm_allbl_h(tm_allbl_h),
     .tm_allbl_l(tm_allbl_l), .ysup_25(ysup_25),
     .tm_allwl_h(tm_allwl_h), .tm_allwl_l(tm_allwl_l),
     .tm_tcol(tm_tcol), .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2],
     fsm_blkadd_b[1], fsm_blkadd[0]}), .tm_testdec_wr(tm_testdec_wr),
     .wr(wr[227:0]), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_multibl_read(fsm_multibl_read), .tm_dma(tm_dma));
ml_core_654x232_top Iblk_0 ( .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .wr(wr[227:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd_b[1],
     fsm_blkadd_b[0]}), .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[0]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_core_654x232_top Iblk_3 ( .tm_allbank_sel(tm_allbank_sel),
     .tm_dma(tm_dma), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .wr(wr[227:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd({fsm_blkadd_b[3], fsm_blkadd_b[2], fsm_blkadd[1],
     fsm_blkadd[0]}), .tm_tcol(tm_tcol), .tm_allwl_l(tm_allwl_l),
     .tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25), .vpxa(vpxa),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .vblinhi_rdo(vblinhi_rdo), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .vblinhi_rde(vblinhi_rde),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .gwl_b_25(gwl_b_25[56:0]), .sbhvsup_hv(sbhvsup_hv),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .sb25sup_25(sb25sup_25),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .ngate_25(ngate_25),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .gwl_b_sup_25(gwl_b_sup_25),
     .fsm_rowadd(fsm_rowadd[1:0]), .bl_pgm_glb(bl_pgm_glb),
     .fsm_rd(fsm_rd), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_tm_trow(fsm_tm_trow), .fsm_pgm(fsm_pgm),
     .fsm_nvcmen(fsm_nvcmen), .nv_dataout(nv_dataout[3]),
     .fsm_coladd(fsm_coladd[9:0]));
ml_gwlwr_top Igwlwr_top_0 ( .tm_testdec_wr(tm_testdec_wr),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wgnden(fsm_wgnden),
     .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_tm_allbl_h(tm_allbl_h),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .fsm_wren(fsm_wren), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_coladd(fsm_coladd[0]), .wr(wr[227:0]),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .testdec_en_b_25(testdec_en_b_25), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]),
     .pgminhi_dmmy_b_25(pgmminhi_dmmy_b_25), .gwp_hv(gwp_hv[56:0]),
     .vpxa(vpxa), .vpp_int(vpp_int), .bl_pgm_glb(bl_pgm_glb),
     .bgr(bgr), .gwl_b_25(gwl_b_25[56:0]), .gwl_b_sup_25(gwl_b_sup_25),
     .tm_testdec(fsm_tm_testdec), .fsm_gwlbdis_b_25(fsm_gwlbdis_b_25),
     .fsm_wpen(fsm_wpen), .fsm_pgmdisc(fsm_pgmdisc),
     .fsm_tm_allwl_l(tm_allwl_l), .fsm_tm_allbl_l(tm_allbl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .fsm_din(fsm_din), .tm_dma(tm_dma));

endmodule
// Library - NVCM, Cell - ml_hv2vddp_sw, View - schematic
// LAST TIME SAVED: May  1 11:01:33 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_hv2vddp_sw ( out_hv, hv2vddp, vddp_tieh );
inout  out_hv;

input  hv2vddp, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_ls_inv_hotsw Iml_hv_ls_inv_vppt ( .sel_b_25(sw_vddp_b),
     .sel_25(net035), .out_b_hv(sw_vpp_b), .in_hv(out_hv),
     .vddp_tieh(vddp_tieh));
pch_25  M1 ( .D(net27), .B(out_hv), .G(sw_vpp_b), .S(out_hv));
pch_25  M0 ( .D(net27), .B(vddp_), .G(sw_vddp_b), .S(vddp_));
inv_25 I62 ( .IN(net37), .OUT(sw_vddp_b), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I71 ( .IN(net060), .OUT(net035), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net060),
     .out_vddio(net37), .in_b(net46));
inv_hvt I65 ( .A(hv2vddp), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));

endmodule
// Library - NVCM, Cell - ml_vpp_ref_sw, View - schematic
// LAST TIME SAVED: Mar 21 16:41:35 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vpp_ref_sw ( in, out, sel_b_25 );
inout  in, out;

input  sel_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I281 ( .IN(sel_b_25), .OUT(net122), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M12 ( .D(out), .B(GND_), .G(net122), .S(in));
pch_25  M14 ( .D(in), .B(vddp_), .G(sel_b_25), .S(out));

endmodule
// Library - NVCM, Cell - ml_vpp_ref, View - schematic
// LAST TIME SAVED: Apr  7 18:49:59 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vpp_ref ( vref_25, bgr, pumpen_25, vppwl_25 );
inout  vref_25;

input  bgr, pumpen_25;

input [2:0]  vppwl_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_b_25;

wire  [7:0]  red_dec_25;



nch_na25  M0 ( .D(net179), .B(GND_), .G(ctrl_gate_25),
     .S(bgr_mirror_25));
nand3_25 I44_7_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[7]),
     .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_6_ ( .B(vppwl_25[1]), .A(vppwl_25[2]), .Y(red_dec_25[6]),
     .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I44_5_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[5]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_4_ ( .B(vppwl_b_25[1]), .A(vppwl_25[2]),
     .Y(red_dec_25[4]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_3_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[3]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_2_ ( .B(vppwl_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[2]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_1_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[1]), .C(vppwl_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
nand3_25 I44_0_ ( .B(vppwl_b_25[1]), .A(vppwl_b_25[2]),
     .Y(red_dec_25[0]), .C(vppwl_b_25[0]), .P(vddp_), .Pb(vddp_),
     .Gb(gnd_), .G(gnd_));
ml_vpp_ref_sw I281 ( .in(net92), .out(vref_25),
     .sel_b_25(red_dec_25[6]));
ml_vpp_ref_sw I287 ( .in(net95), .out(vref_25),
     .sel_b_25(red_dec_25[4]));
ml_vpp_ref_sw I283 ( .in(net98), .out(vref_25),
     .sel_b_25(red_dec_25[7]));
ml_vpp_ref_sw I290 ( .in(net0100), .out(vref_25),
     .sel_b_25(red_dec_25[0]));
ml_vpp_ref_sw I288 ( .in(net104), .out(vref_25),
     .sel_b_25(red_dec_25[3]));
ml_vpp_ref_sw I284 ( .in(net139), .out(vref_25),
     .sel_b_25(red_dec_25[5]));
ml_vpp_ref_sw I291 ( .in(net110), .out(vref_25),
     .sel_b_25(red_dec_25[1]));
ml_vpp_ref_sw I292 ( .in(net113), .out(vref_25),
     .sel_b_25(red_dec_25[2]));
nmoscap_25  C3 ( .MINUS(net0129), .PLUS(net0113));
nmoscap_25  C2 ( .MINUS(gnd_), .PLUS(ctrl_gate_25));
inv_25 I38 ( .IN(pumpen_25), .OUT(vppref_en_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_2_ ( .IN(vppwl_25[2]), .OUT(vppwl_b_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_1_ ( .IN(vppwl_25[1]), .OUT(vppwl_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I305_0_ ( .IN(vppwl_25[0]), .OUT(vppwl_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
rppolywo_m  R11 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R13 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R14 ( .MINUS(net113), .PLUS(net104), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(net110), .PLUS(net113), .BULK(GND_));
rppolywo_m  R15 ( .MINUS(net104), .PLUS(net95), .BULK(GND_));
rppolywo_m  R16 ( .MINUS(net104), .PLUS(net95), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net95), .PLUS(net139), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net95), .PLUS(net139), .BULK(GND_));
rppolywo_m  R19 ( .MINUS(net139), .PLUS(net92), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(net139), .PLUS(net92), .BULK(GND_));
rppolywo_m  R21 ( .MINUS(net92), .PLUS(net98), .BULK(GND_));
rppolywo_m  R22 ( .MINUS(net92), .PLUS(net98), .BULK(GND_));
rppolywo_m  R25 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R24 ( .MINUS(net98), .PLUS(bgr_mirror_25), .BULK(GND_));
rppolywo_m  R8 ( .MINUS(gnd_), .PLUS(net0100), .BULK(GND_));
rppolywo_m  R5 ( .MINUS(net0100), .PLUS(net110), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net0100), .PLUS(net110), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(bgr_mirror_25), .PLUS(net0129), .BULK(GND_));
nch_25  M10 ( .D(net163), .B(GND_), .G(bgr), .S(gnd_));
nch_25  M14 ( .D(net0113), .B(GND_), .G(vppref_en_b_25), .S(gnd_));
nch_25  M15 ( .D(ctrl_gate_25), .B(GND_), .G(vppref_en_b_25),
     .S(gnd_));
nch_25  M8 ( .D(ctrl_gate_25), .B(GND_), .G(bgr_mirror_25),
     .S(net163));
nch_25  M13 ( .D(net0113), .B(GND_), .G(bgr), .S(net163));
pch_25  M18 ( .D(net179), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));
pch_25  M5 ( .D(ctrl_gate_25), .B(vddp_), .G(net0113), .S(net175));
pch_25  M6 ( .D(net0113), .B(vddp_), .G(net0113), .S(net175));
pch_25  M7 ( .D(net175), .B(vddp_), .G(vppref_en_b_25), .S(vddp_));

endmodule
// Library - NVCM, Cell - ml_vpp_ctrl, View - schematic
// LAST TIME SAVED: Apr 30 14:24:32 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vpp_ctrl ( pumpen_25, vpint_en, vpp_2_vdd, vppdisc_25,
     vppwl_25, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_vpgmwl_buf, fsm_wgnden );
output  pumpen_25, vpint_en, vpp_2_vdd, vppdisc_25;

input  fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf,
     fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint, fsm_wgnden;

output [2:0]  vppwl_25;

input [2:0]  fsm_vpgmwl_buf;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:2]  net068;

wire  [0:2]  net038;

wire  [0:2]  net082;

wire  [0:2]  net092;



nand4_hvt I75 ( .D(fsm_pgm_buf), .C(fsm_lshven_buf), .A(net0127),
     .Y(net046), .B(net0127));
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(net0122));
nor2_hvt I111 ( .A(vpp_pumpen_b), .B(net080), .Y(net0133));
nor2_hvt I87 ( .A(vpp_pumpen), .Y(net036), .B(fsm_pgmdisc_buf));
sbtlibn65lp_ml_dff_schematic I77 ( .CLK(net084), .QN(vpp_pumpen_b),
     .R(pgm_dis), .D(vdd_tieh), .Q(vpp_pumpen));
vdd_tiehigh I117 ( .vdd_tieh(vdd_tieh));
nand3_hvt I79 ( .C(net086), .A(fsm_pgm_buf), .Y(pgm_dis),
     .B(fsm_nvcmen_buf));
nand2_hvt I104 ( .A(fsm_tm_xforce), .Y(net049), .B(fsm_tm_xvppint));
inv_25 I95_2_ ( .IN(net068[0]), .OUT(vppwl_25[2]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_1_ ( .IN(net068[1]), .OUT(vppwl_25[1]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I95_0_ ( .IN(net068[2]), .OUT(vppwl_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I81 ( .IN(net073), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(net088), .OUT(vppdisc_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I96_2_ ( .in(net082[0]), .sup(vddp_),
     .out_vddio_b(net068[0]), .out_vddio(net038[0]), .in_b(net092[0]));
ml_ls_vdd2vdd25 I96_1_ ( .in(net082[1]), .sup(vddp_),
     .out_vddio_b(net068[1]), .out_vddio(net038[1]), .in_b(net092[1]));
ml_ls_vdd2vdd25 I96_0_ ( .in(net082[2]), .sup(vddp_),
     .out_vddio_b(net068[2]), .out_vddio(net038[2]), .in_b(net092[2]));
ml_ls_vdd2vdd25 I84 ( .in(net0133), .sup(vddp_), .out_vddio_b(net073),
     .out_vddio(net074), .in_b(net0134));
ml_ls_vdd2vdd25 I173 ( .in(fsm_pgmdisc_buf), .sup(vddp_),
     .out_vddio_b(net088), .out_vddio(net048), .in_b(net0106));
inv_hvt I107 ( .A(net0122), .Y(net0124));
inv_hvt I109 ( .A(fsm_pgmvfy_buf), .Y(net0127));
inv_hvt I131 ( .A(net049), .Y(net080));
inv_hvt I110_2_ ( .A(net092[0]), .Y(net082[0]));
inv_hvt I110_1_ ( .A(net092[1]), .Y(net082[1]));
inv_hvt I110_0_ ( .A(net092[2]), .Y(net082[2]));
inv_hvt I76 ( .A(net046), .Y(net084));
inv_hvt I108 ( .A(fsm_pgmdisc_buf), .Y(net0122));
inv_hvt I78 ( .A(net0124), .Y(net086));
inv_hvt I113 ( .A(vpp_pumpen_b), .Y(vpint_en));
inv_hvt I91 ( .A(net036), .Y(net089));
inv_hvt I90 ( .A(net089), .Y(vpp_2_vdd));
inv_hvt I98_2_ ( .A(fsm_vpgmwl_buf[2]), .Y(net092[0]));
inv_hvt I98_1_ ( .A(fsm_vpgmwl_buf[1]), .Y(net092[1]));
inv_hvt I98_0_ ( .A(fsm_vpgmwl_buf[0]), .Y(net092[2]));
inv_hvt I112 ( .A(net0133), .Y(net0134));
inv_hvt I101 ( .A(fsm_pgmdisc_buf), .Y(net0106));

endmodule
// Library - xpmem, Cell - sg_bufx10, View - schematic
// LAST TIME SAVED: Jul 28 19:09:08 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module sg_bufx10 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - NVCM, Cell - ml_vpp_reg, View - schematic
// LAST TIME SAVED: May  3 15:48:51 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vpp_reg ( slow_25, bgr, pbias_25, pump_in, vpp_int,
     pumpen_25, vppdisc_25, vref_25 );
output  slow_25;

inout  bgr, pbias_25, pump_in, vpp_int;

input  pumpen_25, vppdisc_25, vref_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I261 ( .vddp_tieh(net0208));
nch_na25  M11 ( .D(net0199), .B(GND_), .G(vppdisc_25), .S(VDD_));
nch_na25  M22 ( .D(vpp_int), .B(GND_), .G(pump_gate), .S(pump_in));
nch_na25  M1 ( .D(GND_), .B(GND_), .G(pump_gate), .S(GND_));
nch_na25  M10 ( .D(net0203), .B(GND_), .G(net0208), .S(net0199));
nch_na25  M5 ( .D(pump_opamp_out), .B(GND_), .G(vpp_int),
     .S(pump_opamp_out));
inv_25 I211 ( .IN(en_buf_b_25), .OUT(en_buf_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I212 ( .IN(pumpen_25), .OUT(en_buf_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
pch_25  M31 ( .D(net0203), .B(net0165), .G(dis_pgate_25), .S(net0165));
pch_25  M0 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
pch_25  M9 ( .D(net0166), .B(vddp_), .G(en_buf_b_25), .S(vddp_));
pch_25  M14 ( .D(pump_opamp_out), .B(net125), .G(vref_25), .S(net125));
pch_25  M18 ( .D(net122), .B(vpp_int), .G(net122), .S(vpp_int));
pch_25  M13 ( .D(net124), .B(net125), .G(vdiv), .S(net125));
pch_25  M32 ( .D(dis_pgate_25), .B(vddp_), .G(dis_pgate_25),
     .S(vddp_));
pch_25  M33 ( .D(dis_pgate_25), .B(vddp_), .G(vppdisc_25), .S(vddp_));
pch_25  M12 ( .D(net125), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M19 ( .D(net134), .B(net122), .G(net134), .S(net122));
pch_25  M21 ( .D(net138), .B(net134), .G(net138), .S(net134));
pch_25  M23 ( .D(net142), .B(net138), .G(net142), .S(net138));
pch_25  M24 ( .D(vdiv), .B(net142), .G(vdiv), .S(net142));
pch_25  M25 ( .D(net0224), .B(vdiv), .G(net0224), .S(vdiv));
pch_25  M4_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
pch_25  M4_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net0166));
nch_25  M40 ( .D(dis_pgate_25), .B(GND_), .G(vppdisc_25), .S(gnd_));
nch_25  M8 ( .D(pbias_25), .B(GND_), .G(en_buf_b_25), .S(gnd_));
nch_25  M16 ( .D(net124), .B(GND_), .G(net124), .S(net155));
nch_25  M17 ( .D(net155), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M6 ( .D(vpp_int), .B(GND_), .G(en_buf_25), .S(net168));
nch_25  M20 ( .D(slow_25), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M7 ( .D(net168), .B(GND_), .G(pump_opamp_out), .S(gnd_));
nch_25  M41 ( .D(net0224), .B(GND_), .G(en_buf_25), .S(gnd_));
nch_25  M15 ( .D(pump_opamp_out), .B(GND_), .G(net124), .S(net155));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net0250));
rppolywo_m  R5 ( .MINUS(net0165), .PLUS(vpp_int), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(pump_gate), .PLUS(pump_in), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net0247), .PLUS(net0250), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net0247), .BULK(GND_));

endmodule
// Library - NVCM, Cell - ml_vpp_vco, View - schematic
// LAST TIME SAVED: Apr  8 16:31:55 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vpp_vco ( clk_25_0, pbias_25, slow_25, en_25, freq_25 );
output  clk_25_0;

inout  pbias_25, slow_25;

input  en_25;

input [1:0]  freq_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:1]  freq_b_25;



nch_na25  M4 ( .D(GND_), .B(GND_), .G(net173), .S(GND_));
nch_na25  M15 ( .D(GND_), .B(GND_), .G(net185), .S(GND_));
nch_na25  M16 ( .D(GND_), .B(GND_), .G(net193), .S(GND_));
nch_na25  M2 ( .D(GND_), .B(GND_), .G(net189), .S(GND_));
nch_25  M5 ( .D(net173), .B(GND_), .G(net185), .S(net177));
nch_25  M6 ( .D(net177), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M13 ( .D(net181), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M14 ( .D(net185), .B(GND_), .G(net193), .S(net181));
nch_25  M8 ( .D(net189), .B(GND_), .G(net173), .S(net201));
nch_25  M17 ( .D(net193), .B(GND_), .G(net195), .S(net197));
nch_25  M18 ( .D(net197), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M1 ( .D(net201), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M23 ( .D(pbias_osc_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M24 ( .D(slow_25), .B(GND_), .G(nbias_osc_25), .S(GND_));
nch_25  M25 ( .D(nbias_osc_25), .B(GND_), .G(en_25), .S(slow_25));
pch_25  M7 ( .D(net173), .B(vddp_), .G(net185), .S(net236));
pch_25  M10 ( .D(net236), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M9 ( .D(net248), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M3 ( .D(net189), .B(vddp_), .G(net173), .S(net248));
pch_25  M11 ( .D(net256), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M12 ( .D(net185), .B(vddp_), .G(net193), .S(net256));
pch_25  M19 ( .D(net193), .B(vddp_), .G(net195), .S(net260));
pch_25  M20 ( .D(net260), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
pch_25  M22 ( .D(pbias_osc_25), .B(vddp_), .G(en_b_25), .S(net228));
pch_25  M26_1_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M26_0_ ( .D(nbias_osc_25), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_1_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M27_0_ ( .D(net208), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M28 ( .D(net212), .B(vddp_), .G(pbias_25), .S(vddp_));
pch_25  M29 ( .D(nbias_osc_25), .B(vddp_), .G(freq_25[0]), .S(net212));
pch_25  M30 ( .D(nbias_osc_25), .B(vddp_), .G(freq_b_25[1]),
     .S(net208));
pch_25  M21 ( .D(net228), .B(vddp_), .G(pbias_osc_25), .S(vddp_));
nand2_25 I96 ( .G(GND_), .Pb(vddp_), .A(net189), .Y(net195), .P(vddp_),
     .B(en_25), .Gb(GND_));
inv_25 I201 ( .IN(net195), .OUT(clk_25_0), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I188 ( .IN(en_25), .OUT(en_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I199 ( .IN(freq_25[1]), .OUT(freq_b_25[1]), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));

endmodule
// Library - NVCM, Cell - ml_vpp_pump, View - schematic
// LAST TIME SAVED: Apr  7 18:25:20 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vpp_pump ( pump_in, clkin_25, en_25 );
inout  pump_in;

input  clkin_25, en_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));
nmoscap_25  C1 ( .MINUS(clk_b_25), .PLUS(s_3));
pch_25  M0 ( .D(net23), .B(vddp_), .G(net64), .S(vddp_));
inv_25 I194 ( .IN(clkin_25), .OUT(net70), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(en_25), .OUT(net64), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I210 ( .IN(net28), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I219 ( .IN(net40), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I220 ( .IN(net34), .OUT(net46), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I221 ( .IN(net46), .OUT(net40), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I224 ( .IN(clkin_25), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I209 ( .IN(net70), .OUT(net28), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
nch_na25  M10 ( .D(s_0), .B(GND_), .G(s_0), .S(s_1));
nch_na25  M11 ( .D(s_1), .B(GND_), .G(s_1), .S(s_2));
nch_na25  M12 ( .D(s_2), .B(GND_), .G(s_2), .S(s_3));
nch_na25  M22 ( .D(net23), .B(GND_), .G(net23), .S(s_0));
nch_na25  M1 ( .D(s_3), .B(GND_), .G(s_3), .S(pump_in));

endmodule
// Library - NVCM, Cell - ml_vpp_pumpx3, View - schematic
// LAST TIME SAVED: Apr  8 17:28:05 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vpp_pumpx3 ( pump_in, clkin_0_25, pumpen_25 );
inout  pump_in;

input  clkin_0_25, pumpen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I195 ( .IN(clkin_0_25), .OUT(net13), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I84 ( .IN(net13), .OUT(net024), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
ml_vpp_pump Ivpp_pump_0 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(clkin_0_25));
ml_vpp_pump I79 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net024));
ml_vpp_pump Ivpp_pump_1 ( .pump_in(pump_in), .en_25(pumpen_25),
     .clkin_25(net13));

endmodule
// Library - NVCM, Cell - ml_vppint_top, View - schematic
// LAST TIME SAVED: May  1 11:06:26 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_vppint_top ( vpint_en, vpp_int, bgr, fsm_lshven_buf,
     fsm_nvcmen_buf, fsm_pgm_buf, fsm_pgmdisc_buf, fsm_pgmvfy_buf,
     fsm_tm_xforce, fsm_tm_xvppint, fsm_vpgmwl_buf, fsm_wgnden_buf );
output  vpint_en;

inout  vpp_int;

input  bgr, fsm_lshven_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmvfy_buf, fsm_tm_xforce, fsm_tm_xvppint,
     fsm_wgnden_buf;

input [2:0]  fsm_vpgmwl_buf;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [2:0]  vppwl_25;

wire  [1:0]  freq_25;



ml_hv2vddp_sw Ivpxa_2vddp_sw ( .hv2vddp(vpp_2_vdd),
     .vddp_tieh(vddp_tieh), .out_hv(vpp_int));
inv_25 I38 ( .IN(vddp_tieh), .OUT(freq_25[1]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I86 ( .IN(vddp_tieh), .OUT(freq_25[0]), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
ml_vpp_ref Ivpp_ref ( .vref_25(vref_25), .vppwl_25(vppwl_25[2:0]),
     .pumpen_25(pumpen_25), .bgr(bgr));
ml_vpp_ctrl Ivpp_ctrl ( .vpint_en(vpint_en),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .vppdisc_25(vppdisc_25), .fsm_wgnden(fsm_wgnden_buf),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf), .vppwl_25(vppwl_25[2:0]),
     .vpp_2_vdd(vpp_2_vdd), .pumpen_25(pumpen_25));
ml_vpp_reg Ivpp_reg ( .bgr(bgr), .slow_25(slow_25),
     .pbias_25(pbias_25), .vref_25(vref_25), .vppdisc_25(vppdisc_25),
     .pumpen_25(pumpen_25), .pump_in(pump_in), .vpp_int(vpp_int));
ml_vpp_vco Ivpp_vco ( .pbias_25(pbias_25), .slow_25(slow_25),
     .freq_25(freq_25[1:0]), .en_25(pumpen_25), .clk_25_0(clkin_0_25));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));
nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpp_int));
ml_vpp_pumpx3 Ivpp_pumpx3 ( .pump_in(pump_in), .pumpen_25(pumpen_25),
     .clkin_0_25(clkin_0_25));

endmodule
// Library - NVCM, Cell - UBGR_2511_065_FLAT, View - schematic
// LAST TIME SAVED: Apr  1 15:53:36 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module UBGR_2511_065_FLAT ( VREF, PDN, T0, T1, T2, T3, TEN, VDD25, VSS
     );
output  VREF;

input  PDN, T0, T1, T2, T3, TEN, VDD25, VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_bgr_top, View - schematic
// LAST TIME SAVED: Apr  7 14:19:14 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_bgr_top ( bgr_int, fsm_nvcmen_buf, fsm_trim_vbg_buf );
inout  bgr_int;

input  fsm_nvcmen_buf;

input [3:0]  fsm_trim_vbg_buf;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  bgr_trim_25;

wire  [0:3]  net48;

wire  [0:3]  net53;

wire  [0:3]  net44;



inv_25 I38 ( .IN(net58), .OUT(PDN), .P(vddp_), .Pb(vddp_), .G(gnd_),
     .Gb(gnd_));
vddp_tiehigh I85 ( .vddp_tieh(TEN));
UBGR_2511_065_FLAT Ibgr ( .TEN(TEN), .VSS(gnd_), .VDD25(vddp_),
     .VREF(bgr_int), .T3(bgr_trim_25[3]), .T2(bgr_trim_25[2]),
     .T1(bgr_trim_25[1]), .T0(bgr_trim_25[0]), .PDN(PDN));
inv_hvt I88_3_ ( .A(fsm_trim_vbg_buf[3]), .Y(net48[0]));
inv_hvt I88_2_ ( .A(fsm_trim_vbg_buf[2]), .Y(net48[1]));
inv_hvt I88_1_ ( .A(fsm_trim_vbg_buf[1]), .Y(net48[2]));
inv_hvt I88_0_ ( .A(fsm_trim_vbg_buf[0]), .Y(net48[3]));
inv_hvt I319 ( .A(net50), .Y(net46));
inv_hvt I87_3_ ( .A(net48[0]), .Y(net44[0]));
inv_hvt I87_2_ ( .A(net48[1]), .Y(net44[1]));
inv_hvt I87_1_ ( .A(net48[2]), .Y(net44[2]));
inv_hvt I87_0_ ( .A(net48[3]), .Y(net44[3]));
inv_hvt I323 ( .A(fsm_nvcmen_buf), .Y(net50));
ml_ls_vdd2vdd25 I80_3_ ( .in(net44[0]), .sup(vddp_),
     .out_vddio_b(net53[0]), .out_vddio(bgr_trim_25[3]),
     .in_b(net48[0]));
ml_ls_vdd2vdd25 I80_2_ ( .in(net44[1]), .sup(vddp_),
     .out_vddio_b(net53[1]), .out_vddio(bgr_trim_25[2]),
     .in_b(net48[1]));
ml_ls_vdd2vdd25 I80_1_ ( .in(net44[2]), .sup(vddp_),
     .out_vddio_b(net53[2]), .out_vddio(bgr_trim_25[1]),
     .in_b(net48[2]));
ml_ls_vdd2vdd25 I80_0_ ( .in(net44[3]), .sup(vddp_),
     .out_vddio_b(net53[3]), .out_vddio(bgr_trim_25[0]),
     .in_b(net48[3]));
ml_ls_vdd2vdd25 I335 ( .in(net46), .sup(vddp_), .out_vddio_b(net58),
     .out_vddio(bgr_en_25), .in_b(net50));

endmodule
// Library - NVCM, Cell - ml_pump_vpxa_3.3v, View - schematic
// LAST TIME SAVED: Nov 14 11:57:16 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_pump_vpxa_3_3v ( out, clkin_25, en );
inout  out;

input  clkin_25, en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M10 ( .B(GND_), .D(s_0), .G(s_0), .S(s_1));
nch_na25  M11 ( .B(GND_), .D(s_1), .G(s_1), .S(s_2));
nch_na25  M12 ( .B(GND_), .D(s_2), .G(s_2), .S(out));
nch_na25  M22 ( .B(GND_), .D(net0115), .G(net0115), .S(s_0));
inv_25 I194 ( .IN(clkin_25), .OUT(net064), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I206 ( .IN(en), .OUT(net042), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
inv_25 I210 ( .IN(net076), .OUT(clk_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I219 ( .IN(net040), .OUT(clk_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I220 ( .IN(net034), .OUT(net046), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I221 ( .IN(net046), .OUT(net040), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I224 ( .IN(clkin_25), .OUT(net034), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I209 ( .IN(net064), .OUT(net076), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
pch_25  M0 ( .D(net0115), .B(vddp_), .G(net042), .S(vddp_));
nmoscap_25  C0 ( .MINUS(clk_25), .PLUS(s_0));
nmoscap_25  C4 ( .MINUS(clk_b_25), .PLUS(s_1));
nmoscap_25  C7 ( .MINUS(clk_25), .PLUS(s_2));

endmodule
// Library - sbtlibn65lp, Cell - ml_dlatch_25, View - schematic
// LAST TIME SAVED: Feb 21 13:49:32 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_dlatch_25 ( Q_25, D_25, EN_25, R_25 );
output  Q_25;

input  D_25, EN_25, R_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M9 ( .D(net31), .B(vddp_), .G(EN_25), .S(vddp_));
pch_25  M7 ( .D(net39), .B(vddp_), .G(EN_B_25), .S(vddp_));
pch_25  M3 ( .D(net52), .B(vddp_), .G(D_25), .S(net39));
pch_25  M4 ( .D(net52), .B(vddp_), .G(Q_25), .S(net31));
nch_25  M8 ( .D(net52), .B(GND_), .G(D_25), .S(net48));
nch_25  M1 ( .D(net48), .B(GND_), .G(EN_25), .S(GND_));
nch_25  M5 ( .D(net40), .B(GND_), .G(EN_B_25), .S(GND_));
nch_25  M6 ( .D(net52), .B(GND_), .G(Q_25), .S(net40));
inv_25 I156 ( .IN(EN_25), .OUT(EN_B_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
nor2_25 I161 ( .A(net52), .Y(Q_25), .Gb(GND_), .G(GND_), .Pb(vddp_),
     .P(vddp_), .B(R_25));

endmodule
// Library - NVCM, Cell - ml_pump_clk_reg, View - schematic
// LAST TIME SAVED: Feb 13 16:09:37 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_pump_clk_reg ( clk_out_25, clk_in_25, pump_chrg_25,
     pump_on_25 );
output  clk_out_25;

input  clk_in_25, pump_chrg_25, pump_on_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



exor2_25 I85 ( .A(clk_in_25), .Y(net020), .B(clk_out_25));
nand2_25 I78 ( .G(GND_), .Pb(vddp_), .A(pump_chrg_25), .Y(clk_freeze),
     .P(vddp_), .B(pump_on_25), .Gb(GND_));
inv_25 I72 ( .IN(net020), .OUT(clk_equal), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(vddp_tieh), .OUT(net34), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
vddp_tiehigh I117 ( .vddp_tieh(vddp_tieh));
ml_dlatch_25 I63 ( .D_25(clk_in_25), .EN_25(clk_go), .R_25(net34),
     .Q_25(clk_out_25));
ml_dlatch_25 I64 ( .D_25(vddp_tieh), .EN_25(clk_equal),
     .R_25(clk_freeze), .Q_25(clk_go));

endmodule
// Library - leafcell, Cell - bram_bufferx4, View - schematic
// LAST TIME SAVED: Jun 25 13:46:30 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module bram_bufferx4 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - NVCM, Cell - ml_pump_vpxa_x2, View - schematic
// LAST TIME SAVED: Nov 14 11:57:43 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_pump_vpxa_x2 ( vpxa_int, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, pumpen, pumpen_25, vpxa_clk_25, vpxa_clk_b_25 );
inout  vpxa_int;

input  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25, pumpen,
     pumpen_25, vpxa_clk_25, vpxa_clk_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_pump_vpxa_3_3v Ivpxa_pump_0 ( .en(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_0_25));
ml_pump_vpxa_3_3v Ivpxa_pump_2 ( .en(pumpen_25), .out(vpxa_int),
     .clkin_25(clkin_2_25));
ml_pump_vpxa_3_3v Ivpxa_pump_1 ( .en(pumpen_25), .clkin_25(clkin_1_25),
     .out(vpxa_int));
ml_pump_clk_reg Iclk_reg_0 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_0_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_0_25));
ml_pump_clk_reg Iclk_reg_2 ( .clk_in_25(vpxa_clk_b_25),
     .pump_chrg_25(pump_chrg_2_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_2_25));
ml_pump_clk_reg Iclk_reg_1 ( .clk_in_25(vpxa_clk_25),
     .pump_chrg_25(pump_chrg_1_25), .pump_on_25(pumpen_25),
     .clk_out_25(clkin_1_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_osc, View - schematic
// LAST TIME SAVED: Mar 14 15:11:03 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_vpxa_osc ( vpxa_clk_25, bgr, freq_25, pumpen_25 );
output  vpxa_clk_25;

inout  bgr;

input  pumpen_25;

input [1:0]  freq_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  freq_buf_b_25;



inv_25 I38 ( .IN(pumpen_25), .OUT(pbiasen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I195 ( .IN(freq_25[0]), .OUT(freq_buf_b_25[0]), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
pch_25  M9 ( .D(net64), .B(vddp_), .G(pbiasen_b_25), .S(vddp_));
pch_25  M4_1_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
pch_25  M4_0_ ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
pch_25  M0 ( .D(pbias_25), .B(vddp_), .G(pbias_25), .S(net64));
nch_25  M8 ( .D(pbias_25), .B(GND_), .G(pbiasen_b_25), .S(gnd_));
nch_25  M3 ( .D(pbias_25), .B(GND_), .G(bgr), .S(net74));
rppolywo_m  R2 ( .MINUS(gnd_), .PLUS(gnd_), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(net83), .PLUS(net74), .BULK(GND_));
rppolywo_m  R1 ( .MINUS(gnd_), .PLUS(net83), .BULK(GND_));
ml_vpp_vco Ivpx_vpp_vco ( .pbias_25(pbias_25), .slow_25(net86),
     .freq_25({freq_25[1], freq_buf_b_25[0]}), .en_25(pumpen_25),
     .clk_25_0(vpxa_clk_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_ctrl, View - schematic
// LAST TIME SAVED: Oct 28 15:48:54 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_vpxa_ctrl ( pumpen, pumpen_25, vpxa_2_vdd, fsm_pumpen,
     fsm_tm_xforce, fsm_tm_xvpxaint );
output  pumpen, pumpen_25, vpxa_2_vdd;

input  fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I73 ( .A(fsm_tm_xvpxaint), .B(fsm_tm_xforce), .Y(net042));
inv_25 I38 ( .IN(net045), .OUT(pumpen_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I173 ( .in(net049), .sup(vddp_), .out_vddio_b(net045),
     .out_vddio(net046), .in_b(net075));
nor2_hvt I72 ( .A(vpxa_off), .B(net065), .Y(net049));
nor2_hvt I69 ( .A(vpxa_2_vdd), .B(vpxa_2_vdd), .Y(net043));
inv_hvt I75 ( .A(net049), .Y(net056));
inv_hvt I76 ( .A(net056), .Y(pumpen));
inv_hvt I110 ( .A(net049), .Y(net075));
inv_hvt I74 ( .A(net042), .Y(net065));
inv_hvt I131 ( .A(fsm_pumpen), .Y(vpxa_2_vdd));
inv_hvt I70 ( .A(net043), .Y(vpxa_off));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff_25, View - schematic
// LAST TIME SAVED: Feb 11 11:37:05 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_dff_25 ( Q_25, Q_B_25, CLK_25, D_25, R_25 );
output  Q_25, Q_B_25;

input  CLK_25, D_25, R_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I87 ( .IN(net044), .OUT(net038), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I72 ( .IN(CLK_25), .OUT(net044), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I90 ( .IN(Q_25), .OUT(Q_B_25), .P(vddp_), .Pb(vddp_), .G(GND_),
     .Gb(GND_));
ml_dlatch_25 Ilatch2 ( .D_25(net053), .EN_25(net038), .R_25(R_25),
     .Q_25(Q_25));
ml_dlatch_25 Ilatch1 ( .Q_25(net053), .EN_25(net044), .D_25(D_25),
     .R_25(R_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_n, View - schematic
// LAST TIME SAVED: Feb  5 15:08:44 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp_n ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M0 ( .D(out_div), .B(vddp_), .G(out_ref), .S(vddp_));
pch_25  M4 ( .D(out_ref), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M5 ( .D(out_div), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M7 ( .D(out_ref), .B(vddp_), .G(out_ref), .S(vddp_));
nch_25  M1 ( .D(out_div), .B(GND_), .G(in_div), .S(net049));
nch_25  M2 ( .D(out_ref), .B(GND_), .G(in_ref), .S(net049));
nch_25  M6_1_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net049), .B(GND_), .G(sa_bias), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_top_n, View - schematic
// LAST TIME SAVED: Feb 21 13:55:00 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp_top_n ( pump_chrg_25, in_div, in_ref, sa_bias,
     saen_25 );
output  pump_chrg_25;

input  in_div, in_ref, sa_bias, saen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_25 I103 ( .G(gnd_), .Pb(vddp_), .A(saen_25), .Y(chrg_b_25),
     .P(vddp_), .B(net27), .Gb(gnd_));
nch_25  M6_1_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M6_0_ ( .D(net087), .B(GND_), .G(sa_bias), .S(gnd_));
inv_25 I102 ( .IN(chrg_b_25), .OUT(pump_chrg_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I104 ( .IN(out_div2), .OUT(net27), .P(vddp_), .Pb(vddp_),
     .G(net087), .Gb(gnd_));
ml_core_sa_comp_n Icore_sa_comp_n0 ( .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp_n Iml_core_sa_comp_n1 ( .out_div(out_div2),
     .out_ref(out_ref2), .in_div(in_div2), .in_ref(in_ref2),
     .sa_bias(sa_bias), .saen_25(saen_25));

endmodule
// Library - NVCM, Cell - ml_vpxa_reg, View - schematic
// LAST TIME SAVED: May  3 13:50:36 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_vpxa_reg ( freq_25, pump_chrg_0_25, pump_chrg_1_25,
     pump_chrg_2_25, vpxa_int, bgr, fsm_vrdwl, pumpen, vpxa_clk_25 );
output  pump_chrg_0_25, pump_chrg_1_25, pump_chrg_2_25;

inout  vpxa_int;

input  bgr, pumpen, vpxa_clk_25;

output [1:0]  freq_25;

input [2:0]  fsm_vrdwl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  freq_in_25;

wire  [0:2]  vrdwl_vpxa;

wire  [0:2]  vrdwl_b_vpxa;



nand2_25 I145 ( .G(GND_), .Pb(vddp_), .A(net0171), .Y(freq_in_25[0]),
     .P(vddp_), .B(net0179), .Gb(GND_));
nand2_25 I158 ( .G(GND_), .Pb(vddp_), .A(net0179), .Y(freq_in_25[1]),
     .P(vddp_), .B(net0163), .Gb(GND_));
nand3_25 I44 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0179),
     .C(pump_chrg_0_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I149 ( .B(pump_chrg_1_b_25), .A(pump_chrg_2_25), .Y(net0171),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
nand3_25 I159 ( .B(pump_chrg_1_25), .A(pump_chrg_2_25), .Y(net0163),
     .C(pump_chrg_0_b_25), .P(vddp_), .Pb(vddp_), .Gb(GND_), .G(GND_));
ml_dff_25 I125 ( .Q_B_25(net0187), .R_25(saen_b_25),
     .D_25(freq_in_25[1]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[1]));
ml_dff_25 I126 ( .Q_B_25(net0192), .R_25(saen_b_25),
     .D_25(freq_in_25[0]), .CLK_25(vpxa_clk_25), .Q_25(freq_25[0]));
inv_hvt I85 ( .A(net171), .Y(net175));
inv_hvt I183 ( .A(fsm_vrdwl[2]), .Y(net171));
inv_hvt I83 ( .A(pumpen), .Y(net143));
inv_hvt I82 ( .A(net143), .Y(net145));
inv_hvt I184 ( .A(fsm_vrdwl[1]), .Y(net176));
inv_hvt I187 ( .A(fsm_vrdwl[0]), .Y(net181));
inv_hvt I186 ( .A(net181), .Y(net185));
inv_hvt I185 ( .A(net176), .Y(net180));
inv_25 I155 ( .IN(pump_chrg_0_25), .OUT(pump_chrg_0_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
inv_25 I63 ( .IN(net169), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I75 ( .IN(net168), .OUT(saen_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));
inv_25 I154 ( .IN(pump_chrg_1_25), .OUT(pump_chrg_1_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_ls_vdd2vdd25 I191 ( .in(saen_25), .sup(vpxa_int),
     .out_vddio_b(saen_b_vpxa), .out_vddio(net0210), .in_b(saen_b_25));
ml_ls_vdd2vdd25 I335 ( .in(net145), .sup(vddp_), .out_vddio_b(net168),
     .out_vddio(net169), .in_b(net143));
ml_ls_vdd2vdd25 I87 ( .in(net171), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[2]), .out_vddio(vrdwl_b_vpxa[2]),
     .in_b(net175));
ml_ls_vdd2vdd25 I98 ( .in(net176), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[1]), .out_vddio(vrdwl_b_vpxa[1]),
     .in_b(net180));
ml_ls_vdd2vdd25 I99 ( .in(net181), .sup(vpxa_int),
     .out_vddio_b(vrdwl_vpxa[0]), .out_vddio(vrdwl_b_vpxa[0]),
     .in_b(net185));
ml_core_sa_comp_top_n Icore_sa_comp_top_n2 (
     .pump_chrg_25(pump_chrg_2_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_2));
ml_core_sa_comp_top_n core_sa_comp_top_n0 (
     .pump_chrg_25(pump_chrg_0_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_0));
ml_core_sa_comp_top_n Icore_sa_comp_top_n1 (
     .pump_chrg_25(pump_chrg_1_25), .saen_25(saen_25),
     .sa_bias(sa_bias), .in_ref(bgr), .in_div(in_div_1));
rppolywo_m  R29 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R28 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R20 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R27 ( .MINUS(in_div_2), .PLUS(in_div_1), .BULK(GND_));
rppolywo_m  R26 ( .MINUS(in_div_0), .PLUS(net202), .BULK(GND_));
rppolywo_m  R17 ( .MINUS(net232), .PLUS(net223), .BULK(GND_));
rppolywo_m  R2 ( .MINUS(net270), .PLUS(net226), .BULK(GND_));
rppolywo_m  R18 ( .MINUS(net226), .PLUS(net229), .BULK(GND_));
rppolywo_m  R0 ( .MINUS(sa_bias), .PLUS(net232), .BULK(GND_));
rppolywo_m  R10 ( .MINUS(net202), .PLUS(net237), .BULK(GND_));
rppolywo_m  R3 ( .MINUS(net237), .PLUS(net270), .BULK(GND_));
rppolywo_m  R30 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
rppolywo_m  R12 ( .MINUS(gnd_), .PLUS(in_div_2), .BULK(GND_));
rppolywo_m  R31 ( .MINUS(in_div_1), .PLUS(in_div_0), .BULK(GND_));
pch_25  M3 ( .D(net229), .B(vpxa_int), .G(saen_b_vpxa), .S(vpxa_int));
pch_25  M11_1_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M11_0_ ( .D(in_div_0), .B(in_div_0), .G(vpxa_int),
     .S(in_div_0));
pch_25  M15 ( .D(net237), .B(vpxa_int), .G(vrdwl_vpxa[0]), .S(net270));
pch_25  M37 ( .D(net226), .B(vpxa_int), .G(vrdwl_vpxa[2]), .S(net229));
pch_25  M1 ( .D(net223), .B(vddp_), .G(saen_b_25), .S(vddp_));
pch_25  M14 ( .D(net270), .B(vpxa_int), .G(vrdwl_vpxa[1]), .S(net226));
pch_25  M8_1_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
pch_25  M8_0_ ( .D(net270), .B(net270), .G(vpxa_int), .S(net270));
nch_25  M2 ( .D(sa_bias), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M32 ( .D(net229), .B(GND_), .G(vrdwl_b_vpxa[2]), .S(net226));
nch_25  M0_3_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_2_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_1_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M0_0_ ( .D(sa_bias), .B(GND_), .G(sa_bias), .S(gnd_));
nch_25  M9 ( .D(net270), .B(GND_), .G(vrdwl_b_vpxa[0]), .S(net237));
nch_25  M7 ( .D(net226), .B(GND_), .G(vrdwl_b_vpxa[1]), .S(net270));

endmodule
// Library - NVCM, Cell - ml_hv2vdd_sw, View - schematic
// LAST TIME SAVED: Apr  8 14:27:39 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_hv2vdd_sw ( out_hv, hv2vdd, vddp_tieh );
inout  out_hv;

input  hv2vdd, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M1 ( .D(net27), .B(GND_), .G(vddp_tieh), .S(out_hv));
nch_na25  M2 ( .D(vdd_), .B(GND_), .G(hv2vdd_25), .S(net27));
inv_25 I62 ( .IN(net40), .OUT(hv2vdd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
ml_ls_vdd2vdd25 I64 ( .in(net44), .sup(vddp_), .out_vddio_b(net40),
     .out_vddio(net37), .in_b(net46));
inv_hvt I65 ( .A(hv2vdd), .Y(net46));
inv_hvt I66 ( .A(net46), .Y(net44));

endmodule
// Library - NVCM, Cell - ml_vpxa_top, View - schematic
// LAST TIME SAVED: Sep  3 10:36:27 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_vpxa_top ( vpxa_int, bgr, fsm_pumpen, fsm_tm_xforce,
     fsm_tm_xvpxaint, fsm_vrdwl );
inout  vpxa_int;

input  bgr, fsm_pumpen, fsm_tm_xforce, fsm_tm_xvpxaint;

input [2:0]  fsm_vrdwl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  freq_25;



nmoscap_25  C7 ( .MINUS(gnd_), .PLUS(vpxa_int));
ml_pump_vpxa_x2 Ipump_vpxa_x3 ( .pumpen(pumpen),
     .vpxa_clk_b_25(vpxa_clk_b_25), .vpxa_clk_25(vpxa_clk_25),
     .pumpen_25(pumpen_25), .pump_chrg_2_25(pump_chrg_2_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_0_25(pump_chrg_0_25),
     .vpxa_int(vpxa_int));
inv_25 I73 ( .IN(vpxa_clk_25), .OUT(vpxa_clk_b_25), .P(vddp_),
     .Pb(vddp_), .G(GND_), .Gb(GND_));
ml_vpxa_osc Ivpxa_osc ( .freq_25(freq_25[1:0]), .bgr(bgr),
     .pumpen_25(pumpen_25), .vpxa_clk_25(vpxa_clk_25));
ml_vpxa_ctrl Ivpxa_ctrl ( .fsm_pumpen(fsm_pumpen), .pumpen(pumpen),
     .pumpen_25(pumpen_25), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .vpxa_2_vdd(vpxa_2_vdd));
vddp_tiehigh I118_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I118_0_ ( .vddp_tieh(vddp_tieh));
ml_vpxa_reg Ivpxa_reg ( .pump_chrg_0_25(pump_chrg_0_25),
     .pump_chrg_1_25(pump_chrg_1_25), .pump_chrg_2_25(pump_chrg_2_25),
     .freq_25(freq_25[1:0]), .vpxa_clk_25(vpxa_clk_25),
     .pumpen(pumpen), .fsm_vrdwl(fsm_vrdwl[2:0]), .bgr(bgr),
     .vpxa_int(vpxa_int));
ml_hv2vdd_sw Ivpxa_2vdd_sw ( .vddp_tieh(vddp_tieh),
     .hv2vdd(vpxa_2_vdd), .out_hv(vpxa_int));

endmodule
// Library - NVCM, Cell - ml_hvmux_top_ctrl, View - schematic
// LAST TIME SAVED: May  2 18:30:47 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_hvmux_top_ctrl ( bgrext_en, bgrint_en, en_vblinhi,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp, fsm_lshven,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint, fsm_wgnden,
     fsm_wpen, tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );
output  bgrext_en, bgrint_en, en_vblinhi, ngate_vddp, ngate_vpxa,
     sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint,
     vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint, vpxaint_ext,
     vtmode, ysup25_2vdd, ysup25_2vddp;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_testdec,
     tm_wleqbl, vpint_en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



mux2_hvt I260 ( .in1(fsm_wgnden), .in0(fsm_wpen), .out(net0217),
     .sel(pgmpulse_b));
vdd_tielow I136 ( .gnd_tiel(gnd_tiel));
anor21_hvt I245 ( .A(net0189), .B(net0193), .Y(vppint_ext),
     .C(net0188));
anor21_hvt I109 ( .A(net0201), .B(net0199), .Y(vpxa_ext), .C(net0188));
nand3_hvt I248 ( .Y(net0189), .B(vpint_en), .C(fsm_tm_xvppint),
     .A(fsm_tm_xforce));
nand3_hvt I246 ( .Y(net0201), .B(vddp_rd_b), .C(fsm_tm_xvpxa),
     .A(fsm_tm_xforce));
nand3_hvt I247 ( .Y(net0193), .B(pmprd), .C(pmprd),
     .A(fsm_tm_xvppint));
nand3_hvt I35 ( .C(fsm_lshven), .A(fsm_pgm), .Y(pgmpulse_b),
     .B(net0327));
nand3_hvt I205 ( .Y(net0213), .B(net0321), .C(pgmpulse_b),
     .A(net0321));
nand3_hvt I240 ( .C(pmprd), .A(fsm_tm_xvpxa), .Y(net0199), .B(pmprd));
nor2_hvt I213 ( .A(net0324), .B(fsm_nvcmen_b), .Y(net0251));
nor2_hvt I224 ( .A(vddp_rd_b), .B(net0258), .Y(vpxa_vppd));
nor2_hvt I214 ( .A(net0251), .B(net0266), .Y(sbhvsup_vppint));
nor2_hvt I215 ( .A(net0264), .B(net0311), .Y(sbhvsup_vddp));
nor2_hvt I183 ( .A(net87), .B(net73), .Y(ysup25_2vddp));
nor2_hvt I14 ( .A(net75), .B(net93), .Y(ysup25_2vdd));
nor2_hvt I207 ( .A(net0325), .B(net0260), .Y(sb25sup_vddp));
nor2_hvt I206 ( .A(net0268), .B(net0213), .Y(sb25sup_vpxa));
nor2_hvt I185 ( .A(gnd_tiel), .B(gnd_tiel), .Y(net0240));
nor2_hvt I223 ( .B(net0240), .Y(vddp_rd), .A(net0349));
nor2_hvt I195 ( .A(net0272), .B(rd_vddp), .Y(ngate_vpxa));
nor2_hvt I196 ( .A(net0331), .B(net0270), .Y(ngate_vddp));
nor2_hvt I225 ( .A(net0256), .B(vddp_rd), .Y(vpxa_vpxaint));
ml_pump_a_clkdly I219 ( .in(ysup25_2vddp_b), .out(net75));
ml_pump_a_clkdly I227 ( .in(net0297), .out(net0256));
ml_pump_a_clkdly I226 ( .in(net0319), .out(net0258));
ml_pump_a_clkdly I209 ( .in(net0323), .out(net0260));
ml_pump_a_clkdly I184 ( .in(ysup25_2vdd_b), .out(net73));
ml_pump_a_clkdly I217 ( .in(net0313), .out(net0264));
ml_pump_a_clkdly I216 ( .in(net0309), .out(net0266));
ml_pump_a_clkdly I208 ( .in(net0329), .out(net0268));
ml_pump_a_clkdly I198 ( .in(net0339), .out(net0270));
ml_pump_a_clkdly I197 ( .in(net0335), .out(net0272));
nand2_hvt I254 ( .A(bgrext_en), .Y(bgrint_en), .B(fsm_tm_xforce));
nand2_hvt I104 ( .A(fsm_nvcmen), .Y(net77), .B(tm_wleqbl));
nand2_hvt I179 ( .A(fsm_nvcmen), .Y(net80), .B(net0217));
nand2_hvt I252 ( .A(fsm_nvcmen_buf), .Y(net0277), .B(fsm_tm_xvbg));
nand2_hvt I234 ( .A(fsm_pumpen), .Y(net0286), .B(fsm_tm_xvpxaint));
inv_hvt I259 ( .A(pgmpulse_b), .Y(net0324));
inv_hvt I229 ( .A(vpxa_vppd), .Y(net0297));
inv_hvt I250 ( .A(fsm_pumpen), .Y(net0188));
inv_hvt I182 ( .A(ysup25_2vdd), .Y(ysup25_2vdd_b));
inv_hvt I230 ( .A(vddp_rd), .Y(vddp_rd_b));
inv_hvt I249 ( .A(pgmpulse_b), .Y(pgmpulse));
inv_hvt I131 ( .A(fsm_nvcmen), .Y(fsm_nvcmen_b));
inv_hvt I178 ( .A(net77), .Y(vtmode));
inv_hvt I180 ( .A(net80), .Y(net93));
inv_hvt I253 ( .A(net0277), .Y(bgrext_en));
inv_hvt I218 ( .A(sbhvsup_vddp), .Y(net0309));
inv_hvt I221 ( .A(net0251), .Y(net0311));
inv_hvt I220 ( .A(sbhvsup_vppint), .Y(net0313));
inv_hvt I134 ( .A(net93), .Y(net87));
inv_hvt I181 ( .A(ysup25_2vddp), .Y(ysup25_2vddp_b));
inv_hvt I228 ( .A(vpxa_vpxaint), .Y(net0319));
inv_hvt I204 ( .A(rd_vddp), .Y(net0321));
inv_hvt I212 ( .A(sb25sup_vpxa), .Y(net0323));
inv_hvt I210 ( .A(net0213), .Y(net0325));
inv_hvt I202 ( .A(fsm_pgmvfy), .Y(net0327));
inv_hvt I211 ( .A(sb25sup_vddp), .Y(net0329));
inv_hvt I199 ( .A(rd_vddp), .Y(net0331));
inv_hvt I236 ( .A(fsm_tm_xforce), .Y(pmprd));
inv_hvt I200 ( .A(ngate_vddp), .Y(net0335));
inv_hvt I235 ( .A(net0286), .Y(vpxaint_ext));
inv_hvt I201 ( .A(ngate_vpxa), .Y(net0339));
inv_hvt I233 ( .A(fsm_nvcmen_b), .Y(fsm_nvcmen_buf));
nor3_hvt I105 ( .B(tm_testdec), .Y(en_vblinhi), .A(fsm_nvcmen_b),
     .C(tm_allbl_l));
nor3_hvt I186 ( .C(fsm_rd), .A(fsm_tm_rd_mode), .B(fsm_pgmvfy),
     .Y(net0349));
nor3_hvt I187 ( .B(net0240), .Y(rd_vddp), .A(net0349),
     .C(fsm_nvcmen_b));

endmodule
// Library - misc, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jul  3 16:54:18 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_dff ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));
nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));

endmodule
// Library - NVCM, Cell - ml_hvmux_ls25, View - schematic
// LAST TIME SAVED: Feb 15 14:23:11 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_hvmux_ls25 ( bgrext_en_25, bgrint_en_25, ngate_vddp_25,
     ngate_vpxa_25, sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25, bgrext_en, bgrint_en,
     ngate_vddp, ngate_vpxa, sb25sup_vddp, sb25sup_vpxa, sbhvsup_vddp,
     sbhvsup_vppint, vppint_ext, vpxa_ext, vpxa_vppd, vpxa_vpxaint,
     vpxaint_ext, vtmode, ysup25_2vdd, ysup25_2vddp );
output  bgrext_en_25, bgrint_en_25, ngate_vddp_25, ngate_vpxa_25,
     sb25sup_vddp_25, sb25sup_vpxa_25, sbhvsup_vddp_25,
     sbhvsup_vppint_25, vppint_ext_25, vpxa_ext_25, vpxa_vppd_25,
     vpxa_vpxaint_25, vpxaint_ext_25, vtmode_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25;

input  bgrext_en, bgrint_en, ngate_vddp, ngate_vpxa, sb25sup_vddp,
     sb25sup_vpxa, sbhvsup_vddp, sbhvsup_vppint, vppint_ext, vpxa_ext,
     vpxa_vppd, vpxa_vpxaint, vpxaint_ext, vtmode, ysup25_2vdd,
     ysup25_2vddp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I317 ( .A(net054), .Y(net052));
inv_hvt I314 ( .A(vpxa_vppd), .Y(net054));
inv_hvt I327 ( .A(net066), .Y(net056));
inv_hvt I329 ( .A(bgrint_en), .Y(net058));
inv_hvt I321 ( .A(vpxaint_ext), .Y(net060));
inv_hvt I320 ( .A(net060), .Y(net062));
inv_hvt I325 ( .A(net082), .Y(net064));
inv_hvt I326 ( .A(vppint_ext), .Y(net066));
inv_hvt I312 ( .A(bgrext_en), .Y(net068));
inv_hvt I313 ( .A(net068), .Y(net070));
inv_hvt I328 ( .A(net058), .Y(net0487));
inv_hvt I239 ( .A(sb25sup_vpxa), .Y(net0486));
inv_hvt I319 ( .A(net0112), .Y(net0488));
inv_hvt I240 ( .A(net0486), .Y(net080));
inv_hvt I324 ( .A(vpxa_ext), .Y(net082));
inv_hvt I206 ( .A(vtmode), .Y(net084));
inv_hvt I213 ( .A(ysup25_2vdd), .Y(net086));
inv_hvt I214 ( .A(net086), .Y(net088));
inv_hvt I205 ( .A(net084), .Y(net090));
inv_hvt I216 ( .A(net088), .Y(net092));
inv_hvt I110 ( .A(net072), .Y(net074));
inv_hvt I227 ( .A(net098), .Y(net096));
inv_hvt I228 ( .A(ngate_vddp), .Y(net098));
inv_hvt I217 ( .A(net092), .Y(ysup25_2vdd_buf));
inv_hvt I190 ( .A(ysup25_2vddp), .Y(net072));
inv_hvt I219 ( .A(ngate_vpxa), .Y(net0104));
inv_hvt I220 ( .A(net0104), .Y(net0106));
inv_hvt I232 ( .A(sb25sup_vddp), .Y(net0108));
inv_hvt I231 ( .A(net0108), .Y(net0110));
inv_hvt I323 ( .A(vpxa_vpxaint), .Y(net0112));
inv_hvt I256 ( .A(net0116), .Y(net0114));
inv_hvt I257 ( .A(sbhvsup_vddp), .Y(net0116));
inv_hvt I258 ( .A(net0120), .Y(net0118));
inv_hvt I259 ( .A(sbhvsup_vppint), .Y(net0120));
ml_ls_vdd2vdd25 I336 ( .in(net064), .sup(vddp_), .out_vddio_b(net0123),
     .out_vddio(net0207), .in_b(net082));
ml_ls_vdd2vdd25 I337 ( .in(net056), .sup(vddp_), .out_vddio_b(net0128),
     .out_vddio(net0208), .in_b(net066));
ml_ls_vdd2vdd25 I338 ( .in(net052), .sup(vddp_), .out_vddio_b(net0133),
     .out_vddio(net0211), .in_b(net054));
ml_ls_vdd2vdd25 I339 ( .in(net0487), .sup(vddp_),
     .out_vddio_b(net0138), .out_vddio(net0209), .in_b(net058));
ml_ls_vdd2vdd25 I332 ( .in(net070), .sup(vddp_), .out_vddio_b(net0148),
     .out_vddio(net0149), .in_b(net068));
ml_ls_vdd2vdd25 I238 ( .in(net080), .sup(vddp_), .out_vddio_b(net0153),
     .out_vddio(net0154), .in_b(net0486));
ml_ls_vdd2vdd25 I334 ( .in(net062), .sup(vddp_), .out_vddio_b(net0158),
     .out_vddio(net0214), .in_b(net060));
ml_ls_vdd2vdd25 I335 ( .in(net0488), .sup(vddp_),
     .out_vddio_b(net0163), .out_vddio(net0206), .in_b(net0112));
ml_ls_vdd2vdd25 I212 ( .in(net088), .sup(vddp_), .out_vddio_b(net0168),
     .out_vddio(net0169), .in_b(net086));
ml_ls_vdd2vdd25 I226 ( .in(net096), .sup(vddp_), .out_vddio_b(net0173),
     .out_vddio(net0174), .in_b(net098));
ml_ls_vdd2vdd25 I203 ( .in(net072), .sup(vddp_), .out_vddio_b(net077),
     .out_vddio(net078), .in_b(net074));
ml_ls_vdd2vdd25 I221 ( .in(net0106), .sup(vddp_),
     .out_vddio_b(net0183), .out_vddio(net0184), .in_b(net0104));
ml_ls_vdd2vdd25 I233 ( .in(net0110), .sup(vddp_),
     .out_vddio_b(net0188), .out_vddio(net0219), .in_b(net0108));
ml_ls_vdd2vdd25 I207 ( .in(net090), .sup(vddp_), .out_vddio_b(net0193),
     .out_vddio(net0194), .in_b(net084));
ml_ls_vdd2vdd25 I260 ( .in(net0114), .sup(vddp_),
     .out_vddio_b(net0198), .out_vddio(net0220), .in_b(net0116));
ml_ls_vdd2vdd25 I261 ( .in(net0118), .sup(vddp_),
     .out_vddio_b(net0203), .out_vddio(net0204), .in_b(net0120));
inv_25 I390 ( .IN(net0148), .OUT(bgrext_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I384 ( .IN(net0163), .OUT(vpxa_vpxaint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I386 ( .IN(net0133), .OUT(vpxa_vppd_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I388 ( .IN(net0123), .OUT(vpxa_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I376 ( .IN(net0168), .OUT(ysup25_2vdd_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I387 ( .IN(net0158), .OUT(vpxaint_ext_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I389 ( .IN(net0128), .OUT(vppint_ext_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I362 ( .IN(net077), .OUT(ysup25_2vddp_b_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I383 ( .IN(net0203), .OUT(sbhvsup_vppint_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I379 ( .IN(net0183), .OUT(ngate_vpxa_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I377 ( .IN(net0193), .OUT(vtmode_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I378 ( .IN(net0173), .OUT(ngate_vddp_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I381 ( .IN(net0153), .OUT(sb25sup_vpxa_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I382 ( .IN(net0198), .OUT(sbhvsup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I380 ( .IN(net0188), .OUT(sb25sup_vddp_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I391 ( .IN(net0138), .OUT(bgrint_en_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_bgrxcvr, View - schematic
// LAST TIME SAVED: Apr  8 10:30:41 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_hvmux_bgrxcvr ( bgr, bgr_int, bgrint_en_25, vpp,
     bgrext_en_25, vddp_tieh );
inout  bgr, bgr_int, bgrint_en_25, vpp;

input  bgrext_en_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M0 ( .D(bgr), .B(GND_), .G(bgrint_en_25), .S(bgr_int));
nch_25  M2 ( .D(vpp), .B(GND_), .G(vddp_tieh), .S(net53));
nch_25  M3 ( .D(net53), .B(GND_), .G(bgrext_en_25), .S(bgr));

endmodule
// Library - NVCM, Cell - ml_ysup_25_switch, View - schematic
// LAST TIME SAVED: Apr  8 10:33:54 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_ysup_25_switch ( vdd, vddp, ysup_25, ysup25_2vdd_25,
     ysup25_2vdd_buf, ysup25_2vddp_b_25 );
inout  vdd, vddp, ysup_25;

input  ysup25_2vdd_25, ysup25_2vdd_buf, ysup25_2vddp_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd), .B(GND_), .G(ysup25_2vdd_25), .S(ysup_25));
pch_25  M5 ( .D(net73), .B(vddp), .G(ysup25_2vddp_b_25), .S(vddp));
pch_25  M0 ( .D(ysup_25), .B(ysup_25), .G(ysup25_2vdd_buf), .S(net73));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_vblinhi, View - schematic
// LAST TIME SAVED: Feb  1 08:51:27 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_vblinhi ( vblinhi, vpxa, en_vblinhi, vtmode,
     vtmode_25 );
inout  vblinhi, vpxa;

input  en_vblinhi, vtmode, vtmode_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I191 ( .A(en_vblinhi), .B(vtmode_buf), .Y(ngate_inhi_lv));
nand2_hvt I104 ( .A(net063), .Y(pgate_inhi_lv), .B(en_vblinhi));
inv_hvt I110 ( .A(net063), .Y(vtmode_buf));
inv_hvt I190 ( .A(vtmode), .Y(net063));
nch_25  M9 ( .D(net062), .B(GND_), .G(net062), .S(vblinhi));
nch_25  M8 ( .D(vpxa), .B(GND_), .G(vtmode_25), .S(net062));
pch_hvt  M7_1_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
pch_hvt  M7_0_ ( .D(vblinhi), .B(vdd_), .G(pgate_inhi_lv), .S(vdd_));
nch_hvt  M0_1_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));
nch_hvt  M0_0_ ( .D(vblinhi), .B(GND_), .G(ngate_inhi_lv), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hvmux_top, View - schematic
// LAST TIME SAVED: May  2 18:49:30 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_hvmux_top ( bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv,
     vblinhi, vpp, vpp_int, vpxa, vpxa_int, ysup_25, fsm_lshven,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_tm_rd_mode, fsm_tm_xforce, fsm_tm_xvbg,
     fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint, fsm_wgnden,
     fsm_wpen, tm_allbl_l, tm_testdec, tm_wleqbl, vpint_en );
inout  bgr, bgr_int, ngate_25, sb25sup_25, sbhvsup_hv, vblinhi, vpp,
     vpp_int, vpxa, vpxa_int, ysup_25;

input  fsm_lshven, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_tm_rd_mode,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa,
     fsm_tm_xvpxaint, fsm_wgnden, fsm_wpen, tm_allbl_l, tm_testdec,
     tm_wleqbl, vpint_en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_hv_hotswitch_enhance Ixcvr_vppint ( .vddp_tieh(vddp_tieh),
     .selhv_25(vppint_ext_25), .hv_in_hv(vpp_int), .hv_out_hv(vpp));
ml_hvmux_top_ctrl Ihvmux_top_ctrl ( .vpint_en(vpint_en),
     .fsm_wpen(fsm_wpen), .tm_wleqbl(tm_wleqbl),
     .tm_testdec(tm_testdec), .tm_allbl_l(tm_allbl_l),
     .fsm_wgnden(fsm_wgnden), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvpxa(fsm_tm_xvpxa), .fsm_tm_xvppint(fsm_tm_xvppint),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_rd(fsm_rd),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy),
     .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_lshven(fsm_lshven),
     .ysup25_2vddp(ysup25_2vddp), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vppint(sbhvsup_vppint), .sbhvsup_vddp(sbhvsup_vddp),
     .sb25sup_vpxa(sb25sup_vpxa), .sb25sup_vddp(sb25sup_vddp),
     .ngate_vpxa(ngate_vpxa), .ngate_vddp(ngate_vddp),
     .en_vblinhi(en_vblinhi), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en));
ml_hvmux_ls25 Ihvmux_ls25 ( .ysup25_2vddp(ysup25_2vddp),
     .sbhvsup_vppint(sbhvsup_vppint),
     .sbhvsup_vppint_25(sbhvsup_vppint_25), .ysup25_2vdd(ysup25_2vdd),
     .vtmode(vtmode), .vpxaint_ext(vpxaint_ext),
     .vpxa_vpxaint(vpxa_vpxaint), .vpxa_vppd(vpxa_vppd),
     .vpxa_ext(vpxa_ext), .vppint_ext(vppint_ext),
     .sbhvsup_vddp(sbhvsup_vddp), .sb25sup_vpxa(sb25sup_vpxa),
     .sb25sup_vddp(sb25sup_vddp), .ngate_vpxa(ngate_vpxa),
     .ngate_vddp(ngate_vddp), .bgrint_en(bgrint_en),
     .bgrext_en(bgrext_en), .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vtmode_25(vtmode_25),
     .vpxaint_ext_25(vpxaint_ext_25),
     .vpxa_vpxaint_25(vpxa_vpxaint_25), .vpxa_vppd_25(vpxa_vppd_25),
     .vpxa_ext_25(net164), .vppint_ext_25(vppint_ext_25),
     .sbhvsup_vddp_25(sbhvsup_vddp_25),
     .sb25sup_vpxa_25(sb25sup_vpxa_25),
     .sb25sup_vddp_25(sb25sup_vddp_25), .ngate_vpxa_25(ngate_vpxa_25),
     .ngate_vddp_25(ngate_vddp_25), .bgrint_en_25(bgrint_en_25),
     .bgrext_en_25(bgrext_en_25));
ml_hvmux_bgrxcvr Ixcvr_bgr ( .vddp_tieh(vddp_tieh),
     .bgrext_en_25(bgrext_en_25), .vpp(vpp),
     .bgrint_en_25(bgrint_en_25), .bgr_int(bgr_int), .bgr(bgr));
ml_hv_hotswitch Ixcvr_vpxa_int ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa_int), .hv_out_hv(vpp));
ml_hv_hotswitch Ixcvr_vpxa ( .vddp_tieh(vddp_tieh),
     .selhv_25(vpxaint_ext_25), .hv_in_hv(vpxa), .hv_out_hv(vpp));
ml_hvmux_hotswitch Isw_sbhvsup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sbhvsup_vppint_25), .sel_hv_a_25(sbhvsup_vddp_25),
     .out_hv(sbhvsup_hv), .hvin_b_hv(vpp_int), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_sb25sup ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(sb25sup_vpxa_25), .sel_hv_a_25(sb25sup_vddp_25),
     .out_hv(sb25sup_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_ngate ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(ngate_vpxa_25), .sel_hv_a_25(ngate_vddp_25),
     .out_hv(ngate_25), .hvin_b_hv(vpxa), .hvin_a_hv(vddp_));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_1_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vpxa_int), .hvin_a_hv(vpxa_int));
ml_hvmux_hotswitch Isw_vpxa_int_vddp_0_ ( .vddp_tieh(vddp_tieh),
     .sel_hv_b_25(vpxa_vppd_25), .sel_hv_a_25(vpxa_vpxaint_25),
     .out_hv(vpxa), .hvin_b_hv(vpxa_int), .hvin_a_hv(vpxa_int));
ml_ysup_25_switch Isw_ysup25_1_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
ml_ysup_25_switch Isw_ysup25_0_ (
     .ysup25_2vddp_b_25(ysup25_2vddp_b_25),
     .ysup25_2vdd_buf(ysup25_2vdd_buf),
     .ysup25_2vdd_25(ysup25_2vdd_25), .vdd(vdd_), .ysup_25(ysup_25),
     .vddp(vddp_));
vddp_tiehigh I188_9_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_8_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I188_0_ ( .vddp_tieh(vddp_tieh));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_1_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));
ml_ymux_ctrl_vblinhi Isw_ymux_ctrl_vblinhi_0_ ( .vtmode(vtmode),
     .vtmode_25(vtmode_25), .en_vblinhi(en_vblinhi), .vpxa(vpxa),
     .vblinhi(vblinhi));

endmodule
// Library - NVCM, Cell - ml_chip_nvcm_8f, View - schematic
// LAST TIME SAVED: Sep 11 17:55:36 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_chip_nvcm_8f ( nv_dataout, vpp, fsm_blkadd, fsm_blkadd_b,
     fsm_coladd, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rowadd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint,
     fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_trim_vbg,
     fsm_vpgmwl, fsm_vpxaset, fsm_vrdwl, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl
     );

inout  vpp;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_rst_b, fsm_sample,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvppint, fsm_tm_xvpxa, fsm_tm_xvpxaint,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     tm_allbank_sel, tm_allbl_h, tm_allbl_l, tm_allwl_h, tm_allwl_l,
     tm_dma, tm_tcol, tm_testdec_wr, tm_wleqbl;

output [8:0]  nv_dataout;

input [7:0]  fsm_rowadd;
input [3:0]  fsm_trim_vbg;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_vpgmwl;
input [3:0]  fsm_trim_ipp;
input [2:0]  fsm_vrdwl;
input [3:0]  fsm_blkadd_b;
input [9:0]  fsm_coladd;
input [2:0]  fsm_trim_rrefpgm;
input [2:0]  fsm_trim_rrefrd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  fsm_trim_ipp_buf;

wire  [2:0]  fsm_trim_rrefpgm_buf;

wire  [7:0]  fsm_rowadd_buf;

wire  [3:0]  fsm_blkadd_b_buf;

wire  [3:0]  fsm_blkadd_buf;

wire  [2:0]  fsm_trim_rrefred_buf;

wire  [9:0]  fsm_coladd_buf;

wire  [3:0]  fsm_trim_vbg_buf;

wire  [3:0]  nv_dataout_unbuf;

wire  [2:0]  fsm_vpgmwl_buf;



ml_chip_spare Ich_spare_1 ( );
ml_chip_spare Ich_spare_2 ( );
ml_chip_buf_top_8f Ichip_buf_top ( .fsm_rst_b_buf(fsm_rst_b_buf),
     .tm_allbank_sel_buf(tm_allbank_sel_buf),
     .tm_allbank_sel(tm_allbank_sel), .nv_dataout_buf(nv_dataout[3:0]),
     .nv_dataout(nv_dataout_unbuf[3:0]), .tm_dma_buf(tm_dma_buf),
     .fsm_wren_buf(fsm_wren_buf), .fsm_pgmhv_buf(fsm_pgmhv_buf),
     .fsm_gwlbdis_buf(fsm_gwlbdis_buf),
     .fsm_nv_bstream_buf(fsm_nv_bstream_buf),
     .fsm_pgmien_buf(fsm_pgmien_buf), .fsm_din_buf(fsm_din_buf),
     .fsm_rd_buf(fsm_rd_buf), .fsm_rowadd_buf(fsm_rowadd_buf[7:0]),
     .fsm_tm_trow_buf(fsm_tm_trow_buf),
     .fsm_sample_buf(fsm_sample_buf),
     .fsm_blkadd_b_buf(fsm_blkadd_b_buf[3:0]),
     .fsm_tm_rd_mode_buf(fsm_tm_rd_mode_buf),
     .fsm_trim_ipp_buf(fsm_trim_ipp_buf[3:0]),
     .fsm_tm_testdec_buf(fsm_tm_testdec_buf),
     .fsm_trim_rrefpgm_buf(fsm_trim_rrefpgm_buf[2:0]),
     .fsm_trim_rrefrd_buf(fsm_trim_rrefred_buf[2:0]),
     .fsm_vpxaset_buf(fsm_vpxaset_buf), .fsm_wpen_buf(fsm_wpen_buf),
     .fsm_ymuxdis_buf(fsm_ymuxdis_buf),
     .tm_allbl_h_buf(tm_allbl_h_buf), .tm_allbl_l_buf(tm_allbl_l_buf),
     .tm_allwl_h_buf(tm_allwl_h_buf), .tm_allwl_l_buf(tm_allwl_l_buf),
     .tm_tcol_buf(tm_tcol_buf), .fsm_blkadd_buf(fsm_blkadd_buf[3:0]),
     .tm_testdec_wr_buf(tm_testdec_wr_buf),
     .fsm_coladd_buf(fsm_coladd_buf[9:0]),
     .fsm_nv_rrow_buf(fsm_nv_rrow_buf),
     .fsm_nv_sisi_ui_buf(fsm_nv_sisi_ui_buf),
     .fsm_nv_rri_trim_buf(fsm_nv_rri_trim_buf),
     .fsm_multibl_read_buf(fsm_multibl_read_buf), .tm_dma(tm_dma),
     .fsm_multibl_read(fsm_multibl_read),
     .fsm_nv_rri_trim(fsm_nv_rri_trim),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_coladd(fsm_coladd[9:0]), .tm_testdec_wr(tm_testdec_wr),
     .fsm_blkadd(fsm_blkadd[3:0]), .tm_tcol(tm_tcol),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_trim_ipp(fsm_trim_ipp[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode), .fsm_blkadd_b(fsm_blkadd_b[3:0]),
     .fsm_sample(fsm_sample), .fsm_tm_trow(fsm_tm_trow),
     .fsm_rst_b(fsm_rst_b), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_rd(fsm_rd), .fsm_din(fsm_din), .fsm_pgmien(fsm_pgmien),
     .fsm_nv_bstream(fsm_nv_bstream), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_pgmhv(fsm_pgmhv), .fsm_wren(fsm_wren),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmvfy_buf(fsm_pgmvfy_buf),
     .fsm_pgm(fsm_pgm), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_wgnden_buf(fsm_wgnden_buf), .fsm_wgnden(fsm_wgnden),
     .fsm_vpgmwl(fsm_vpgmwl[2:0]), .fsm_trim_vbg(fsm_trim_vbg[3:0]),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_nvcmen(fsm_nvcmen),
     .fsm_lshven(fsm_lshven), .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .fsm_lshven_buf(fsm_lshven_buf));
ml_core_bank_1_8f Ibank_1 ( .tm_allbank_sel(tm_allbank_sel),
     .nv_dataout(nv_dataout[8:4]), .fsm_coladd(fsm_coladd[9:0]),
     .fsm_pgmdisc(fsm_pgmdisc), .fsm_din(fsm_din),
     .tm_testdec_wr(tm_testdec_wr), .tm_tcol(tm_tcol), .tm_dma(tm_dma),
     .tm_allwl_l(tm_allwl_l), .tm_allwl_h(tm_allwl_h),
     .tm_allbl_l(tm_allbl_l), .tm_allbl_h(tm_allbl_h),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wren(fsm_wren),
     .fsm_wpen(fsm_wpen), .fsm_wgnden(fsm_wgnden),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_trim_ipp(fsm_trim_ipp[3:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_sample(fsm_sample), .fsm_rst_b(fsm_rst_b), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_pgmhv(fsm_pgmhv), .fsm_pgm(fsm_pgm), .fsm_nvcmen(fsm_nvcmen),
     .fsm_nv_rrow(fsm_nv_rrow), .fsm_gwlbdis(fsm_gwlbdis),
     .fsm_nv_bstream(fsm_nv_bstream),
     .fsm_multibl_read(fsm_multibl_read), .fsm_lshven(fsm_lshven),
     .fsm_blkadd_b(fsm_blkadd_b[3:0]), .fsm_blkadd(fsm_blkadd[3:0]),
     .bgr(bgr), .ngate_25(ngate_25), .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .vblinhi_rde(vblinhi),
     .vblinhi_rdo(vblinhi), .vpp_int(vpp_int), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_rowadd(fsm_rowadd[7:0]),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim));
ml_core_bank_0_8f Ibank_0 ( .tm_allbank_sel(tm_allbank_sel_buf),
     .fsm_gwlbdis(fsm_gwlbdis_buf), .vpp_int(vpp_int),
     .fsm_nvcmen(fsm_nvcmen_buf), .fsm_pgm(fsm_pgm_buf),
     .fsm_pgmien(fsm_pgmien_buf), .fsm_pgmvfy(fsm_pgmvfy_buf),
     .fsm_rd(fsm_rd_buf), .fsm_rowadd(fsm_rowadd_buf[7:0]),
     .fsm_rst_b(fsm_rst_b_buf), .fsm_sample(fsm_sample_buf),
     .fsm_blkadd_b(fsm_blkadd_b_buf[3:0]),
     .fsm_tm_rd_mode(fsm_tm_rd_mode_buf),
     .fsm_tm_testdec(fsm_tm_testdec_buf),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm_buf[2:0]),
     .fsm_trim_rrefrd(fsm_trim_rrefred_buf[2:0]),
     .fsm_vpxaset(fsm_vpxaset_buf), .fsm_wpen(fsm_wpen_buf),
     .fsm_ymuxdis(fsm_ymuxdis_buf), .tm_allbl_h(tm_allbl_h_buf),
     .tm_allbl_l(tm_allbl_l_buf), .tm_allwl_h(tm_allwl_h_buf),
     .tm_allwl_l(tm_allwl_l_buf), .tm_tcol(tm_tcol_buf),
     .fsm_blkadd(fsm_blkadd_buf[3:0]),
     .tm_testdec_wr(tm_testdec_wr_buf),
     .fsm_coladd(fsm_coladd_buf[9:0]), .fsm_nv_rrow(fsm_nv_rrow_buf),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui_buf),
     .fsm_nv_rri_trim(fsm_nv_rri_trim_buf),
     .fsm_lshven(fsm_lshven_buf),
     .fsm_multibl_read(fsm_multibl_read_buf), .tm_dma(tm_dma_buf),
     .sb25sup_25(sb25sup_25), .sbhvsup_hv(sbhvsup_hv),
     .vblinhi_rde(vblinhi), .vblinhi_rdo(vblinhi), .vpxa(vpxa),
     .ysup_25(ysup_25), .fsm_wren(fsm_wren_buf),
     .fsm_pgmhv(fsm_pgmhv_buf), .fsm_nv_bstream(fsm_nv_bstream_buf),
     .fsm_din(fsm_din_buf), .fsm_tm_trow(fsm_tm_trow_buf),
     .fsm_trim_ipp(fsm_trim_ipp_buf[3:0]), .fsm_wgnden(fsm_wgnden_buf),
     .fsm_pgmdisc(fsm_pgmdisc_buf), .ngate_25(ngate_25), .bgr(bgr),
     .nv_dataout(nv_dataout_unbuf[3:0]));
nmoscap_25  C7 ( .MINUS(GND_), .PLUS(vddp_));
ml_vppint_top Ivppint_top ( .vpint_en(vpint_en),
     .fsm_pgmvfy_buf(fsm_pgmvfy_buf), .fsm_nvcmen_buf(fsm_nvcmen_buf),
     .vpp_int(vpp_int), .fsm_wgnden_buf(fsm_wgnden_buf), .bgr(bgr),
     .fsm_tm_xvppint(fsm_tm_xvppint), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_vpgmwl_buf(fsm_vpgmwl_buf[2:0]),
     .fsm_pgmdisc_buf(fsm_pgmdisc_buf), .fsm_pgm_buf(fsm_pgm_buf),
     .fsm_lshven_buf(fsm_lshven_buf));
ml_bgr_top Ibgr_top ( .fsm_trim_vbg_buf(fsm_trim_vbg_buf[3:0]),
     .fsm_nvcmen_buf(fsm_nvcmen_buf), .bgr_int(bgr_int));
ml_vpxa_top Ivpxa_top ( .fsm_pumpen(fsm_pumpen),
     .fsm_vrdwl(fsm_vrdwl[2:0]), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xforce(fsm_tm_xforce), .bgr(bgr), .vpxa_int(vpxa));
ml_hvmux_top Ihvmux_top ( .vpint_en(vpint_en), .fsm_wpen(fsm_wpen_buf),
     .tm_wleqbl(tm_wleqbl), .tm_allbl_l(tm_allbl_l_buf),
     .fsm_wgnden(fsm_wgnden_buf), .fsm_tm_xvpxaint(fsm_tm_xvpxaint),
     .fsm_tm_xvpxa(fsm_tm_xvpxa), .fsm_tm_xvppint(fsm_tm_xvppint),
     .fsm_tm_xvbg(fsm_tm_xvbg), .fsm_tm_xforce(fsm_tm_xforce),
     .fsm_tm_rd_mode(fsm_tm_rd_mode_buf), .fsm_rd(fsm_rd_buf),
     .fsm_pumpen(fsm_pumpen), .fsm_pgmvfy(fsm_pgmvfy_buf),
     .fsm_pgm(fsm_pgm_buf), .fsm_nvcmen(fsm_nvcmen_buf),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui_buf),
     .fsm_nv_rri_trim(fsm_nv_rri_trim_buf),
     .fsm_lshven(fsm_lshven_buf), .bgr(bgr), .bgr_int(bgr_int),
     .ngate_25(ngate_25), .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .vpp(vpp), .vpp_int(vpp_int),
     .vpxa(vpxa), .vpxa_int(vpxa), .ysup_25(ysup_25),
     .vblinhi(vblinhi), .tm_testdec(fsm_tm_testdec_buf));

endmodule
// Library - misc, Cell - nvcm_top, View - schematic
// LAST TIME SAVED: Sep 17 16:05:54 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module nvcm_top ( bp0, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_nv_bstream, fsm_nv_redrow,
     fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmdisc,
     fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_pumpen, fsm_rd, fsm_recall,
     fsm_rowadd, fsm_sample, fsm_tm_allbank_sel, fsm_tm_allbl_h,
     fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l, fsm_tm_dma,
     fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_tcol, fsm_tm_testdec,
     fsm_tm_testdec_wr, fsm_tm_trow, fsm_tm_vwleqbl, fsm_tm_xforce,
     fsm_tm_xvbg, fsm_tm_xvpp, fsm_tm_xvpxa, fsm_tm_xvpxa_int,
     fsm_trim_ipp, fsm_trim_multibl_read, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_trim_vbg, fsm_trim_vpgmwl, fsm_trim_vrdwl,
     fsm_vpxaset, fsm_wgnden, fsm_wpen, fsm_wren, fsm_ymuxdis,
     nvcm_boot, nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b, clk,
     icef_member_sel, nv_dataout, nvcm_ce_b, rst_b,
     smc_load_nvcm_bstream, spi_sdi, spi_ss_b );
output  bp0, fsm_din, fsm_gwlbdis, fsm_lshven, fsm_nv_bstream,
     fsm_nv_redrow, fsm_nv_rri_trim, fsm_nv_sisi_ui, fsm_nvcmen,
     fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy,
     fsm_pumpen, fsm_rd, fsm_recall, fsm_sample, fsm_tm_allbank_sel,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_dma, fsm_tm_margin0_read, fsm_tm_rd_mode, fsm_tm_tcol,
     fsm_tm_testdec, fsm_tm_testdec_wr, fsm_tm_trow, fsm_tm_vwleqbl,
     fsm_tm_xforce, fsm_tm_xvbg, fsm_tm_xvpp, fsm_tm_xvpxa,
     fsm_tm_xvpxa_int, fsm_trim_multibl_read, fsm_vpxaset, fsm_wgnden,
     fsm_wpen, fsm_wren, fsm_ymuxdis, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

output [3:0]  fsm_trim_vbg;
output [8:0]  fsm_rowadd;
output [9:0]  fsm_coladd;
output [2:0]  fsm_trim_vpgmwl;
output [3:0]  fsm_trim_ipp;
output [2:0]  fsm_trim_rrefpgm;
output [2:0]  fsm_trim_rrefrd;
output [3:0]  fsm_blkadd;
output [2:0]  fsm_trim_vrdwl;
output [3:0]  fsm_blkadd_b;

input [1:0]  icef_member_sel;
input [8:0]  nv_dataout;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - misc, Cell - nvcm_ml_block, View - schematic
// LAST TIME SAVED: Sep 17 16:06:07 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module nvcm_ml_block ( bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, spi_sdo, spi_sdo_oe_b, vpp, clk,
     icef_member_sel, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi,
     spi_ss_b );
output  bp0, fsm_recall, fsm_tm_margin0_read, nvcm_boot, nvcm_rdy,
     nvcm_relextspi, spi_sdo, spi_sdo_oe_b;

inout  vpp;

input  clk, nvcm_ce_b, rst_b, smc_load_nvcm_bstream, spi_sdi, spi_ss_b;

input [1:0]  icef_member_sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [8:0]  fsm_rowadd;

wire  [0:2]  net209;

wire  [0:3]  net212;

wire  [0:3]  net249;

wire  [0:8]  net0144;

wire  [0:2]  net207;

wire  [0:2]  net206;

wire  [0:2]  net210;

wire  [0:9]  net0140;

wire  [0:3]  net248;

wire  [0:3]  net208;


/*
ml_chip_nvcm_8f Iml_chip_nvcm ( .tm_allbank_sel(net0145),
     .fsm_coladd(net0140[0:9]), .tm_wleqbl(net217),
     .tm_testdec_wr(net219), .tm_tcol(net221), .tm_dma(net224),
     .tm_allwl_l(net225), .tm_allwl_h(net226), .tm_allbl_l(net227),
     .tm_allbl_h(net228), .fsm_ymuxdis(net200), .fsm_wren(net201),
     .fsm_wpen(net202), .fsm_wgnden(net203), .fsm_vrdwl(net206[0:2]),
     .fsm_vpxaset(net204), .fsm_vpgmwl(net207[0:2]),
     .fsm_trim_vbg(net208[0:3]), .fsm_trim_rrefrd(net209[0:2]),
     .fsm_trim_rrefpgm(net210[0:2]), .fsm_trim_ipp(net212[0:3]),
     .fsm_tm_xvpxaint(net213), .fsm_tm_xvpxa(net214),
     .fsm_tm_xvppint(net272), .fsm_tm_xvbg(net205),
     .fsm_tm_xforce(net216), .fsm_tm_trow(net218),
     .fsm_tm_testdec(net220), .fsm_tm_rd_mode(net222),
     .fsm_sample(net229), .fsm_rst_b(rst_bd),
     .fsm_rowadd(fsm_rowadd[7:0]), .fsm_rd(net232),
     .fsm_pumpen(net233), .fsm_pgmvfy(net234), .fsm_pgmien(net235),
     .fsm_pgmhv(net236), .fsm_pgmdisc(net237), .fsm_pgm(net238),
     .fsm_nvcmen(net239), .fsm_nv_sisi_ui(net240),
     .fsm_nv_rrow(net242), .fsm_nv_rri_trim(net241),
     .fsm_nv_bstream(net243), .fsm_multibl_read(net211),
     .fsm_lshven(net244), .fsm_gwlbdis(net245), .fsm_din(net246),
     .fsm_blkadd_b(net248[0:3]), .fsm_blkadd(net249[0:3]),
     .nv_dataout(net0144[0:8]), .vpp(vpp));
sg_bufx10 I217 ( .in(rst_b), .out(rst_bd));
nvcm_top Invcm_top ( .fsm_tm_allbank_sel(net0145),
     .nvcm_boot(nvcm_boot), .fsm_coladd(net0140[0:9]),
     .spi_ss_b(spi_ss_b), .spi_sdi(spi_sdi),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_ce_b(nvcm_ce_b), .nv_dataout(net0144[0:8]),
     .icef_member_sel(icef_member_sel[1:0]), .clk(clk),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .nvcm_relextspi(nvcm_relextspi), .nvcm_rdy(nvcm_rdy),
     .fsm_ymuxdis(net200), .fsm_wren(net201), .fsm_wpen(net202),
     .fsm_wgnden(net203), .fsm_vpxaset(net204), .fsm_tm_xvbg(net205),
     .fsm_trim_vrdwl(net206[0:2]), .fsm_trim_vpgmwl(net207[0:2]),
     .fsm_trim_vbg(net208[0:3]), .fsm_trim_rrefrd(net209[0:2]),
     .fsm_trim_rrefpgm(net210[0:2]), .fsm_trim_multibl_read(net211),
     .fsm_trim_ipp(net212[0:3]), .fsm_tm_xvpxa_int(net213),
     .fsm_tm_xvpxa(net214), .fsm_tm_xvpp(net272),
     .fsm_tm_xforce(net216), .fsm_tm_vwleqbl(net217),
     .fsm_tm_trow(net218), .fsm_tm_testdec_wr(net219),
     .fsm_tm_testdec(net220), .fsm_tm_tcol(net221),
     .fsm_tm_rd_mode(net222),
     .fsm_tm_margin0_read(fsm_tm_margin0_read), .fsm_tm_dma(net224),
     .fsm_tm_allwl_l(net225), .fsm_tm_allwl_h(net226),
     .fsm_tm_allbl_l(net227), .fsm_tm_allbl_h(net228),
     .fsm_sample(net229), .fsm_rowadd(fsm_rowadd[8:0]),
     .fsm_recall(fsm_recall), .fsm_rd(net232), .fsm_pumpen(net233),
     .fsm_pgmvfy(net234), .fsm_pgmien(net235), .fsm_pgmhv(net236),
     .fsm_pgmdisc(net237), .fsm_pgm(net238), .fsm_nvcmen(net239),
     .fsm_nv_sisi_ui(net240), .fsm_nv_rri_trim(net241),
     .fsm_nv_redrow(net242), .fsm_nv_bstream(net243),
     .fsm_lshven(net244), .fsm_gwlbdis(net245), .fsm_din(net246),
     .fsm_blkadd_b(net248[0:3]), .fsm_blkadd(net249[0:3]), .bp0(bp0));
*/
endmodule
// Library - io, Cell - PMEMIO, View - schematic
// LAST TIME SAVED: Aug 18 15:53:39 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PMEMIO ( C, NET107, PAD, VREF, A2, A6, DS, I, LVCMOS, OEN, PWD,
     S0, S1 );
output  C;

inout  NET107, PAD, VREF;

input  A2, A6, DS, I, LVCMOS, OEN, PWD, S0, S1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PMEMIO_pair_ice8, View - schematic
// LAST TIME SAVED: May 20 13:28:05 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PMEMIO_pair_ice8 ( c_n, c_p, PAD_n, PAD_p, VREFSSTL, cbit, i_n,
     i_p, oen_n, oen_p );
output  c_n, c_p;

inout  PAD_n, PAD_p, VREFSSTL;

input  i_n, i_p, oen_n, oen_p;

input [14:0]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PMEMIO I50 ( .PAD(PAD_p), .VREF(VREFSSTL), .NET107(net107),
     .A6(cbit[8]), .A2(cbit[9]), .DS(cbit[10]), .LVCMOS(cbit[11]),
     .S1(cbit[12]), .S0(cbit[13]), .PWD(cbit[14]), .C(c_p),
     .OEN(oen_p), .I(i_p));
PMEMIO I54 ( .PAD(PAD_n), .VREF(input_), .NET107(net_056),
     .A6(cbit[0]), .A2(cbit[1]), .DS(cbit[2]), .LVCMOS(cbit[3]),
     .S1(cbit[4]), .S0(cbit[5]), .PWD(cbit[6]), .C(c_n), .OEN(oen_n),
     .I(i_n));
LVDS_con I52 ( .VREF(VREFSSTL), .input_(input_), .cbit_7(cbit[7]),
     .Top_Pad_input(net107));

endmodule
// Library - xpmem, Cell - sg_dffbuf_modified, View - schematic
// LAST TIME SAVED: Aug 28 14:33:30 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module sg_dffbuf_modified ( dffout, clk, d, r );
output  dffout;

input  clk, d, r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I2 ( .in(net10), .out(dffout));
ml_dff I0 ( .R(r), .D(d), .CLK(clk), .QN(net9), .Q(net10));

endmodule
// Library - io, Cell - PVSSRSSTL, View - schematic
// LAST TIME SAVED: Sep  4 18:59:25 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVSSRSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVD25SSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:14:18 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVD25SSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDDSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:16:16 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVDDSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDDSSTLE, View - schematic
// LAST TIME SAVED: Jul 28 17:16:16 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVDDSSTLE (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVSSSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:17:35 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVSSSSTL ( VSSC );
input  VSSC;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDDSSTLD, View - schematic
// LAST TIME SAVED: Jul 28 17:15:51 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVDDSSTLD ( VDDD, VDDSSTLD );
input  VDDD, VDDSSTLD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVDDPSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:15:34 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVDDPSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVSSPSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:17:20 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVSSPSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVREFSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:16:31 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVREFSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVSSSSTLD, View - schematic
// LAST TIME SAVED: Jul 28 17:17:58 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVSSSSTLD ( VSSD );
input  VSSD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - misc, Cell - smc_and_jtag_ice8f, View - schematic
// LAST TIME SAVED: Aug  8 16:20:55 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module smc_and_jtag_ice8f ( bm_bank_sdi, bm_banksel, bm_clk, bm_init,
     bm_rcapmux_en, bm_sa, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_banksel, cm_clk, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2, cm_sdi_u3, data_muxsel, data_muxsel1,
     en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0, j_hiz_b,
     j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck, j_tdi,
     j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, psdo, rst_b,
     smc_load_nvcm_bstream, smc_osc_fsel, smc_oscoff_b, smc_podt_off,
     smc_podt_rst, smc_read, smc_row_inc, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rsr_rst, smc_rwl_en, smc_seq_rst,
     smc_wcram_rst, smc_wdis_dclk, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out,
     spi_sdo, spi_sdo_oe_b, spi_ss_out_b, tdo_oe_pad, tdo_pad,
     bm_bank_sdo, boot, bp0, bschain_sdo, cdone_in, cm_last_rsr,
     cm_monitor_cell, cm_sdo_u0, cm_sdo_u1, cm_sdo_u2, cm_sdo_u3,
     cnt_podt_out, coldboot_sel, creset_b, idcode_msb20bits, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     osc_clk, por_b, psdi, spi_clk_in, spi_sdi, spi_ss_in_b, tck_pad,
     tdi_pad, tms_pad, trst_pad, warmboot_sel );
output  bm_clk, bm_init, bm_rcapmux_en, bm_sclkrw, bm_sreb, bm_sweb,
     bm_wdummymux_en, bs_en, cdone_out, cm_clk, data_muxsel,
     data_muxsel1, en_8bconfig_b, end_of_startup, gint_hz, gsr, j_ceb0,
     j_hiz_b, j_mode, j_row_test, j_rst_b, j_sft_dr, j_shift0, j_tck,
     j_tdi, j_upd_dr, md_spi_b, nvcm_spi_sdi, nvcm_spi_ss_b, rst_b,
     smc_load_nvcm_bstream, smc_oscoff_b, smc_podt_off, smc_podt_rst,
     smc_read, smc_row_inc, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rsr_rst, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_wdis_dclk, smc_write, smc_wset_prec, smc_wset_precgnd,
     smc_wwlwrt_dis, smc_wwlwrt_en, spi_clk_out, spi_sdo, spi_sdo_oe_b,
     spi_ss_out_b, tdo_oe_pad, tdo_pad;

input  boot, bp0, bschain_sdo, cdone_in, cm_last_rsr, cnt_podt_out,
     creset_b, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, osc_clk, por_b, spi_clk_in, spi_sdi,
     spi_ss_in_b, tck_pad, tdi_pad, tms_pad, trst_pad;

output [3:0]  bm_bank_sdi;
output [3:0]  bm_banksel;
output [3:0]  cm_banksel;
output [1:0]  cm_sdi_u2;
output [1:0]  cm_sdi_u1;
output [7:1]  psdo;
output [1:0]  smc_osc_fsel;
output [7:0]  bm_sa;
output [1:0]  cm_sdi_u0;
output [1:0]  cm_sdi_u3;

input [3:0]  cm_monitor_cell;
input [1:0]  cm_sdo_u3;
input [1:0]  cm_sdo_u0;
input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdo_u2;
input [1:0]  warmboot_sel;
input [19:0]  idcode_msb20bits;
input [3:0]  bm_bank_sdo;
input [7:1]  psdi;
input [1:0]  coldboot_sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PVD25POCSSTL, View - schematic
// LAST TIME SAVED: Jul 28 17:14:18 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PVD25POCSSTL (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - lefbank_rev, View - schematic
// LAST TIME SAVED: May 20 13:37:32 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module lefbank_rev ( in, VREFSSTL, pad, cbit, oen, out );

inout  VREFSSTL;


output [49:0]  in;

inout [49:0]  pad;

input [374:0]  cbit;
input [49:0]  oen;
input [49:0]  out;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net274;

wire  [0:1]  net273;



PMEMIO_pair_ice8 I46_15_ ( .oen_p(oen[31]), .oen_n(oen[30]),
     .PAD_n(pad[30]), .VREFSSTL(VREFSSTL), .c_p(in[31]), .c_n(in[30]),
     .PAD_p(pad[31]), .i_n(out[30]), .i_p(out[31]),
     .cbit(cbit[239:225]));
PMEMIO_pair_ice8 I46_14_ ( .oen_p(oen[29]), .oen_n(oen[28]),
     .PAD_n(pad[28]), .VREFSSTL(VREFSSTL), .c_p(in[29]), .c_n(in[28]),
     .PAD_p(pad[29]), .i_n(out[28]), .i_p(out[29]),
     .cbit(cbit[224:210]));
PMEMIO_pair_ice8 I46_13_ ( .oen_p(oen[27]), .oen_n(oen[26]),
     .PAD_n(pad[26]), .VREFSSTL(VREFSSTL), .c_p(in[27]), .c_n(in[26]),
     .PAD_p(pad[27]), .i_n(out[26]), .i_p(out[27]),
     .cbit(cbit[209:195]));
PMEMIO_pair_ice8 I47_22_ ( .oen_p(oen[45]), .oen_n(oen[44]),
     .PAD_n(pad[44]), .VREFSSTL(VREFSSTL), .c_p(in[45]), .c_n(in[44]),
     .PAD_p(pad[45]), .i_n(out[44]), .i_p(out[45]),
     .cbit(cbit[344:330]));
PMEMIO_pair_ice8 I47_21_ ( .oen_p(oen[43]), .oen_n(oen[42]),
     .PAD_n(pad[42]), .VREFSSTL(VREFSSTL), .c_p(in[43]), .c_n(in[42]),
     .PAD_p(pad[43]), .i_n(out[42]), .i_p(out[43]),
     .cbit(cbit[329:315]));
PMEMIO_pair_ice8 I48_12_ ( .oen_p(oen[25]), .oen_n(oen[24]),
     .PAD_n(pad[24]), .VREFSSTL(VREFSSTL), .c_p(in[25]), .c_n(in[24]),
     .PAD_p(pad[25]), .i_n(out[24]), .i_p(out[25]),
     .cbit(cbit[194:180]));
PMEMIO_pair_ice8 I49_20_ ( .oen_p(oen[41]), .oen_n(oen[40]),
     .PAD_n(pad[40]), .VREFSSTL(VREFSSTL), .c_p(in[41]), .c_n(in[40]),
     .PAD_p(pad[41]), .i_n(out[40]), .i_p(out[41]),
     .cbit(cbit[314:300]));
PMEMIO_pair_ice8 I49_19_ ( .oen_p(oen[39]), .oen_n(oen[38]),
     .PAD_n(pad[38]), .VREFSSTL(VREFSSTL), .c_p(in[39]), .c_n(in[38]),
     .PAD_p(pad[39]), .i_n(out[38]), .i_p(out[39]),
     .cbit(cbit[299:285]));
PMEMIO_pair_ice8 I50_11_ ( .oen_p(oen[23]), .oen_n(oen[22]),
     .PAD_n(pad[22]), .VREFSSTL(VREFSSTL), .c_p(in[23]), .c_n(in[22]),
     .PAD_p(pad[23]), .i_n(out[22]), .i_p(out[23]),
     .cbit(cbit[179:165]));
PMEMIO_pair_ice8 I50_10_ ( .oen_p(oen[21]), .oen_n(oen[20]),
     .PAD_n(pad[20]), .VREFSSTL(VREFSSTL), .c_p(in[21]), .c_n(in[20]),
     .PAD_p(pad[21]), .i_n(out[20]), .i_p(out[21]),
     .cbit(cbit[164:150]));
PMEMIO_pair_ice8 I50_9_ ( .oen_p(oen[19]), .oen_n(oen[18]),
     .PAD_n(pad[18]), .VREFSSTL(VREFSSTL), .c_p(in[19]), .c_n(in[18]),
     .PAD_p(pad[19]), .i_n(out[18]), .i_p(out[19]),
     .cbit(cbit[149:135]));
PMEMIO_pair_ice8 I51_18_ ( .oen_p(oen[37]), .oen_n(oen[36]),
     .PAD_n(pad[36]), .VREFSSTL(VREFSSTL), .c_p(in[37]), .c_n(in[36]),
     .PAD_p(pad[37]), .i_n(out[36]), .i_p(out[37]),
     .cbit(cbit[284:270]));
PMEMIO_pair_ice8 I53_17_ ( .oen_p(oen[35]), .oen_n(oen[34]),
     .PAD_n(pad[34]), .VREFSSTL(VREFSSTL), .c_p(in[35]), .c_n(in[34]),
     .PAD_p(pad[35]), .i_n(out[34]), .i_p(out[35]),
     .cbit(cbit[269:255]));
PMEMIO_pair_ice8 I54_7_ ( .oen_p(oen[15]), .oen_n(oen[14]),
     .PAD_n(pad[14]), .VREFSSTL(VREFSSTL), .c_p(in[15]), .c_n(in[14]),
     .PAD_p(pad[15]), .i_n(out[14]), .i_p(out[15]),
     .cbit(cbit[119:105]));
PMEMIO_pair_ice8 I54_6_ ( .oen_p(oen[13]), .oen_n(oen[12]),
     .PAD_n(pad[12]), .VREFSSTL(VREFSSTL), .c_p(in[13]), .c_n(in[12]),
     .PAD_p(pad[13]), .i_n(out[12]), .i_p(out[13]),
     .cbit(cbit[104:90]));
PMEMIO_pair_ice8 I54_5_ ( .oen_p(oen[11]), .oen_n(oen[10]),
     .PAD_n(pad[10]), .VREFSSTL(VREFSSTL), .c_p(in[11]), .c_n(in[10]),
     .PAD_p(pad[11]), .i_n(out[10]), .i_p(out[11]),
     .cbit(cbit[89:75]));
PMEMIO_pair_ice8 I54_4_ ( .oen_p(oen[9]), .oen_n(oen[8]),
     .PAD_n(pad[8]), .VREFSSTL(VREFSSTL), .c_p(in[9]), .c_n(in[8]),
     .PAD_p(pad[9]), .i_n(out[8]), .i_p(out[9]), .cbit(cbit[74:60]));
PMEMIO_pair_ice8 I45_24_ ( .oen_p(oen[49]), .oen_n(oen[48]),
     .PAD_n(pad[48]), .VREFSSTL(VREFSSTL), .c_p(in[49]), .c_n(in[48]),
     .PAD_p(pad[49]), .i_n(out[48]), .i_p(out[49]),
     .cbit(cbit[374:360]));
PMEMIO_pair_ice8 I45_23_ ( .oen_p(oen[47]), .oen_n(oen[46]),
     .PAD_n(pad[46]), .VREFSSTL(VREFSSTL), .c_p(in[47]), .c_n(in[46]),
     .PAD_p(pad[47]), .i_n(out[46]), .i_p(out[47]),
     .cbit(cbit[359:345]));
PMEMIO_pair_ice8 I58_16_ ( .oen_p(oen[33]), .oen_n(oen[32]),
     .PAD_n(pad[32]), .VREFSSTL(VREFSSTL), .c_p(in[33]), .c_n(in[32]),
     .PAD_p(pad[33]), .i_n(out[32]), .i_p(out[33]),
     .cbit(cbit[254:240]));
PMEMIO_pair_ice8 I59_2_ ( .oen_p(oen[5]), .oen_n(oen[4]),
     .PAD_n(pad[4]), .VREFSSTL(VREFSSTL), .c_p(in[5]), .c_n(in[4]),
     .PAD_p(pad[5]), .i_n(out[4]), .i_p(out[5]), .cbit(cbit[44:30]));
PMEMIO_pair_ice8 I59_1_ ( .oen_p(oen[3]), .oen_n(oen[2]),
     .PAD_n(pad[2]), .VREFSSTL(VREFSSTL), .c_p(in[3]), .c_n(in[2]),
     .PAD_p(pad[3]), .i_n(out[2]), .i_p(out[3]), .cbit(cbit[29:15]));
PMEMIO_pair_ice8 I59_0_ ( .oen_p(oen[1]), .oen_n(oen[0]),
     .PAD_n(pad[0]), .VREFSSTL(VREFSSTL), .c_p(in[1]), .c_n(in[0]),
     .PAD_p(pad[1]), .i_n(out[0]), .i_p(out[1]), .cbit(cbit[14:0]));
PMEMIO_pair_ice8 I57_3_ ( .oen_p(oen[7]), .oen_n(oen[6]),
     .PAD_n(pad[6]), .VREFSSTL(VREFSSTL), .c_p(in[7]), .c_n(in[6]),
     .PAD_p(pad[7]), .i_n(out[6]), .i_p(out[7]), .cbit(cbit[59:45]));
PMEMIO_pair_ice8 I52_8_ ( .oen_p(oen[17]), .oen_n(oen[16]),
     .PAD_n(pad[16]), .VREFSSTL(VREFSSTL), .c_p(in[17]), .c_n(in[16]),
     .PAD_p(pad[17]), .i_n(out[16]), .i_p(out[17]),
     .cbit(cbit[134:120]));
PVSSRSSTL I83 ( );
PVD25SSTL I32 ( );
PVD25SSTL I81_1_ ( );
PVD25SSTL I81_0_ ( );
PVDDSSTL I72 ( );
PVDDSSTL I68 ( );
PVDDSSTL I62 ( );
PVDDSSTLE I69 ( );
PVSSSSTL I39_1_ ( .VSSC(net274[0]));
PVSSSSTL I39_0_ ( .VSSC(net274[1]));
PVSSSSTL I82_1_ ( .VSSC(net273[0]));
PVSSSSTL I82_0_ ( .VSSC(net273[1]));
PVSSSSTL I79 ( .VSSC(net272));
PVSSSSTL I65 ( .VSSC(net275));
PVDDSSTLD I73 ( .VDDSSTLD(net276), .VDDD(net277));
PVDDSSTLD I63 ( .VDDSSTLD(net280), .VDDD(net281));
PVDDPSSTL I61_1_ ( );
PVDDPSSTL I61_0_ ( );
PVDDPSSTL I77_1_ ( );
PVDDPSSTL I77_0_ ( );
PVDDPSSTL I74_1_ ( );
PVDDPSSTL I74_0_ ( );
PVDDPSSTL I70_1_ ( );
PVDDPSSTL I70_0_ ( );
PVDDPSSTL I67_1_ ( );
PVDDPSSTL I67_0_ ( );
PVSSPSSTL I60_1_ ( );
PVSSPSSTL I60_0_ ( );
PVSSPSSTL I78_1_ ( );
PVSSPSSTL I78_0_ ( );
PVSSPSSTL I75_1_ ( );
PVSSPSSTL I75_0_ ( );
PVSSPSSTL I71_1_ ( );
PVSSPSSTL I71_0_ ( );
PVSSPSSTL I66_1_ ( );
PVSSPSSTL I66_0_ ( );
PVREFSSTL I35_1_ ( );
PVREFSSTL I35_0_ ( );
PVSSSSTLD I76 ( .VSSD(net282));
PVSSSSTLD I64 ( .VSSD(net0277));
PVD25POCSSTL I80 ( );

endmodule
// Library - io, Cell - PDU08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 17:45:09 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PDU08DGZ ( C, PAD, I, OEN );
output  C;

inout  PAD;

input  I, OEN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - botbank, View - schematic
// LAST TIME SAVED: Dec 13 15:20:47 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module botbank ( cdone_int, ctst_b_int, in, done, pad, cdone_out,
     ctst_b, oen, out, ren );
output  cdone_int, ctst_b_int;

inout  done;

input  cdone_out, ctst_b;

output [56:0]  in;

inout [56:0]  pad;

input [56:0]  out;
input [56:0]  oen;
input [56:0]  ren;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDIDGZ I41 ( .PAD(ctst_b), .C(ctst_b_int));
PDU08DGZ I39 ( .PAD(done), .C(cdone_int), .OEN(cdone_out), .I(gnd_));
PDUW08DGZ I46_30_ ( .PAD(pad[30]), .C(in[30]), .OEN(oen[30]),
     .I(out[30]), .REN(ren[30]));
PDUW08DGZ I46_29_ ( .PAD(pad[29]), .C(in[29]), .OEN(oen[29]),
     .I(out[29]), .REN(ren[29]));
PDUW08DGZ I46_28_ ( .PAD(pad[28]), .C(in[28]), .OEN(oen[28]),
     .I(out[28]), .REN(ren[28]));
PDUW08DGZ I38_10_ ( .PAD(pad[10]), .C(in[10]), .OEN(oen[10]),
     .I(out[10]), .REN(ren[10]));
PDUW08DGZ I38_9_ ( .PAD(pad[9]), .C(in[9]), .OEN(oen[9]), .I(out[9]),
     .REN(ren[9]));
PDUW08DGZ I32_46_ ( .PAD(pad[46]), .C(in[46]), .OEN(oen[46]),
     .I(out[46]), .REN(ren[46]));
PDUW08DGZ I32_45_ ( .PAD(pad[45]), .C(in[45]), .OEN(oen[45]),
     .I(out[45]), .REN(ren[45]));
PDUW08DGZ I40_18_ ( .PAD(pad[18]), .C(in[18]), .OEN(oen[18]),
     .I(out[18]), .REN(ren[18]));
PDUW08DGZ I40_17_ ( .PAD(pad[17]), .C(in[17]), .OEN(oen[17]),
     .I(out[17]), .REN(ren[17]));
PDUW08DGZ I40_16_ ( .PAD(pad[16]), .C(in[16]), .OEN(oen[16]),
     .I(out[16]), .REN(ren[16]));
PDUW08DGZ I40_15_ ( .PAD(pad[15]), .C(in[15]), .OEN(oen[15]),
     .I(out[15]), .REN(ren[15]));
PDUW08DGZ I40_14_ ( .PAD(pad[14]), .C(in[14]), .OEN(oen[14]),
     .I(out[14]), .REN(ren[14]));
PDUW08DGZ I40_13_ ( .PAD(pad[13]), .C(in[13]), .OEN(oen[13]),
     .I(out[13]), .REN(ren[13]));
PDUW08DGZ I40_12_ ( .PAD(pad[12]), .C(in[12]), .OEN(oen[12]),
     .I(out[12]), .REN(ren[12]));
PDUW08DGZ I40_11_ ( .PAD(pad[11]), .C(in[11]), .OEN(oen[11]),
     .I(out[11]), .REN(ren[11]));
PDUW08DGZ I60_52_ ( .PAD(pad[52]), .C(in[52]), .OEN(oen[52]),
     .I(out[52]), .REN(ren[52]));
PDUW08DGZ I60_51_ ( .PAD(pad[51]), .C(in[51]), .OEN(oen[51]),
     .I(out[51]), .REN(ren[51]));
PDUW08DGZ I60_50_ ( .PAD(pad[50]), .C(in[50]), .OEN(oen[50]),
     .I(out[50]), .REN(ren[50]));
PDUW08DGZ I60_49_ ( .PAD(pad[49]), .C(in[49]), .OEN(oen[49]),
     .I(out[49]), .REN(ren[49]));
PDUW08DGZ I60_48_ ( .PAD(pad[48]), .C(in[48]), .OEN(oen[48]),
     .I(out[48]), .REN(ren[48]));
PDUW08DGZ I34_47_ ( .PAD(pad[47]), .C(in[47]), .OEN(oen[47]),
     .I(out[47]), .REN(ren[47]));
PDUW08DGZ I30_44_ ( .PAD(pad[44]), .C(in[44]), .OEN(oen[44]),
     .I(out[44]), .REN(ren[44]));
PDUW08DGZ I30_43_ ( .PAD(pad[43]), .C(in[43]), .OEN(oen[43]),
     .I(out[43]), .REN(ren[43]));
PDUW08DGZ I30_42_ ( .PAD(pad[42]), .C(in[42]), .OEN(oen[42]),
     .I(out[42]), .REN(ren[42]));
PDUW08DGZ I30_41_ ( .PAD(pad[41]), .C(in[41]), .OEN(oen[41]),
     .I(out[41]), .REN(ren[41]));
PDUW08DGZ I30_40_ ( .PAD(pad[40]), .C(in[40]), .OEN(oen[40]),
     .I(out[40]), .REN(ren[40]));
PDUW08DGZ I30_39_ ( .PAD(pad[39]), .C(in[39]), .OEN(oen[39]),
     .I(out[39]), .REN(ren[39]));
PDUW08DGZ I30_38_ ( .PAD(pad[38]), .C(in[38]), .OEN(oen[38]),
     .I(out[38]), .REN(ren[38]));
PDUW08DGZ I30_37_ ( .PAD(pad[37]), .C(in[37]), .OEN(oen[37]),
     .I(out[37]), .REN(ren[37]));
PDUW08DGZ I30_36_ ( .PAD(pad[36]), .C(in[36]), .OEN(oen[36]),
     .I(out[36]), .REN(ren[36]));
PDUW08DGZ I30_35_ ( .PAD(pad[35]), .C(in[35]), .OEN(oen[35]),
     .I(out[35]), .REN(ren[35]));
PDUW08DGZ I30_34_ ( .PAD(pad[34]), .C(in[34]), .OEN(oen[34]),
     .I(out[34]), .REN(ren[34]));
PDUW08DGZ I30_33_ ( .PAD(pad[33]), .C(in[33]), .OEN(oen[33]),
     .I(out[33]), .REN(ren[33]));
PDUW08DGZ I30_32_ ( .PAD(pad[32]), .C(in[32]), .OEN(oen[32]),
     .I(out[32]), .REN(ren[32]));
PDUW08DGZ I30_31_ ( .PAD(pad[31]), .C(in[31]), .OEN(oen[31]),
     .I(out[31]), .REN(ren[31]));
PDUW08DGZ I37_8_ ( .PAD(pad[8]), .C(in[8]), .OEN(oen[8]), .I(out[8]),
     .REN(ren[8]));
PDUW08DGZ I37_7_ ( .PAD(pad[7]), .C(in[7]), .OEN(oen[7]), .I(out[7]),
     .REN(ren[7]));
PDUW08DGZ I37_6_ ( .PAD(pad[6]), .C(in[6]), .OEN(oen[6]), .I(out[6]),
     .REN(ren[6]));
PDUW08DGZ I37_5_ ( .PAD(pad[5]), .C(in[5]), .OEN(oen[5]), .I(out[5]),
     .REN(ren[5]));
PDUW08DGZ I37_4_ ( .PAD(pad[4]), .C(in[4]), .OEN(oen[4]), .I(out[4]),
     .REN(ren[4]));
PDUW08DGZ I37_3_ ( .PAD(pad[3]), .C(in[3]), .OEN(oen[3]), .I(out[3]),
     .REN(ren[3]));
PDUW08DGZ I42_20_ ( .PAD(pad[20]), .C(in[20]), .OEN(oen[20]),
     .I(out[20]), .REN(ren[20]));
PDUW08DGZ I42_19_ ( .PAD(pad[19]), .C(in[19]), .OEN(oen[19]),
     .I(out[19]), .REN(ren[19]));
PDUW08DGZ I43_54_ ( .PAD(pad[54]), .C(in[54]), .OEN(oen[54]),
     .I(out[54]), .REN(ren[54]));
PDUW08DGZ I43_53_ ( .PAD(pad[53]), .C(in[53]), .OEN(oen[53]),
     .I(out[53]), .REN(ren[53]));
PDUW08DGZ I44_27_ ( .PAD(pad[27]), .C(in[27]), .OEN(oen[27]),
     .I(out[27]), .REN(ren[27]));
PDUW08DGZ I44_26_ ( .PAD(pad[26]), .C(in[26]), .OEN(oen[26]),
     .I(out[26]), .REN(ren[26]));
PDUW08DGZ I44_25_ ( .PAD(pad[25]), .C(in[25]), .OEN(oen[25]),
     .I(out[25]), .REN(ren[25]));
PDUW08DGZ I44_24_ ( .PAD(pad[24]), .C(in[24]), .OEN(oen[24]),
     .I(out[24]), .REN(ren[24]));
PDUW08DGZ I44_23_ ( .PAD(pad[23]), .C(in[23]), .OEN(oen[23]),
     .I(out[23]), .REN(ren[23]));
PDUW08DGZ I44_22_ ( .PAD(pad[22]), .C(in[22]), .OEN(oen[22]),
     .I(out[22]), .REN(ren[22]));
PDUW08DGZ I44_21_ ( .PAD(pad[21]), .C(in[21]), .OEN(oen[21]),
     .I(out[21]), .REN(ren[21]));
PDUW08DGZ I36_2_ ( .PAD(pad[2]), .C(in[2]), .OEN(oen[2]), .I(out[2]),
     .REN(ren[2]));
PDUW08DGZ I36_1_ ( .PAD(pad[1]), .C(in[1]), .OEN(oen[1]), .I(out[1]),
     .REN(ren[1]));
PDUW08DGZ I36_0_ ( .PAD(pad[0]), .C(in[0]), .OEN(oen[0]), .I(out[0]),
     .REN(ren[0]));
PDUW08DGZ I45_56_ ( .PAD(pad[56]), .C(in[56]), .OEN(oen[56]),
     .I(out[56]), .REN(ren[56]));
PDUW08DGZ I45_55_ ( .PAD(pad[55]), .C(in[55]), .OEN(oen[55]),
     .I(out[55]), .REN(ren[55]));
PVDD1DGZ I58_1_ ( .VDD(vdd_));
PVDD1DGZ I58_0_ ( .VDD(vdd_));
PVDD1DGZ I50_1_ ( .VDD(vdd_));
PVDD1DGZ I50_0_ ( .VDD(vdd_));
PVDD1DGZ I52_1_ ( .VDD(vdd_));
PVDD1DGZ I52_0_ ( .VDD(vdd_));
PVDD2DGZ I56 ( .VDDPST(vddio_spi));
PVDD2DGZ I48_1_ ( .VDDPST(vddio_bottombank));
PVDD2DGZ I48_0_ ( .VDDPST(vddio_bottombank));
PVDD2DGZ I54 ( .VDDPST(vddio_bottombank));
PVDD2DGZ I61_1_ ( .VDDPST(vddio_bottombank));
PVDD2DGZ I61_0_ ( .VDDPST(vddio_bottombank));
PVDD2POC I57 ( .VDDPST(vddio_spi));
PVDD2POC I53 ( .VDDPST(vddio_bottombank));
PVSS3DGZ I37_1_ ( .VSS(gnd_));
PVSS3DGZ I37_0_ ( .VSS(gnd_));
PVSS3DGZ I47_1_ ( .VSS(gnd_));
PVSS3DGZ I47_0_ ( .VSS(gnd_));
PVSS3DGZ I55_1_ ( .VSS(gnd_));
PVSS3DGZ I55_0_ ( .VSS(gnd_));
PVSS3DGZ I59_1_ ( .VSS(gnd_));
PVSS3DGZ I59_0_ ( .VSS(gnd_));
PVSS3DGZ I49_1_ ( .VSS(gnd_));
PVSS3DGZ I49_0_ ( .VSS(gnd_));
PVSS3DGZ I51_1_ ( .VSS(gnd_));
PVSS3DGZ I51_0_ ( .VSS(gnd_));

endmodule
// Library - chip, Cell - CHIP_route_left10k, View - schematic
// LAST TIME SAVED: Oct  7 17:53:09 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module CHIP_route_left10k ( cm_banksel_bltld3_1_, cm_clk_bltld3,
     cm_sdi_u1d3[1:0], cm_sdo_u1d1[1:0], core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, last_rsr[1:0],
     monitor_celld2[1:0], pgate_l[543:0], reset_l[543:0],
     smc_wdis_dclk_bltld3, vdd_cntl_l[543:0], wl_l[543:0],
     cf_lbank[300], cf_lbank[479], cm_banksel_blbld1[0],
     cm_banksel_blbld[1], cm_clk_blbld, cm_sdi_u1d[1:0],
     cm_sdo_u1[1:0], core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0 );
output  cm_banksel_bltld3_1_, cm_clk_bltld3, core_por_b_rowu0,
     core_por_b_rowu1, cram_prec_bltld3, cram_pullup_bltld3,
     cram_write_bltld3, data_muxsel1_bltld3, data_muxsel_bltld3,
     en_8bconfig_b_bltld3, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, last_rsr0, smc_wdis_dclk_bltld3;

input  cm_clk_blbld, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0;

output [1:0]  cm_sdo_u1d1;
output [1:0]  last_rsr;
output [543:0]  reset_l;
output [1:0]  monitor_celld2;
output [543:0]  wl_l;
output [1:0]  cm_sdi_u1d3;
output [543:0]  vdd_cntl_l;
output [543:0]  pgate_l;

input [1:1]  cm_banksel_blbld;
input [1:0]  cm_sdo_u1;
input [1:0]  cm_sdi_u1d;
input [0:0]  cm_banksel_blbld1;
input [300:479]  cf_lbank;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u1d;

wire  [1:0]  cm_sdi_u1d0;

wire  [1:1]  monitor_celld;

wire  [0:1]  net081;

wire  [1:1]  cm_banksel_bltld;

wire  [1:1]  monitor_celld1;

wire  [1:0]  cm_sdo_u1d0;

wire  [1:0]  dff_out;



tielo I451_1_ ( .tielo(net081[0]));
tielo I451_0_ ( .tielo(net081[1]));
tielo I452 ( .tielo(net080));
sg_dffbuf_modified I261_1_ ( .r(net081[0]), .dffout(dff_out[1]),
     .d(cm_sdo_u1d[1]), .clk(net148));
sg_dffbuf_modified I261_0_ ( .r(net081[1]), .dffout(dff_out[0]),
     .d(cm_sdo_u1d[0]), .clk(net148));
sg_dffbuf_modified I289 ( .r(net080), .d(last_rsr[0]), .clk(net146),
     .dffout(last_rsr0));
ml_rowdrv_bank10k Irowul ( .vddctrl({vdd_cntl_l[272], vdd_cntl_l[273],
     vdd_cntl_l[274], vdd_cntl_l[275], vdd_cntl_l[276],
     vdd_cntl_l[277], vdd_cntl_l[278], vdd_cntl_l[279],
     vdd_cntl_l[280], vdd_cntl_l[281], vdd_cntl_l[282],
     vdd_cntl_l[283], vdd_cntl_l[284], vdd_cntl_l[285],
     vdd_cntl_l[286], vdd_cntl_l[287], vdd_cntl_l[288],
     vdd_cntl_l[289], vdd_cntl_l[290], vdd_cntl_l[291],
     vdd_cntl_l[292], vdd_cntl_l[293], vdd_cntl_l[294],
     vdd_cntl_l[295], vdd_cntl_l[296], vdd_cntl_l[297],
     vdd_cntl_l[298], vdd_cntl_l[299], vdd_cntl_l[300],
     vdd_cntl_l[301], vdd_cntl_l[302], vdd_cntl_l[303],
     vdd_cntl_l[304], vdd_cntl_l[305], vdd_cntl_l[306],
     vdd_cntl_l[307], vdd_cntl_l[308], vdd_cntl_l[309],
     vdd_cntl_l[310], vdd_cntl_l[311], vdd_cntl_l[312],
     vdd_cntl_l[313], vdd_cntl_l[314], vdd_cntl_l[315],
     vdd_cntl_l[316], vdd_cntl_l[317], vdd_cntl_l[318],
     vdd_cntl_l[319], vdd_cntl_l[320], vdd_cntl_l[321],
     vdd_cntl_l[322], vdd_cntl_l[323], vdd_cntl_l[324],
     vdd_cntl_l[325], vdd_cntl_l[326], vdd_cntl_l[327],
     vdd_cntl_l[328], vdd_cntl_l[329], vdd_cntl_l[330],
     vdd_cntl_l[331], vdd_cntl_l[332], vdd_cntl_l[333],
     vdd_cntl_l[334], vdd_cntl_l[335], vdd_cntl_l[336],
     vdd_cntl_l[337], vdd_cntl_l[338], vdd_cntl_l[339],
     vdd_cntl_l[340], vdd_cntl_l[341], vdd_cntl_l[342],
     vdd_cntl_l[343], vdd_cntl_l[344], vdd_cntl_l[345],
     vdd_cntl_l[346], vdd_cntl_l[347], vdd_cntl_l[348],
     vdd_cntl_l[349], vdd_cntl_l[350], vdd_cntl_l[351],
     vdd_cntl_l[352], vdd_cntl_l[353], vdd_cntl_l[354],
     vdd_cntl_l[355], vdd_cntl_l[356], vdd_cntl_l[357],
     vdd_cntl_l[358], vdd_cntl_l[359], vdd_cntl_l[360],
     vdd_cntl_l[361], vdd_cntl_l[362], vdd_cntl_l[363],
     vdd_cntl_l[364], vdd_cntl_l[365], vdd_cntl_l[366],
     vdd_cntl_l[367], vdd_cntl_l[368], vdd_cntl_l[369],
     vdd_cntl_l[370], vdd_cntl_l[371], vdd_cntl_l[372],
     vdd_cntl_l[373], vdd_cntl_l[374], vdd_cntl_l[375],
     vdd_cntl_l[376], vdd_cntl_l[377], vdd_cntl_l[378],
     vdd_cntl_l[379], vdd_cntl_l[380], vdd_cntl_l[381],
     vdd_cntl_l[382], vdd_cntl_l[383], vdd_cntl_l[384],
     vdd_cntl_l[385], vdd_cntl_l[386], vdd_cntl_l[387],
     vdd_cntl_l[388], vdd_cntl_l[389], vdd_cntl_l[390],
     vdd_cntl_l[391], vdd_cntl_l[392], vdd_cntl_l[393],
     vdd_cntl_l[394], vdd_cntl_l[395], vdd_cntl_l[396],
     vdd_cntl_l[397], vdd_cntl_l[398], vdd_cntl_l[399],
     vdd_cntl_l[400], vdd_cntl_l[401], vdd_cntl_l[402],
     vdd_cntl_l[403], vdd_cntl_l[404], vdd_cntl_l[405],
     vdd_cntl_l[406], vdd_cntl_l[407], vdd_cntl_l[408],
     vdd_cntl_l[409], vdd_cntl_l[410], vdd_cntl_l[411],
     vdd_cntl_l[412], vdd_cntl_l[413], vdd_cntl_l[414],
     vdd_cntl_l[415], vdd_cntl_l[416], vdd_cntl_l[417],
     vdd_cntl_l[418], vdd_cntl_l[419], vdd_cntl_l[420],
     vdd_cntl_l[421], vdd_cntl_l[422], vdd_cntl_l[423],
     vdd_cntl_l[424], vdd_cntl_l[425], vdd_cntl_l[426],
     vdd_cntl_l[427], vdd_cntl_l[428], vdd_cntl_l[429],
     vdd_cntl_l[430], vdd_cntl_l[431], vdd_cntl_l[432],
     vdd_cntl_l[433], vdd_cntl_l[434], vdd_cntl_l[435],
     vdd_cntl_l[436], vdd_cntl_l[437], vdd_cntl_l[438],
     vdd_cntl_l[439], vdd_cntl_l[440], vdd_cntl_l[441],
     vdd_cntl_l[442], vdd_cntl_l[443], vdd_cntl_l[444],
     vdd_cntl_l[445], vdd_cntl_l[446], vdd_cntl_l[447],
     vdd_cntl_l[448], vdd_cntl_l[449], vdd_cntl_l[450],
     vdd_cntl_l[451], vdd_cntl_l[452], vdd_cntl_l[453],
     vdd_cntl_l[454], vdd_cntl_l[455], vdd_cntl_l[456],
     vdd_cntl_l[457], vdd_cntl_l[458], vdd_cntl_l[459],
     vdd_cntl_l[460], vdd_cntl_l[461], vdd_cntl_l[462],
     vdd_cntl_l[463], vdd_cntl_l[464], vdd_cntl_l[465],
     vdd_cntl_l[466], vdd_cntl_l[467], vdd_cntl_l[468],
     vdd_cntl_l[469], vdd_cntl_l[470], vdd_cntl_l[471],
     vdd_cntl_l[472], vdd_cntl_l[473], vdd_cntl_l[474],
     vdd_cntl_l[475], vdd_cntl_l[476], vdd_cntl_l[477],
     vdd_cntl_l[478], vdd_cntl_l[479], vdd_cntl_l[480],
     vdd_cntl_l[481], vdd_cntl_l[482], vdd_cntl_l[483],
     vdd_cntl_l[484], vdd_cntl_l[485], vdd_cntl_l[486],
     vdd_cntl_l[487], vdd_cntl_l[488], vdd_cntl_l[489],
     vdd_cntl_l[490], vdd_cntl_l[491], vdd_cntl_l[492],
     vdd_cntl_l[493], vdd_cntl_l[494], vdd_cntl_l[495],
     vdd_cntl_l[496], vdd_cntl_l[497], vdd_cntl_l[498],
     vdd_cntl_l[499], vdd_cntl_l[500], vdd_cntl_l[501],
     vdd_cntl_l[502], vdd_cntl_l[503], vdd_cntl_l[504],
     vdd_cntl_l[505], vdd_cntl_l[506], vdd_cntl_l[507],
     vdd_cntl_l[508], vdd_cntl_l[509], vdd_cntl_l[510],
     vdd_cntl_l[511], vdd_cntl_l[512], vdd_cntl_l[513],
     vdd_cntl_l[514], vdd_cntl_l[515], vdd_cntl_l[516],
     vdd_cntl_l[517], vdd_cntl_l[518], vdd_cntl_l[519],
     vdd_cntl_l[520], vdd_cntl_l[521], vdd_cntl_l[522],
     vdd_cntl_l[523], vdd_cntl_l[524], vdd_cntl_l[525],
     vdd_cntl_l[526], vdd_cntl_l[527], vdd_cntl_l[528],
     vdd_cntl_l[529], vdd_cntl_l[530], vdd_cntl_l[531],
     vdd_cntl_l[532], vdd_cntl_l[533], vdd_cntl_l[534],
     vdd_cntl_l[535], vdd_cntl_l[536], vdd_cntl_l[537],
     vdd_cntl_l[538], vdd_cntl_l[539], vdd_cntl_l[540],
     vdd_cntl_l[541], vdd_cntl_l[542], vdd_cntl_l[543]}),
     .pgate({pgate_l[272], pgate_l[273], pgate_l[274], pgate_l[275],
     pgate_l[276], pgate_l[277], pgate_l[278], pgate_l[279],
     pgate_l[280], pgate_l[281], pgate_l[282], pgate_l[283],
     pgate_l[284], pgate_l[285], pgate_l[286], pgate_l[287],
     pgate_l[288], pgate_l[289], pgate_l[290], pgate_l[291],
     pgate_l[292], pgate_l[293], pgate_l[294], pgate_l[295],
     pgate_l[296], pgate_l[297], pgate_l[298], pgate_l[299],
     pgate_l[300], pgate_l[301], pgate_l[302], pgate_l[303],
     pgate_l[304], pgate_l[305], pgate_l[306], pgate_l[307],
     pgate_l[308], pgate_l[309], pgate_l[310], pgate_l[311],
     pgate_l[312], pgate_l[313], pgate_l[314], pgate_l[315],
     pgate_l[316], pgate_l[317], pgate_l[318], pgate_l[319],
     pgate_l[320], pgate_l[321], pgate_l[322], pgate_l[323],
     pgate_l[324], pgate_l[325], pgate_l[326], pgate_l[327],
     pgate_l[328], pgate_l[329], pgate_l[330], pgate_l[331],
     pgate_l[332], pgate_l[333], pgate_l[334], pgate_l[335],
     pgate_l[336], pgate_l[337], pgate_l[338], pgate_l[339],
     pgate_l[340], pgate_l[341], pgate_l[342], pgate_l[343],
     pgate_l[344], pgate_l[345], pgate_l[346], pgate_l[347],
     pgate_l[348], pgate_l[349], pgate_l[350], pgate_l[351],
     pgate_l[352], pgate_l[353], pgate_l[354], pgate_l[355],
     pgate_l[356], pgate_l[357], pgate_l[358], pgate_l[359],
     pgate_l[360], pgate_l[361], pgate_l[362], pgate_l[363],
     pgate_l[364], pgate_l[365], pgate_l[366], pgate_l[367],
     pgate_l[368], pgate_l[369], pgate_l[370], pgate_l[371],
     pgate_l[372], pgate_l[373], pgate_l[374], pgate_l[375],
     pgate_l[376], pgate_l[377], pgate_l[378], pgate_l[379],
     pgate_l[380], pgate_l[381], pgate_l[382], pgate_l[383],
     pgate_l[384], pgate_l[385], pgate_l[386], pgate_l[387],
     pgate_l[388], pgate_l[389], pgate_l[390], pgate_l[391],
     pgate_l[392], pgate_l[393], pgate_l[394], pgate_l[395],
     pgate_l[396], pgate_l[397], pgate_l[398], pgate_l[399],
     pgate_l[400], pgate_l[401], pgate_l[402], pgate_l[403],
     pgate_l[404], pgate_l[405], pgate_l[406], pgate_l[407],
     pgate_l[408], pgate_l[409], pgate_l[410], pgate_l[411],
     pgate_l[412], pgate_l[413], pgate_l[414], pgate_l[415],
     pgate_l[416], pgate_l[417], pgate_l[418], pgate_l[419],
     pgate_l[420], pgate_l[421], pgate_l[422], pgate_l[423],
     pgate_l[424], pgate_l[425], pgate_l[426], pgate_l[427],
     pgate_l[428], pgate_l[429], pgate_l[430], pgate_l[431],
     pgate_l[432], pgate_l[433], pgate_l[434], pgate_l[435],
     pgate_l[436], pgate_l[437], pgate_l[438], pgate_l[439],
     pgate_l[440], pgate_l[441], pgate_l[442], pgate_l[443],
     pgate_l[444], pgate_l[445], pgate_l[446], pgate_l[447],
     pgate_l[448], pgate_l[449], pgate_l[450], pgate_l[451],
     pgate_l[452], pgate_l[453], pgate_l[454], pgate_l[455],
     pgate_l[456], pgate_l[457], pgate_l[458], pgate_l[459],
     pgate_l[460], pgate_l[461], pgate_l[462], pgate_l[463],
     pgate_l[464], pgate_l[465], pgate_l[466], pgate_l[467],
     pgate_l[468], pgate_l[469], pgate_l[470], pgate_l[471],
     pgate_l[472], pgate_l[473], pgate_l[474], pgate_l[475],
     pgate_l[476], pgate_l[477], pgate_l[478], pgate_l[479],
     pgate_l[480], pgate_l[481], pgate_l[482], pgate_l[483],
     pgate_l[484], pgate_l[485], pgate_l[486], pgate_l[487],
     pgate_l[488], pgate_l[489], pgate_l[490], pgate_l[491],
     pgate_l[492], pgate_l[493], pgate_l[494], pgate_l[495],
     pgate_l[496], pgate_l[497], pgate_l[498], pgate_l[499],
     pgate_l[500], pgate_l[501], pgate_l[502], pgate_l[503],
     pgate_l[504], pgate_l[505], pgate_l[506], pgate_l[507],
     pgate_l[508], pgate_l[509], pgate_l[510], pgate_l[511],
     pgate_l[512], pgate_l[513], pgate_l[514], pgate_l[515],
     pgate_l[516], pgate_l[517], pgate_l[518], pgate_l[519],
     pgate_l[520], pgate_l[521], pgate_l[522], pgate_l[523],
     pgate_l[524], pgate_l[525], pgate_l[526], pgate_l[527],
     pgate_l[528], pgate_l[529], pgate_l[530], pgate_l[531],
     pgate_l[532], pgate_l[533], pgate_l[534], pgate_l[535],
     pgate_l[536], pgate_l[537], pgate_l[538], pgate_l[539],
     pgate_l[540], pgate_l[541], pgate_l[542], pgate_l[543]}),
     .reset({reset_l[272], reset_l[273], reset_l[274], reset_l[275],
     reset_l[276], reset_l[277], reset_l[278], reset_l[279],
     reset_l[280], reset_l[281], reset_l[282], reset_l[283],
     reset_l[284], reset_l[285], reset_l[286], reset_l[287],
     reset_l[288], reset_l[289], reset_l[290], reset_l[291],
     reset_l[292], reset_l[293], reset_l[294], reset_l[295],
     reset_l[296], reset_l[297], reset_l[298], reset_l[299],
     reset_l[300], reset_l[301], reset_l[302], reset_l[303],
     reset_l[304], reset_l[305], reset_l[306], reset_l[307],
     reset_l[308], reset_l[309], reset_l[310], reset_l[311],
     reset_l[312], reset_l[313], reset_l[314], reset_l[315],
     reset_l[316], reset_l[317], reset_l[318], reset_l[319],
     reset_l[320], reset_l[321], reset_l[322], reset_l[323],
     reset_l[324], reset_l[325], reset_l[326], reset_l[327],
     reset_l[328], reset_l[329], reset_l[330], reset_l[331],
     reset_l[332], reset_l[333], reset_l[334], reset_l[335],
     reset_l[336], reset_l[337], reset_l[338], reset_l[339],
     reset_l[340], reset_l[341], reset_l[342], reset_l[343],
     reset_l[344], reset_l[345], reset_l[346], reset_l[347],
     reset_l[348], reset_l[349], reset_l[350], reset_l[351],
     reset_l[352], reset_l[353], reset_l[354], reset_l[355],
     reset_l[356], reset_l[357], reset_l[358], reset_l[359],
     reset_l[360], reset_l[361], reset_l[362], reset_l[363],
     reset_l[364], reset_l[365], reset_l[366], reset_l[367],
     reset_l[368], reset_l[369], reset_l[370], reset_l[371],
     reset_l[372], reset_l[373], reset_l[374], reset_l[375],
     reset_l[376], reset_l[377], reset_l[378], reset_l[379],
     reset_l[380], reset_l[381], reset_l[382], reset_l[383],
     reset_l[384], reset_l[385], reset_l[386], reset_l[387],
     reset_l[388], reset_l[389], reset_l[390], reset_l[391],
     reset_l[392], reset_l[393], reset_l[394], reset_l[395],
     reset_l[396], reset_l[397], reset_l[398], reset_l[399],
     reset_l[400], reset_l[401], reset_l[402], reset_l[403],
     reset_l[404], reset_l[405], reset_l[406], reset_l[407],
     reset_l[408], reset_l[409], reset_l[410], reset_l[411],
     reset_l[412], reset_l[413], reset_l[414], reset_l[415],
     reset_l[416], reset_l[417], reset_l[418], reset_l[419],
     reset_l[420], reset_l[421], reset_l[422], reset_l[423],
     reset_l[424], reset_l[425], reset_l[426], reset_l[427],
     reset_l[428], reset_l[429], reset_l[430], reset_l[431],
     reset_l[432], reset_l[433], reset_l[434], reset_l[435],
     reset_l[436], reset_l[437], reset_l[438], reset_l[439],
     reset_l[440], reset_l[441], reset_l[442], reset_l[443],
     reset_l[444], reset_l[445], reset_l[446], reset_l[447],
     reset_l[448], reset_l[449], reset_l[450], reset_l[451],
     reset_l[452], reset_l[453], reset_l[454], reset_l[455],
     reset_l[456], reset_l[457], reset_l[458], reset_l[459],
     reset_l[460], reset_l[461], reset_l[462], reset_l[463],
     reset_l[464], reset_l[465], reset_l[466], reset_l[467],
     reset_l[468], reset_l[469], reset_l[470], reset_l[471],
     reset_l[472], reset_l[473], reset_l[474], reset_l[475],
     reset_l[476], reset_l[477], reset_l[478], reset_l[479],
     reset_l[480], reset_l[481], reset_l[482], reset_l[483],
     reset_l[484], reset_l[485], reset_l[486], reset_l[487],
     reset_l[488], reset_l[489], reset_l[490], reset_l[491],
     reset_l[492], reset_l[493], reset_l[494], reset_l[495],
     reset_l[496], reset_l[497], reset_l[498], reset_l[499],
     reset_l[500], reset_l[501], reset_l[502], reset_l[503],
     reset_l[504], reset_l[505], reset_l[506], reset_l[507],
     reset_l[508], reset_l[509], reset_l[510], reset_l[511],
     reset_l[512], reset_l[513], reset_l[514], reset_l[515],
     reset_l[516], reset_l[517], reset_l[518], reset_l[519],
     reset_l[520], reset_l[521], reset_l[522], reset_l[523],
     reset_l[524], reset_l[525], reset_l[526], reset_l[527],
     reset_l[528], reset_l[529], reset_l[530], reset_l[531],
     reset_l[532], reset_l[533], reset_l[534], reset_l[535],
     reset_l[536], reset_l[537], reset_l[538], reset_l[539],
     reset_l[540], reset_l[541], reset_l[542], reset_l[543]}),
     .wl({wl_l[272], wl_l[273], wl_l[274], wl_l[275], wl_l[276],
     wl_l[277], wl_l[278], wl_l[279], wl_l[280], wl_l[281], wl_l[282],
     wl_l[283], wl_l[284], wl_l[285], wl_l[286], wl_l[287], wl_l[288],
     wl_l[289], wl_l[290], wl_l[291], wl_l[292], wl_l[293], wl_l[294],
     wl_l[295], wl_l[296], wl_l[297], wl_l[298], wl_l[299], wl_l[300],
     wl_l[301], wl_l[302], wl_l[303], wl_l[304], wl_l[305], wl_l[306],
     wl_l[307], wl_l[308], wl_l[309], wl_l[310], wl_l[311], wl_l[312],
     wl_l[313], wl_l[314], wl_l[315], wl_l[316], wl_l[317], wl_l[318],
     wl_l[319], wl_l[320], wl_l[321], wl_l[322], wl_l[323], wl_l[324],
     wl_l[325], wl_l[326], wl_l[327], wl_l[328], wl_l[329], wl_l[330],
     wl_l[331], wl_l[332], wl_l[333], wl_l[334], wl_l[335], wl_l[336],
     wl_l[337], wl_l[338], wl_l[339], wl_l[340], wl_l[341], wl_l[342],
     wl_l[343], wl_l[344], wl_l[345], wl_l[346], wl_l[347], wl_l[348],
     wl_l[349], wl_l[350], wl_l[351], wl_l[352], wl_l[353], wl_l[354],
     wl_l[355], wl_l[356], wl_l[357], wl_l[358], wl_l[359], wl_l[360],
     wl_l[361], wl_l[362], wl_l[363], wl_l[364], wl_l[365], wl_l[366],
     wl_l[367], wl_l[368], wl_l[369], wl_l[370], wl_l[371], wl_l[372],
     wl_l[373], wl_l[374], wl_l[375], wl_l[376], wl_l[377], wl_l[378],
     wl_l[379], wl_l[380], wl_l[381], wl_l[382], wl_l[383], wl_l[384],
     wl_l[385], wl_l[386], wl_l[387], wl_l[388], wl_l[389], wl_l[390],
     wl_l[391], wl_l[392], wl_l[393], wl_l[394], wl_l[395], wl_l[396],
     wl_l[397], wl_l[398], wl_l[399], wl_l[400], wl_l[401], wl_l[402],
     wl_l[403], wl_l[404], wl_l[405], wl_l[406], wl_l[407], wl_l[408],
     wl_l[409], wl_l[410], wl_l[411], wl_l[412], wl_l[413], wl_l[414],
     wl_l[415], wl_l[416], wl_l[417], wl_l[418], wl_l[419], wl_l[420],
     wl_l[421], wl_l[422], wl_l[423], wl_l[424], wl_l[425], wl_l[426],
     wl_l[427], wl_l[428], wl_l[429], wl_l[430], wl_l[431], wl_l[432],
     wl_l[433], wl_l[434], wl_l[435], wl_l[436], wl_l[437], wl_l[438],
     wl_l[439], wl_l[440], wl_l[441], wl_l[442], wl_l[443], wl_l[444],
     wl_l[445], wl_l[446], wl_l[447], wl_l[448], wl_l[449], wl_l[450],
     wl_l[451], wl_l[452], wl_l[453], wl_l[454], wl_l[455], wl_l[456],
     wl_l[457], wl_l[458], wl_l[459], wl_l[460], wl_l[461], wl_l[462],
     wl_l[463], wl_l[464], wl_l[465], wl_l[466], wl_l[467], wl_l[468],
     wl_l[469], wl_l[470], wl_l[471], wl_l[472], wl_l[473], wl_l[474],
     wl_l[475], wl_l[476], wl_l[477], wl_l[478], wl_l[479], wl_l[480],
     wl_l[481], wl_l[482], wl_l[483], wl_l[484], wl_l[485], wl_l[486],
     wl_l[487], wl_l[488], wl_l[489], wl_l[490], wl_l[491], wl_l[492],
     wl_l[493], wl_l[494], wl_l[495], wl_l[496], wl_l[497], wl_l[498],
     wl_l[499], wl_l[500], wl_l[501], wl_l[502], wl_l[503], wl_l[504],
     wl_l[505], wl_l[506], wl_l[507], wl_l[508], wl_l[509], wl_l[510],
     wl_l[511], wl_l[512], wl_l[513], wl_l[514], wl_l[515], wl_l[516],
     wl_l[517], wl_l[518], wl_l[519], wl_l[520], wl_l[521], wl_l[522],
     wl_l[523], wl_l[524], wl_l[525], wl_l[526], wl_l[527], wl_l[528],
     wl_l[529], wl_l[530], wl_l[531], wl_l[532], wl_l[533], wl_l[534],
     wl_l[535], wl_l[536], wl_l[537], wl_l[538], wl_l[539], wl_l[540],
     wl_l[541], wl_l[542], wl_l[543]}),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu1_b),
     .smc_write(smc_write_rowu1), .smc_rsr_inc(smc_row_inc_rowu1),
     .rsr_rst(smc_rsr_rst_rowu1), .por_rst(core_por_b_rowu1),
     .cram_wl_en(cram_wl_en_rowu1), .cram_vddoff(cram_vddoff_rowu1),
     .cram_rst(cram_rst_rowu1), .cram_pgateoff(cram_pgateoff_rowu1),
     .banksel(cm_banksel_bltld3_1_), .last_rsr(last_rsr[1]),
     .trst_b(trst_rowu1), .jtag_rowtest_rst(row_test_rowu1),
     .jtag_clk(tck_pad_rowu1));
ml_rowdrv_bank10k Irowbl ( .vddctrl(vdd_cntl_l[271:0]),
     .pgate(pgate_l[271:0]), .reset(reset_l[271:0]), .wl(wl_l[271:0]),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu0_b),
     .smc_write(smc_write_rowu0), .smc_rsr_inc(smc_row_inc_rowu0),
     .rsr_rst(smc_rsr_rst_rowu0), .por_rst(core_por_b_rowu0),
     .cram_wl_en(cram_wl_en_rowu0), .cram_vddoff(cram_vddoff_rowu0),
     .cram_rst(cram_rst_rowu0), .cram_pgateoff(cram_pgateoff_rowu0),
     .banksel(cm_banksel_blbld1[0]), .last_rsr(last_rsr[0]),
     .trst_b(trst_rowu0), .jtag_rowtest_rst(row_test_rowu0),
     .jtag_clk(tck_pad_rowu0));
bram_bufferx16 I381 ( .in(j_rst_bl1), .out(trst_rowu0));
bram_bufferx16 I391 ( .in(j_rst_bl2), .out(trst_rowu1));
bram_bufferx16 I392 ( .in(row_testl3), .out(row_test_rowu1));
bram_bufferx16 I393 ( .in(cram_pgateoffl2), .out(cram_pgateoff_rowu1));
bram_bufferx16 I394 ( .in(cram_rstl2), .out(cram_rst_rowu1));
bram_bufferx16 I395 ( .in(cram_wl_enl2), .out(cram_wl_en_rowu1));
bram_bufferx16 I396 ( .in(smc_writel2), .out(smc_write_rowu1));
bram_bufferx16 I397 ( .in(cram_vddoffl2), .out(cram_vddoff_rowu1));
bram_bufferx16 I398 ( .in(smc_row_incl2), .out(smc_row_inc_rowu1));
bram_bufferx16 I400 ( .in(smc_rsr_rstl2), .out(smc_rsr_rst_rowu1));
bram_bufferx16 I390 ( .in(smc_rsr_rstl1), .out(smc_rsr_rst_rowu0));
bram_bufferx16 I435 ( .in(tck_padl2), .out(tck_pad_rowu1));
bram_bufferx16 I384 ( .in(cram_rstl1), .out(cram_rst_rowu0));
bram_bufferx16 I290 ( .in(cm_clk_blbld), .out(net146));
bram_bufferx16 I260 ( .in(cm_clk_blbld), .out(net148));
bram_bufferx16 I385 ( .in(cram_vddoffl1), .out(cram_vddoff_rowu0));
bram_bufferx16 I386 ( .in(cram_wl_enl1), .out(cram_wl_en_rowu0));
bram_bufferx16 I387 ( .in(smc_row_incl1), .out(smc_row_inc_rowu0));
bram_bufferx16 I388 ( .in(smc_writel1), .out(smc_write_rowu0));
bram_bufferx16 I389 ( .in(core_por_bbl1), .out(core_por_b_rowu0));
bram_bufferx16 I383 ( .in(cram_pgateoffl1), .out(cram_pgateoff_rowu0));
bram_bufferx16 I437 ( .in(tck_padl1), .out(tck_pad_rowu0));
bram_bufferx16 I382 ( .in(row_testl2), .out(row_test_rowu0));
sg_bufx10 I421 ( .in(cf_lbank[479]), .out(monitor_celld[1]));
sg_bufx10 I235 ( .in(data_muxsel_bltld), .out(data_muxsel_bltld3));
sg_bufx10 I425 ( .in(monitor_celld[1]), .out(monitor_celld1[1]));
sg_bufx10 I424 ( .in(cf_lbank[300]), .out(monitor_celld2[0]));
sg_bufx10 I426 ( .in(monitor_celld1[1]), .out(monitor_celld2[1]));
sg_bufx10 I450_1_ ( .in(dff_out[1]), .out(cm_sdo_u1d1[1]));
sg_bufx10 I450_0_ ( .in(dff_out[0]), .out(cm_sdo_u1d1[0]));
sg_bufx10 I106_1_ ( .in(cm_sdo_u1[1]), .out(cm_sdo_u1d0[1]));
sg_bufx10 I106_0_ ( .in(cm_sdo_u1[0]), .out(cm_sdo_u1d0[0]));
sg_bufx10 I337 ( .in(core_por_bbl0), .out(core_por_bbl1));
sg_bufx10 I338 ( .in(smc_rsr_rstl0), .out(smc_rsr_rstl1));
sg_bufx10 I339 ( .in(row_testl1), .out(row_testl2));
sg_bufx10 I340 ( .in(j_rst_bl0), .out(j_rst_bl1));
sg_bufx10 I342 ( .in(smc_writel0), .out(smc_writel1));
sg_bufx10 I343 ( .in(smc_row_incl0), .out(smc_row_incl1));
sg_bufx10 I344 ( .in(cram_wl_enl0), .out(cram_wl_enl1));
sg_bufx10 I345 ( .in(cram_vddoffl0), .out(cram_vddoffl1));
sg_bufx10 I346 ( .in(cram_rstl0), .out(cram_rstl1));
sg_bufx10 I347 ( .in(cram_pgateoffl0), .out(cram_pgateoffl1));
sg_bufx10 I355 ( .in(cram_pgateoffl1), .out(cram_pgateoffl2));
sg_bufx10 I438 ( .in(tck_padl0), .out(tck_padl1));
sg_bufx10 I237 ( .in(data_muxsel1_bltld), .out(data_muxsel1_bltld3));
sg_bufx10 I351 ( .in(smc_row_incl1), .out(smc_row_incl2));
sg_bufx10 I368 ( .in(cram_pullup_bltld), .out(cram_pullup_bltld3));
sg_bufx10 I277 ( .in(cm_banksel_blbld[1]), .out(cm_banksel_bltld[1]));
sg_bufx10 I348 ( .in(smc_rsr_rstl1), .out(smc_rsr_rstl2));
sg_bufx10 I278_1_ ( .in(cm_sdo_u1d0[1]), .out(cm_sdo_u1d[1]));
sg_bufx10 I278_0_ ( .in(cm_sdo_u1d0[0]), .out(cm_sdo_u1d[0]));
sg_bufx10 I354 ( .in(cram_rstl1), .out(cram_rstl2));
sg_bufx10 I271 ( .in(data_muxsel1_blbld), .out(data_muxsel1_bltld));
sg_bufx10 I275 ( .in(cram_prec_blbld), .out(cram_prec_bltld));
sg_bufx10 I241 ( .in(en_8bconfig_b_bltld), .out(en_8bconfig_b_bltld3));
sg_bufx10 I353 ( .in(cram_vddoffl1), .out(cram_vddoffl2));
sg_bufx10 I357 ( .in(j_rst_bl1), .out(j_rst_bl2));
sg_bufx10 I356 ( .in(row_testl2), .out(row_testl3));
sg_bufx10 I273 ( .in(smc_wdis_dclk_blbld), .out(smc_wdis_dclk_bltld));
sg_bufx10 I279_1_ ( .in(cm_sdi_u1d[1]), .out(cm_sdi_u1d0[1]));
sg_bufx10 I279_0_ ( .in(cm_sdi_u1d[0]), .out(cm_sdi_u1d0[0]));
sg_bufx10 I272 ( .in(en_8bconfig_b_blbld), .out(en_8bconfig_b_bltld));
sg_bufx10 I274 ( .in(cram_write_blbld), .out(cram_write_bltld));
sg_bufx10 I239 ( .in(smc_wdis_dclk_bltld), .out(smc_wdis_dclk_bltld3));
sg_bufx10 I270 ( .in(data_muxsel_blbld), .out(data_muxsel_bltld));
sg_bufx10 I240 ( .in(cram_write_bltld), .out(cram_write_bltld3));
sg_bufx10 I238 ( .in(cram_prec_bltld), .out(cram_prec_bltld3));
sg_bufx10 I242 ( .in(cm_clk_bltld), .out(cm_clk_bltld3));
sg_bufx10 I236 ( .in(cm_banksel_bltld[1]), .out(cm_banksel_bltld3_1_));
sg_bufx10 I276 ( .in(cm_clk_blbld), .out(cm_clk_bltld));
sg_bufx10 I352 ( .in(cram_wl_enl1), .out(cram_wl_enl2));
sg_bufx10 I280_1_ ( .in(cm_sdi_u1d0[1]), .out(cm_sdi_u1d3[1]));
sg_bufx10 I280_0_ ( .in(cm_sdi_u1d0[0]), .out(cm_sdi_u1d3[0]));
sg_bufx10 I350 ( .in(smc_writel1), .out(smc_writel2));
sg_bufx10 I349 ( .in(core_por_bbl1), .out(core_por_b_rowu1));
sg_bufx10 I369 ( .in(cram_pullup_blbld), .out(cram_pullup_bltld));
sg_bufx10 I436 ( .in(tck_padl1), .out(tck_padl2));

endmodule
// Library - xpmem, Cell - ml_dff_bl, View - schematic
// LAST TIME SAVED: Sep  6 14:18:45 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_dff_bl ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - xpmem, Cell - ml_blsa_clk_buf, View - schematic
// LAST TIME SAVED: Sep  5 15:09:27 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_clk_buf ( o, in );
output  o;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net77), .Y(o));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_powersurg_buf, View - schematic
// LAST TIME SAVED: Jul 31 18:29:48 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_powersurg_buf ( o, in );
output  o;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I404 ( .A(net016), .Y(net012));
inv_hvt I405 ( .A(net012), .Y(o));
inv_hvt I391 ( .A(net77), .Y(net016));
inv_hvt I392 ( .A(in), .Y(net77));

endmodule
// Library - xpmem, Cell - ml_blsa_sch, View - schematic
// LAST TIME SAVED: Sep  6 14:30:13 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_sch ( dataout, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, datain, latch_clock, latch_reset, smc_wdic_clk );
output  dataout;

inout  bl;

input  cram_prec, cram_pullup_b, cram_write, data_muxsel, datain,
     latch_clock, latch_reset, smc_wdic_clk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_dff_bl Idff ( .R(latch_reset), .D(dff_in), .CLK(latch_clock),
     .QN(write_data_b), .Q(dff_data));
nor2_hvt I223 ( .A(net084), .B(write_data_b), .Y(n_gate));
inv_hvt I163 ( .A(write_data_b), .Y(dataout));
inv_hvt I159 ( .A(cram_prec), .Y(net0161));
inv_hvt I160 ( .A(cram_write), .Y(net084));
mux2_hvt I161 ( .in1(sa_out), .in0(datain), .out(latch_in),
     .sel(data_muxsel));
mux2_hvt I164 ( .in1(dff_data), .in0(latch_in), .out(dff_in),
     .sel(smc_wdic_clk));
nch_hvt  MN12 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN8 ( .D(sa_out), .B(gnd_), .G(cram_pullup_b), .S(gnd_));
nch_hvt  MN10 ( .D(net0166), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN13 ( .D(net0184), .B(gnd_), .G(n_gate), .S(gnd_));
nch_hvt  MN3 ( .D(sa_out), .B(gnd_), .G(bl), .S(gnd_));
nch_hvt  MN6 ( .D(bl), .B(gnd_), .G(n_gate), .S(gnd_));
pch_hvt  MP8 ( .D(net0148), .B(vdd_), .G(dataout), .S(vdd_));
pch_hvt  MP9 ( .D(bl), .B(vdd_), .G(net084), .S(net0148));
pch_hvt  MP13 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP12 ( .D(bl), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP14 ( .D(net0208), .B(vdd_), .G(net0161), .S(vdd_));
pch_hvt  MP4 ( .D(net0143), .B(vdd_), .G(cram_pullup_b), .S(vdd_));
pch_hvt  MP5 ( .D(sa_out), .B(vdd_), .G(bl), .S(net0143));
pch_hvt  MP15 ( .D(net0204), .B(vdd_), .G(net0161), .S(vdd_));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_bram10k, View - schematic
// LAST TIME SAVED: Mar 20 10:20:41 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tile_bram10k ( cram_prec_out, cram_write_out, data_out,
     para_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock, latch_reset, para_en, para_in,
     smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out, para_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, para_en, para_in, smc_wdic_clk;

inout [41:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:4]  data_dummy_in;

wire  [0:41]  dataout;

wire  [0:14]  ck;

wire  [0:5]  data_in;



ml_dff_bl I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net97), .Q(net119));
ml_dff_bl I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net92), .Q(data_dummy_in[4]));
ml_dff_bl I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net87), .Q(data_dummy_in[2]));
ml_dff_bl I179 ( .R(latch_reset), .D(data_in[0]), .CLK(ck[14]),
     .QN(net82), .Q(data_dummy_in[1]));
ml_dff_bl I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net77), .Q(data_dummy_in[3]));
ml_blsa_clk_buf I192_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I192_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I192_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I192_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I192_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I192_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I192_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I192_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I192_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I192_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I192_0_ ( .in(latch_clock), .o(ck[0]));
mux2_hvt I194 ( .in1(data_dummy_in[2]), .in0(dataout[3]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I161 ( .in1(para_in), .in0(dataout[1]), .out(data_out_mux),
     .sel(para_en));
mux2_hvt I199 ( .in1(net119), .in0(dataout[6]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I198 ( .in1(data_dummy_in[4]), .in0(dataout[5]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I196 ( .in1(data_dummy_in[1]), .in0(dataout[2]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I197 ( .in1(data_dummy_in[3]), .in0(dataout[4]),
     .out(data_in[3]), .sel(data_muxsel1));
inv_hvt I262 ( .A(data_out_mux), .Y(net151));
inv_hvt I261 ( .A(net151), .Y(data_in[0]));
inv_hvt I175 ( .A(dataout[1]), .Y(net154));
inv_hvt I176 ( .A(net154), .Y(para_out));
inv_hvt I172 ( .A(net160), .Y(data_out));
inv_hvt I171 ( .A(dataout[41]), .Y(net160));
inv_hvt I200 ( .A(net133), .Y(net0132));
inv_hvt I201 ( .A(net0132), .Y(net0133));
inv_hvt I202 ( .A(net0133), .Y(net0131));
inv_hvt I229 ( .A(latch_clock), .Y(net133));
inv_hvt I203 ( .A(net0131), .Y(net0126));
inv_hvt I204 ( .A(net0126), .Y(ck[14]));
ml_powersurg_buf I165 ( .in(cram_prec), .o(net162));
ml_powersurg_buf I163 ( .in(net162), .o(net164));
ml_powersurg_buf I162 ( .in(net170), .o(net166));
ml_powersurg_buf I169 ( .in(net166), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(cram_write), .o(net170));
ml_powersurg_buf I168 ( .in(net164), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[7]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[8]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[9]),
     .datain(data_in[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(data_in[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_41_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_40_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_39_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_38_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_37_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_36_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_35_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_34_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_33_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_32_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_31_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_30_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_29_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_28_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_27_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_26_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net170), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net162));
ml_blsa_sch Iml_blsa_sch_25_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_24_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_23_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_22_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_21_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_20_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_19_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_18_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[14]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[15]),
     .dataout(dataout[15]), .cram_prec(net164));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[13]),
     .data_muxsel(data_muxsel), .cram_write(net166), .bl(bl[14]),
     .dataout(dataout[14]), .cram_prec(net164));

endmodule
// Library - xpmem, Cell - ml_buf_ice5_2, View - schematic
// LAST TIME SAVED: Aug 15 18:07:29 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_buf_ice5_2 ( o, in, sel );
output  o;

input  in, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));
inv_hvt I391 ( .A(net77), .Y(o));

endmodule
// Library - xpmem, Cell - ml_blsa_tile, View - schematic
// LAST TIME SAVED: Sep  5 14:53:52 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tile ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [53:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [53:0]  dataout;

wire  [13:0]  ck;



ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
inv_hvt I172 ( .A(net48), .Y(data_out));
inv_hvt I171 ( .A(dataout[53]), .Y(net48));
ml_powersurg_buf I161 ( .in(cram_write), .o(net53));
ml_powersurg_buf I165 ( .in(net57), .o(net55));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net57));
ml_powersurg_buf I163 ( .in(net55), .o(net59));
ml_powersurg_buf I162 ( .in(net65), .o(net61));
ml_powersurg_buf I169 ( .in(net61), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net53), .o(net65));
ml_powersurg_buf I168 ( .in(net59), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[10]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[11]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[12]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[13]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));
ml_blsa_sch Iml_blsa_sch_47_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[47]),
     .dataout(dataout[47]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_46_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[46]),
     .dataout(dataout[46]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_45_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[45]),
     .dataout(dataout[45]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_44_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[44]),
     .dataout(dataout[44]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_43_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[43]),
     .dataout(dataout[43]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_42_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[42]),
     .dataout(dataout[42]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_41_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[41]),
     .dataout(dataout[41]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_40_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[40]),
     .dataout(dataout[40]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_39_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[39]),
     .dataout(dataout[39]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_38_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[38]),
     .dataout(dataout[38]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_37_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[37]),
     .dataout(dataout[37]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_36_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[36]),
     .dataout(dataout[36]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_35_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[35]),
     .dataout(dataout[35]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_34_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[34]),
     .dataout(dataout[34]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_33_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[33]),
     .dataout(dataout[33]), .cram_prec(net55));
ml_blsa_sch Iml_blsa_sch_32_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]),
     .data_muxsel(data_muxsel), .cram_write(net65), .bl(bl[32]),
     .dataout(dataout[32]), .cram_prec(net55));
ml_blsa_sch I170_53_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[52]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[53]),
     .dataout(dataout[53]), .cram_prec(net57));
ml_blsa_sch I170_52_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[0]), .datain(dataout[51]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[52]),
     .dataout(dataout[52]), .cram_prec(net57));
ml_blsa_sch I170_51_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[50]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[51]),
     .dataout(dataout[51]), .cram_prec(net57));
ml_blsa_sch I170_50_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[49]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[50]),
     .dataout(dataout[50]), .cram_prec(net57));
ml_blsa_sch I170_49_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[48]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[49]),
     .dataout(dataout[49]), .cram_prec(net57));
ml_blsa_sch I170_48_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[1]), .datain(dataout[47]),
     .data_muxsel(data_muxsel), .cram_write(net53), .bl(bl[48]),
     .dataout(dataout[48]), .cram_prec(net57));
ml_blsa_sch Iml_blsa_sch_31_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[31]),
     .dataout(dataout[31]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_30_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[30]),
     .dataout(dataout[30]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_29_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[29]),
     .dataout(dataout[29]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_28_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[28]),
     .dataout(dataout[28]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_27_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[27]),
     .dataout(dataout[27]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_26_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[26]),
     .dataout(dataout[26]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_25_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[25]),
     .dataout(dataout[25]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_24_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[24]),
     .dataout(dataout[24]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_23_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[23]),
     .dataout(dataout[23]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_22_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[22]),
     .dataout(dataout[22]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_21_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[21]),
     .dataout(dataout[21]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_20_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[20]),
     .dataout(dataout[20]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_19_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[19]),
     .dataout(dataout[19]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_18_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[18]),
     .dataout(dataout[18]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[17]),
     .dataout(dataout[17]), .cram_prec(net59));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]),
     .data_muxsel(data_muxsel), .cram_write(net61), .bl(bl[16]),
     .dataout(dataout[16]), .cram_prec(net59));

endmodule
// Library - xpmem, Cell - ml_blprecwrt_en, View - schematic
// LAST TIME SAVED: May 16 10:09:58 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blprecwrt_en ( data_out, action, clkin, data_in, rst );
output  data_out;

input  action, clkin, data_in, rst;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I161 ( .A(net89), .Y(net88));
inv_hvt I162 ( .A(action), .Y(net86));
inv_hvt I165 ( .A(net98), .Y(data_out));
nand3_hvt I160 ( .Y(net89), .B(data_in), .C(action), .A(clkin));
nor2_hvt I385 ( .A(net88), .B(net94), .Y(net98));
nor3_hvt I387 ( .B(net86), .Y(net94), .A(net98), .C(rst));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_bram10k, View - schematic
// LAST TIME SAVED: Nov 30 09:32:34 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2_bram10k ( data_out, latch_clock_out, para_out,
     prec_out, wrt_out, bl, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, datain, latch_clock_in, latch_reset,
     para_en, para_in, prec_in, smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, para_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, para_en, para_in, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in;

inout [95:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile_bram10k Iml_blsa_tile_0 ( .para_en(para_en),
     .para_in(para_in), .para_out(para_out), .bl(bl[41:0]),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[95:42]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
inv_hvt I183 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I184 ( .A(smc_wdic_clk), .Y(net088));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_buf_ice5, View - schematic
// LAST TIME SAVED: Aug 13 13:53:01 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_buf_ice5 ( o, in, sel );
output  o;

input  in, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(sel), .B(in), .Y(net77));
inv_hvt I391 ( .A(net77), .Y(o));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_last, View - schematic
// LAST TIME SAVED: Aug 28 08:58:43 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tile_last ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [17:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [17:0]  dataout;

wire  [4:0]  ck;



tiehi I186 ( .tiehi(net040));
ml_dff_bl Idff ( .R(latch_reset), .D(dataout[16]), .CLK(ck[0]),
     .QN(net50), .Q(net45));
ml_dff_bl I179 ( .R(latch_reset), .D(net58), .CLK(ck[0]), .QN(net49),
     .Q(net61));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_buf_ice5 I205 ( .in(net61), .o(data_out), .sel(net040));
mux2_hvt I174 ( .in1(net45), .in0(dataout[17]), .out(net58),
     .sel(data_muxsel));
ml_powersurg_buf I169 ( .in(cram_write), .o(cram_write_out));
ml_powersurg_buf I168 ( .in(cram_prec), .o(cram_prec_out));
ml_blsa_sch Iml_blsa_sch_17_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[16]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[17]), .dataout(dataout[17]));
ml_blsa_sch Iml_blsa_sch_16_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[15]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[16]), .dataout(dataout[16]));
ml_blsa_sch Iml_blsa_sch_15_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[14]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]));
ml_blsa_sch Iml_blsa_sch_14_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[13]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]));
ml_blsa_sch Iml_blsa_sch_13_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[12]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]));
ml_blsa_sch Iml_blsa_sch_12_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[11]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]));
ml_blsa_sch Iml_blsa_sch_11_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[10]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]));
ml_blsa_sch Iml_blsa_sch_10_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[9]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]));
ml_blsa_sch Iml_blsa_sch_9_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[8]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]));
ml_blsa_sch Iml_blsa_sch_8_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[2]),
     .datain(dataout[7]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]));
ml_blsa_sch Iml_blsa_sch_7_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[6]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]));
ml_blsa_sch Iml_blsa_sch_6_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[5]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]));
ml_blsa_sch Iml_blsa_sch_5_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[4]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]));
ml_blsa_sch Iml_blsa_sch_4_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[3]),
     .datain(dataout[3]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]));
ml_blsa_sch Iml_blsa_sch_3_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[2]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]));
ml_blsa_sch Iml_blsa_sch_2_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[1]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]));
ml_blsa_sch Iml_blsa_sch_1_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]),
     .datain(dataout[0]), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]));
ml_blsa_sch Iml_blsa_sch_0_ ( .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk), .cram_prec(cram_prec_out),
     .latch_reset(latch_reset), .latch_clock(ck[4]), .datain(datain),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_last, View - schematic
// LAST TIME SAVED: Nov 27 11:54:15 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2_last ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [125:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_1 ( .latch_reset(latch_reset_buf),
     .datain(data_tile), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_1st),
     .cram_prec(prec_en_1st), .data_out(datain_io),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[107:54]), .latch_clock(latch_clock_out),
     .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blsa_tile Iml_blsa_tile_0 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_dic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
ml_blsa_tile_last Iml_blsa_tile_last ( .bl(bl[125:108]),
     .latch_reset(latch_reset_buf), .datain(datain_io),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_1st), .cram_prec_out(prec_en_1st),
     .latch_clock(latch_clock_out), .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_dic_clk_buf));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
inv_hvt I185 ( .A(smc_wdic_clk), .Y(net091));
inv_hvt I184 ( .A(net091), .Y(smc_dic_clk_buf));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_blsa_tile_1st, View - schematic
// LAST TIME SAVED: Sep  6 14:29:58 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tile_1st ( cram_prec_out, cram_write_out, data_out, bl,
     cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk );
output  cram_prec_out, cram_write_out, data_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock, latch_reset, smc_wdic_clk;

inout [55:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:4]  data_dummy_in;

wire  [1:5]  data_in;

wire  [0:55]  dataout;

wire  [0:14]  ck;



ml_dff_bl I195 ( .R(latch_reset), .D(data_dummy_in[4]), .CLK(ck[14]),
     .QN(net132), .Q(net154));
ml_dff_bl I191 ( .R(latch_reset), .D(data_dummy_in[3]), .CLK(ck[14]),
     .QN(net137), .Q(data_dummy_in[4]));
ml_dff_bl I183 ( .R(latch_reset), .D(data_dummy_in[1]), .CLK(ck[14]),
     .QN(net142), .Q(data_dummy_in[2]));
ml_dff_bl I179 ( .R(latch_reset), .D(datain), .CLK(ck[14]),
     .QN(net147), .Q(data_dummy_in[1]));
ml_dff_bl I190 ( .R(latch_reset), .D(data_dummy_in[2]), .CLK(ck[14]),
     .QN(net152), .Q(data_dummy_in[3]));
ml_blsa_clk_buf I178_13_ ( .in(latch_clock), .o(ck[13]));
ml_blsa_clk_buf I178_12_ ( .in(latch_clock), .o(ck[12]));
ml_blsa_clk_buf I178_11_ ( .in(latch_clock), .o(ck[11]));
ml_blsa_clk_buf I178_10_ ( .in(latch_clock), .o(ck[10]));
ml_blsa_clk_buf I178_9_ ( .in(latch_clock), .o(ck[9]));
ml_blsa_clk_buf I178_8_ ( .in(latch_clock), .o(ck[8]));
ml_blsa_clk_buf I178_7_ ( .in(latch_clock), .o(ck[7]));
ml_blsa_clk_buf I178_6_ ( .in(latch_clock), .o(ck[6]));
ml_blsa_clk_buf I178_5_ ( .in(latch_clock), .o(ck[5]));
ml_blsa_clk_buf I178_4_ ( .in(latch_clock), .o(ck[4]));
ml_blsa_clk_buf I178_3_ ( .in(latch_clock), .o(ck[3]));
ml_blsa_clk_buf I178_2_ ( .in(latch_clock), .o(ck[2]));
ml_blsa_clk_buf I178_1_ ( .in(latch_clock), .o(ck[1]));
ml_blsa_clk_buf I178_0_ ( .in(latch_clock), .o(ck[0]));
ml_blsa_sch Iml_blsa_sch_15_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[14]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[15]), .dataout(dataout[15]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_14_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[13]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[14]), .dataout(dataout[14]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_13_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[12]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[13]), .dataout(dataout[13]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_12_ ( .latch_reset(latch_reset),
     .latch_clock(ck[10]), .datain(dataout[11]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[12]), .dataout(dataout[12]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_11_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[10]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[11]), .dataout(dataout[11]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_10_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[9]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[10]), .dataout(dataout[10]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_9_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[8]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[9]), .dataout(dataout[9]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_8_ ( .latch_reset(latch_reset),
     .latch_clock(ck[11]), .datain(dataout[7]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[8]), .dataout(dataout[8]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_7_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[6]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[7]), .dataout(dataout[7]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_6_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(dataout[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[6]), .dataout(dataout[6]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_5_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[5]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[5]), .dataout(dataout[5]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_4_ ( .latch_reset(latch_reset),
     .latch_clock(ck[12]), .datain(data_in[4]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[4]), .dataout(dataout[4]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_3_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[3]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[3]), .dataout(dataout[3]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_2_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[2]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[2]), .dataout(dataout[2]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_1_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(data_in[1]),
     .cram_prec(cram_prec_out), .data_muxsel(data_muxsel),
     .cram_write(cram_write_out), .bl(bl[1]), .dataout(dataout[1]),
     .cram_pullup_b(cram_pullup_b), .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_0_ ( .latch_reset(latch_reset),
     .latch_clock(ck[13]), .datain(datain), .cram_prec(cram_prec_out),
     .data_muxsel(data_muxsel), .cram_write(cram_write_out),
     .bl(bl[0]), .dataout(dataout[0]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_47_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[46]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[47]),
     .dataout(dataout[47]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_46_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[45]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[46]),
     .dataout(dataout[46]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_45_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[44]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[45]),
     .dataout(dataout[45]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_44_ ( .latch_reset(latch_reset),
     .latch_clock(ck[2]), .datain(dataout[43]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[44]),
     .dataout(dataout[44]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_43_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[42]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[43]),
     .dataout(dataout[43]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_42_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[41]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[42]),
     .dataout(dataout[42]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_41_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[40]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[41]),
     .dataout(dataout[41]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_40_ ( .latch_reset(latch_reset),
     .latch_clock(ck[3]), .datain(dataout[39]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[40]),
     .dataout(dataout[40]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_39_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[38]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[39]),
     .dataout(dataout[39]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_38_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[37]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[38]),
     .dataout(dataout[38]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_37_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[36]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[37]),
     .dataout(dataout[37]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_36_ ( .latch_reset(latch_reset),
     .latch_clock(ck[4]), .datain(dataout[35]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[36]),
     .dataout(dataout[36]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_35_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[34]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[35]),
     .dataout(dataout[35]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_34_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[33]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[34]),
     .dataout(dataout[34]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_33_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[32]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[33]),
     .dataout(dataout[33]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_32_ ( .latch_reset(latch_reset),
     .latch_clock(ck[5]), .datain(dataout[31]), .cram_prec(net106),
     .data_muxsel(data_muxsel), .cram_write(net116), .bl(bl[32]),
     .dataout(dataout[32]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_55_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[54]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[55]),
     .dataout(dataout[55]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_54_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[53]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[54]),
     .dataout(dataout[54]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_53_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[52]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[53]),
     .dataout(dataout[53]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_52_ ( .latch_reset(latch_reset), .latch_clock(ck[0]),
     .datain(dataout[51]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[52]),
     .dataout(dataout[52]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_51_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[50]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[51]),
     .dataout(dataout[51]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_50_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[49]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[50]),
     .dataout(dataout[50]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_49_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[48]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[49]),
     .dataout(dataout[49]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch I170_48_ ( .latch_reset(latch_reset), .latch_clock(ck[1]),
     .datain(dataout[47]), .cram_prec(net108),
     .data_muxsel(data_muxsel), .cram_write(net104), .bl(bl[48]),
     .dataout(dataout[48]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_31_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[30]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[31]),
     .dataout(dataout[31]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_30_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[29]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[30]),
     .dataout(dataout[30]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_29_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[28]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[29]),
     .dataout(dataout[29]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_28_ ( .latch_reset(latch_reset),
     .latch_clock(ck[6]), .datain(dataout[27]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[28]),
     .dataout(dataout[28]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_27_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[26]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[27]),
     .dataout(dataout[27]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_26_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[25]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[26]),
     .dataout(dataout[26]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_25_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[24]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[25]),
     .dataout(dataout[25]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_24_ ( .latch_reset(latch_reset),
     .latch_clock(ck[7]), .datain(dataout[23]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[24]),
     .dataout(dataout[24]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_23_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[22]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[23]),
     .dataout(dataout[23]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_22_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[21]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[22]),
     .dataout(dataout[22]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_21_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[20]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[21]),
     .dataout(dataout[21]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_20_ ( .latch_reset(latch_reset),
     .latch_clock(ck[8]), .datain(dataout[19]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[20]),
     .dataout(dataout[20]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_19_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[18]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[19]),
     .dataout(dataout[19]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_18_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[17]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[18]),
     .dataout(dataout[18]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_17_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[16]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[17]),
     .dataout(dataout[17]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_blsa_sch Iml_blsa_sch_16_ ( .latch_reset(latch_reset),
     .latch_clock(ck[9]), .datain(dataout[15]), .cram_prec(net110),
     .data_muxsel(data_muxsel), .cram_write(net112), .bl(bl[16]),
     .dataout(dataout[16]), .cram_pullup_b(cram_pullup_b),
     .smc_wdic_clk(smc_wdic_clk));
ml_powersurg_buf I161 ( .in(cram_write), .o(net104));
ml_powersurg_buf I165 ( .in(net108), .o(net106));
ml_powersurg_buf I160 ( .in(cram_prec), .o(net108));
ml_powersurg_buf I163 ( .in(net106), .o(net110));
ml_powersurg_buf I162 ( .in(net116), .o(net112));
ml_powersurg_buf I169 ( .in(net112), .o(cram_write_out));
ml_powersurg_buf I166 ( .in(net104), .o(net116));
ml_powersurg_buf I168 ( .in(net110), .o(cram_prec_out));
inv_hvt I171 ( .A(dataout[55]), .Y(net121));
inv_hvt I172 ( .A(net121), .Y(data_out));
inv_hvt I224 ( .A(net0130), .Y(ck[14]));
inv_hvt I225 ( .A(net0129), .Y(net0130));
inv_hvt I226 ( .A(net0126), .Y(net0129));
inv_hvt I229 ( .A(latch_clock), .Y(net0122));
inv_hvt I227 ( .A(net0124), .Y(net0126));
inv_hvt I228 ( .A(net0122), .Y(net0124));
mux2_hvt I197 ( .in1(net154), .in0(dataout[4]), .out(data_in[5]),
     .sel(data_muxsel1));
mux2_hvt I185 ( .in1(data_dummy_in[2]), .in0(dataout[1]),
     .out(data_in[2]), .sel(data_muxsel1));
mux2_hvt I193 ( .in1(data_dummy_in[4]), .in0(dataout[3]),
     .out(data_in[4]), .sel(data_muxsel1));
mux2_hvt I180 ( .in1(data_dummy_in[1]), .in0(dataout[0]),
     .out(data_in[1]), .sel(data_muxsel1));
mux2_hvt I188 ( .in1(data_dummy_in[3]), .in0(dataout[2]),
     .out(data_in[3]), .sel(data_muxsel1));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2_1st, View - schematic
// LAST TIME SAVED: Aug 13 13:56:25 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2_1st ( data_out, latch_clock_out, prec_out,
     wrt_out, bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [109:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I186 ( .A(data_muxsel), .Y(net55));
inv_hvt I187 ( .A(net55), .Y(data_muxsel_buf));
inv_hvt I190 ( .A(net61), .Y(cram_pullup_buf));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net61));
inv_hvt I198 ( .A(smc_wdic_clk), .Y(net63));
inv_hvt I199 ( .A(net63), .Y(smc_wdic_clk_buf));
inv_hvt I197 ( .A(latch_clock_in), .Y(net67));
inv_hvt I196 ( .A(net67), .Y(latch_clock_out));
inv_hvt I194 ( .A(latch_reset), .Y(net71));
inv_hvt I195 ( .A(net71), .Y(latch_reset_buf));
ml_blsa_tile_1st Iml_blsa_tile_1st_0 ( .bl(bl[55:0]),
     .cram_pullup_b(cram_pullup_buf), .latch_clock(latch_clock_out),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .datain(datain), .data_muxsel1(data_muxsel1),
     .data_muxsel(data_muxsel_buf), .cram_write(wrt_en_mid),
     .cram_prec(prec_en_mid), .data_out(data_tile),
     .cram_write_out(wrt_en_last), .cram_prec_out(prec_en_last));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_buf),
     .latch_clock(latch_clock_out), .smc_wdic_clk(smc_wdic_clk_buf),
     .latch_reset(latch_reset_buf), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[109:56]));

endmodule
// Library - xpmem, Cell - ml_blsa_tilex2, View - schematic
// LAST TIME SAVED: Jun 29 11:04:00 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_tilex2 ( data_out, latch_clock_out, prec_out, wrt_out,
     bl, cram_prec, cram_pullup_b, cram_write, data_muxsel,
     data_muxsel1, datain, latch_clock_in, latch_reset, prec_in,
     smc_clk_dpr, smc_wdic_clk, wrt_in );
output  data_out, latch_clock_out, prec_out, wrt_out;


input  cram_prec, cram_pullup_b, cram_write, data_muxsel, data_muxsel1,
     datain, latch_clock_in, latch_reset, prec_in, smc_clk_dpr,
     smc_wdic_clk, wrt_in;

inout [107:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tile Iml_blsa_tile_0 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(datain),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_en_mid), .cram_prec(prec_en_mid),
     .data_out(data_tile), .cram_write_out(wrt_en_last),
     .cram_prec_out(prec_en_last), .bl(bl[53:0]));
ml_blsa_tile Iml_blsa_tile_1 ( .cram_pullup_b(cram_pullup_b_buf),
     .smc_wdic_clk(smc_wdic_clk_buf), .latch_reset(latch_reset_buf),
     .latch_clock(latch_clock_out), .datain(data_tile),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel_buf),
     .cram_write(wrt_out), .cram_prec(prec_out), .data_out(data_out),
     .cram_write_out(wrt_en_mid), .cram_prec_out(prec_en_mid),
     .bl(bl[107:54]));
ml_blprecwrt_en Iml_blprecwrt_en_wrt ( .rst(latch_reset),
     .data_in(wrt_in), .clkin(smc_clk_dpr), .action(cram_write),
     .data_out(wrt_out));
ml_blprecwrt_en Iml_blprecwrt_en_rd ( .rst(latch_reset),
     .data_in(prec_in), .clkin(smc_clk_dpr), .action(cram_prec),
     .data_out(prec_out));
inv_hvt I183 ( .A(net088), .Y(smc_wdic_clk_buf));
inv_hvt I184 ( .A(smc_wdic_clk), .Y(net088));
inv_hvt I197 ( .A(latch_clock_in), .Y(net100));
inv_hvt I190 ( .A(net92), .Y(cram_pullup_b_buf));
inv_hvt I196 ( .A(net100), .Y(latch_clock_out));
inv_hvt I195 ( .A(net94), .Y(latch_reset_buf));
inv_hvt I194 ( .A(latch_reset), .Y(net94));
inv_hvt I191 ( .A(cram_pullup_b), .Y(net92));
inv_hvt I187 ( .A(net86), .Y(data_muxsel_buf));
inv_hvt I186 ( .A(data_muxsel), .Y(net86));

endmodule
// Library - xpmem, Cell - ml_blsa_bank10k, View - schematic
// LAST TIME SAVED: Nov 30 09:26:09 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module ml_blsa_bank10k ( cm_sdo_u, bl, banksel, cm_sdi_u,
     cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk );


input  banksel, cor_en_8bpcfg_b, cram_prec, cram_pullup_b, cram_write,
     data_muxsel, data_muxsel1, latch_reset, smc_clk, smc_wdic_clk;

output [1:0]  cm_sdo_u;

inout [871:0]  bl;

input [1:0]  cm_sdi_u;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_tilex2_bram10k Ilt_0809 ( .para_en(cor_en_8bpcfg_buf),
     .para_in(sdi1_buf), .para_out(para_out), .bl(bl[529:434]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net370),
     .latch_clock_out(net164), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret), .wrt_in(wrt_out_1011),
     .prec_in(prec_out_1011), .latch_reset(latch_reset_buf),
     .datain(data_out_67), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_89),
     .prec_out(prec_out_89), .data_out(data_out_89));
tiehi I267 ( .tiehi(net272));
tiehi I268 ( .tiehi(net147));
tiehi I272 ( .tiehi(net148));
tiehi I271 ( .tiehi(net149));
tiehi I273 ( .tiehi(net150));
tiehi I270 ( .tiehi(net151));
tiehi I269 ( .tiehi(net152));
ml_dff_bl I146 ( .R(latch_reset_buf), .D(para_out), .CLK(smc_clk),
     .QN(net156), .Q(net197));
nor2_hvt I254 ( .B(net184), .Y(net185), .A(cram_pullup_b));
inv_hvt I253 ( .A(cor_en_8bpcfg_b), .Y(net182));
inv_hvt I256 ( .A(banksel), .Y(net184));
inv_hvt I255 ( .A(net185), .Y(cram_pullup_logic_b));
inv_hvt I189 ( .A(smc_clk), .Y(net188));
ml_buf_ice5 I247 ( .in(cm_sdi_u[1]), .o(sdi1_buf), .sel(net148));
ml_buf_ice5 I249 ( .in(net182), .o(cor_en_8bpcfg_buf), .sel(net148));
ml_buf_ice5 I265 ( .in(net148), .o(cm_sdo_u[0]), .sel(net197));
ml_buf_ice5 I257 ( .in(smc_wdic_clk), .o(smc_wdic_clk_buf),
     .sel(banksel));
ml_buf_ice5 I203 ( .in(data_muxsel1), .o(data_muxsel1_buf),
     .sel(banksel));
ml_buf_ice5 I205 ( .in(latch_reset), .o(latch_reset_buf),
     .sel(net150));
ml_buf_ice5 I207 ( .in(cram_write), .o(cram_write_buf), .sel(banksel));
ml_buf_ice5 I208 ( .in(cram_pullup_logic_b), .o(cram_pullup_b_buf),
     .sel(cram_pullup_logic_b));
ml_buf_ice5 I201 ( .in(cram_prec), .o(cram_prec_buf), .sel(banksel));
ml_buf_ice5 I216 ( .in(net149), .o(net217), .sel(net149));
ml_buf_ice5 I245 ( .in(cm_sdi_u[0]), .o(sdi0_buf), .sel(net148));
ml_buf_ice5 I187 ( .in(smc_clk), .o(smc_clk_buf), .sel(smc_clk));
ml_buf_ice5 I188 ( .in(net188), .o(smc_clk_buf_b_ret), .sel(net188));
ml_buf_ice5 I204 ( .in(data_muxsel), .o(data_muxsel_buf),
     .sel(banksel));
ml_buf_ice5 I227 ( .in(net152), .o(net232), .sel(net152));
nor3_hvt I217 ( .B(net151), .Y(net235), .A(net151), .C(net151));
nor3_hvt I220 ( .B(net243), .Y(net239), .A(net243), .C(net243));
nor3_hvt I218 ( .B(net235), .Y(net243), .A(net235), .C(net235));
nand3_hvt I231 ( .Y(net246), .B(net250), .C(net250), .A(net250));
nand3_hvt I230 ( .Y(net250), .B(net254), .C(net254), .A(net254));
nand3_hvt I224 ( .Y(net254), .B(net147), .C(net147), .A(net147));
ml_blsa_tilex2_last Ilt_1415 ( .bl(bl[871:746]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(smc_clk),
     .latch_clock_out(net269), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf), .wrt_in(net272), .prec_in(net272),
     .latch_reset(latch_reset_buf), .datain(data_out_1213),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_1415), .prec_out(prec_out_1415),
     .data_out(cm_sdo_u[1]));
ml_blsa_tilex2_1st ilt_0001 ( .wrt_in(wrt_out_23),
     .prec_in(prec_out_23), .latch_reset(latch_reset_buf),
     .datain(sdi0_buf), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .bl(bl[109:0]), .cram_prec(cram_prec_buf), .wrt_out(wrt_out_01),
     .prec_out(prec_out_01), .data_out(data_out_01),
     .latch_clock_in(net303), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_out(net297), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret));
ml_blsa_tilex2 Ilt_0203 ( .bl(bl[217:110]),
     .cram_pullup_b(cram_pullup_b_buf), .latch_clock_in(net353),
     .latch_clock_out(net303), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf), .wrt_in(wrt_out_45),
     .prec_in(prec_out_45), .latch_reset(latch_reset_buf),
     .datain(data_out_01), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_23),
     .prec_out(prec_out_23), .data_out(data_out_23));
ml_blsa_tilex2 Ilt_0607 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(net164), .latch_clock_out(net319),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf),
     .wrt_in(wrt_out_89), .prec_in(prec_out_89),
     .latch_reset(latch_reset_buf), .datain(data_out_45),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_67), .prec_out(prec_out_67),
     .data_out(data_out_67), .bl(bl[433:326]));
ml_blsa_tilex2 Ilt_1213 ( .wrt_in(wrt_out_1415),
     .prec_in(prec_out_1415), .latch_reset(latch_reset_buf),
     .datain(data_out_1011), .data_muxsel1(data_muxsel1_buf),
     .data_muxsel(data_muxsel_buf), .cram_write(cram_write_buf),
     .cram_prec(cram_prec_buf), .wrt_out(wrt_out_1213),
     .prec_out(prec_out_1213), .data_out(data_out_1213),
     .latch_clock_in(net269), .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_out(net347), .smc_wdic_clk(smc_wdic_clk_buf),
     .smc_clk_dpr(smc_clk_buf_b_ret), .bl(bl[745:638]));
ml_blsa_tilex2 Ilt_0405 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(net319), .latch_clock_out(net353),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf_b_ret),
     .wrt_in(wrt_out_67), .prec_in(prec_out_67),
     .latch_reset(latch_reset_buf), .datain(data_out_23),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_45), .prec_out(prec_out_45),
     .data_out(data_out_45), .bl(bl[325:218]));
ml_blsa_tilex2 Ilt_1011 ( .cram_pullup_b(cram_pullup_b_buf),
     .latch_clock_in(net347), .latch_clock_out(net370),
     .smc_wdic_clk(smc_wdic_clk_buf), .smc_clk_dpr(smc_clk_buf),
     .wrt_in(wrt_out_1213), .prec_in(prec_out_1213),
     .latch_reset(latch_reset_buf), .datain(data_out_89),
     .data_muxsel1(data_muxsel1_buf), .data_muxsel(data_muxsel_buf),
     .cram_write(cram_write_buf), .cram_prec(cram_prec_buf),
     .wrt_out(wrt_out_1011), .prec_out(prec_out_1011),
     .data_out(data_out_1011), .bl(bl[637:530]));

endmodule
// Library - xpmem, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jun  5 11:34:46 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - io, Cell - PDT08DGZ, View - schematic
// LAST TIME SAVED: Aug 13 15:32:26 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module PDT08DGZ ( PAD, I, OEN );
inout  PAD;

input  I, OEN;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - xpmem, Cell - sg_bufx10bot, View - schematic
// LAST TIME SAVED: Sep 18 11:01:27 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module sg_bufx10bot ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - chip, Cell - CHIP_route_bot10k, View - schematic
// LAST TIME SAVED: Oct  6 15:01:12 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module CHIP_route_bot10k ( cm_banksel_blbld1_0_, cm_banksel_blbld_1_,
     cm_clk_blbld, cm_sdi_u1d, cm_sdo_u0d1, cm_sdo_u1d3, cm_sdo_u2d1,
     core_por_b2, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, crst_filterout, data_muxsel1_blbld,
     data_muxsel_blbld, en_8bconfig_b_blbld, j_rst_bl0, last_rsr3,
     monitor_celld4, row_testl1, smc_core_por_bottom1,
     smc_core_por_bottom2, smc_row_incl0, smc_rsr_rstl0,
     smc_wdis_dclk_blbld, smc_writel0, spi_ss_in_bbankd, tck_padl0,
     bl_bot, cm_banksel, cm_banksel_blbrd_2_, cm_clk_blbrd, cm_sdi_u0,
     cm_sdi_u1, cm_sdi_u2d, cm_sdo_u1d1, core_por_b0, core_por_b_rowu2,
     core_por_bb, core_por_rowu0, cram_pgateoff, cram_prec,
     cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en, cram_write,
     creset_b_int, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, monitor_celld2,
     row_test0, smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd,
     smc_write, spi_ss_in_bbank, vddio_botbank, vddio_spi );
output  cm_banksel_blbld1_0_, cm_banksel_blbld_1_, cm_clk_blbld,
     core_por_b2, core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, crst_filterout, data_muxsel1_blbld,
     data_muxsel_blbld, en_8bconfig_b_blbld, j_rst_bl0, last_rsr3,
     row_testl1, smc_core_por_bottom1, smc_core_por_bottom2,
     smc_row_incl0, smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0,
     tck_padl0;


input  cm_banksel_blbrd_2_, cm_clk_blbrd, core_por_b0,
     core_por_b_rowu2, core_por_bb, core_por_rowu0, cram_pgateoff,
     cram_prec, cram_pullup_b, cram_rst, cram_vddoff, cram_wl_en,
     cram_write, creset_b_int, data_muxsel1_blbrd, data_muxsel_blbrd,
     en_8bconfig_b_blbrd, j_rst_b, j_tck, last_rsr1, row_test0,
     smc_row_inc, smc_rsr_rst, smc_wdis_dclk_blbrd, smc_write,
     vddio_botbank, vddio_spi;

output [4:0]  spi_ss_in_bbankd;
output [1:0]  cm_sdo_u2d1;
output [1:0]  cm_sdo_u0d1;
output [1:0]  cm_sdi_u1d;
output [1:0]  monitor_celld4;
output [1:0]  cm_sdo_u1d3;

inout [1743:0]  bl_bot;

input [1:0]  cm_sdi_u1;
input [4:0]  spi_ss_in_bbank;
input [1:0]  cm_sdi_u2d;
input [1:0]  cm_sdo_u1d1;
input [1:0]  cm_banksel;
input [1:0]  monitor_celld2;
input [1:0]  cm_sdi_u0;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u2;

wire  [1:0]  dff_u2_d1;

wire  [1:0]  monitor_celld3;

wire  [0:1]  net0195;

wire  [0:1]  net0200;

wire  [0:1]  net0194;

wire  [1:0]  dff_u1_d1;

wire  [1:0]  cm_sdo_u1_buf;

wire  [1:0]  cm_sdo_u0_buf;

wire  [1:0]  dff_u0_d1;

wire  [1:0]  cm_sdo_u0;

wire  [1:0]  dff_u0_d0;

wire  [1:0]  cm_sdi_u0d1;

wire  [2:2]  cm_banksel_blbrd1;

wire  [1:0]  dff_u2_d0;

wire  [1:0]  cm_sdi_u2d_buf;

wire  [0:1]  net0254;

wire  [0:1]  net0197;

wire  [0:1]  net0193;

wire  [0:1]  net0260;

wire  [0:1]  net0192;

wire  [0:1]  net0278;



eh_io_pup_2_new I4 ( .core_por_b(core_por_b0), .vdd_io(vddio_botbank),
     .por_b(smc_core_por_bottom1));
eh_io_pup_2_new I5 ( .core_por_b(core_por_b0), .vdd_io(vddio_spi),
     .por_b(smc_core_por_bottom2));
tielo I559_1_ ( .tielo(net0197[0]));
tielo I559_0_ ( .tielo(net0197[1]));
tielo I560_1_ ( .tielo(net0192[0]));
tielo I560_0_ ( .tielo(net0192[1]));
tielo I561_1_ ( .tielo(net0193[0]));
tielo I561_0_ ( .tielo(net0193[1]));
tielo I562_1_ ( .tielo(net0194[0]));
tielo I562_0_ ( .tielo(net0194[1]));
tielo I563_1_ ( .tielo(net0195[0]));
tielo I563_0_ ( .tielo(net0195[1]));
tielo I564 ( .tielo(net0196));
sg_dffbuf_modified I535_1_ ( .r(net0197[0]), .d(cm_sdo_u0[1]),
     .clk(net395), .dffout(dff_u0_d0[1]));
sg_dffbuf_modified I535_0_ ( .r(net0197[1]), .d(cm_sdo_u0[0]),
     .clk(net395), .dffout(dff_u0_d0[0]));
sg_dffbuf_modified I546_1_ ( .r(net0194[0]), .d(cm_sdo_u2[1]),
     .clk(net400), .dffout(dff_u2_d0[1]));
sg_dffbuf_modified I546_0_ ( .r(net0194[1]), .d(cm_sdo_u2[0]),
     .clk(net400), .dffout(dff_u2_d0[0]));
sg_dffbuf_modified I537_1_ ( .r(net0192[0]), .d(cm_sdo_u1_buf[1]),
     .clk(net393), .dffout(dff_u1_d1[1]));
sg_dffbuf_modified I537_0_ ( .r(net0192[1]), .d(cm_sdo_u1_buf[0]),
     .clk(net393), .dffout(dff_u1_d1[0]));
sg_dffbuf_modified I545_1_ ( .r(net0195[0]), .d(dff_u2_d0[1]),
     .clk(net401), .dffout(dff_u2_d1[1]));
sg_dffbuf_modified I545_0_ ( .r(net0195[1]), .d(dff_u2_d0[0]),
     .clk(net401), .dffout(dff_u2_d1[0]));
sg_dffbuf_modified I462_1_ ( .r(net0193[0]), .d(cm_sdo_u0_buf[1]),
     .clk(net393), .dffout(dff_u0_d1[1]));
sg_dffbuf_modified I462_0_ ( .r(net0193[1]), .d(cm_sdo_u0_buf[0]),
     .clk(net393), .dffout(dff_u0_d1[0]));
sg_dffbuf_modified I512 ( .r(net0196), .d(last_rsr2), .clk(net393),
     .dffout(net374));
ml_blsa_bank10k Iblbr ( .bl(bl_bot[1743:872]),
     .smc_wdic_clk(predata_smc_wdis_dclk),
     .smc_clk(predata_smc_clk_out), .cm_sdi_u(cm_sdi_u2d_buf[1:0]),
     .latch_reset(core_por_b_rowu2), .cm_sdo_u(cm_sdo_u2[1:0]),
     .data_muxsel1(predata_muxsel1), .data_muxsel(predata_muxsel),
     .cram_write(predata_cram_write), .cram_prec(predata_cram_prec),
     .cor_en_8bpcfg_b(predata_en_8bconfig_b),
     .cram_pullup_b(predata_cram_pullup_b),
     .banksel(cm_banksel_blbrd1[2]));
ml_blsa_bank10k Iblbl ( .bl({bl_bot[0], bl_bot[1], bl_bot[2],
     bl_bot[3], bl_bot[4], bl_bot[5], bl_bot[6], bl_bot[7], bl_bot[8],
     bl_bot[9], bl_bot[10], bl_bot[11], bl_bot[12], bl_bot[13],
     bl_bot[14], bl_bot[15], bl_bot[16], bl_bot[17], bl_bot[18],
     bl_bot[19], bl_bot[20], bl_bot[21], bl_bot[22], bl_bot[23],
     bl_bot[24], bl_bot[25], bl_bot[26], bl_bot[27], bl_bot[28],
     bl_bot[29], bl_bot[30], bl_bot[31], bl_bot[32], bl_bot[33],
     bl_bot[34], bl_bot[35], bl_bot[36], bl_bot[37], bl_bot[38],
     bl_bot[39], bl_bot[40], bl_bot[41], bl_bot[42], bl_bot[43],
     bl_bot[44], bl_bot[45], bl_bot[46], bl_bot[47], bl_bot[48],
     bl_bot[49], bl_bot[50], bl_bot[51], bl_bot[52], bl_bot[53],
     bl_bot[54], bl_bot[55], bl_bot[56], bl_bot[57], bl_bot[58],
     bl_bot[59], bl_bot[60], bl_bot[61], bl_bot[62], bl_bot[63],
     bl_bot[64], bl_bot[65], bl_bot[66], bl_bot[67], bl_bot[68],
     bl_bot[69], bl_bot[70], bl_bot[71], bl_bot[72], bl_bot[73],
     bl_bot[74], bl_bot[75], bl_bot[76], bl_bot[77], bl_bot[78],
     bl_bot[79], bl_bot[80], bl_bot[81], bl_bot[82], bl_bot[83],
     bl_bot[84], bl_bot[85], bl_bot[86], bl_bot[87], bl_bot[88],
     bl_bot[89], bl_bot[90], bl_bot[91], bl_bot[92], bl_bot[93],
     bl_bot[94], bl_bot[95], bl_bot[96], bl_bot[97], bl_bot[98],
     bl_bot[99], bl_bot[100], bl_bot[101], bl_bot[102], bl_bot[103],
     bl_bot[104], bl_bot[105], bl_bot[106], bl_bot[107], bl_bot[108],
     bl_bot[109], bl_bot[110], bl_bot[111], bl_bot[112], bl_bot[113],
     bl_bot[114], bl_bot[115], bl_bot[116], bl_bot[117], bl_bot[118],
     bl_bot[119], bl_bot[120], bl_bot[121], bl_bot[122], bl_bot[123],
     bl_bot[124], bl_bot[125], bl_bot[126], bl_bot[127], bl_bot[128],
     bl_bot[129], bl_bot[130], bl_bot[131], bl_bot[132], bl_bot[133],
     bl_bot[134], bl_bot[135], bl_bot[136], bl_bot[137], bl_bot[138],
     bl_bot[139], bl_bot[140], bl_bot[141], bl_bot[142], bl_bot[143],
     bl_bot[144], bl_bot[145], bl_bot[146], bl_bot[147], bl_bot[148],
     bl_bot[149], bl_bot[150], bl_bot[151], bl_bot[152], bl_bot[153],
     bl_bot[154], bl_bot[155], bl_bot[156], bl_bot[157], bl_bot[158],
     bl_bot[159], bl_bot[160], bl_bot[161], bl_bot[162], bl_bot[163],
     bl_bot[164], bl_bot[165], bl_bot[166], bl_bot[167], bl_bot[168],
     bl_bot[169], bl_bot[170], bl_bot[171], bl_bot[172], bl_bot[173],
     bl_bot[174], bl_bot[175], bl_bot[176], bl_bot[177], bl_bot[178],
     bl_bot[179], bl_bot[180], bl_bot[181], bl_bot[182], bl_bot[183],
     bl_bot[184], bl_bot[185], bl_bot[186], bl_bot[187], bl_bot[188],
     bl_bot[189], bl_bot[190], bl_bot[191], bl_bot[192], bl_bot[193],
     bl_bot[194], bl_bot[195], bl_bot[196], bl_bot[197], bl_bot[198],
     bl_bot[199], bl_bot[200], bl_bot[201], bl_bot[202], bl_bot[203],
     bl_bot[204], bl_bot[205], bl_bot[206], bl_bot[207], bl_bot[208],
     bl_bot[209], bl_bot[210], bl_bot[211], bl_bot[212], bl_bot[213],
     bl_bot[214], bl_bot[215], bl_bot[216], bl_bot[217], bl_bot[218],
     bl_bot[219], bl_bot[220], bl_bot[221], bl_bot[222], bl_bot[223],
     bl_bot[224], bl_bot[225], bl_bot[226], bl_bot[227], bl_bot[228],
     bl_bot[229], bl_bot[230], bl_bot[231], bl_bot[232], bl_bot[233],
     bl_bot[234], bl_bot[235], bl_bot[236], bl_bot[237], bl_bot[238],
     bl_bot[239], bl_bot[240], bl_bot[241], bl_bot[242], bl_bot[243],
     bl_bot[244], bl_bot[245], bl_bot[246], bl_bot[247], bl_bot[248],
     bl_bot[249], bl_bot[250], bl_bot[251], bl_bot[252], bl_bot[253],
     bl_bot[254], bl_bot[255], bl_bot[256], bl_bot[257], bl_bot[258],
     bl_bot[259], bl_bot[260], bl_bot[261], bl_bot[262], bl_bot[263],
     bl_bot[264], bl_bot[265], bl_bot[266], bl_bot[267], bl_bot[268],
     bl_bot[269], bl_bot[270], bl_bot[271], bl_bot[272], bl_bot[273],
     bl_bot[274], bl_bot[275], bl_bot[276], bl_bot[277], bl_bot[278],
     bl_bot[279], bl_bot[280], bl_bot[281], bl_bot[282], bl_bot[283],
     bl_bot[284], bl_bot[285], bl_bot[286], bl_bot[287], bl_bot[288],
     bl_bot[289], bl_bot[290], bl_bot[291], bl_bot[292], bl_bot[293],
     bl_bot[294], bl_bot[295], bl_bot[296], bl_bot[297], bl_bot[298],
     bl_bot[299], bl_bot[300], bl_bot[301], bl_bot[302], bl_bot[303],
     bl_bot[304], bl_bot[305], bl_bot[306], bl_bot[307], bl_bot[308],
     bl_bot[309], bl_bot[310], bl_bot[311], bl_bot[312], bl_bot[313],
     bl_bot[314], bl_bot[315], bl_bot[316], bl_bot[317], bl_bot[318],
     bl_bot[319], bl_bot[320], bl_bot[321], bl_bot[322], bl_bot[323],
     bl_bot[324], bl_bot[325], bl_bot[326], bl_bot[327], bl_bot[328],
     bl_bot[329], bl_bot[330], bl_bot[331], bl_bot[332], bl_bot[333],
     bl_bot[334], bl_bot[335], bl_bot[336], bl_bot[337], bl_bot[338],
     bl_bot[339], bl_bot[340], bl_bot[341], bl_bot[342], bl_bot[343],
     bl_bot[344], bl_bot[345], bl_bot[346], bl_bot[347], bl_bot[348],
     bl_bot[349], bl_bot[350], bl_bot[351], bl_bot[352], bl_bot[353],
     bl_bot[354], bl_bot[355], bl_bot[356], bl_bot[357], bl_bot[358],
     bl_bot[359], bl_bot[360], bl_bot[361], bl_bot[362], bl_bot[363],
     bl_bot[364], bl_bot[365], bl_bot[366], bl_bot[367], bl_bot[368],
     bl_bot[369], bl_bot[370], bl_bot[371], bl_bot[372], bl_bot[373],
     bl_bot[374], bl_bot[375], bl_bot[376], bl_bot[377], bl_bot[378],
     bl_bot[379], bl_bot[380], bl_bot[381], bl_bot[382], bl_bot[383],
     bl_bot[384], bl_bot[385], bl_bot[386], bl_bot[387], bl_bot[388],
     bl_bot[389], bl_bot[390], bl_bot[391], bl_bot[392], bl_bot[393],
     bl_bot[394], bl_bot[395], bl_bot[396], bl_bot[397], bl_bot[398],
     bl_bot[399], bl_bot[400], bl_bot[401], bl_bot[402], bl_bot[403],
     bl_bot[404], bl_bot[405], bl_bot[406], bl_bot[407], bl_bot[408],
     bl_bot[409], bl_bot[410], bl_bot[411], bl_bot[412], bl_bot[413],
     bl_bot[414], bl_bot[415], bl_bot[416], bl_bot[417], bl_bot[418],
     bl_bot[419], bl_bot[420], bl_bot[421], bl_bot[422], bl_bot[423],
     bl_bot[424], bl_bot[425], bl_bot[426], bl_bot[427], bl_bot[428],
     bl_bot[429], bl_bot[430], bl_bot[431], bl_bot[432], bl_bot[433],
     bl_bot[434], bl_bot[435], bl_bot[436], bl_bot[437], bl_bot[438],
     bl_bot[439], bl_bot[440], bl_bot[441], bl_bot[442], bl_bot[443],
     bl_bot[444], bl_bot[445], bl_bot[446], bl_bot[447], bl_bot[448],
     bl_bot[449], bl_bot[450], bl_bot[451], bl_bot[452], bl_bot[453],
     bl_bot[454], bl_bot[455], bl_bot[456], bl_bot[457], bl_bot[458],
     bl_bot[459], bl_bot[460], bl_bot[461], bl_bot[462], bl_bot[463],
     bl_bot[464], bl_bot[465], bl_bot[466], bl_bot[467], bl_bot[468],
     bl_bot[469], bl_bot[470], bl_bot[471], bl_bot[472], bl_bot[473],
     bl_bot[474], bl_bot[475], bl_bot[476], bl_bot[477], bl_bot[478],
     bl_bot[479], bl_bot[480], bl_bot[481], bl_bot[482], bl_bot[483],
     bl_bot[484], bl_bot[485], bl_bot[486], bl_bot[487], bl_bot[488],
     bl_bot[489], bl_bot[490], bl_bot[491], bl_bot[492], bl_bot[493],
     bl_bot[494], bl_bot[495], bl_bot[496], bl_bot[497], bl_bot[498],
     bl_bot[499], bl_bot[500], bl_bot[501], bl_bot[502], bl_bot[503],
     bl_bot[504], bl_bot[505], bl_bot[506], bl_bot[507], bl_bot[508],
     bl_bot[509], bl_bot[510], bl_bot[511], bl_bot[512], bl_bot[513],
     bl_bot[514], bl_bot[515], bl_bot[516], bl_bot[517], bl_bot[518],
     bl_bot[519], bl_bot[520], bl_bot[521], bl_bot[522], bl_bot[523],
     bl_bot[524], bl_bot[525], bl_bot[526], bl_bot[527], bl_bot[528],
     bl_bot[529], bl_bot[530], bl_bot[531], bl_bot[532], bl_bot[533],
     bl_bot[534], bl_bot[535], bl_bot[536], bl_bot[537], bl_bot[538],
     bl_bot[539], bl_bot[540], bl_bot[541], bl_bot[542], bl_bot[543],
     bl_bot[544], bl_bot[545], bl_bot[546], bl_bot[547], bl_bot[548],
     bl_bot[549], bl_bot[550], bl_bot[551], bl_bot[552], bl_bot[553],
     bl_bot[554], bl_bot[555], bl_bot[556], bl_bot[557], bl_bot[558],
     bl_bot[559], bl_bot[560], bl_bot[561], bl_bot[562], bl_bot[563],
     bl_bot[564], bl_bot[565], bl_bot[566], bl_bot[567], bl_bot[568],
     bl_bot[569], bl_bot[570], bl_bot[571], bl_bot[572], bl_bot[573],
     bl_bot[574], bl_bot[575], bl_bot[576], bl_bot[577], bl_bot[578],
     bl_bot[579], bl_bot[580], bl_bot[581], bl_bot[582], bl_bot[583],
     bl_bot[584], bl_bot[585], bl_bot[586], bl_bot[587], bl_bot[588],
     bl_bot[589], bl_bot[590], bl_bot[591], bl_bot[592], bl_bot[593],
     bl_bot[594], bl_bot[595], bl_bot[596], bl_bot[597], bl_bot[598],
     bl_bot[599], bl_bot[600], bl_bot[601], bl_bot[602], bl_bot[603],
     bl_bot[604], bl_bot[605], bl_bot[606], bl_bot[607], bl_bot[608],
     bl_bot[609], bl_bot[610], bl_bot[611], bl_bot[612], bl_bot[613],
     bl_bot[614], bl_bot[615], bl_bot[616], bl_bot[617], bl_bot[618],
     bl_bot[619], bl_bot[620], bl_bot[621], bl_bot[622], bl_bot[623],
     bl_bot[624], bl_bot[625], bl_bot[626], bl_bot[627], bl_bot[628],
     bl_bot[629], bl_bot[630], bl_bot[631], bl_bot[632], bl_bot[633],
     bl_bot[634], bl_bot[635], bl_bot[636], bl_bot[637], bl_bot[638],
     bl_bot[639], bl_bot[640], bl_bot[641], bl_bot[642], bl_bot[643],
     bl_bot[644], bl_bot[645], bl_bot[646], bl_bot[647], bl_bot[648],
     bl_bot[649], bl_bot[650], bl_bot[651], bl_bot[652], bl_bot[653],
     bl_bot[654], bl_bot[655], bl_bot[656], bl_bot[657], bl_bot[658],
     bl_bot[659], bl_bot[660], bl_bot[661], bl_bot[662], bl_bot[663],
     bl_bot[664], bl_bot[665], bl_bot[666], bl_bot[667], bl_bot[668],
     bl_bot[669], bl_bot[670], bl_bot[671], bl_bot[672], bl_bot[673],
     bl_bot[674], bl_bot[675], bl_bot[676], bl_bot[677], bl_bot[678],
     bl_bot[679], bl_bot[680], bl_bot[681], bl_bot[682], bl_bot[683],
     bl_bot[684], bl_bot[685], bl_bot[686], bl_bot[687], bl_bot[688],
     bl_bot[689], bl_bot[690], bl_bot[691], bl_bot[692], bl_bot[693],
     bl_bot[694], bl_bot[695], bl_bot[696], bl_bot[697], bl_bot[698],
     bl_bot[699], bl_bot[700], bl_bot[701], bl_bot[702], bl_bot[703],
     bl_bot[704], bl_bot[705], bl_bot[706], bl_bot[707], bl_bot[708],
     bl_bot[709], bl_bot[710], bl_bot[711], bl_bot[712], bl_bot[713],
     bl_bot[714], bl_bot[715], bl_bot[716], bl_bot[717], bl_bot[718],
     bl_bot[719], bl_bot[720], bl_bot[721], bl_bot[722], bl_bot[723],
     bl_bot[724], bl_bot[725], bl_bot[726], bl_bot[727], bl_bot[728],
     bl_bot[729], bl_bot[730], bl_bot[731], bl_bot[732], bl_bot[733],
     bl_bot[734], bl_bot[735], bl_bot[736], bl_bot[737], bl_bot[738],
     bl_bot[739], bl_bot[740], bl_bot[741], bl_bot[742], bl_bot[743],
     bl_bot[744], bl_bot[745], bl_bot[746], bl_bot[747], bl_bot[748],
     bl_bot[749], bl_bot[750], bl_bot[751], bl_bot[752], bl_bot[753],
     bl_bot[754], bl_bot[755], bl_bot[756], bl_bot[757], bl_bot[758],
     bl_bot[759], bl_bot[760], bl_bot[761], bl_bot[762], bl_bot[763],
     bl_bot[764], bl_bot[765], bl_bot[766], bl_bot[767], bl_bot[768],
     bl_bot[769], bl_bot[770], bl_bot[771], bl_bot[772], bl_bot[773],
     bl_bot[774], bl_bot[775], bl_bot[776], bl_bot[777], bl_bot[778],
     bl_bot[779], bl_bot[780], bl_bot[781], bl_bot[782], bl_bot[783],
     bl_bot[784], bl_bot[785], bl_bot[786], bl_bot[787], bl_bot[788],
     bl_bot[789], bl_bot[790], bl_bot[791], bl_bot[792], bl_bot[793],
     bl_bot[794], bl_bot[795], bl_bot[796], bl_bot[797], bl_bot[798],
     bl_bot[799], bl_bot[800], bl_bot[801], bl_bot[802], bl_bot[803],
     bl_bot[804], bl_bot[805], bl_bot[806], bl_bot[807], bl_bot[808],
     bl_bot[809], bl_bot[810], bl_bot[811], bl_bot[812], bl_bot[813],
     bl_bot[814], bl_bot[815], bl_bot[816], bl_bot[817], bl_bot[818],
     bl_bot[819], bl_bot[820], bl_bot[821], bl_bot[822], bl_bot[823],
     bl_bot[824], bl_bot[825], bl_bot[826], bl_bot[827], bl_bot[828],
     bl_bot[829], bl_bot[830], bl_bot[831], bl_bot[832], bl_bot[833],
     bl_bot[834], bl_bot[835], bl_bot[836], bl_bot[837], bl_bot[838],
     bl_bot[839], bl_bot[840], bl_bot[841], bl_bot[842], bl_bot[843],
     bl_bot[844], bl_bot[845], bl_bot[846], bl_bot[847], bl_bot[848],
     bl_bot[849], bl_bot[850], bl_bot[851], bl_bot[852], bl_bot[853],
     bl_bot[854], bl_bot[855], bl_bot[856], bl_bot[857], bl_bot[858],
     bl_bot[859], bl_bot[860], bl_bot[861], bl_bot[862], bl_bot[863],
     bl_bot[864], bl_bot[865], bl_bot[866], bl_bot[867], bl_bot[868],
     bl_bot[869], bl_bot[870], bl_bot[871]}),
     .smc_wdic_clk(smc_wdis_dclk_blbld), .smc_clk(cm_clk_blbld),
     .cm_sdi_u(cm_sdi_u0d1[1:0]), .latch_reset(core_por_rowu0),
     .cm_sdo_u(cm_sdo_u0[1:0]), .data_muxsel1(data_muxsel1_blbld),
     .data_muxsel(data_muxsel_blbld), .cram_write(cram_write_blbld),
     .cram_prec(cram_prec_blbld),
     .cor_en_8bpcfg_b(en_8bconfig_b_blbld),
     .cram_pullup_b(cram_pullup_blbld),
     .banksel(cm_banksel_blbld1_0_));
sg_bufx10bot I531_1_ ( .in(net0200[0]), .out(net0278[0]));
sg_bufx10bot I531_0_ ( .in(net0200[1]), .out(net0278[1]));
sg_bufx10bot I175 ( .in(net272), .out(data_muxsel_blbld));
sg_bufx10bot I333 ( .in(j_rst_b), .out(j_rst_bl0));
sg_bufx10bot I486 ( .in(net270), .out(cram_prec_blbld));
sg_bufx10bot I492 ( .in(net268), .out(cram_write_blbld));
sg_bufx10bot I474 ( .in(net302), .out(net312));
sg_bufx10bot I496 ( .in(en_8bconfig_b_blbrd),
     .out(predata_en_8bconfig_b));
sg_bufx10bot I481 ( .in(net318), .out(cram_rstl0));
sg_bufx10bot I495 ( .in(net264), .out(en_8bconfig_b_blbld));
sg_bufx10bot I467 ( .in(predata_muxsel1), .out(net260));
sg_bufx10bot I466 ( .in(net260), .out(data_muxsel1_blbld));
sg_bufx10bot I429_1_ ( .in(monitor_celld3[1]),
     .out(monitor_celld4[1]));
sg_bufx10bot I429_0_ ( .in(monitor_celld3[0]),
     .out(monitor_celld4[0]));
sg_bufx10bot I523 ( .in(smc_clk_mid), .out(cm_clk_blbld));
sg_bufx10bot I489 ( .in(net256), .out(cram_pullup_blbld));
sg_bufx10bot I485 ( .in(cram_prec), .out(predata_cram_prec));
sg_bufx10bot I487 ( .in(predata_cram_prec), .out(net270));
sg_bufx10bot I533_1_ ( .in(cm_sdi_u1[1]), .out(net0200[0]));
sg_bufx10bot I533_0_ ( .in(cm_sdi_u1[0]), .out(net0200[1]));
sg_bufx10bot I527_1_ ( .in(cm_sdi_u0[1]), .out(net0260[0]));
sg_bufx10bot I527_0_ ( .in(cm_sdi_u0[0]), .out(net0260[1]));
sg_bufx10bot I520 ( .in(net282), .out(net280));
sg_bufx10bot I517 ( .in(net250), .out(net206));
sg_bufx10bot I493 ( .in(predata_cram_write), .out(net268));
sg_bufx10bot I505 ( .in(net248), .out(smc_rsr_rstl0));
sg_bufx10bot I509 ( .in(net246), .out(row_testl1));
sg_bufx10bot I519 ( .in(cm_banksel[0]), .out(net282));
sg_bufx10bot I491 ( .in(cram_write), .out(predata_cram_write));
sg_bufx10bot I504 ( .in(smc_rsr_rst), .out(net298));
sg_bufx10bot I494 ( .in(predata_en_8bconfig_b), .out(net264));
sg_bufx10bot I529_1_ ( .in(net0254[0]), .out(cm_sdi_u0d1[1]));
sg_bufx10bot I529_0_ ( .in(net0254[1]), .out(cm_sdi_u0d1[0]));
sg_bufx10bot I476 ( .in(net236), .out(cram_vddoffl0));
sg_bufx10bot I479 ( .in(cram_rst), .out(net214));
sg_bufx10bot I530_1_ ( .in(net0260[0]), .out(net0254[0]));
sg_bufx10bot I530_0_ ( .in(net0260[1]), .out(net0254[1]));
sg_bufx10bot I439 ( .in(j_tck), .out(tck_padl0));
sg_bufx10bot I510 ( .in(net276), .out(net246));
sg_bufx10bot I482 ( .in(net228), .out(cram_pgateoffl0));
sg_bufx10bot I483 ( .in(net226), .out(net228));
sg_bufx10bot I464 ( .in(predata_muxsel), .out(net272));
sg_bufx10bot I525 ( .in(cm_clk_blbrd), .out(predata_smc_clk_out));
sg_bufx10bot I503 ( .in(net298), .out(net248));
sg_bufx10bot I490 ( .in(cram_pullup_b), .out(predata_cram_pullup_b));
sg_bufx10bot I532_1_ ( .in(net0278[0]), .out(cm_sdi_u1d[1]));
sg_bufx10bot I532_0_ ( .in(net0278[1]), .out(cm_sdi_u1d[0]));
sg_bufx10bot I521 ( .in(net280), .out(cm_banksel_blbld1_0_));
sg_bufx10bot I465 ( .in(data_muxsel1_blbrd), .out(predata_muxsel1));
sg_bufx10bot I484 ( .in(cram_pgateoff), .out(net226));
sg_bufx10bot I480 ( .in(net214), .out(net318));
sg_bufx10bot I518 ( .in(cm_banksel[1]), .out(net250));
sg_bufx10bot I488 ( .in(predata_cram_pullup_b), .out(net256));
sg_bufx10bot I524 ( .in(predata_smc_clk_out), .out(smc_clk_mid));
sg_bufx10bot I516 ( .in(net206), .out(cm_banksel_blbld_1_));
sg_bufx10bot I470 ( .in(net204), .out(cram_wl_enl0));
sg_bufx10bot I293 ( .in(last_rsr1), .out(last_rsr2));
sg_bufx10bot I541_1_ ( .in(dff_u0_d1[1]), .out(cm_sdo_u0d1[1]));
sg_bufx10bot I541_0_ ( .in(dff_u0_d1[0]), .out(cm_sdo_u0d1[0]));
sg_bufx10bot I539_1_ ( .in(cm_sdo_u1d1[1]), .out(cm_sdo_u1_buf[1]));
sg_bufx10bot I539_0_ ( .in(cm_sdo_u1d1[0]), .out(cm_sdo_u1_buf[0]));
sg_bufx10bot I455 ( .in(data_muxsel_blbrd), .out(predata_muxsel));
sg_bufx10bot I475 ( .in(net312), .out(smc_writel0));
sg_bufx10bot I526_1_ ( .in(cm_sdi_u2d[1]), .out(cm_sdi_u2d_buf[1]));
sg_bufx10bot I526_0_ ( .in(cm_sdi_u2d[0]), .out(cm_sdi_u2d_buf[0]));
sg_bufx10bot I459 ( .in(smc_row_inc), .out(net316));
sg_bufx10bot I477 ( .in(net292), .out(net236));
sg_bufx10bot I543_1_ ( .in(dff_u0_d0[1]), .out(cm_sdo_u0_buf[1]));
sg_bufx10bot I543_0_ ( .in(dff_u0_d0[0]), .out(cm_sdo_u0_buf[0]));
sg_bufx10bot I469 ( .in(net274), .out(smc_row_incl0));
sg_bufx10bot I522 ( .in(cm_banksel_blbrd_2_),
     .out(cm_banksel_blbrd1[2]));
sg_bufx10bot I427_1_ ( .in(monitor_celld2[1]),
     .out(monitor_celld3[1]));
sg_bufx10bot I427_0_ ( .in(monitor_celld2[0]),
     .out(monitor_celld3[0]));
sg_bufx10bot I540_1_ ( .in(dff_u1_d1[1]), .out(cm_sdo_u1d3[1]));
sg_bufx10bot I540_0_ ( .in(dff_u1_d1[0]), .out(cm_sdo_u1d3[0]));
sg_bufx10bot I473 ( .in(smc_write), .out(net302));
sg_bufx10bot I542 ( .in(net374), .out(last_rsr3));
sg_bufx10bot I497 ( .in(smc_wdis_dclk_blbrd),
     .out(predata_smc_wdis_dclk));
sg_bufx10bot I511 ( .in(row_test0), .out(net276));
sg_bufx10bot I498 ( .in(net324), .out(smc_wdis_dclk_blbld));
sg_bufx10bot I471 ( .in(net278), .out(net204));
sg_bufx10bot I499 ( .in(predata_smc_wdis_dclk), .out(net324));
sg_bufx10bot I330 ( .in(net316), .out(net274));
sg_bufx10bot I478 ( .in(cram_vddoff), .out(net292));
sg_bufx10bot I336 ( .in(core_por_bb), .out(core_por_bbl0));
sg_bufx10bot I472 ( .in(cram_wl_en), .out(net278));
creset_filter I141 ( .in(creset_b_int), .out(crst_filterout));
bram_bufferx16 I534 ( .in(smc_clk_mid), .out(net393));
bram_bufferx16 I550_1_ ( .in(dff_u2_d1[1]), .out(cm_sdo_u2d1[1]));
bram_bufferx16 I550_0_ ( .in(dff_u2_d1[0]), .out(cm_sdo_u2d1[0]));
bram_bufferx16 I549 ( .in(net400), .out(net401));
bram_bufferx16 I450_4_ ( .in(spi_ss_in_bbank[4]),
     .out(spi_ss_in_bbankd[4]));
bram_bufferx16 I450_3_ ( .in(spi_ss_in_bbank[3]),
     .out(spi_ss_in_bbankd[3]));
bram_bufferx16 I450_2_ ( .in(spi_ss_in_bbank[2]),
     .out(spi_ss_in_bbankd[2]));
bram_bufferx16 I450_1_ ( .in(spi_ss_in_bbank[1]),
     .out(spi_ss_in_bbankd[1]));
bram_bufferx16 I450_0_ ( .in(spi_ss_in_bbank[0]),
     .out(spi_ss_in_bbankd[0]));
bram_bufferx16 I548 ( .in(predata_smc_clk_out), .out(net400));
bram_bufferx16 I536 ( .in(cm_clk_blbld), .out(net395));
bram_bufferx16 I186 ( .in(core_por_b0), .out(core_por_b2));

endmodule
// Library - chip, Cell - CHIP_route_top10k, View - schematic
// LAST TIME SAVED: Oct  7 17:49:11 2008
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module CHIP_route_top10k ( cm_sdo_u1, cm_sdo_u3, bl_top,
     cm_banksel_bltld3, cm_banksel_bltrd1, cm_clk_bltld3,
     cm_clk_bltrd1, .cm_prec_bltld3(cram_prec_bltld3), cm_sdi_u1d3,
     cm_sdi_u3d2, core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3,
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1) );


input  cm_clk_bltld3, cm_clk_bltrd1, cram_prec_bltld3,
     core_por_b_rowu1, core_por_b_rowu3, cram_prec_bltrd1,
     cram_pullup_b_bltrd1, cram_pullup_bltld3, cram_write_bltld3,
     cram_write_bltrd1, data_muxsel1_bltld3, data_muxsel1_bltrd1,
     data_muxsel_bltld3, data_muxsel_bltrd1, en_8bconfig_b_bltld3,
     en_8bconfig_b_bltrd1, smc_wdis_dclk_bltld3, smc_wdis_dclk_bltrd1;

output [1:0]  cm_sdo_u1;
output [1:0]  cm_sdo_u3;

inout [1743:0]  bl_top;

input [1:0]  cm_sdi_u1d3;
input [1:0]  cm_sdi_u3d2;
input [3:3]  cm_banksel_bltrd1;
input [1:1]  cm_banksel_bltld3;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_blsa_bank10k Ibltr ( .bl(bl_top[1743:872]),
     .smc_wdic_clk(smc_wdis_dclk_bltrd1), .smc_clk(cm_clk_bltrd1),
     .cm_sdi_u(cm_sdi_u3d2[1:0]), .latch_reset(core_por_b_rowu3),
     .cm_sdo_u(cm_sdo_u3[1:0]), .data_muxsel1(data_muxsel1_bltrd1),
     .data_muxsel(data_muxsel_bltrd1), .cram_write(cram_write_bltrd1),
     .cram_prec(cram_prec_bltrd1),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltrd1),
     .cram_pullup_b(cram_pullup_b_bltrd1),
     .banksel(cm_banksel_bltrd1[3]));
ml_blsa_bank10k Ibltlu1 ( .bl({bl_top[0], bl_top[1], bl_top[2],
     bl_top[3], bl_top[4], bl_top[5], bl_top[6], bl_top[7], bl_top[8],
     bl_top[9], bl_top[10], bl_top[11], bl_top[12], bl_top[13],
     bl_top[14], bl_top[15], bl_top[16], bl_top[17], bl_top[18],
     bl_top[19], bl_top[20], bl_top[21], bl_top[22], bl_top[23],
     bl_top[24], bl_top[25], bl_top[26], bl_top[27], bl_top[28],
     bl_top[29], bl_top[30], bl_top[31], bl_top[32], bl_top[33],
     bl_top[34], bl_top[35], bl_top[36], bl_top[37], bl_top[38],
     bl_top[39], bl_top[40], bl_top[41], bl_top[42], bl_top[43],
     bl_top[44], bl_top[45], bl_top[46], bl_top[47], bl_top[48],
     bl_top[49], bl_top[50], bl_top[51], bl_top[52], bl_top[53],
     bl_top[54], bl_top[55], bl_top[56], bl_top[57], bl_top[58],
     bl_top[59], bl_top[60], bl_top[61], bl_top[62], bl_top[63],
     bl_top[64], bl_top[65], bl_top[66], bl_top[67], bl_top[68],
     bl_top[69], bl_top[70], bl_top[71], bl_top[72], bl_top[73],
     bl_top[74], bl_top[75], bl_top[76], bl_top[77], bl_top[78],
     bl_top[79], bl_top[80], bl_top[81], bl_top[82], bl_top[83],
     bl_top[84], bl_top[85], bl_top[86], bl_top[87], bl_top[88],
     bl_top[89], bl_top[90], bl_top[91], bl_top[92], bl_top[93],
     bl_top[94], bl_top[95], bl_top[96], bl_top[97], bl_top[98],
     bl_top[99], bl_top[100], bl_top[101], bl_top[102], bl_top[103],
     bl_top[104], bl_top[105], bl_top[106], bl_top[107], bl_top[108],
     bl_top[109], bl_top[110], bl_top[111], bl_top[112], bl_top[113],
     bl_top[114], bl_top[115], bl_top[116], bl_top[117], bl_top[118],
     bl_top[119], bl_top[120], bl_top[121], bl_top[122], bl_top[123],
     bl_top[124], bl_top[125], bl_top[126], bl_top[127], bl_top[128],
     bl_top[129], bl_top[130], bl_top[131], bl_top[132], bl_top[133],
     bl_top[134], bl_top[135], bl_top[136], bl_top[137], bl_top[138],
     bl_top[139], bl_top[140], bl_top[141], bl_top[142], bl_top[143],
     bl_top[144], bl_top[145], bl_top[146], bl_top[147], bl_top[148],
     bl_top[149], bl_top[150], bl_top[151], bl_top[152], bl_top[153],
     bl_top[154], bl_top[155], bl_top[156], bl_top[157], bl_top[158],
     bl_top[159], bl_top[160], bl_top[161], bl_top[162], bl_top[163],
     bl_top[164], bl_top[165], bl_top[166], bl_top[167], bl_top[168],
     bl_top[169], bl_top[170], bl_top[171], bl_top[172], bl_top[173],
     bl_top[174], bl_top[175], bl_top[176], bl_top[177], bl_top[178],
     bl_top[179], bl_top[180], bl_top[181], bl_top[182], bl_top[183],
     bl_top[184], bl_top[185], bl_top[186], bl_top[187], bl_top[188],
     bl_top[189], bl_top[190], bl_top[191], bl_top[192], bl_top[193],
     bl_top[194], bl_top[195], bl_top[196], bl_top[197], bl_top[198],
     bl_top[199], bl_top[200], bl_top[201], bl_top[202], bl_top[203],
     bl_top[204], bl_top[205], bl_top[206], bl_top[207], bl_top[208],
     bl_top[209], bl_top[210], bl_top[211], bl_top[212], bl_top[213],
     bl_top[214], bl_top[215], bl_top[216], bl_top[217], bl_top[218],
     bl_top[219], bl_top[220], bl_top[221], bl_top[222], bl_top[223],
     bl_top[224], bl_top[225], bl_top[226], bl_top[227], bl_top[228],
     bl_top[229], bl_top[230], bl_top[231], bl_top[232], bl_top[233],
     bl_top[234], bl_top[235], bl_top[236], bl_top[237], bl_top[238],
     bl_top[239], bl_top[240], bl_top[241], bl_top[242], bl_top[243],
     bl_top[244], bl_top[245], bl_top[246], bl_top[247], bl_top[248],
     bl_top[249], bl_top[250], bl_top[251], bl_top[252], bl_top[253],
     bl_top[254], bl_top[255], bl_top[256], bl_top[257], bl_top[258],
     bl_top[259], bl_top[260], bl_top[261], bl_top[262], bl_top[263],
     bl_top[264], bl_top[265], bl_top[266], bl_top[267], bl_top[268],
     bl_top[269], bl_top[270], bl_top[271], bl_top[272], bl_top[273],
     bl_top[274], bl_top[275], bl_top[276], bl_top[277], bl_top[278],
     bl_top[279], bl_top[280], bl_top[281], bl_top[282], bl_top[283],
     bl_top[284], bl_top[285], bl_top[286], bl_top[287], bl_top[288],
     bl_top[289], bl_top[290], bl_top[291], bl_top[292], bl_top[293],
     bl_top[294], bl_top[295], bl_top[296], bl_top[297], bl_top[298],
     bl_top[299], bl_top[300], bl_top[301], bl_top[302], bl_top[303],
     bl_top[304], bl_top[305], bl_top[306], bl_top[307], bl_top[308],
     bl_top[309], bl_top[310], bl_top[311], bl_top[312], bl_top[313],
     bl_top[314], bl_top[315], bl_top[316], bl_top[317], bl_top[318],
     bl_top[319], bl_top[320], bl_top[321], bl_top[322], bl_top[323],
     bl_top[324], bl_top[325], bl_top[326], bl_top[327], bl_top[328],
     bl_top[329], bl_top[330], bl_top[331], bl_top[332], bl_top[333],
     bl_top[334], bl_top[335], bl_top[336], bl_top[337], bl_top[338],
     bl_top[339], bl_top[340], bl_top[341], bl_top[342], bl_top[343],
     bl_top[344], bl_top[345], bl_top[346], bl_top[347], bl_top[348],
     bl_top[349], bl_top[350], bl_top[351], bl_top[352], bl_top[353],
     bl_top[354], bl_top[355], bl_top[356], bl_top[357], bl_top[358],
     bl_top[359], bl_top[360], bl_top[361], bl_top[362], bl_top[363],
     bl_top[364], bl_top[365], bl_top[366], bl_top[367], bl_top[368],
     bl_top[369], bl_top[370], bl_top[371], bl_top[372], bl_top[373],
     bl_top[374], bl_top[375], bl_top[376], bl_top[377], bl_top[378],
     bl_top[379], bl_top[380], bl_top[381], bl_top[382], bl_top[383],
     bl_top[384], bl_top[385], bl_top[386], bl_top[387], bl_top[388],
     bl_top[389], bl_top[390], bl_top[391], bl_top[392], bl_top[393],
     bl_top[394], bl_top[395], bl_top[396], bl_top[397], bl_top[398],
     bl_top[399], bl_top[400], bl_top[401], bl_top[402], bl_top[403],
     bl_top[404], bl_top[405], bl_top[406], bl_top[407], bl_top[408],
     bl_top[409], bl_top[410], bl_top[411], bl_top[412], bl_top[413],
     bl_top[414], bl_top[415], bl_top[416], bl_top[417], bl_top[418],
     bl_top[419], bl_top[420], bl_top[421], bl_top[422], bl_top[423],
     bl_top[424], bl_top[425], bl_top[426], bl_top[427], bl_top[428],
     bl_top[429], bl_top[430], bl_top[431], bl_top[432], bl_top[433],
     bl_top[434], bl_top[435], bl_top[436], bl_top[437], bl_top[438],
     bl_top[439], bl_top[440], bl_top[441], bl_top[442], bl_top[443],
     bl_top[444], bl_top[445], bl_top[446], bl_top[447], bl_top[448],
     bl_top[449], bl_top[450], bl_top[451], bl_top[452], bl_top[453],
     bl_top[454], bl_top[455], bl_top[456], bl_top[457], bl_top[458],
     bl_top[459], bl_top[460], bl_top[461], bl_top[462], bl_top[463],
     bl_top[464], bl_top[465], bl_top[466], bl_top[467], bl_top[468],
     bl_top[469], bl_top[470], bl_top[471], bl_top[472], bl_top[473],
     bl_top[474], bl_top[475], bl_top[476], bl_top[477], bl_top[478],
     bl_top[479], bl_top[480], bl_top[481], bl_top[482], bl_top[483],
     bl_top[484], bl_top[485], bl_top[486], bl_top[487], bl_top[488],
     bl_top[489], bl_top[490], bl_top[491], bl_top[492], bl_top[493],
     bl_top[494], bl_top[495], bl_top[496], bl_top[497], bl_top[498],
     bl_top[499], bl_top[500], bl_top[501], bl_top[502], bl_top[503],
     bl_top[504], bl_top[505], bl_top[506], bl_top[507], bl_top[508],
     bl_top[509], bl_top[510], bl_top[511], bl_top[512], bl_top[513],
     bl_top[514], bl_top[515], bl_top[516], bl_top[517], bl_top[518],
     bl_top[519], bl_top[520], bl_top[521], bl_top[522], bl_top[523],
     bl_top[524], bl_top[525], bl_top[526], bl_top[527], bl_top[528],
     bl_top[529], bl_top[530], bl_top[531], bl_top[532], bl_top[533],
     bl_top[534], bl_top[535], bl_top[536], bl_top[537], bl_top[538],
     bl_top[539], bl_top[540], bl_top[541], bl_top[542], bl_top[543],
     bl_top[544], bl_top[545], bl_top[546], bl_top[547], bl_top[548],
     bl_top[549], bl_top[550], bl_top[551], bl_top[552], bl_top[553],
     bl_top[554], bl_top[555], bl_top[556], bl_top[557], bl_top[558],
     bl_top[559], bl_top[560], bl_top[561], bl_top[562], bl_top[563],
     bl_top[564], bl_top[565], bl_top[566], bl_top[567], bl_top[568],
     bl_top[569], bl_top[570], bl_top[571], bl_top[572], bl_top[573],
     bl_top[574], bl_top[575], bl_top[576], bl_top[577], bl_top[578],
     bl_top[579], bl_top[580], bl_top[581], bl_top[582], bl_top[583],
     bl_top[584], bl_top[585], bl_top[586], bl_top[587], bl_top[588],
     bl_top[589], bl_top[590], bl_top[591], bl_top[592], bl_top[593],
     bl_top[594], bl_top[595], bl_top[596], bl_top[597], bl_top[598],
     bl_top[599], bl_top[600], bl_top[601], bl_top[602], bl_top[603],
     bl_top[604], bl_top[605], bl_top[606], bl_top[607], bl_top[608],
     bl_top[609], bl_top[610], bl_top[611], bl_top[612], bl_top[613],
     bl_top[614], bl_top[615], bl_top[616], bl_top[617], bl_top[618],
     bl_top[619], bl_top[620], bl_top[621], bl_top[622], bl_top[623],
     bl_top[624], bl_top[625], bl_top[626], bl_top[627], bl_top[628],
     bl_top[629], bl_top[630], bl_top[631], bl_top[632], bl_top[633],
     bl_top[634], bl_top[635], bl_top[636], bl_top[637], bl_top[638],
     bl_top[639], bl_top[640], bl_top[641], bl_top[642], bl_top[643],
     bl_top[644], bl_top[645], bl_top[646], bl_top[647], bl_top[648],
     bl_top[649], bl_top[650], bl_top[651], bl_top[652], bl_top[653],
     bl_top[654], bl_top[655], bl_top[656], bl_top[657], bl_top[658],
     bl_top[659], bl_top[660], bl_top[661], bl_top[662], bl_top[663],
     bl_top[664], bl_top[665], bl_top[666], bl_top[667], bl_top[668],
     bl_top[669], bl_top[670], bl_top[671], bl_top[672], bl_top[673],
     bl_top[674], bl_top[675], bl_top[676], bl_top[677], bl_top[678],
     bl_top[679], bl_top[680], bl_top[681], bl_top[682], bl_top[683],
     bl_top[684], bl_top[685], bl_top[686], bl_top[687], bl_top[688],
     bl_top[689], bl_top[690], bl_top[691], bl_top[692], bl_top[693],
     bl_top[694], bl_top[695], bl_top[696], bl_top[697], bl_top[698],
     bl_top[699], bl_top[700], bl_top[701], bl_top[702], bl_top[703],
     bl_top[704], bl_top[705], bl_top[706], bl_top[707], bl_top[708],
     bl_top[709], bl_top[710], bl_top[711], bl_top[712], bl_top[713],
     bl_top[714], bl_top[715], bl_top[716], bl_top[717], bl_top[718],
     bl_top[719], bl_top[720], bl_top[721], bl_top[722], bl_top[723],
     bl_top[724], bl_top[725], bl_top[726], bl_top[727], bl_top[728],
     bl_top[729], bl_top[730], bl_top[731], bl_top[732], bl_top[733],
     bl_top[734], bl_top[735], bl_top[736], bl_top[737], bl_top[738],
     bl_top[739], bl_top[740], bl_top[741], bl_top[742], bl_top[743],
     bl_top[744], bl_top[745], bl_top[746], bl_top[747], bl_top[748],
     bl_top[749], bl_top[750], bl_top[751], bl_top[752], bl_top[753],
     bl_top[754], bl_top[755], bl_top[756], bl_top[757], bl_top[758],
     bl_top[759], bl_top[760], bl_top[761], bl_top[762], bl_top[763],
     bl_top[764], bl_top[765], bl_top[766], bl_top[767], bl_top[768],
     bl_top[769], bl_top[770], bl_top[771], bl_top[772], bl_top[773],
     bl_top[774], bl_top[775], bl_top[776], bl_top[777], bl_top[778],
     bl_top[779], bl_top[780], bl_top[781], bl_top[782], bl_top[783],
     bl_top[784], bl_top[785], bl_top[786], bl_top[787], bl_top[788],
     bl_top[789], bl_top[790], bl_top[791], bl_top[792], bl_top[793],
     bl_top[794], bl_top[795], bl_top[796], bl_top[797], bl_top[798],
     bl_top[799], bl_top[800], bl_top[801], bl_top[802], bl_top[803],
     bl_top[804], bl_top[805], bl_top[806], bl_top[807], bl_top[808],
     bl_top[809], bl_top[810], bl_top[811], bl_top[812], bl_top[813],
     bl_top[814], bl_top[815], bl_top[816], bl_top[817], bl_top[818],
     bl_top[819], bl_top[820], bl_top[821], bl_top[822], bl_top[823],
     bl_top[824], bl_top[825], bl_top[826], bl_top[827], bl_top[828],
     bl_top[829], bl_top[830], bl_top[831], bl_top[832], bl_top[833],
     bl_top[834], bl_top[835], bl_top[836], bl_top[837], bl_top[838],
     bl_top[839], bl_top[840], bl_top[841], bl_top[842], bl_top[843],
     bl_top[844], bl_top[845], bl_top[846], bl_top[847], bl_top[848],
     bl_top[849], bl_top[850], bl_top[851], bl_top[852], bl_top[853],
     bl_top[854], bl_top[855], bl_top[856], bl_top[857], bl_top[858],
     bl_top[859], bl_top[860], bl_top[861], bl_top[862], bl_top[863],
     bl_top[864], bl_top[865], bl_top[866], bl_top[867], bl_top[868],
     bl_top[869], bl_top[870], bl_top[871]}),
     .smc_wdic_clk(smc_wdis_dclk_bltld3), .smc_clk(cm_clk_bltld3),
     .cm_sdi_u(cm_sdi_u1d3[1:0]), .latch_reset(core_por_b_rowu1),
     .cm_sdo_u(cm_sdo_u1[1:0]), .data_muxsel1(data_muxsel1_bltld3),
     .data_muxsel(data_muxsel_bltld3), .cram_write(cram_write_bltld3),
     .cram_prec(cram_prec_bltld3),
     .cor_en_8bpcfg_b(en_8bconfig_b_bltld3),
     .cram_pullup_b(cram_pullup_bltld3),
     .banksel(cm_banksel_bltld3[1]));

endmodule
// Library - io, Cell - PRCUTSSTLSTDR, View - schematic
// LAST TIME SAVED: Oct 24 13:01:45 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PRCUTSSTLSTDR ( VSS, VSSPST );
input  VSS, VSSPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - PRCUTSSTLSTDL, View - schematic
// LAST TIME SAVED: Oct 24 13:01:45 2007
// NETLIST TIME: Nov 14 16:17:13 2008
`timescale 1ns / 1ns 

module PRCUTSSTLSTDL ( VSS, VSSPST );
input  VSS, VSSPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - chip, Cell - ring_route8k_f, View - schematic
// LAST TIME SAVED: Oct  7 17:54:08 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module ring_route8k_f ( bm_banksel_i, bm_init_i, bm_rcapmux_en_i,
     bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bs_en0, ceb0, en_8bconfig_b, end_of_startup,
     gint_hz, gsr, hiz_b0, in_bbank, in_lbank, in_rbank, in_tbank,
     j_tck, j_tdi, jtag_rowtest_mode_rowu0_b,
     jtag_rowtest_mode_rowu1_b, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr, md_spi_b, mode0, pgate_l,
     pgate_r, psdo, reset_l, reset_r, shift0, spi_clk_out, spi_sdo,
     spi_sdo_oe_b, spi_ss_out_b, tdo, update0, vdd_cntl_l, vdd_cntl_r,
     wl_l, wl_r, bl_bot, bl_top, cdone, uio_bbank, uio_lbank,
     uio_rbank, uio_tbank, vpp, VREFSSTL, bm_sdo_o, cf_bbank, cf_lbank,
     cf_r_ext, cf_rbank, cf_tbank, creset_b, fabric_out_32_00,
     fabric_out_33_01, fabric_out_33_02, fromsdo, oen_bbank, oen_lbank,
     oen_rbank, oen_tbank, out_bbank, out_lbank, out_rbank, out_tbank,
     spi_ss_in_bbank, spi_ss_in_r, tck, tdi, tiegnd, tievdd, tms, trstb
     );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, ceb0, en_8bconfig_b,
     end_of_startup, gint_hz, gsr, hiz_b0, j_tck, j_tdi,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b,
     jtag_rowtest_mode_rowu2_b, jtag_rowtest_mode_rowu3_b, md_spi_b,
     mode0, shift0, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out_b,
     tdo, update0;

inout  cdone, vpp;

input  VREFSSTL, creset_b, fabric_out_32_00, fabric_out_33_01,
     fabric_out_33_02, fromsdo, tck, tdi, tiegnd, tievdd, tms, trstb;

output [7:0]  bm_sa_i;
output [543:0]  vdd_cntl_r;
output [3:0]  bm_banksel_i;
output [543:0]  wl_r;
output [54:0]  in_rbank;
output [543:0]  pgate_r;
output [543:0]  reset_r;
output [7:1]  psdo;
output [3:0]  bm_sdi_i;
output [543:0]  pgate_l;
output [56:0]  in_bbank;
output [59:0]  in_tbank;
output [3:0]  last_rsr;
output [543:0]  reset_l;
output [543:0]  vdd_cntl_l;
output [49:0]  in_lbank;
output [543:0]  wl_l;

inout [49:0]  uio_lbank;
inout [56:0]  uio_bbank;
inout [59:0]  uio_tbank;
inout [1743:0]  bl_bot;
inout [54:0]  uio_rbank;
inout [1743:0]  bl_top;

input [59:0]  cf_tbank;
input [3:0]  bm_sdo_o;
input [54:0]  out_rbank;
input [7:1]  spi_ss_in_r;
input [59:0]  out_tbank;
input [54:0]  cf_rbank;
input [54:0]  oen_rbank;
input [1:0]  cf_r_ext;
input [61:56]  spi_ss_in_bbank;
input [56:0]  oen_bbank;
input [56:0]  cf_bbank;
input [59:0]  oen_tbank;
input [56:0]  out_bbank;
input [49:0]  out_lbank;
input [49:0]  oen_lbank;
input [376:0]  cf_lbank;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  cm_sdo_u3;

wire  [3:3]  cm_banksel_bltrd1;

wire  [1:0]  cm_sdi_u3d2;

wire  [2:2]  cm_banksel_blbrd;

wire  [1:0]  cm_sdo_u1;

wire  [1:0]  cm_sdi_u1d3;

wire  [1:0]  monitor_celld2;

wire  [1:0]  cm_sdi_u1d;

wire  [1:0]  cm_sdi_u1;

wire  [1:0]  cm_sdi_u0;

wire  [1:0]  cm_sdi_u2d;

wire  [1:0]  cm_banksel;

wire  [1:1]  cm_banksel_bltld3;

wire  [1:0]  cm_sdo_u0d1;

wire  [1:0]  cm_sdo_u1d3;

wire  [1:1]  cm_banksel_blbld;

wire  [1:0]  cm_sdo_u2d1;

wire  [0:0]  cm_banksel_blbld1;

wire  [1:0]  cm_sdo_u1d1;

wire  [42:47]  spi_ss_in_bbankd;

wire  [1:0]  monitor_celld4;



rgtbank_f Iright_bank ( .tdi_int(tdi_pad), .tck_int(tck_pad),
     .tms_int(tms_pad), .tdo_int(totdopad), .tdo_en(sdo_enable),
     .trstb_int(trst_pad), .pad(uio_rbank[54:0]),
     .oen(oen_rbank[54:0]), .out(out_rbank[54:0]), .in(in_rbank[54:0]),
     .ren(cf_rbank[54:0]), .Tdo(tdo), .TRSTb(trstb), .Tdi(tdi),
     .Tms(tms), .Tck(tck));
topbank_f Iio_topcell ( .vppin(vppin), .vpp(vpp),
     .out(out_tbank[59:0]), .oen(oen_tbank[59:0]),
     .ren(cf_tbank[59:0]), .in(in_tbank[59:0]), .pad(uio_tbank[59:0]));
sg_bufx10 I465 ( .in(spi_clk_out), .out(spi_clk_out2fsm));
CHIP_route_right_ice8f Ismc_chip_rout_right (
     .idcode_msb20bits({tiegnd, tiegnd, tiegnd, tievdd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tievdd, tiegnd, tiegnd, tiegnd}),
     .pgate_r(pgate_r[543:0]), .reset_b_r(reset_r[543:0]),
     .vdd_cntl_r(vdd_cntl_r[543:0]), .wl_r(wl_r[543:0]),
     .fabric_out_33_01(fabric_out_33_01),
     .fabric_out_32_00(fabric_out_32_00),
     .fabric_out_33_02(fabric_out_33_02), .nvcm_spi_sdo(nvcm_spi_sdo),
     .bp0(bp0), .nvcm_boot(nvcm_boot), .nvcm_rdy(nvcm_rdy),
     .nvcm_relextspi(nvcm_relextspi),
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b), .rst_b(rst_b_4smc2nvcm),
     .nvcm_spi_ss_b(nvcm_spi_ss_b), .nvcm_spi_sdi(nvcm_spi_sdi),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .ceb0(ceb0),
     .en_8bconfig_b(en_8bconfig_b), .spi_ss_in_r(spi_ss_in_r[7:1]),
     .smc_write0(smc_write), .cm_banksel_bldld(cm_banksel[1:0]),
     .cm_banksel_bltrd1_3_(cm_banksel_bltrd1[3]),
     .cm_banksel_blbrd_2_(cm_banksel_blbrd[2]),
     .last_rsr(last_rsr[3:2]), .spi_ss_in_bbank({spi_ss_in_bbankd[47],
     spi_ss_in_bbankd[46], spi_ss_in_bbankd[45], spi_ss_in_bbankd[43],
     spi_ss_in_bbankd[42]}), .cf_r(cf_r_ext[1:0]),
     .core_por_b_rowu2(core_por_b_rowu2), .core_por_b0(core_por_b0),
     .row_test0(row_test0), .smc_row_inc(smc_row_inc),
     .cram_pgateoff(cram_pgateoff), .core_por_bb(core_por_bb),
     .cram_wl_en(cram_wl_en), .cram_vddoff(cram_vddoff),
     .cram_rst(cram_rst), .smc_rsr_rst(smc_rsr_rst), .j_rst_b(j_rst_b),
     .smc_wdis_dclk_bltrd1(smc_wdis_dclk_bltrd1),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .cm_clk_blbrd(cm_clk_blbrd),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .cram_write(cram_write), .cram_prec(cram_prec),
     .cram_pullup_b(cram_pullup_b), .last_rsr3(last_rsr3),
     .core_por_b_rowu3(core_por_b_rowu3),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .cm_sdo_u3(cm_sdo_u3[1:0]), .vddio_rightbank(vddp_),
     .trst_pad(trst_pad), .tms_pad(tms_pad), .tdi_pad(tdi_pad),
     .tck_pad(tck_pad), .monitor_celld4(monitor_celld4[1:0]),
     .fromsdo(fromsdo), .crst_filterout(crst_filterout),
     .cm_sdo_u2d1(cm_sdo_u2d1[1:0]), .cm_sdo_u1d3(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0d1(cm_sdo_u0d1[1:0]), .cdone_in(cdone_in),
     .bm_sdo_o(bm_sdo_o[3:0]), .update0(update0), .totdopad(totdopad),
     .spi_ss_out_b(spi_ss_out_b), .spi_sdo_oe_b(spi_sdo_oe_b),
     .spi_sdo(spi_sdo), .spi_clk_out(spi_clk_out), .shift0(shift0),
     .sdo_enable(sdo_enable), .psdo(psdo[7:1]), .mode0(mode0),
     .md_spi_b(md_spi_b),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .j_tdi(j_tdi), .j_tck(j_tck), .hiz_b0(hiz_b0), .gsr(gsr),
     .gint_hz(gint_hz), .end_of_startup(end_of_startup),
     .en_8bcibfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel1_bltrd1(data_muxsel1_bltrd1),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1), .core_por_b1(core_por_b1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .cm_sdi_u1(cm_sdi_u1[1:0]), .cm_sdi_u0(cm_sdi_u0[1:0]),
     .cm_clk_bltrd1(cm_clk_bltrd1), .cdone_out(cdone_out),
     .bs_en0(bs_en0), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sweb_i(bm_sweb_i), .bm_sreb_i(bm_sreb_i),
     .bm_sdi_i(bm_sdi_i[3:0]), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bm_banksel_i(bm_banksel_i[3:0]),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b));
nvcm_ml_block I464 ( .spi_ss_b(nvcm_spi_ss_b), .spi_sdi(nvcm_spi_sdi),
     .rst_b(rst_b_4smc2nvcm), .nvcm_ce_b(end_of_startup),
     .icef_member_sel({tievdd, tiegnd}), .clk(spi_clk_out2fsm),
     .spi_sdo_oe_b(nvcm_spi_sdo_oe_b), .spi_sdo(nvcm_spi_sdo),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream),
     .fsm_tm_margin0_read(net269), .fsm_recall(net270), .bp0(bp0),
     .nvcm_relextspi(nvcm_relextspi), .vpp(vppin));
lefbank_rev Iio_lftcell ( .oen(oen_lbank[49:0]), .out(out_lbank[49:0]),
     .in(in_lbank[49:0]), .pad(uio_lbank[49:0]),
     .cbit(cf_lbank[374:0]), .VREFSSTL(VREFSSTL));
botbank Iio_botcell ( .oen(oen_bbank[56:0]), .ren(cf_bbank[56:0]),
     .cdone_int(cdone_in), .pad(uio_bbank[56:0]), .in(in_bbank[56:0]),
     .out(out_bbank[56:0]), .cdone_out(cdone_out), .done(cdone),
     .ctst_b(creset_b), .ctst_b_int(creset_b_int));
CHIP_route_left10k Ichip_route_left ( cm_banksel_bltld3[1],
     cm_clk_bltld3, cm_sdi_u1d3[1:0], cm_sdo_u1d1[1:0],
     core_por_b_rowu0, core_por_b_rowu1, cram_prec_bltld3,
     cram_pullup_b_bltld3, cram_write_bltld3, data_muxsel1_bltld3,
     data_muxsel_bltld3, en_8bconfig_b_bltld3,
     jtag_rowtest_mode_rowu0_b, jtag_rowtest_mode_rowu1_b, last_rsr0,
     last_rsr[1:0], monitor_celld2[1:0], pgate_l[543:0],
     reset_l[543:0], smc_wdis_dclk_bltld3r, vdd_cntl_l[543:0],
     wl_l[543:0], cf_lbank[375], cf_lbank[376], cm_banksel_blbld1[0],
     cm_banksel_blbld[1], cm_clk_blbld, cm_sdi_u1d[1:0],
     cm_sdo_u1[1:0], core_por_bbl0, cram_pgateoffl0, cram_prec_blbld,
     cram_pullup_blbld, cram_rstl0, cram_vddoffl0, cram_wl_enl0,
     cram_write_blbld, data_muxsel1_blbld, data_muxsel_blbld,
     en_8bconfig_b_blbld, j_rst_bl0, row_testl1, smc_row_incl0,
     smc_rsr_rstl0, smc_wdis_dclk_blbld, smc_writel0, tck_padl0);
CHIP_route_bot10k Ichip_route_bot (
     .cm_banksel_blbrd_2_(cm_banksel_blbrd[2]),
     .bl_bot(bl_bot[1743:0]),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2),
     .vddio_spi(vddio_spi), .vddio_botbank(vddio_bottombank),
     .cm_banksel_blbld1_0_(cm_banksel_blbld1[0]),
     .cm_banksel_blbld_1_(cm_banksel_blbld[1]), .j_rst_b(j_rst_b),
     .spi_ss_in_bbankd({spi_ss_in_bbankd[47], spi_ss_in_bbankd[46],
     spi_ss_in_bbankd[45], spi_ss_in_bbankd[43],
     spi_ss_in_bbankd[42]}), .spi_ss_in_bbank({spi_ss_in_bbank[61],
     spi_ss_in_bbank[60], spi_ss_in_bbank[59], spi_ss_in_bbank[57],
     spi_ss_in_bbank[56]}), .cm_banksel(cm_banksel[1:0]),
     .monitor_celld2(monitor_celld2[1:0]),
     .data_muxsel1_blbld(data_muxsel1_blbld),
     .data_muxsel_blbld(data_muxsel_blbld),
     .smc_wdis_dclk_blbld(smc_wdis_dclk_blbld),
     .en_8bconfig_b_blbld(en_8bconfig_b_blbld),
     .cram_write_blbld(cram_write_blbld),
     .cram_pullup_blbld(cram_pullup_blbld),
     .cram_prec_blbld(cram_prec_blbld), .cm_clk_blbld(cm_clk_blbld),
     .cram_pullup_b(cram_pullup_b), .cram_write(cram_write),
     .cm_sdi_u2d(cm_sdi_u2d[1:0]),
     .data_muxsel1_blbrd(data_muxsel1_blbrd),
     .data_muxsel_blbrd(data_muxsel_blbrd),
     .en_8bconfig_b_blbrd(en_8bconfig_b_blbrd),
     .smc_wdis_dclk_blbrd(smc_wdis_dclk_blbrd),
     .cm_clk_blbrd(cm_clk_blbrd), .smc_write(smc_write),
     .smc_rsr_rst(smc_rsr_rst), .smc_row_inc(smc_row_inc),
     .row_test0(row_test0), .last_rsr1(last_rsr0), .j_tck(j_tck),
     .creset_b_int(creset_b_int), .cram_wl_en(cram_wl_en),
     .cram_vddoff(cram_vddoff), .cram_rst(cram_rst),
     .cram_prec(cram_prec), .cram_pgateoff(cram_pgateoff),
     .core_por_rowu0(core_por_b_rowu0), .core_por_bb(core_por_bb),
     .core_por_b_rowu2(core_por_b_rowu2), .core_por_b0(core_por_b0),
     .cm_sdo_u1d1(cm_sdo_u1d1[1:0]), .cm_sdi_u1(cm_sdi_u1[1:0]),
     .cm_sdi_u0(cm_sdi_u0[1:0]), .tck_padl0(tck_padl0),
     .smc_writel0(smc_writel0), .smc_rsr_rstl0(smc_rsr_rstl0),
     .smc_row_incl0(smc_row_incl0), .row_testl1(row_testl1),
     .monitor_celld4(monitor_celld4[1:0]), .last_rsr3(last_rsr3),
     .j_rst_bl0(j_rst_bl0), .crst_filterout(crst_filterout),
     .cram_wl_enl0(cram_wl_enl0), .cram_vddoffl0(cram_vddoffl0),
     .cram_rstl0(cram_rstl0), .cram_pgateoffl0(cram_pgateoffl0),
     .core_por_bbl0(core_por_bbl0), .core_por_b2(core_por_b2),
     .cm_sdo_u2d1(cm_sdo_u2d1[1:0]), .cm_sdo_u1d3(cm_sdo_u1d3[1:0]),
     .cm_sdo_u0d1(cm_sdo_u0d1[1:0]), .cm_sdi_u1d(cm_sdi_u1d[1:0]));
CHIP_route_top10k Ichip_route_top ( .bl_top(bl_top[1743:0]),
     .data_muxsel1_bltrd1(data_muxsel1_bltrd1),
     .smc_wdis_dclk_bltrd1r(smc_wdis_dclk_bltrd1),
     .smc_wdis_dclk_bltld3(smc_wdis_dclk_bltld3r),
     .en_8bconfig_b_bltrd1(en_8bconfig_b_bltrd1),
     .en_8bconfig_b_bltld3(en_8bconfig_b_bltld3),
     .data_muxsel_bltrd1(data_muxsel_bltrd1),
     .data_muxsel_bltld3(data_muxsel_bltld3),
     .data_muxsel1_bltld3(data_muxsel1_bltld3),
     .cram_write_bltrd1(cram_write_bltrd1),
     .cram_write_bltld3(cram_write_bltld3),
     .cram_pullup_bltld3(cram_pullup_b_bltld3),
     .cram_pullup_b_bltrd1(cram_pullup_b_bltrd1),
     .cram_prec_bltrd1(cram_prec_bltrd1),
     .core_por_b_rowu3(core_por_b_rowu3),
     .core_por_b_rowu1(core_por_b_rowu1),
     .cm_sdi_u3d2(cm_sdi_u3d2[1:0]), .cm_sdi_u1d3(cm_sdi_u1d3[1:0]),
     .cm_prec_bltld3(cram_prec_bltld3), .cm_clk_bltrd1(cm_clk_bltrd1),
     .cm_clk_bltld3(cm_clk_bltld3),
     .cm_banksel_bltrd1(cm_banksel_bltrd1[3]),
     .cm_banksel_bltld3(cm_banksel_bltld3[1]),
     .cm_sdo_u3(cm_sdo_u3[1:0]), .cm_sdo_u1(cm_sdo_u1[1:0]));
//PRCUTSSTLSTDR I40cutr ( .VSS(gnd_), .VSSPST(gnd_));
//PRCUTSSTLSTDL I40cutl ( .VSS(gnd_), .VSSPST(gnd_));

endmodule
// Library - leafcell, Cell - clk_mux2to18k, View - schematic
// LAST TIME SAVED: Apr 24 16:46:58 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module clk_mux2to18k ( clk, cbit, cbitb, min, prog );
output  clk;

input  cbit, cbitb, prog;

input [1:0]  min;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I289 ( .A(net29), .Y(clk));
inv_hvt I288 ( .A(prog), .Y(net27));
nand2_hvt I287 ( .A(net27), .Y(net29), .B(st2));
txgate_hvt I249 ( .in(min[1]), .out(st2), .pp(cbitb), .nn(cbit));
txgate_hvt I248 ( .in(min[0]), .out(st2), .pp(cbit), .nn(cbitb));

endmodule
// Library - xpmem, Cell - cram2x2, View - schematic
// LAST TIME SAVED: Jul 28 08:23:43 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module cram2x2 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [3:0]  q;
output [3:0]  q_b;

inout [1:0]  bl;

input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  r_vdd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



eh_cram_cell_4 Icram_cellb831r255 ( .q_b(q_b[1]), .q(q[1]), .wl(wl[0]),
     .bl(bl[1]), .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I20 ( .q_b(q_b[2]), .q(q[2]), .wl(wl[1]), .bl(bl[0]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));
eh_cram_cell_4 I15 ( .q_b(q_b[0]), .q(q[0]), .wl(wl[0]), .bl(bl[0]),
     .r_vdd(r_vdd[0]), .pgate(pgate[0]), .reset(reset[0]));
eh_cram_cell_4 I19 ( .q_b(q_b[3]), .q(q[3]), .wl(wl[1]), .bl(bl[1]),
     .r_vdd(r_vdd[1]), .pgate(pgate[1]), .reset(reset[1]));

endmodule
// Library - leafcell, Cell - clk_mux2to1x48k, View - schematic
// LAST TIME SAVED: Jan 15 15:45:32 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module clk_mux2to1x48k ( gnet, bl, min0, min1, min2, min3, pgate_l,
     pgate_r, prog, reset_l, reset_r, vdd_cntl_l, vdd_cntl_r, wl_l,
     wl_r );


input  prog;

output [3:0]  gnet;

inout [3:0]  bl;

input [1:0]  min2;
input [1:0]  pgate_l;
input [1:0]  reset_r;
input [1:0]  min0;
input [1:0]  wl_r;
input [1:0]  reset_l;
input [1:0]  pgate_r;
input [1:0]  vdd_cntl_r;
input [1:0]  min1;
input [1:0]  wl_l;
input [1:0]  vdd_cntl_l;
input [1:0]  min3;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [7:0]  cbitb;

wire  [0:1]  l_vdd;

wire  [7:0]  cbit;



clk_mux2to18k I295 ( .prog(prog), .cbit(cbit[3]), .cbitb(cbitb[3]),
     .min(min3[1:0]), .clk(gnet[3]));
clk_mux2to18k I293 ( .prog(prog), .cbit(cbit[1]), .cbitb(cbitb[1]),
     .min(min1[1:0]), .clk(gnet[1]));
clk_mux2to18k I294 ( .prog(prog), .cbit(cbit[2]), .cbitb(cbitb[2]),
     .min(min2[1:0]), .clk(gnet[2]));
clk_mux2to18k I291 ( .prog(prog), .cbit(cbit[0]), .cbitb(cbitb[0]),
     .min(min0[1:0]), .clk(gnet[0]));
pch_hvt  vdd_cntrl_1_ ( .D(l_vdd[0]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(l_vdd[1]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));
pch_hvt  M1_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl_r[1]), .S(vdd_));
pch_hvt  M1_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl_r[0]), .S(vdd_));
cram2x2 I292 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset_l[1:0]),
     .q(cbit[3:0]), .wl(wl_l[1:0]), .r_vdd(l_vdd[0:1]),
     .pgate(pgate_l[1:0]));
cram2x2 I298 ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset_r[1:0]),
     .q(cbit[7:4]), .wl(wl_r[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate_r[1:0]));

endmodule
// Library - xpmem, Cell - cram2x2x2, View - schematic
// LAST TIME SAVED: Apr 14 10:22:48 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module cram2x2x2 ( q, q_b, bl, pgate_l, pgate_r, r_gnd_l, r_gnd_r,
     reset_b_l, reset_b_r, wl_l, wl_r );



output [7:0]  q_b;
output [7:0]  q;

inout [3:0]  bl;

input [1:0]  reset_b_r;
input [1:0]  pgate_l;
input [1:0]  r_gnd_r;
input [1:0]  r_gnd_l;
input [1:0]  pgate_r;
input [1:0]  wl_l;
input [1:0]  reset_b_l;
input [1:0]  wl_r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imrgt ( .bl(bl[3:2]), .q_b(q_b[7:4]), .reset(reset_b_r[1:0]),
     .q(q[7:4]), .wl(wl_r[1:0]), .r_vdd(r_gnd_r[1:0]),
     .pgate(pgate_r[1:0]));
cram2x2 Imleft ( .reset(reset_b_l[1:0]), .r_vdd(r_gnd_l[1:0]),
     .pgate(pgate_l[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl_l[1:0]));

endmodule
// Library - xpmem, Cell - ml_rowdrv2_last, View - schematic
// LAST TIME SAVED: Sep 26 14:07:07 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_rowdrv2_last ( pgate, reset, smc_rsr_out, vddctrl, wl,
     wl_rd_sup, wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write
     );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  NM0 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
ml_dff_schematic I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));

endmodule
// Library - leafcell, Cell - cram_row270col4, View - schematic
// LAST TIME SAVED: Dec  6 09:25:12 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module cram_row270col4 ( bl, pgate_l, pgate_r, reset_l, reset_r,
     vdd_cntl_l, vdd_cntl_r, wl_l, wl_r );


inout [3:0]  bl;

input [269:0]  reset_r;
input [269:0]  wl_l;
input [269:0]  pgate_r;
input [269:0]  pgate_l;
input [269:0]  vdd_cntl_l;
input [269:0]  vdd_cntl_r;
input [269:0]  wl_r;
input [269:0]  reset_l;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1079]  net37;

wire  [0:1079]  net36;

wire  [0:269]  net32;

wire  [0:269]  net43;



cram2x2x2 xcram_134_ ( .pgate_l(pgate_l[269:268]),
     .wl_l(wl_l[269:268]), .reset_b_l(reset_l[269:268]),
     .r_gnd_l(net43[0:1]), .r_gnd_r(net32[0:1]),
     .pgate_r(pgate_r[269:268]), .wl_r(wl_r[269:268]),
     .reset_b_r(reset_r[269:268]), .q(net36[0:7]), .q_b(net37[0:7]),
     .bl(bl[3:0]));
cram2x2x2 xcram_133_ ( .pgate_l(pgate_l[267:266]),
     .wl_l(wl_l[267:266]), .reset_b_l(reset_l[267:266]),
     .r_gnd_l(net43[2:3]), .r_gnd_r(net32[2:3]),
     .pgate_r(pgate_r[267:266]), .wl_r(wl_r[267:266]),
     .reset_b_r(reset_r[267:266]), .q(net36[8:15]), .q_b(net37[8:15]),
     .bl(bl[3:0]));
cram2x2x2 xcram_132_ ( .pgate_l(pgate_l[265:264]),
     .wl_l(wl_l[265:264]), .reset_b_l(reset_l[265:264]),
     .r_gnd_l(net43[4:5]), .r_gnd_r(net32[4:5]),
     .pgate_r(pgate_r[265:264]), .wl_r(wl_r[265:264]),
     .reset_b_r(reset_r[265:264]), .q(net36[16:23]),
     .q_b(net37[16:23]), .bl(bl[3:0]));
cram2x2x2 xcram_131_ ( .pgate_l(pgate_l[263:262]),
     .wl_l(wl_l[263:262]), .reset_b_l(reset_l[263:262]),
     .r_gnd_l(net43[6:7]), .r_gnd_r(net32[6:7]),
     .pgate_r(pgate_r[263:262]), .wl_r(wl_r[263:262]),
     .reset_b_r(reset_r[263:262]), .q(net36[24:31]),
     .q_b(net37[24:31]), .bl(bl[3:0]));
cram2x2x2 xcram_130_ ( .pgate_l(pgate_l[261:260]),
     .wl_l(wl_l[261:260]), .reset_b_l(reset_l[261:260]),
     .r_gnd_l(net43[8:9]), .r_gnd_r(net32[8:9]),
     .pgate_r(pgate_r[261:260]), .wl_r(wl_r[261:260]),
     .reset_b_r(reset_r[261:260]), .q(net36[32:39]),
     .q_b(net37[32:39]), .bl(bl[3:0]));
cram2x2x2 xcram_129_ ( .pgate_l(pgate_l[259:258]),
     .wl_l(wl_l[259:258]), .reset_b_l(reset_l[259:258]),
     .r_gnd_l(net43[10:11]), .r_gnd_r(net32[10:11]),
     .pgate_r(pgate_r[259:258]), .wl_r(wl_r[259:258]),
     .reset_b_r(reset_r[259:258]), .q(net36[40:47]),
     .q_b(net37[40:47]), .bl(bl[3:0]));
cram2x2x2 xcram_128_ ( .pgate_l(pgate_l[257:256]),
     .wl_l(wl_l[257:256]), .reset_b_l(reset_l[257:256]),
     .r_gnd_l(net43[12:13]), .r_gnd_r(net32[12:13]),
     .pgate_r(pgate_r[257:256]), .wl_r(wl_r[257:256]),
     .reset_b_r(reset_r[257:256]), .q(net36[48:55]),
     .q_b(net37[48:55]), .bl(bl[3:0]));
cram2x2x2 xcram_127_ ( .pgate_l(pgate_l[255:254]),
     .wl_l(wl_l[255:254]), .reset_b_l(reset_l[255:254]),
     .r_gnd_l(net43[14:15]), .r_gnd_r(net32[14:15]),
     .pgate_r(pgate_r[255:254]), .wl_r(wl_r[255:254]),
     .reset_b_r(reset_r[255:254]), .q(net36[56:63]),
     .q_b(net37[56:63]), .bl(bl[3:0]));
cram2x2x2 xcram_126_ ( .pgate_l(pgate_l[253:252]),
     .wl_l(wl_l[253:252]), .reset_b_l(reset_l[253:252]),
     .r_gnd_l(net43[16:17]), .r_gnd_r(net32[16:17]),
     .pgate_r(pgate_r[253:252]), .wl_r(wl_r[253:252]),
     .reset_b_r(reset_r[253:252]), .q(net36[64:71]),
     .q_b(net37[64:71]), .bl(bl[3:0]));
cram2x2x2 xcram_125_ ( .pgate_l(pgate_l[251:250]),
     .wl_l(wl_l[251:250]), .reset_b_l(reset_l[251:250]),
     .r_gnd_l(net43[18:19]), .r_gnd_r(net32[18:19]),
     .pgate_r(pgate_r[251:250]), .wl_r(wl_r[251:250]),
     .reset_b_r(reset_r[251:250]), .q(net36[72:79]),
     .q_b(net37[72:79]), .bl(bl[3:0]));
cram2x2x2 xcram_124_ ( .pgate_l(pgate_l[249:248]),
     .wl_l(wl_l[249:248]), .reset_b_l(reset_l[249:248]),
     .r_gnd_l(net43[20:21]), .r_gnd_r(net32[20:21]),
     .pgate_r(pgate_r[249:248]), .wl_r(wl_r[249:248]),
     .reset_b_r(reset_r[249:248]), .q(net36[80:87]),
     .q_b(net37[80:87]), .bl(bl[3:0]));
cram2x2x2 xcram_123_ ( .pgate_l(pgate_l[247:246]),
     .wl_l(wl_l[247:246]), .reset_b_l(reset_l[247:246]),
     .r_gnd_l(net43[22:23]), .r_gnd_r(net32[22:23]),
     .pgate_r(pgate_r[247:246]), .wl_r(wl_r[247:246]),
     .reset_b_r(reset_r[247:246]), .q(net36[88:95]),
     .q_b(net37[88:95]), .bl(bl[3:0]));
cram2x2x2 xcram_122_ ( .pgate_l(pgate_l[245:244]),
     .wl_l(wl_l[245:244]), .reset_b_l(reset_l[245:244]),
     .r_gnd_l(net43[24:25]), .r_gnd_r(net32[24:25]),
     .pgate_r(pgate_r[245:244]), .wl_r(wl_r[245:244]),
     .reset_b_r(reset_r[245:244]), .q(net36[96:103]),
     .q_b(net37[96:103]), .bl(bl[3:0]));
cram2x2x2 xcram_121_ ( .pgate_l(pgate_l[243:242]),
     .wl_l(wl_l[243:242]), .reset_b_l(reset_l[243:242]),
     .r_gnd_l(net43[26:27]), .r_gnd_r(net32[26:27]),
     .pgate_r(pgate_r[243:242]), .wl_r(wl_r[243:242]),
     .reset_b_r(reset_r[243:242]), .q(net36[104:111]),
     .q_b(net37[104:111]), .bl(bl[3:0]));
cram2x2x2 xcram_120_ ( .pgate_l(pgate_l[241:240]),
     .wl_l(wl_l[241:240]), .reset_b_l(reset_l[241:240]),
     .r_gnd_l(net43[28:29]), .r_gnd_r(net32[28:29]),
     .pgate_r(pgate_r[241:240]), .wl_r(wl_r[241:240]),
     .reset_b_r(reset_r[241:240]), .q(net36[112:119]),
     .q_b(net37[112:119]), .bl(bl[3:0]));
cram2x2x2 xcram_119_ ( .pgate_l(pgate_l[239:238]),
     .wl_l(wl_l[239:238]), .reset_b_l(reset_l[239:238]),
     .r_gnd_l(net43[30:31]), .r_gnd_r(net32[30:31]),
     .pgate_r(pgate_r[239:238]), .wl_r(wl_r[239:238]),
     .reset_b_r(reset_r[239:238]), .q(net36[120:127]),
     .q_b(net37[120:127]), .bl(bl[3:0]));
cram2x2x2 xcram_118_ ( .pgate_l(pgate_l[237:236]),
     .wl_l(wl_l[237:236]), .reset_b_l(reset_l[237:236]),
     .r_gnd_l(net43[32:33]), .r_gnd_r(net32[32:33]),
     .pgate_r(pgate_r[237:236]), .wl_r(wl_r[237:236]),
     .reset_b_r(reset_r[237:236]), .q(net36[128:135]),
     .q_b(net37[128:135]), .bl(bl[3:0]));
cram2x2x2 xcram_117_ ( .pgate_l(pgate_l[235:234]),
     .wl_l(wl_l[235:234]), .reset_b_l(reset_l[235:234]),
     .r_gnd_l(net43[34:35]), .r_gnd_r(net32[34:35]),
     .pgate_r(pgate_r[235:234]), .wl_r(wl_r[235:234]),
     .reset_b_r(reset_r[235:234]), .q(net36[136:143]),
     .q_b(net37[136:143]), .bl(bl[3:0]));
cram2x2x2 xcram_116_ ( .pgate_l(pgate_l[233:232]),
     .wl_l(wl_l[233:232]), .reset_b_l(reset_l[233:232]),
     .r_gnd_l(net43[36:37]), .r_gnd_r(net32[36:37]),
     .pgate_r(pgate_r[233:232]), .wl_r(wl_r[233:232]),
     .reset_b_r(reset_r[233:232]), .q(net36[144:151]),
     .q_b(net37[144:151]), .bl(bl[3:0]));
cram2x2x2 xcram_115_ ( .pgate_l(pgate_l[231:230]),
     .wl_l(wl_l[231:230]), .reset_b_l(reset_l[231:230]),
     .r_gnd_l(net43[38:39]), .r_gnd_r(net32[38:39]),
     .pgate_r(pgate_r[231:230]), .wl_r(wl_r[231:230]),
     .reset_b_r(reset_r[231:230]), .q(net36[152:159]),
     .q_b(net37[152:159]), .bl(bl[3:0]));
cram2x2x2 xcram_114_ ( .pgate_l(pgate_l[229:228]),
     .wl_l(wl_l[229:228]), .reset_b_l(reset_l[229:228]),
     .r_gnd_l(net43[40:41]), .r_gnd_r(net32[40:41]),
     .pgate_r(pgate_r[229:228]), .wl_r(wl_r[229:228]),
     .reset_b_r(reset_r[229:228]), .q(net36[160:167]),
     .q_b(net37[160:167]), .bl(bl[3:0]));
cram2x2x2 xcram_113_ ( .pgate_l(pgate_l[227:226]),
     .wl_l(wl_l[227:226]), .reset_b_l(reset_l[227:226]),
     .r_gnd_l(net43[42:43]), .r_gnd_r(net32[42:43]),
     .pgate_r(pgate_r[227:226]), .wl_r(wl_r[227:226]),
     .reset_b_r(reset_r[227:226]), .q(net36[168:175]),
     .q_b(net37[168:175]), .bl(bl[3:0]));
cram2x2x2 xcram_112_ ( .pgate_l(pgate_l[225:224]),
     .wl_l(wl_l[225:224]), .reset_b_l(reset_l[225:224]),
     .r_gnd_l(net43[44:45]), .r_gnd_r(net32[44:45]),
     .pgate_r(pgate_r[225:224]), .wl_r(wl_r[225:224]),
     .reset_b_r(reset_r[225:224]), .q(net36[176:183]),
     .q_b(net37[176:183]), .bl(bl[3:0]));
cram2x2x2 xcram_111_ ( .pgate_l(pgate_l[223:222]),
     .wl_l(wl_l[223:222]), .reset_b_l(reset_l[223:222]),
     .r_gnd_l(net43[46:47]), .r_gnd_r(net32[46:47]),
     .pgate_r(pgate_r[223:222]), .wl_r(wl_r[223:222]),
     .reset_b_r(reset_r[223:222]), .q(net36[184:191]),
     .q_b(net37[184:191]), .bl(bl[3:0]));
cram2x2x2 xcram_110_ ( .pgate_l(pgate_l[221:220]),
     .wl_l(wl_l[221:220]), .reset_b_l(reset_l[221:220]),
     .r_gnd_l(net43[48:49]), .r_gnd_r(net32[48:49]),
     .pgate_r(pgate_r[221:220]), .wl_r(wl_r[221:220]),
     .reset_b_r(reset_r[221:220]), .q(net36[192:199]),
     .q_b(net37[192:199]), .bl(bl[3:0]));
cram2x2x2 xcram_109_ ( .pgate_l(pgate_l[219:218]),
     .wl_l(wl_l[219:218]), .reset_b_l(reset_l[219:218]),
     .r_gnd_l(net43[50:51]), .r_gnd_r(net32[50:51]),
     .pgate_r(pgate_r[219:218]), .wl_r(wl_r[219:218]),
     .reset_b_r(reset_r[219:218]), .q(net36[200:207]),
     .q_b(net37[200:207]), .bl(bl[3:0]));
cram2x2x2 xcram_108_ ( .pgate_l(pgate_l[217:216]),
     .wl_l(wl_l[217:216]), .reset_b_l(reset_l[217:216]),
     .r_gnd_l(net43[52:53]), .r_gnd_r(net32[52:53]),
     .pgate_r(pgate_r[217:216]), .wl_r(wl_r[217:216]),
     .reset_b_r(reset_r[217:216]), .q(net36[208:215]),
     .q_b(net37[208:215]), .bl(bl[3:0]));
cram2x2x2 xcram_107_ ( .pgate_l(pgate_l[215:214]),
     .wl_l(wl_l[215:214]), .reset_b_l(reset_l[215:214]),
     .r_gnd_l(net43[54:55]), .r_gnd_r(net32[54:55]),
     .pgate_r(pgate_r[215:214]), .wl_r(wl_r[215:214]),
     .reset_b_r(reset_r[215:214]), .q(net36[216:223]),
     .q_b(net37[216:223]), .bl(bl[3:0]));
cram2x2x2 xcram_106_ ( .pgate_l(pgate_l[213:212]),
     .wl_l(wl_l[213:212]), .reset_b_l(reset_l[213:212]),
     .r_gnd_l(net43[56:57]), .r_gnd_r(net32[56:57]),
     .pgate_r(pgate_r[213:212]), .wl_r(wl_r[213:212]),
     .reset_b_r(reset_r[213:212]), .q(net36[224:231]),
     .q_b(net37[224:231]), .bl(bl[3:0]));
cram2x2x2 xcram_105_ ( .pgate_l(pgate_l[211:210]),
     .wl_l(wl_l[211:210]), .reset_b_l(reset_l[211:210]),
     .r_gnd_l(net43[58:59]), .r_gnd_r(net32[58:59]),
     .pgate_r(pgate_r[211:210]), .wl_r(wl_r[211:210]),
     .reset_b_r(reset_r[211:210]), .q(net36[232:239]),
     .q_b(net37[232:239]), .bl(bl[3:0]));
cram2x2x2 xcram_104_ ( .pgate_l(pgate_l[209:208]),
     .wl_l(wl_l[209:208]), .reset_b_l(reset_l[209:208]),
     .r_gnd_l(net43[60:61]), .r_gnd_r(net32[60:61]),
     .pgate_r(pgate_r[209:208]), .wl_r(wl_r[209:208]),
     .reset_b_r(reset_r[209:208]), .q(net36[240:247]),
     .q_b(net37[240:247]), .bl(bl[3:0]));
cram2x2x2 xcram_103_ ( .pgate_l(pgate_l[207:206]),
     .wl_l(wl_l[207:206]), .reset_b_l(reset_l[207:206]),
     .r_gnd_l(net43[62:63]), .r_gnd_r(net32[62:63]),
     .pgate_r(pgate_r[207:206]), .wl_r(wl_r[207:206]),
     .reset_b_r(reset_r[207:206]), .q(net36[248:255]),
     .q_b(net37[248:255]), .bl(bl[3:0]));
cram2x2x2 xcram_102_ ( .pgate_l(pgate_l[205:204]),
     .wl_l(wl_l[205:204]), .reset_b_l(reset_l[205:204]),
     .r_gnd_l(net43[64:65]), .r_gnd_r(net32[64:65]),
     .pgate_r(pgate_r[205:204]), .wl_r(wl_r[205:204]),
     .reset_b_r(reset_r[205:204]), .q(net36[256:263]),
     .q_b(net37[256:263]), .bl(bl[3:0]));
cram2x2x2 xcram_101_ ( .pgate_l(pgate_l[203:202]),
     .wl_l(wl_l[203:202]), .reset_b_l(reset_l[203:202]),
     .r_gnd_l(net43[66:67]), .r_gnd_r(net32[66:67]),
     .pgate_r(pgate_r[203:202]), .wl_r(wl_r[203:202]),
     .reset_b_r(reset_r[203:202]), .q(net36[264:271]),
     .q_b(net37[264:271]), .bl(bl[3:0]));
cram2x2x2 xcram_100_ ( .pgate_l(pgate_l[201:200]),
     .wl_l(wl_l[201:200]), .reset_b_l(reset_l[201:200]),
     .r_gnd_l(net43[68:69]), .r_gnd_r(net32[68:69]),
     .pgate_r(pgate_r[201:200]), .wl_r(wl_r[201:200]),
     .reset_b_r(reset_r[201:200]), .q(net36[272:279]),
     .q_b(net37[272:279]), .bl(bl[3:0]));
cram2x2x2 xcram_99_ ( .pgate_l(pgate_l[199:198]), .wl_l(wl_l[199:198]),
     .reset_b_l(reset_l[199:198]), .r_gnd_l(net43[70:71]),
     .r_gnd_r(net32[70:71]), .pgate_r(pgate_r[199:198]),
     .wl_r(wl_r[199:198]), .reset_b_r(reset_r[199:198]),
     .q(net36[280:287]), .q_b(net37[280:287]), .bl(bl[3:0]));
cram2x2x2 xcram_98_ ( .pgate_l(pgate_l[197:196]), .wl_l(wl_l[197:196]),
     .reset_b_l(reset_l[197:196]), .r_gnd_l(net43[72:73]),
     .r_gnd_r(net32[72:73]), .pgate_r(pgate_r[197:196]),
     .wl_r(wl_r[197:196]), .reset_b_r(reset_r[197:196]),
     .q(net36[288:295]), .q_b(net37[288:295]), .bl(bl[3:0]));
cram2x2x2 xcram_97_ ( .pgate_l(pgate_l[195:194]), .wl_l(wl_l[195:194]),
     .reset_b_l(reset_l[195:194]), .r_gnd_l(net43[74:75]),
     .r_gnd_r(net32[74:75]), .pgate_r(pgate_r[195:194]),
     .wl_r(wl_r[195:194]), .reset_b_r(reset_r[195:194]),
     .q(net36[296:303]), .q_b(net37[296:303]), .bl(bl[3:0]));
cram2x2x2 xcram_96_ ( .pgate_l(pgate_l[193:192]), .wl_l(wl_l[193:192]),
     .reset_b_l(reset_l[193:192]), .r_gnd_l(net43[76:77]),
     .r_gnd_r(net32[76:77]), .pgate_r(pgate_r[193:192]),
     .wl_r(wl_r[193:192]), .reset_b_r(reset_r[193:192]),
     .q(net36[304:311]), .q_b(net37[304:311]), .bl(bl[3:0]));
cram2x2x2 xcram_95_ ( .pgate_l(pgate_l[191:190]), .wl_l(wl_l[191:190]),
     .reset_b_l(reset_l[191:190]), .r_gnd_l(net43[78:79]),
     .r_gnd_r(net32[78:79]), .pgate_r(pgate_r[191:190]),
     .wl_r(wl_r[191:190]), .reset_b_r(reset_r[191:190]),
     .q(net36[312:319]), .q_b(net37[312:319]), .bl(bl[3:0]));
cram2x2x2 xcram_94_ ( .pgate_l(pgate_l[189:188]), .wl_l(wl_l[189:188]),
     .reset_b_l(reset_l[189:188]), .r_gnd_l(net43[80:81]),
     .r_gnd_r(net32[80:81]), .pgate_r(pgate_r[189:188]),
     .wl_r(wl_r[189:188]), .reset_b_r(reset_r[189:188]),
     .q(net36[320:327]), .q_b(net37[320:327]), .bl(bl[3:0]));
cram2x2x2 xcram_93_ ( .pgate_l(pgate_l[187:186]), .wl_l(wl_l[187:186]),
     .reset_b_l(reset_l[187:186]), .r_gnd_l(net43[82:83]),
     .r_gnd_r(net32[82:83]), .pgate_r(pgate_r[187:186]),
     .wl_r(wl_r[187:186]), .reset_b_r(reset_r[187:186]),
     .q(net36[328:335]), .q_b(net37[328:335]), .bl(bl[3:0]));
cram2x2x2 xcram_92_ ( .pgate_l(pgate_l[185:184]), .wl_l(wl_l[185:184]),
     .reset_b_l(reset_l[185:184]), .r_gnd_l(net43[84:85]),
     .r_gnd_r(net32[84:85]), .pgate_r(pgate_r[185:184]),
     .wl_r(wl_r[185:184]), .reset_b_r(reset_r[185:184]),
     .q(net36[336:343]), .q_b(net37[336:343]), .bl(bl[3:0]));
cram2x2x2 xcram_91_ ( .pgate_l(pgate_l[183:182]), .wl_l(wl_l[183:182]),
     .reset_b_l(reset_l[183:182]), .r_gnd_l(net43[86:87]),
     .r_gnd_r(net32[86:87]), .pgate_r(pgate_r[183:182]),
     .wl_r(wl_r[183:182]), .reset_b_r(reset_r[183:182]),
     .q(net36[344:351]), .q_b(net37[344:351]), .bl(bl[3:0]));
cram2x2x2 xcram_90_ ( .pgate_l(pgate_l[181:180]), .wl_l(wl_l[181:180]),
     .reset_b_l(reset_l[181:180]), .r_gnd_l(net43[88:89]),
     .r_gnd_r(net32[88:89]), .pgate_r(pgate_r[181:180]),
     .wl_r(wl_r[181:180]), .reset_b_r(reset_r[181:180]),
     .q(net36[352:359]), .q_b(net37[352:359]), .bl(bl[3:0]));
cram2x2x2 xcram_89_ ( .pgate_l(pgate_l[179:178]), .wl_l(wl_l[179:178]),
     .reset_b_l(reset_l[179:178]), .r_gnd_l(net43[90:91]),
     .r_gnd_r(net32[90:91]), .pgate_r(pgate_r[179:178]),
     .wl_r(wl_r[179:178]), .reset_b_r(reset_r[179:178]),
     .q(net36[360:367]), .q_b(net37[360:367]), .bl(bl[3:0]));
cram2x2x2 xcram_88_ ( .pgate_l(pgate_l[177:176]), .wl_l(wl_l[177:176]),
     .reset_b_l(reset_l[177:176]), .r_gnd_l(net43[92:93]),
     .r_gnd_r(net32[92:93]), .pgate_r(pgate_r[177:176]),
     .wl_r(wl_r[177:176]), .reset_b_r(reset_r[177:176]),
     .q(net36[368:375]), .q_b(net37[368:375]), .bl(bl[3:0]));
cram2x2x2 xcram_87_ ( .pgate_l(pgate_l[175:174]), .wl_l(wl_l[175:174]),
     .reset_b_l(reset_l[175:174]), .r_gnd_l(net43[94:95]),
     .r_gnd_r(net32[94:95]), .pgate_r(pgate_r[175:174]),
     .wl_r(wl_r[175:174]), .reset_b_r(reset_r[175:174]),
     .q(net36[376:383]), .q_b(net37[376:383]), .bl(bl[3:0]));
cram2x2x2 xcram_86_ ( .pgate_l(pgate_l[173:172]), .wl_l(wl_l[173:172]),
     .reset_b_l(reset_l[173:172]), .r_gnd_l(net43[96:97]),
     .r_gnd_r(net32[96:97]), .pgate_r(pgate_r[173:172]),
     .wl_r(wl_r[173:172]), .reset_b_r(reset_r[173:172]),
     .q(net36[384:391]), .q_b(net37[384:391]), .bl(bl[3:0]));
cram2x2x2 xcram_85_ ( .pgate_l(pgate_l[171:170]), .wl_l(wl_l[171:170]),
     .reset_b_l(reset_l[171:170]), .r_gnd_l(net43[98:99]),
     .r_gnd_r(net32[98:99]), .pgate_r(pgate_r[171:170]),
     .wl_r(wl_r[171:170]), .reset_b_r(reset_r[171:170]),
     .q(net36[392:399]), .q_b(net37[392:399]), .bl(bl[3:0]));
cram2x2x2 xcram_84_ ( .pgate_l(pgate_l[169:168]), .wl_l(wl_l[169:168]),
     .reset_b_l(reset_l[169:168]), .r_gnd_l(net43[100:101]),
     .r_gnd_r(net32[100:101]), .pgate_r(pgate_r[169:168]),
     .wl_r(wl_r[169:168]), .reset_b_r(reset_r[169:168]),
     .q(net36[400:407]), .q_b(net37[400:407]), .bl(bl[3:0]));
cram2x2x2 xcram_83_ ( .pgate_l(pgate_l[167:166]), .wl_l(wl_l[167:166]),
     .reset_b_l(reset_l[167:166]), .r_gnd_l(net43[102:103]),
     .r_gnd_r(net32[102:103]), .pgate_r(pgate_r[167:166]),
     .wl_r(wl_r[167:166]), .reset_b_r(reset_r[167:166]),
     .q(net36[408:415]), .q_b(net37[408:415]), .bl(bl[3:0]));
cram2x2x2 xcram_82_ ( .pgate_l(pgate_l[165:164]), .wl_l(wl_l[165:164]),
     .reset_b_l(reset_l[165:164]), .r_gnd_l(net43[104:105]),
     .r_gnd_r(net32[104:105]), .pgate_r(pgate_r[165:164]),
     .wl_r(wl_r[165:164]), .reset_b_r(reset_r[165:164]),
     .q(net36[416:423]), .q_b(net37[416:423]), .bl(bl[3:0]));
cram2x2x2 xcram_81_ ( .pgate_l(pgate_l[163:162]), .wl_l(wl_l[163:162]),
     .reset_b_l(reset_l[163:162]), .r_gnd_l(net43[106:107]),
     .r_gnd_r(net32[106:107]), .pgate_r(pgate_r[163:162]),
     .wl_r(wl_r[163:162]), .reset_b_r(reset_r[163:162]),
     .q(net36[424:431]), .q_b(net37[424:431]), .bl(bl[3:0]));
cram2x2x2 xcram_80_ ( .pgate_l(pgate_l[161:160]), .wl_l(wl_l[161:160]),
     .reset_b_l(reset_l[161:160]), .r_gnd_l(net43[108:109]),
     .r_gnd_r(net32[108:109]), .pgate_r(pgate_r[161:160]),
     .wl_r(wl_r[161:160]), .reset_b_r(reset_r[161:160]),
     .q(net36[432:439]), .q_b(net37[432:439]), .bl(bl[3:0]));
cram2x2x2 xcram_79_ ( .pgate_l(pgate_l[159:158]), .wl_l(wl_l[159:158]),
     .reset_b_l(reset_l[159:158]), .r_gnd_l(net43[110:111]),
     .r_gnd_r(net32[110:111]), .pgate_r(pgate_r[159:158]),
     .wl_r(wl_r[159:158]), .reset_b_r(reset_r[159:158]),
     .q(net36[440:447]), .q_b(net37[440:447]), .bl(bl[3:0]));
cram2x2x2 xcram_78_ ( .pgate_l(pgate_l[157:156]), .wl_l(wl_l[157:156]),
     .reset_b_l(reset_l[157:156]), .r_gnd_l(net43[112:113]),
     .r_gnd_r(net32[112:113]), .pgate_r(pgate_r[157:156]),
     .wl_r(wl_r[157:156]), .reset_b_r(reset_r[157:156]),
     .q(net36[448:455]), .q_b(net37[448:455]), .bl(bl[3:0]));
cram2x2x2 xcram_77_ ( .pgate_l(pgate_l[155:154]), .wl_l(wl_l[155:154]),
     .reset_b_l(reset_l[155:154]), .r_gnd_l(net43[114:115]),
     .r_gnd_r(net32[114:115]), .pgate_r(pgate_r[155:154]),
     .wl_r(wl_r[155:154]), .reset_b_r(reset_r[155:154]),
     .q(net36[456:463]), .q_b(net37[456:463]), .bl(bl[3:0]));
cram2x2x2 xcram_76_ ( .pgate_l(pgate_l[153:152]), .wl_l(wl_l[153:152]),
     .reset_b_l(reset_l[153:152]), .r_gnd_l(net43[116:117]),
     .r_gnd_r(net32[116:117]), .pgate_r(pgate_r[153:152]),
     .wl_r(wl_r[153:152]), .reset_b_r(reset_r[153:152]),
     .q(net36[464:471]), .q_b(net37[464:471]), .bl(bl[3:0]));
cram2x2x2 xcram_75_ ( .pgate_l(pgate_l[151:150]), .wl_l(wl_l[151:150]),
     .reset_b_l(reset_l[151:150]), .r_gnd_l(net43[118:119]),
     .r_gnd_r(net32[118:119]), .pgate_r(pgate_r[151:150]),
     .wl_r(wl_r[151:150]), .reset_b_r(reset_r[151:150]),
     .q(net36[472:479]), .q_b(net37[472:479]), .bl(bl[3:0]));
cram2x2x2 xcram_74_ ( .pgate_l(pgate_l[149:148]), .wl_l(wl_l[149:148]),
     .reset_b_l(reset_l[149:148]), .r_gnd_l(net43[120:121]),
     .r_gnd_r(net32[120:121]), .pgate_r(pgate_r[149:148]),
     .wl_r(wl_r[149:148]), .reset_b_r(reset_r[149:148]),
     .q(net36[480:487]), .q_b(net37[480:487]), .bl(bl[3:0]));
cram2x2x2 xcram_73_ ( .pgate_l(pgate_l[147:146]), .wl_l(wl_l[147:146]),
     .reset_b_l(reset_l[147:146]), .r_gnd_l(net43[122:123]),
     .r_gnd_r(net32[122:123]), .pgate_r(pgate_r[147:146]),
     .wl_r(wl_r[147:146]), .reset_b_r(reset_r[147:146]),
     .q(net36[488:495]), .q_b(net37[488:495]), .bl(bl[3:0]));
cram2x2x2 xcram_72_ ( .pgate_l(pgate_l[145:144]), .wl_l(wl_l[145:144]),
     .reset_b_l(reset_l[145:144]), .r_gnd_l(net43[124:125]),
     .r_gnd_r(net32[124:125]), .pgate_r(pgate_r[145:144]),
     .wl_r(wl_r[145:144]), .reset_b_r(reset_r[145:144]),
     .q(net36[496:503]), .q_b(net37[496:503]), .bl(bl[3:0]));
cram2x2x2 xcram_71_ ( .pgate_l(pgate_l[143:142]), .wl_l(wl_l[143:142]),
     .reset_b_l(reset_l[143:142]), .r_gnd_l(net43[126:127]),
     .r_gnd_r(net32[126:127]), .pgate_r(pgate_r[143:142]),
     .wl_r(wl_r[143:142]), .reset_b_r(reset_r[143:142]),
     .q(net36[504:511]), .q_b(net37[504:511]), .bl(bl[3:0]));
cram2x2x2 xcram_70_ ( .pgate_l(pgate_l[141:140]), .wl_l(wl_l[141:140]),
     .reset_b_l(reset_l[141:140]), .r_gnd_l(net43[128:129]),
     .r_gnd_r(net32[128:129]), .pgate_r(pgate_r[141:140]),
     .wl_r(wl_r[141:140]), .reset_b_r(reset_r[141:140]),
     .q(net36[512:519]), .q_b(net37[512:519]), .bl(bl[3:0]));
cram2x2x2 xcram_69_ ( .pgate_l(pgate_l[139:138]), .wl_l(wl_l[139:138]),
     .reset_b_l(reset_l[139:138]), .r_gnd_l(net43[130:131]),
     .r_gnd_r(net32[130:131]), .pgate_r(pgate_r[139:138]),
     .wl_r(wl_r[139:138]), .reset_b_r(reset_r[139:138]),
     .q(net36[520:527]), .q_b(net37[520:527]), .bl(bl[3:0]));
cram2x2x2 xcram_68_ ( .pgate_l(pgate_l[137:136]), .wl_l(wl_l[137:136]),
     .reset_b_l(reset_l[137:136]), .r_gnd_l(net43[132:133]),
     .r_gnd_r(net32[132:133]), .pgate_r(pgate_r[137:136]),
     .wl_r(wl_r[137:136]), .reset_b_r(reset_r[137:136]),
     .q(net36[528:535]), .q_b(net37[528:535]), .bl(bl[3:0]));
cram2x2x2 xcram_67_ ( .pgate_l(pgate_l[135:134]), .wl_l(wl_l[135:134]),
     .reset_b_l(reset_l[135:134]), .r_gnd_l(net43[134:135]),
     .r_gnd_r(net32[134:135]), .pgate_r(pgate_r[135:134]),
     .wl_r(wl_r[135:134]), .reset_b_r(reset_r[135:134]),
     .q(net36[536:543]), .q_b(net37[536:543]), .bl(bl[3:0]));
cram2x2x2 xcram_66_ ( .pgate_l(pgate_l[133:132]), .wl_l(wl_l[133:132]),
     .reset_b_l(reset_l[133:132]), .r_gnd_l(net43[136:137]),
     .r_gnd_r(net32[136:137]), .pgate_r(pgate_r[133:132]),
     .wl_r(wl_r[133:132]), .reset_b_r(reset_r[133:132]),
     .q(net36[544:551]), .q_b(net37[544:551]), .bl(bl[3:0]));
cram2x2x2 xcram_65_ ( .pgate_l(pgate_l[131:130]), .wl_l(wl_l[131:130]),
     .reset_b_l(reset_l[131:130]), .r_gnd_l(net43[138:139]),
     .r_gnd_r(net32[138:139]), .pgate_r(pgate_r[131:130]),
     .wl_r(wl_r[131:130]), .reset_b_r(reset_r[131:130]),
     .q(net36[552:559]), .q_b(net37[552:559]), .bl(bl[3:0]));
cram2x2x2 xcram_64_ ( .pgate_l(pgate_l[129:128]), .wl_l(wl_l[129:128]),
     .reset_b_l(reset_l[129:128]), .r_gnd_l(net43[140:141]),
     .r_gnd_r(net32[140:141]), .pgate_r(pgate_r[129:128]),
     .wl_r(wl_r[129:128]), .reset_b_r(reset_r[129:128]),
     .q(net36[560:567]), .q_b(net37[560:567]), .bl(bl[3:0]));
cram2x2x2 xcram_63_ ( .pgate_l(pgate_l[127:126]), .wl_l(wl_l[127:126]),
     .reset_b_l(reset_l[127:126]), .r_gnd_l(net43[142:143]),
     .r_gnd_r(net32[142:143]), .pgate_r(pgate_r[127:126]),
     .wl_r(wl_r[127:126]), .reset_b_r(reset_r[127:126]),
     .q(net36[568:575]), .q_b(net37[568:575]), .bl(bl[3:0]));
cram2x2x2 xcram_62_ ( .pgate_l(pgate_l[125:124]), .wl_l(wl_l[125:124]),
     .reset_b_l(reset_l[125:124]), .r_gnd_l(net43[144:145]),
     .r_gnd_r(net32[144:145]), .pgate_r(pgate_r[125:124]),
     .wl_r(wl_r[125:124]), .reset_b_r(reset_r[125:124]),
     .q(net36[576:583]), .q_b(net37[576:583]), .bl(bl[3:0]));
cram2x2x2 xcram_61_ ( .pgate_l(pgate_l[123:122]), .wl_l(wl_l[123:122]),
     .reset_b_l(reset_l[123:122]), .r_gnd_l(net43[146:147]),
     .r_gnd_r(net32[146:147]), .pgate_r(pgate_r[123:122]),
     .wl_r(wl_r[123:122]), .reset_b_r(reset_r[123:122]),
     .q(net36[584:591]), .q_b(net37[584:591]), .bl(bl[3:0]));
cram2x2x2 xcram_60_ ( .pgate_l(pgate_l[121:120]), .wl_l(wl_l[121:120]),
     .reset_b_l(reset_l[121:120]), .r_gnd_l(net43[148:149]),
     .r_gnd_r(net32[148:149]), .pgate_r(pgate_r[121:120]),
     .wl_r(wl_r[121:120]), .reset_b_r(reset_r[121:120]),
     .q(net36[592:599]), .q_b(net37[592:599]), .bl(bl[3:0]));
cram2x2x2 xcram_59_ ( .pgate_l(pgate_l[119:118]), .wl_l(wl_l[119:118]),
     .reset_b_l(reset_l[119:118]), .r_gnd_l(net43[150:151]),
     .r_gnd_r(net32[150:151]), .pgate_r(pgate_r[119:118]),
     .wl_r(wl_r[119:118]), .reset_b_r(reset_r[119:118]),
     .q(net36[600:607]), .q_b(net37[600:607]), .bl(bl[3:0]));
cram2x2x2 xcram_58_ ( .pgate_l(pgate_l[117:116]), .wl_l(wl_l[117:116]),
     .reset_b_l(reset_l[117:116]), .r_gnd_l(net43[152:153]),
     .r_gnd_r(net32[152:153]), .pgate_r(pgate_r[117:116]),
     .wl_r(wl_r[117:116]), .reset_b_r(reset_r[117:116]),
     .q(net36[608:615]), .q_b(net37[608:615]), .bl(bl[3:0]));
cram2x2x2 xcram_57_ ( .pgate_l(pgate_l[115:114]), .wl_l(wl_l[115:114]),
     .reset_b_l(reset_l[115:114]), .r_gnd_l(net43[154:155]),
     .r_gnd_r(net32[154:155]), .pgate_r(pgate_r[115:114]),
     .wl_r(wl_r[115:114]), .reset_b_r(reset_r[115:114]),
     .q(net36[616:623]), .q_b(net37[616:623]), .bl(bl[3:0]));
cram2x2x2 xcram_56_ ( .pgate_l(pgate_l[113:112]), .wl_l(wl_l[113:112]),
     .reset_b_l(reset_l[113:112]), .r_gnd_l(net43[156:157]),
     .r_gnd_r(net32[156:157]), .pgate_r(pgate_r[113:112]),
     .wl_r(wl_r[113:112]), .reset_b_r(reset_r[113:112]),
     .q(net36[624:631]), .q_b(net37[624:631]), .bl(bl[3:0]));
cram2x2x2 xcram_55_ ( .pgate_l(pgate_l[111:110]), .wl_l(wl_l[111:110]),
     .reset_b_l(reset_l[111:110]), .r_gnd_l(net43[158:159]),
     .r_gnd_r(net32[158:159]), .pgate_r(pgate_r[111:110]),
     .wl_r(wl_r[111:110]), .reset_b_r(reset_r[111:110]),
     .q(net36[632:639]), .q_b(net37[632:639]), .bl(bl[3:0]));
cram2x2x2 xcram_54_ ( .pgate_l(pgate_l[109:108]), .wl_l(wl_l[109:108]),
     .reset_b_l(reset_l[109:108]), .r_gnd_l(net43[160:161]),
     .r_gnd_r(net32[160:161]), .pgate_r(pgate_r[109:108]),
     .wl_r(wl_r[109:108]), .reset_b_r(reset_r[109:108]),
     .q(net36[640:647]), .q_b(net37[640:647]), .bl(bl[3:0]));
cram2x2x2 xcram_53_ ( .pgate_l(pgate_l[107:106]), .wl_l(wl_l[107:106]),
     .reset_b_l(reset_l[107:106]), .r_gnd_l(net43[162:163]),
     .r_gnd_r(net32[162:163]), .pgate_r(pgate_r[107:106]),
     .wl_r(wl_r[107:106]), .reset_b_r(reset_r[107:106]),
     .q(net36[648:655]), .q_b(net37[648:655]), .bl(bl[3:0]));
cram2x2x2 xcram_52_ ( .pgate_l(pgate_l[105:104]), .wl_l(wl_l[105:104]),
     .reset_b_l(reset_l[105:104]), .r_gnd_l(net43[164:165]),
     .r_gnd_r(net32[164:165]), .pgate_r(pgate_r[105:104]),
     .wl_r(wl_r[105:104]), .reset_b_r(reset_r[105:104]),
     .q(net36[656:663]), .q_b(net37[656:663]), .bl(bl[3:0]));
cram2x2x2 xcram_51_ ( .pgate_l(pgate_l[103:102]), .wl_l(wl_l[103:102]),
     .reset_b_l(reset_l[103:102]), .r_gnd_l(net43[166:167]),
     .r_gnd_r(net32[166:167]), .pgate_r(pgate_r[103:102]),
     .wl_r(wl_r[103:102]), .reset_b_r(reset_r[103:102]),
     .q(net36[664:671]), .q_b(net37[664:671]), .bl(bl[3:0]));
cram2x2x2 xcram_50_ ( .pgate_l(pgate_l[101:100]), .wl_l(wl_l[101:100]),
     .reset_b_l(reset_l[101:100]), .r_gnd_l(net43[168:169]),
     .r_gnd_r(net32[168:169]), .pgate_r(pgate_r[101:100]),
     .wl_r(wl_r[101:100]), .reset_b_r(reset_r[101:100]),
     .q(net36[672:679]), .q_b(net37[672:679]), .bl(bl[3:0]));
cram2x2x2 xcram_49_ ( .pgate_l(pgate_l[99:98]), .wl_l(wl_l[99:98]),
     .reset_b_l(reset_l[99:98]), .r_gnd_l(net43[170:171]),
     .r_gnd_r(net32[170:171]), .pgate_r(pgate_r[99:98]),
     .wl_r(wl_r[99:98]), .reset_b_r(reset_r[99:98]),
     .q(net36[680:687]), .q_b(net37[680:687]), .bl(bl[3:0]));
cram2x2x2 xcram_48_ ( .pgate_l(pgate_l[97:96]), .wl_l(wl_l[97:96]),
     .reset_b_l(reset_l[97:96]), .r_gnd_l(net43[172:173]),
     .r_gnd_r(net32[172:173]), .pgate_r(pgate_r[97:96]),
     .wl_r(wl_r[97:96]), .reset_b_r(reset_r[97:96]),
     .q(net36[688:695]), .q_b(net37[688:695]), .bl(bl[3:0]));
cram2x2x2 xcram_47_ ( .pgate_l(pgate_l[95:94]), .wl_l(wl_l[95:94]),
     .reset_b_l(reset_l[95:94]), .r_gnd_l(net43[174:175]),
     .r_gnd_r(net32[174:175]), .pgate_r(pgate_r[95:94]),
     .wl_r(wl_r[95:94]), .reset_b_r(reset_r[95:94]),
     .q(net36[696:703]), .q_b(net37[696:703]), .bl(bl[3:0]));
cram2x2x2 xcram_46_ ( .pgate_l(pgate_l[93:92]), .wl_l(wl_l[93:92]),
     .reset_b_l(reset_l[93:92]), .r_gnd_l(net43[176:177]),
     .r_gnd_r(net32[176:177]), .pgate_r(pgate_r[93:92]),
     .wl_r(wl_r[93:92]), .reset_b_r(reset_r[93:92]),
     .q(net36[704:711]), .q_b(net37[704:711]), .bl(bl[3:0]));
cram2x2x2 xcram_45_ ( .pgate_l(pgate_l[91:90]), .wl_l(wl_l[91:90]),
     .reset_b_l(reset_l[91:90]), .r_gnd_l(net43[178:179]),
     .r_gnd_r(net32[178:179]), .pgate_r(pgate_r[91:90]),
     .wl_r(wl_r[91:90]), .reset_b_r(reset_r[91:90]),
     .q(net36[712:719]), .q_b(net37[712:719]), .bl(bl[3:0]));
cram2x2x2 xcram_44_ ( .pgate_l(pgate_l[89:88]), .wl_l(wl_l[89:88]),
     .reset_b_l(reset_l[89:88]), .r_gnd_l(net43[180:181]),
     .r_gnd_r(net32[180:181]), .pgate_r(pgate_r[89:88]),
     .wl_r(wl_r[89:88]), .reset_b_r(reset_r[89:88]),
     .q(net36[720:727]), .q_b(net37[720:727]), .bl(bl[3:0]));
cram2x2x2 xcram_43_ ( .pgate_l(pgate_l[87:86]), .wl_l(wl_l[87:86]),
     .reset_b_l(reset_l[87:86]), .r_gnd_l(net43[182:183]),
     .r_gnd_r(net32[182:183]), .pgate_r(pgate_r[87:86]),
     .wl_r(wl_r[87:86]), .reset_b_r(reset_r[87:86]),
     .q(net36[728:735]), .q_b(net37[728:735]), .bl(bl[3:0]));
cram2x2x2 xcram_42_ ( .pgate_l(pgate_l[85:84]), .wl_l(wl_l[85:84]),
     .reset_b_l(reset_l[85:84]), .r_gnd_l(net43[184:185]),
     .r_gnd_r(net32[184:185]), .pgate_r(pgate_r[85:84]),
     .wl_r(wl_r[85:84]), .reset_b_r(reset_r[85:84]),
     .q(net36[736:743]), .q_b(net37[736:743]), .bl(bl[3:0]));
cram2x2x2 xcram_41_ ( .pgate_l(pgate_l[83:82]), .wl_l(wl_l[83:82]),
     .reset_b_l(reset_l[83:82]), .r_gnd_l(net43[186:187]),
     .r_gnd_r(net32[186:187]), .pgate_r(pgate_r[83:82]),
     .wl_r(wl_r[83:82]), .reset_b_r(reset_r[83:82]),
     .q(net36[744:751]), .q_b(net37[744:751]), .bl(bl[3:0]));
cram2x2x2 xcram_40_ ( .pgate_l(pgate_l[81:80]), .wl_l(wl_l[81:80]),
     .reset_b_l(reset_l[81:80]), .r_gnd_l(net43[188:189]),
     .r_gnd_r(net32[188:189]), .pgate_r(pgate_r[81:80]),
     .wl_r(wl_r[81:80]), .reset_b_r(reset_r[81:80]),
     .q(net36[752:759]), .q_b(net37[752:759]), .bl(bl[3:0]));
cram2x2x2 xcram_39_ ( .pgate_l(pgate_l[79:78]), .wl_l(wl_l[79:78]),
     .reset_b_l(reset_l[79:78]), .r_gnd_l(net43[190:191]),
     .r_gnd_r(net32[190:191]), .pgate_r(pgate_r[79:78]),
     .wl_r(wl_r[79:78]), .reset_b_r(reset_r[79:78]),
     .q(net36[760:767]), .q_b(net37[760:767]), .bl(bl[3:0]));
cram2x2x2 xcram_38_ ( .pgate_l(pgate_l[77:76]), .wl_l(wl_l[77:76]),
     .reset_b_l(reset_l[77:76]), .r_gnd_l(net43[192:193]),
     .r_gnd_r(net32[192:193]), .pgate_r(pgate_r[77:76]),
     .wl_r(wl_r[77:76]), .reset_b_r(reset_r[77:76]),
     .q(net36[768:775]), .q_b(net37[768:775]), .bl(bl[3:0]));
cram2x2x2 xcram_37_ ( .pgate_l(pgate_l[75:74]), .wl_l(wl_l[75:74]),
     .reset_b_l(reset_l[75:74]), .r_gnd_l(net43[194:195]),
     .r_gnd_r(net32[194:195]), .pgate_r(pgate_r[75:74]),
     .wl_r(wl_r[75:74]), .reset_b_r(reset_r[75:74]),
     .q(net36[776:783]), .q_b(net37[776:783]), .bl(bl[3:0]));
cram2x2x2 xcram_36_ ( .pgate_l(pgate_l[73:72]), .wl_l(wl_l[73:72]),
     .reset_b_l(reset_l[73:72]), .r_gnd_l(net43[196:197]),
     .r_gnd_r(net32[196:197]), .pgate_r(pgate_r[73:72]),
     .wl_r(wl_r[73:72]), .reset_b_r(reset_r[73:72]),
     .q(net36[784:791]), .q_b(net37[784:791]), .bl(bl[3:0]));
cram2x2x2 xcram_35_ ( .pgate_l(pgate_l[71:70]), .wl_l(wl_l[71:70]),
     .reset_b_l(reset_l[71:70]), .r_gnd_l(net43[198:199]),
     .r_gnd_r(net32[198:199]), .pgate_r(pgate_r[71:70]),
     .wl_r(wl_r[71:70]), .reset_b_r(reset_r[71:70]),
     .q(net36[792:799]), .q_b(net37[792:799]), .bl(bl[3:0]));
cram2x2x2 xcram_34_ ( .pgate_l(pgate_l[69:68]), .wl_l(wl_l[69:68]),
     .reset_b_l(reset_l[69:68]), .r_gnd_l(net43[200:201]),
     .r_gnd_r(net32[200:201]), .pgate_r(pgate_r[69:68]),
     .wl_r(wl_r[69:68]), .reset_b_r(reset_r[69:68]),
     .q(net36[800:807]), .q_b(net37[800:807]), .bl(bl[3:0]));
cram2x2x2 xcram_33_ ( .pgate_l(pgate_l[67:66]), .wl_l(wl_l[67:66]),
     .reset_b_l(reset_l[67:66]), .r_gnd_l(net43[202:203]),
     .r_gnd_r(net32[202:203]), .pgate_r(pgate_r[67:66]),
     .wl_r(wl_r[67:66]), .reset_b_r(reset_r[67:66]),
     .q(net36[808:815]), .q_b(net37[808:815]), .bl(bl[3:0]));
cram2x2x2 xcram_32_ ( .pgate_l(pgate_l[65:64]), .wl_l(wl_l[65:64]),
     .reset_b_l(reset_l[65:64]), .r_gnd_l(net43[204:205]),
     .r_gnd_r(net32[204:205]), .pgate_r(pgate_r[65:64]),
     .wl_r(wl_r[65:64]), .reset_b_r(reset_r[65:64]),
     .q(net36[816:823]), .q_b(net37[816:823]), .bl(bl[3:0]));
cram2x2x2 xcram_31_ ( .pgate_l(pgate_l[63:62]), .wl_l(wl_l[63:62]),
     .reset_b_l(reset_l[63:62]), .r_gnd_l(net43[206:207]),
     .r_gnd_r(net32[206:207]), .pgate_r(pgate_r[63:62]),
     .wl_r(wl_r[63:62]), .reset_b_r(reset_r[63:62]),
     .q(net36[824:831]), .q_b(net37[824:831]), .bl(bl[3:0]));
cram2x2x2 xcram_30_ ( .pgate_l(pgate_l[61:60]), .wl_l(wl_l[61:60]),
     .reset_b_l(reset_l[61:60]), .r_gnd_l(net43[208:209]),
     .r_gnd_r(net32[208:209]), .pgate_r(pgate_r[61:60]),
     .wl_r(wl_r[61:60]), .reset_b_r(reset_r[61:60]),
     .q(net36[832:839]), .q_b(net37[832:839]), .bl(bl[3:0]));
cram2x2x2 xcram_29_ ( .pgate_l(pgate_l[59:58]), .wl_l(wl_l[59:58]),
     .reset_b_l(reset_l[59:58]), .r_gnd_l(net43[210:211]),
     .r_gnd_r(net32[210:211]), .pgate_r(pgate_r[59:58]),
     .wl_r(wl_r[59:58]), .reset_b_r(reset_r[59:58]),
     .q(net36[840:847]), .q_b(net37[840:847]), .bl(bl[3:0]));
cram2x2x2 xcram_28_ ( .pgate_l(pgate_l[57:56]), .wl_l(wl_l[57:56]),
     .reset_b_l(reset_l[57:56]), .r_gnd_l(net43[212:213]),
     .r_gnd_r(net32[212:213]), .pgate_r(pgate_r[57:56]),
     .wl_r(wl_r[57:56]), .reset_b_r(reset_r[57:56]),
     .q(net36[848:855]), .q_b(net37[848:855]), .bl(bl[3:0]));
cram2x2x2 xcram_27_ ( .pgate_l(pgate_l[55:54]), .wl_l(wl_l[55:54]),
     .reset_b_l(reset_l[55:54]), .r_gnd_l(net43[214:215]),
     .r_gnd_r(net32[214:215]), .pgate_r(pgate_r[55:54]),
     .wl_r(wl_r[55:54]), .reset_b_r(reset_r[55:54]),
     .q(net36[856:863]), .q_b(net37[856:863]), .bl(bl[3:0]));
cram2x2x2 xcram_26_ ( .pgate_l(pgate_l[53:52]), .wl_l(wl_l[53:52]),
     .reset_b_l(reset_l[53:52]), .r_gnd_l(net43[216:217]),
     .r_gnd_r(net32[216:217]), .pgate_r(pgate_r[53:52]),
     .wl_r(wl_r[53:52]), .reset_b_r(reset_r[53:52]),
     .q(net36[864:871]), .q_b(net37[864:871]), .bl(bl[3:0]));
cram2x2x2 xcram_25_ ( .pgate_l(pgate_l[51:50]), .wl_l(wl_l[51:50]),
     .reset_b_l(reset_l[51:50]), .r_gnd_l(net43[218:219]),
     .r_gnd_r(net32[218:219]), .pgate_r(pgate_r[51:50]),
     .wl_r(wl_r[51:50]), .reset_b_r(reset_r[51:50]),
     .q(net36[872:879]), .q_b(net37[872:879]), .bl(bl[3:0]));
cram2x2x2 xcram_24_ ( .pgate_l(pgate_l[49:48]), .wl_l(wl_l[49:48]),
     .reset_b_l(reset_l[49:48]), .r_gnd_l(net43[220:221]),
     .r_gnd_r(net32[220:221]), .pgate_r(pgate_r[49:48]),
     .wl_r(wl_r[49:48]), .reset_b_r(reset_r[49:48]),
     .q(net36[880:887]), .q_b(net37[880:887]), .bl(bl[3:0]));
cram2x2x2 xcram_23_ ( .pgate_l(pgate_l[47:46]), .wl_l(wl_l[47:46]),
     .reset_b_l(reset_l[47:46]), .r_gnd_l(net43[222:223]),
     .r_gnd_r(net32[222:223]), .pgate_r(pgate_r[47:46]),
     .wl_r(wl_r[47:46]), .reset_b_r(reset_r[47:46]),
     .q(net36[888:895]), .q_b(net37[888:895]), .bl(bl[3:0]));
cram2x2x2 xcram_22_ ( .pgate_l(pgate_l[45:44]), .wl_l(wl_l[45:44]),
     .reset_b_l(reset_l[45:44]), .r_gnd_l(net43[224:225]),
     .r_gnd_r(net32[224:225]), .pgate_r(pgate_r[45:44]),
     .wl_r(wl_r[45:44]), .reset_b_r(reset_r[45:44]),
     .q(net36[896:903]), .q_b(net37[896:903]), .bl(bl[3:0]));
cram2x2x2 xcram_21_ ( .pgate_l(pgate_l[43:42]), .wl_l(wl_l[43:42]),
     .reset_b_l(reset_l[43:42]), .r_gnd_l(net43[226:227]),
     .r_gnd_r(net32[226:227]), .pgate_r(pgate_r[43:42]),
     .wl_r(wl_r[43:42]), .reset_b_r(reset_r[43:42]),
     .q(net36[904:911]), .q_b(net37[904:911]), .bl(bl[3:0]));
cram2x2x2 xcram_20_ ( .pgate_l(pgate_l[41:40]), .wl_l(wl_l[41:40]),
     .reset_b_l(reset_l[41:40]), .r_gnd_l(net43[228:229]),
     .r_gnd_r(net32[228:229]), .pgate_r(pgate_r[41:40]),
     .wl_r(wl_r[41:40]), .reset_b_r(reset_r[41:40]),
     .q(net36[912:919]), .q_b(net37[912:919]), .bl(bl[3:0]));
cram2x2x2 xcram_19_ ( .pgate_l(pgate_l[39:38]), .wl_l(wl_l[39:38]),
     .reset_b_l(reset_l[39:38]), .r_gnd_l(net43[230:231]),
     .r_gnd_r(net32[230:231]), .pgate_r(pgate_r[39:38]),
     .wl_r(wl_r[39:38]), .reset_b_r(reset_r[39:38]),
     .q(net36[920:927]), .q_b(net37[920:927]), .bl(bl[3:0]));
cram2x2x2 xcram_18_ ( .pgate_l(pgate_l[37:36]), .wl_l(wl_l[37:36]),
     .reset_b_l(reset_l[37:36]), .r_gnd_l(net43[232:233]),
     .r_gnd_r(net32[232:233]), .pgate_r(pgate_r[37:36]),
     .wl_r(wl_r[37:36]), .reset_b_r(reset_r[37:36]),
     .q(net36[928:935]), .q_b(net37[928:935]), .bl(bl[3:0]));
cram2x2x2 xcram_17_ ( .pgate_l(pgate_l[35:34]), .wl_l(wl_l[35:34]),
     .reset_b_l(reset_l[35:34]), .r_gnd_l(net43[234:235]),
     .r_gnd_r(net32[234:235]), .pgate_r(pgate_r[35:34]),
     .wl_r(wl_r[35:34]), .reset_b_r(reset_r[35:34]),
     .q(net36[936:943]), .q_b(net37[936:943]), .bl(bl[3:0]));
cram2x2x2 xcram_16_ ( .pgate_l(pgate_l[33:32]), .wl_l(wl_l[33:32]),
     .reset_b_l(reset_l[33:32]), .r_gnd_l(net43[236:237]),
     .r_gnd_r(net32[236:237]), .pgate_r(pgate_r[33:32]),
     .wl_r(wl_r[33:32]), .reset_b_r(reset_r[33:32]),
     .q(net36[944:951]), .q_b(net37[944:951]), .bl(bl[3:0]));
cram2x2x2 xcram_15_ ( .pgate_l(pgate_l[31:30]), .wl_l(wl_l[31:30]),
     .reset_b_l(reset_l[31:30]), .r_gnd_l(net43[238:239]),
     .r_gnd_r(net32[238:239]), .pgate_r(pgate_r[31:30]),
     .wl_r(wl_r[31:30]), .reset_b_r(reset_r[31:30]),
     .q(net36[952:959]), .q_b(net37[952:959]), .bl(bl[3:0]));
cram2x2x2 xcram_14_ ( .pgate_l(pgate_l[29:28]), .wl_l(wl_l[29:28]),
     .reset_b_l(reset_l[29:28]), .r_gnd_l(net43[240:241]),
     .r_gnd_r(net32[240:241]), .pgate_r(pgate_r[29:28]),
     .wl_r(wl_r[29:28]), .reset_b_r(reset_r[29:28]),
     .q(net36[960:967]), .q_b(net37[960:967]), .bl(bl[3:0]));
cram2x2x2 xcram_13_ ( .pgate_l(pgate_l[27:26]), .wl_l(wl_l[27:26]),
     .reset_b_l(reset_l[27:26]), .r_gnd_l(net43[242:243]),
     .r_gnd_r(net32[242:243]), .pgate_r(pgate_r[27:26]),
     .wl_r(wl_r[27:26]), .reset_b_r(reset_r[27:26]),
     .q(net36[968:975]), .q_b(net37[968:975]), .bl(bl[3:0]));
cram2x2x2 xcram_12_ ( .pgate_l(pgate_l[25:24]), .wl_l(wl_l[25:24]),
     .reset_b_l(reset_l[25:24]), .r_gnd_l(net43[244:245]),
     .r_gnd_r(net32[244:245]), .pgate_r(pgate_r[25:24]),
     .wl_r(wl_r[25:24]), .reset_b_r(reset_r[25:24]),
     .q(net36[976:983]), .q_b(net37[976:983]), .bl(bl[3:0]));
cram2x2x2 xcram_11_ ( .pgate_l(pgate_l[23:22]), .wl_l(wl_l[23:22]),
     .reset_b_l(reset_l[23:22]), .r_gnd_l(net43[246:247]),
     .r_gnd_r(net32[246:247]), .pgate_r(pgate_r[23:22]),
     .wl_r(wl_r[23:22]), .reset_b_r(reset_r[23:22]),
     .q(net36[984:991]), .q_b(net37[984:991]), .bl(bl[3:0]));
cram2x2x2 xcram_10_ ( .pgate_l(pgate_l[21:20]), .wl_l(wl_l[21:20]),
     .reset_b_l(reset_l[21:20]), .r_gnd_l(net43[248:249]),
     .r_gnd_r(net32[248:249]), .pgate_r(pgate_r[21:20]),
     .wl_r(wl_r[21:20]), .reset_b_r(reset_r[21:20]),
     .q(net36[992:999]), .q_b(net37[992:999]), .bl(bl[3:0]));
cram2x2x2 xcram_9_ ( .pgate_l(pgate_l[19:18]), .wl_l(wl_l[19:18]),
     .reset_b_l(reset_l[19:18]), .r_gnd_l(net43[250:251]),
     .r_gnd_r(net32[250:251]), .pgate_r(pgate_r[19:18]),
     .wl_r(wl_r[19:18]), .reset_b_r(reset_r[19:18]),
     .q(net36[1000:1007]), .q_b(net37[1000:1007]), .bl(bl[3:0]));
cram2x2x2 xcram_8_ ( .pgate_l(pgate_l[17:16]), .wl_l(wl_l[17:16]),
     .reset_b_l(reset_l[17:16]), .r_gnd_l(net43[252:253]),
     .r_gnd_r(net32[252:253]), .pgate_r(pgate_r[17:16]),
     .wl_r(wl_r[17:16]), .reset_b_r(reset_r[17:16]),
     .q(net36[1008:1015]), .q_b(net37[1008:1015]), .bl(bl[3:0]));
cram2x2x2 xcram_7_ ( .pgate_l(pgate_l[15:14]), .wl_l(wl_l[15:14]),
     .reset_b_l(reset_l[15:14]), .r_gnd_l(net43[254:255]),
     .r_gnd_r(net32[254:255]), .pgate_r(pgate_r[15:14]),
     .wl_r(wl_r[15:14]), .reset_b_r(reset_r[15:14]),
     .q(net36[1016:1023]), .q_b(net37[1016:1023]), .bl(bl[3:0]));
cram2x2x2 xcram_6_ ( .pgate_l(pgate_l[13:12]), .wl_l(wl_l[13:12]),
     .reset_b_l(reset_l[13:12]), .r_gnd_l(net43[256:257]),
     .r_gnd_r(net32[256:257]), .pgate_r(pgate_r[13:12]),
     .wl_r(wl_r[13:12]), .reset_b_r(reset_r[13:12]),
     .q(net36[1024:1031]), .q_b(net37[1024:1031]), .bl(bl[3:0]));
cram2x2x2 xcram_5_ ( .pgate_l(pgate_l[11:10]), .wl_l(wl_l[11:10]),
     .reset_b_l(reset_l[11:10]), .r_gnd_l(net43[258:259]),
     .r_gnd_r(net32[258:259]), .pgate_r(pgate_r[11:10]),
     .wl_r(wl_r[11:10]), .reset_b_r(reset_r[11:10]),
     .q(net36[1032:1039]), .q_b(net37[1032:1039]), .bl(bl[3:0]));
cram2x2x2 xcram_4_ ( .pgate_l(pgate_l[9:8]), .wl_l(wl_l[9:8]),
     .reset_b_l(reset_l[9:8]), .r_gnd_l(net43[260:261]),
     .r_gnd_r(net32[260:261]), .pgate_r(pgate_r[9:8]),
     .wl_r(wl_r[9:8]), .reset_b_r(reset_r[9:8]), .q(net36[1040:1047]),
     .q_b(net37[1040:1047]), .bl(bl[3:0]));
cram2x2x2 xcram_3_ ( .pgate_l(pgate_l[7:6]), .wl_l(wl_l[7:6]),
     .reset_b_l(reset_l[7:6]), .r_gnd_l(net43[262:263]),
     .r_gnd_r(net32[262:263]), .pgate_r(pgate_r[7:6]),
     .wl_r(wl_r[7:6]), .reset_b_r(reset_r[7:6]), .q(net36[1048:1055]),
     .q_b(net37[1048:1055]), .bl(bl[3:0]));
cram2x2x2 xcram_2_ ( .pgate_l(pgate_l[5:4]), .wl_l(wl_l[5:4]),
     .reset_b_l(reset_l[5:4]), .r_gnd_l(net43[264:265]),
     .r_gnd_r(net32[264:265]), .pgate_r(pgate_r[5:4]),
     .wl_r(wl_r[5:4]), .reset_b_r(reset_r[5:4]), .q(net36[1056:1063]),
     .q_b(net37[1056:1063]), .bl(bl[3:0]));
cram2x2x2 xcram_1_ ( .pgate_l(pgate_l[3:2]), .wl_l(wl_l[3:2]),
     .reset_b_l(reset_l[3:2]), .r_gnd_l(net43[266:267]),
     .r_gnd_r(net32[266:267]), .pgate_r(pgate_r[3:2]),
     .wl_r(wl_r[3:2]), .reset_b_r(reset_r[3:2]), .q(net36[1064:1071]),
     .q_b(net37[1064:1071]), .bl(bl[3:0]));
cram2x2x2 xcram_0_ ( .pgate_l(pgate_l[1:0]), .wl_l(wl_l[1:0]),
     .reset_b_l(reset_l[1:0]), .r_gnd_l(net43[268:269]),
     .r_gnd_r(net32[268:269]), .pgate_r(pgate_r[1:0]),
     .wl_r(wl_r[1:0]), .reset_b_r(reset_r[1:0]), .q(net36[1072:1079]),
     .q_b(net37[1072:1079]), .bl(bl[3:0]));
pch_hvt  M0_269_ ( .D(net32[0]), .B(vdd_), .G(vdd_cntl_r[269]),
     .S(vdd_));
pch_hvt  M0_268_ ( .D(net32[1]), .B(vdd_), .G(vdd_cntl_r[268]),
     .S(vdd_));
pch_hvt  M0_267_ ( .D(net32[2]), .B(vdd_), .G(vdd_cntl_r[267]),
     .S(vdd_));
pch_hvt  M0_266_ ( .D(net32[3]), .B(vdd_), .G(vdd_cntl_r[266]),
     .S(vdd_));
pch_hvt  M0_265_ ( .D(net32[4]), .B(vdd_), .G(vdd_cntl_r[265]),
     .S(vdd_));
pch_hvt  M0_264_ ( .D(net32[5]), .B(vdd_), .G(vdd_cntl_r[264]),
     .S(vdd_));
pch_hvt  M0_263_ ( .D(net32[6]), .B(vdd_), .G(vdd_cntl_r[263]),
     .S(vdd_));
pch_hvt  M0_262_ ( .D(net32[7]), .B(vdd_), .G(vdd_cntl_r[262]),
     .S(vdd_));
pch_hvt  M0_261_ ( .D(net32[8]), .B(vdd_), .G(vdd_cntl_r[261]),
     .S(vdd_));
pch_hvt  M0_260_ ( .D(net32[9]), .B(vdd_), .G(vdd_cntl_r[260]),
     .S(vdd_));
pch_hvt  M0_259_ ( .D(net32[10]), .B(vdd_), .G(vdd_cntl_r[259]),
     .S(vdd_));
pch_hvt  M0_258_ ( .D(net32[11]), .B(vdd_), .G(vdd_cntl_r[258]),
     .S(vdd_));
pch_hvt  M0_257_ ( .D(net32[12]), .B(vdd_), .G(vdd_cntl_r[257]),
     .S(vdd_));
pch_hvt  M0_256_ ( .D(net32[13]), .B(vdd_), .G(vdd_cntl_r[256]),
     .S(vdd_));
pch_hvt  M0_255_ ( .D(net32[14]), .B(vdd_), .G(vdd_cntl_r[255]),
     .S(vdd_));
pch_hvt  M0_254_ ( .D(net32[15]), .B(vdd_), .G(vdd_cntl_r[254]),
     .S(vdd_));
pch_hvt  M0_253_ ( .D(net32[16]), .B(vdd_), .G(vdd_cntl_r[253]),
     .S(vdd_));
pch_hvt  M0_252_ ( .D(net32[17]), .B(vdd_), .G(vdd_cntl_r[252]),
     .S(vdd_));
pch_hvt  M0_251_ ( .D(net32[18]), .B(vdd_), .G(vdd_cntl_r[251]),
     .S(vdd_));
pch_hvt  M0_250_ ( .D(net32[19]), .B(vdd_), .G(vdd_cntl_r[250]),
     .S(vdd_));
pch_hvt  M0_249_ ( .D(net32[20]), .B(vdd_), .G(vdd_cntl_r[249]),
     .S(vdd_));
pch_hvt  M0_248_ ( .D(net32[21]), .B(vdd_), .G(vdd_cntl_r[248]),
     .S(vdd_));
pch_hvt  M0_247_ ( .D(net32[22]), .B(vdd_), .G(vdd_cntl_r[247]),
     .S(vdd_));
pch_hvt  M0_246_ ( .D(net32[23]), .B(vdd_), .G(vdd_cntl_r[246]),
     .S(vdd_));
pch_hvt  M0_245_ ( .D(net32[24]), .B(vdd_), .G(vdd_cntl_r[245]),
     .S(vdd_));
pch_hvt  M0_244_ ( .D(net32[25]), .B(vdd_), .G(vdd_cntl_r[244]),
     .S(vdd_));
pch_hvt  M0_243_ ( .D(net32[26]), .B(vdd_), .G(vdd_cntl_r[243]),
     .S(vdd_));
pch_hvt  M0_242_ ( .D(net32[27]), .B(vdd_), .G(vdd_cntl_r[242]),
     .S(vdd_));
pch_hvt  M0_241_ ( .D(net32[28]), .B(vdd_), .G(vdd_cntl_r[241]),
     .S(vdd_));
pch_hvt  M0_240_ ( .D(net32[29]), .B(vdd_), .G(vdd_cntl_r[240]),
     .S(vdd_));
pch_hvt  M0_239_ ( .D(net32[30]), .B(vdd_), .G(vdd_cntl_r[239]),
     .S(vdd_));
pch_hvt  M0_238_ ( .D(net32[31]), .B(vdd_), .G(vdd_cntl_r[238]),
     .S(vdd_));
pch_hvt  M0_237_ ( .D(net32[32]), .B(vdd_), .G(vdd_cntl_r[237]),
     .S(vdd_));
pch_hvt  M0_236_ ( .D(net32[33]), .B(vdd_), .G(vdd_cntl_r[236]),
     .S(vdd_));
pch_hvt  M0_235_ ( .D(net32[34]), .B(vdd_), .G(vdd_cntl_r[235]),
     .S(vdd_));
pch_hvt  M0_234_ ( .D(net32[35]), .B(vdd_), .G(vdd_cntl_r[234]),
     .S(vdd_));
pch_hvt  M0_233_ ( .D(net32[36]), .B(vdd_), .G(vdd_cntl_r[233]),
     .S(vdd_));
pch_hvt  M0_232_ ( .D(net32[37]), .B(vdd_), .G(vdd_cntl_r[232]),
     .S(vdd_));
pch_hvt  M0_231_ ( .D(net32[38]), .B(vdd_), .G(vdd_cntl_r[231]),
     .S(vdd_));
pch_hvt  M0_230_ ( .D(net32[39]), .B(vdd_), .G(vdd_cntl_r[230]),
     .S(vdd_));
pch_hvt  M0_229_ ( .D(net32[40]), .B(vdd_), .G(vdd_cntl_r[229]),
     .S(vdd_));
pch_hvt  M0_228_ ( .D(net32[41]), .B(vdd_), .G(vdd_cntl_r[228]),
     .S(vdd_));
pch_hvt  M0_227_ ( .D(net32[42]), .B(vdd_), .G(vdd_cntl_r[227]),
     .S(vdd_));
pch_hvt  M0_226_ ( .D(net32[43]), .B(vdd_), .G(vdd_cntl_r[226]),
     .S(vdd_));
pch_hvt  M0_225_ ( .D(net32[44]), .B(vdd_), .G(vdd_cntl_r[225]),
     .S(vdd_));
pch_hvt  M0_224_ ( .D(net32[45]), .B(vdd_), .G(vdd_cntl_r[224]),
     .S(vdd_));
pch_hvt  M0_223_ ( .D(net32[46]), .B(vdd_), .G(vdd_cntl_r[223]),
     .S(vdd_));
pch_hvt  M0_222_ ( .D(net32[47]), .B(vdd_), .G(vdd_cntl_r[222]),
     .S(vdd_));
pch_hvt  M0_221_ ( .D(net32[48]), .B(vdd_), .G(vdd_cntl_r[221]),
     .S(vdd_));
pch_hvt  M0_220_ ( .D(net32[49]), .B(vdd_), .G(vdd_cntl_r[220]),
     .S(vdd_));
pch_hvt  M0_219_ ( .D(net32[50]), .B(vdd_), .G(vdd_cntl_r[219]),
     .S(vdd_));
pch_hvt  M0_218_ ( .D(net32[51]), .B(vdd_), .G(vdd_cntl_r[218]),
     .S(vdd_));
pch_hvt  M0_217_ ( .D(net32[52]), .B(vdd_), .G(vdd_cntl_r[217]),
     .S(vdd_));
pch_hvt  M0_216_ ( .D(net32[53]), .B(vdd_), .G(vdd_cntl_r[216]),
     .S(vdd_));
pch_hvt  M0_215_ ( .D(net32[54]), .B(vdd_), .G(vdd_cntl_r[215]),
     .S(vdd_));
pch_hvt  M0_214_ ( .D(net32[55]), .B(vdd_), .G(vdd_cntl_r[214]),
     .S(vdd_));
pch_hvt  M0_213_ ( .D(net32[56]), .B(vdd_), .G(vdd_cntl_r[213]),
     .S(vdd_));
pch_hvt  M0_212_ ( .D(net32[57]), .B(vdd_), .G(vdd_cntl_r[212]),
     .S(vdd_));
pch_hvt  M0_211_ ( .D(net32[58]), .B(vdd_), .G(vdd_cntl_r[211]),
     .S(vdd_));
pch_hvt  M0_210_ ( .D(net32[59]), .B(vdd_), .G(vdd_cntl_r[210]),
     .S(vdd_));
pch_hvt  M0_209_ ( .D(net32[60]), .B(vdd_), .G(vdd_cntl_r[209]),
     .S(vdd_));
pch_hvt  M0_208_ ( .D(net32[61]), .B(vdd_), .G(vdd_cntl_r[208]),
     .S(vdd_));
pch_hvt  M0_207_ ( .D(net32[62]), .B(vdd_), .G(vdd_cntl_r[207]),
     .S(vdd_));
pch_hvt  M0_206_ ( .D(net32[63]), .B(vdd_), .G(vdd_cntl_r[206]),
     .S(vdd_));
pch_hvt  M0_205_ ( .D(net32[64]), .B(vdd_), .G(vdd_cntl_r[205]),
     .S(vdd_));
pch_hvt  M0_204_ ( .D(net32[65]), .B(vdd_), .G(vdd_cntl_r[204]),
     .S(vdd_));
pch_hvt  M0_203_ ( .D(net32[66]), .B(vdd_), .G(vdd_cntl_r[203]),
     .S(vdd_));
pch_hvt  M0_202_ ( .D(net32[67]), .B(vdd_), .G(vdd_cntl_r[202]),
     .S(vdd_));
pch_hvt  M0_201_ ( .D(net32[68]), .B(vdd_), .G(vdd_cntl_r[201]),
     .S(vdd_));
pch_hvt  M0_200_ ( .D(net32[69]), .B(vdd_), .G(vdd_cntl_r[200]),
     .S(vdd_));
pch_hvt  M0_199_ ( .D(net32[70]), .B(vdd_), .G(vdd_cntl_r[199]),
     .S(vdd_));
pch_hvt  M0_198_ ( .D(net32[71]), .B(vdd_), .G(vdd_cntl_r[198]),
     .S(vdd_));
pch_hvt  M0_197_ ( .D(net32[72]), .B(vdd_), .G(vdd_cntl_r[197]),
     .S(vdd_));
pch_hvt  M0_196_ ( .D(net32[73]), .B(vdd_), .G(vdd_cntl_r[196]),
     .S(vdd_));
pch_hvt  M0_195_ ( .D(net32[74]), .B(vdd_), .G(vdd_cntl_r[195]),
     .S(vdd_));
pch_hvt  M0_194_ ( .D(net32[75]), .B(vdd_), .G(vdd_cntl_r[194]),
     .S(vdd_));
pch_hvt  M0_193_ ( .D(net32[76]), .B(vdd_), .G(vdd_cntl_r[193]),
     .S(vdd_));
pch_hvt  M0_192_ ( .D(net32[77]), .B(vdd_), .G(vdd_cntl_r[192]),
     .S(vdd_));
pch_hvt  M0_191_ ( .D(net32[78]), .B(vdd_), .G(vdd_cntl_r[191]),
     .S(vdd_));
pch_hvt  M0_190_ ( .D(net32[79]), .B(vdd_), .G(vdd_cntl_r[190]),
     .S(vdd_));
pch_hvt  M0_189_ ( .D(net32[80]), .B(vdd_), .G(vdd_cntl_r[189]),
     .S(vdd_));
pch_hvt  M0_188_ ( .D(net32[81]), .B(vdd_), .G(vdd_cntl_r[188]),
     .S(vdd_));
pch_hvt  M0_187_ ( .D(net32[82]), .B(vdd_), .G(vdd_cntl_r[187]),
     .S(vdd_));
pch_hvt  M0_186_ ( .D(net32[83]), .B(vdd_), .G(vdd_cntl_r[186]),
     .S(vdd_));
pch_hvt  M0_185_ ( .D(net32[84]), .B(vdd_), .G(vdd_cntl_r[185]),
     .S(vdd_));
pch_hvt  M0_184_ ( .D(net32[85]), .B(vdd_), .G(vdd_cntl_r[184]),
     .S(vdd_));
pch_hvt  M0_183_ ( .D(net32[86]), .B(vdd_), .G(vdd_cntl_r[183]),
     .S(vdd_));
pch_hvt  M0_182_ ( .D(net32[87]), .B(vdd_), .G(vdd_cntl_r[182]),
     .S(vdd_));
pch_hvt  M0_181_ ( .D(net32[88]), .B(vdd_), .G(vdd_cntl_r[181]),
     .S(vdd_));
pch_hvt  M0_180_ ( .D(net32[89]), .B(vdd_), .G(vdd_cntl_r[180]),
     .S(vdd_));
pch_hvt  M0_179_ ( .D(net32[90]), .B(vdd_), .G(vdd_cntl_r[179]),
     .S(vdd_));
pch_hvt  M0_178_ ( .D(net32[91]), .B(vdd_), .G(vdd_cntl_r[178]),
     .S(vdd_));
pch_hvt  M0_177_ ( .D(net32[92]), .B(vdd_), .G(vdd_cntl_r[177]),
     .S(vdd_));
pch_hvt  M0_176_ ( .D(net32[93]), .B(vdd_), .G(vdd_cntl_r[176]),
     .S(vdd_));
pch_hvt  M0_175_ ( .D(net32[94]), .B(vdd_), .G(vdd_cntl_r[175]),
     .S(vdd_));
pch_hvt  M0_174_ ( .D(net32[95]), .B(vdd_), .G(vdd_cntl_r[174]),
     .S(vdd_));
pch_hvt  M0_173_ ( .D(net32[96]), .B(vdd_), .G(vdd_cntl_r[173]),
     .S(vdd_));
pch_hvt  M0_172_ ( .D(net32[97]), .B(vdd_), .G(vdd_cntl_r[172]),
     .S(vdd_));
pch_hvt  M0_171_ ( .D(net32[98]), .B(vdd_), .G(vdd_cntl_r[171]),
     .S(vdd_));
pch_hvt  M0_170_ ( .D(net32[99]), .B(vdd_), .G(vdd_cntl_r[170]),
     .S(vdd_));
pch_hvt  M0_169_ ( .D(net32[100]), .B(vdd_), .G(vdd_cntl_r[169]),
     .S(vdd_));
pch_hvt  M0_168_ ( .D(net32[101]), .B(vdd_), .G(vdd_cntl_r[168]),
     .S(vdd_));
pch_hvt  M0_167_ ( .D(net32[102]), .B(vdd_), .G(vdd_cntl_r[167]),
     .S(vdd_));
pch_hvt  M0_166_ ( .D(net32[103]), .B(vdd_), .G(vdd_cntl_r[166]),
     .S(vdd_));
pch_hvt  M0_165_ ( .D(net32[104]), .B(vdd_), .G(vdd_cntl_r[165]),
     .S(vdd_));
pch_hvt  M0_164_ ( .D(net32[105]), .B(vdd_), .G(vdd_cntl_r[164]),
     .S(vdd_));
pch_hvt  M0_163_ ( .D(net32[106]), .B(vdd_), .G(vdd_cntl_r[163]),
     .S(vdd_));
pch_hvt  M0_162_ ( .D(net32[107]), .B(vdd_), .G(vdd_cntl_r[162]),
     .S(vdd_));
pch_hvt  M0_161_ ( .D(net32[108]), .B(vdd_), .G(vdd_cntl_r[161]),
     .S(vdd_));
pch_hvt  M0_160_ ( .D(net32[109]), .B(vdd_), .G(vdd_cntl_r[160]),
     .S(vdd_));
pch_hvt  M0_159_ ( .D(net32[110]), .B(vdd_), .G(vdd_cntl_r[159]),
     .S(vdd_));
pch_hvt  M0_158_ ( .D(net32[111]), .B(vdd_), .G(vdd_cntl_r[158]),
     .S(vdd_));
pch_hvt  M0_157_ ( .D(net32[112]), .B(vdd_), .G(vdd_cntl_r[157]),
     .S(vdd_));
pch_hvt  M0_156_ ( .D(net32[113]), .B(vdd_), .G(vdd_cntl_r[156]),
     .S(vdd_));
pch_hvt  M0_155_ ( .D(net32[114]), .B(vdd_), .G(vdd_cntl_r[155]),
     .S(vdd_));
pch_hvt  M0_154_ ( .D(net32[115]), .B(vdd_), .G(vdd_cntl_r[154]),
     .S(vdd_));
pch_hvt  M0_153_ ( .D(net32[116]), .B(vdd_), .G(vdd_cntl_r[153]),
     .S(vdd_));
pch_hvt  M0_152_ ( .D(net32[117]), .B(vdd_), .G(vdd_cntl_r[152]),
     .S(vdd_));
pch_hvt  M0_151_ ( .D(net32[118]), .B(vdd_), .G(vdd_cntl_r[151]),
     .S(vdd_));
pch_hvt  M0_150_ ( .D(net32[119]), .B(vdd_), .G(vdd_cntl_r[150]),
     .S(vdd_));
pch_hvt  M0_149_ ( .D(net32[120]), .B(vdd_), .G(vdd_cntl_r[149]),
     .S(vdd_));
pch_hvt  M0_148_ ( .D(net32[121]), .B(vdd_), .G(vdd_cntl_r[148]),
     .S(vdd_));
pch_hvt  M0_147_ ( .D(net32[122]), .B(vdd_), .G(vdd_cntl_r[147]),
     .S(vdd_));
pch_hvt  M0_146_ ( .D(net32[123]), .B(vdd_), .G(vdd_cntl_r[146]),
     .S(vdd_));
pch_hvt  M0_145_ ( .D(net32[124]), .B(vdd_), .G(vdd_cntl_r[145]),
     .S(vdd_));
pch_hvt  M0_144_ ( .D(net32[125]), .B(vdd_), .G(vdd_cntl_r[144]),
     .S(vdd_));
pch_hvt  M0_143_ ( .D(net32[126]), .B(vdd_), .G(vdd_cntl_r[143]),
     .S(vdd_));
pch_hvt  M0_142_ ( .D(net32[127]), .B(vdd_), .G(vdd_cntl_r[142]),
     .S(vdd_));
pch_hvt  M0_141_ ( .D(net32[128]), .B(vdd_), .G(vdd_cntl_r[141]),
     .S(vdd_));
pch_hvt  M0_140_ ( .D(net32[129]), .B(vdd_), .G(vdd_cntl_r[140]),
     .S(vdd_));
pch_hvt  M0_139_ ( .D(net32[130]), .B(vdd_), .G(vdd_cntl_r[139]),
     .S(vdd_));
pch_hvt  M0_138_ ( .D(net32[131]), .B(vdd_), .G(vdd_cntl_r[138]),
     .S(vdd_));
pch_hvt  M0_137_ ( .D(net32[132]), .B(vdd_), .G(vdd_cntl_r[137]),
     .S(vdd_));
pch_hvt  M0_136_ ( .D(net32[133]), .B(vdd_), .G(vdd_cntl_r[136]),
     .S(vdd_));
pch_hvt  M0_135_ ( .D(net32[134]), .B(vdd_), .G(vdd_cntl_r[135]),
     .S(vdd_));
pch_hvt  M0_134_ ( .D(net32[135]), .B(vdd_), .G(vdd_cntl_r[134]),
     .S(vdd_));
pch_hvt  M0_133_ ( .D(net32[136]), .B(vdd_), .G(vdd_cntl_r[133]),
     .S(vdd_));
pch_hvt  M0_132_ ( .D(net32[137]), .B(vdd_), .G(vdd_cntl_r[132]),
     .S(vdd_));
pch_hvt  M0_131_ ( .D(net32[138]), .B(vdd_), .G(vdd_cntl_r[131]),
     .S(vdd_));
pch_hvt  M0_130_ ( .D(net32[139]), .B(vdd_), .G(vdd_cntl_r[130]),
     .S(vdd_));
pch_hvt  M0_129_ ( .D(net32[140]), .B(vdd_), .G(vdd_cntl_r[129]),
     .S(vdd_));
pch_hvt  M0_128_ ( .D(net32[141]), .B(vdd_), .G(vdd_cntl_r[128]),
     .S(vdd_));
pch_hvt  M0_127_ ( .D(net32[142]), .B(vdd_), .G(vdd_cntl_r[127]),
     .S(vdd_));
pch_hvt  M0_126_ ( .D(net32[143]), .B(vdd_), .G(vdd_cntl_r[126]),
     .S(vdd_));
pch_hvt  M0_125_ ( .D(net32[144]), .B(vdd_), .G(vdd_cntl_r[125]),
     .S(vdd_));
pch_hvt  M0_124_ ( .D(net32[145]), .B(vdd_), .G(vdd_cntl_r[124]),
     .S(vdd_));
pch_hvt  M0_123_ ( .D(net32[146]), .B(vdd_), .G(vdd_cntl_r[123]),
     .S(vdd_));
pch_hvt  M0_122_ ( .D(net32[147]), .B(vdd_), .G(vdd_cntl_r[122]),
     .S(vdd_));
pch_hvt  M0_121_ ( .D(net32[148]), .B(vdd_), .G(vdd_cntl_r[121]),
     .S(vdd_));
pch_hvt  M0_120_ ( .D(net32[149]), .B(vdd_), .G(vdd_cntl_r[120]),
     .S(vdd_));
pch_hvt  M0_119_ ( .D(net32[150]), .B(vdd_), .G(vdd_cntl_r[119]),
     .S(vdd_));
pch_hvt  M0_118_ ( .D(net32[151]), .B(vdd_), .G(vdd_cntl_r[118]),
     .S(vdd_));
pch_hvt  M0_117_ ( .D(net32[152]), .B(vdd_), .G(vdd_cntl_r[117]),
     .S(vdd_));
pch_hvt  M0_116_ ( .D(net32[153]), .B(vdd_), .G(vdd_cntl_r[116]),
     .S(vdd_));
pch_hvt  M0_115_ ( .D(net32[154]), .B(vdd_), .G(vdd_cntl_r[115]),
     .S(vdd_));
pch_hvt  M0_114_ ( .D(net32[155]), .B(vdd_), .G(vdd_cntl_r[114]),
     .S(vdd_));
pch_hvt  M0_113_ ( .D(net32[156]), .B(vdd_), .G(vdd_cntl_r[113]),
     .S(vdd_));
pch_hvt  M0_112_ ( .D(net32[157]), .B(vdd_), .G(vdd_cntl_r[112]),
     .S(vdd_));
pch_hvt  M0_111_ ( .D(net32[158]), .B(vdd_), .G(vdd_cntl_r[111]),
     .S(vdd_));
pch_hvt  M0_110_ ( .D(net32[159]), .B(vdd_), .G(vdd_cntl_r[110]),
     .S(vdd_));
pch_hvt  M0_109_ ( .D(net32[160]), .B(vdd_), .G(vdd_cntl_r[109]),
     .S(vdd_));
pch_hvt  M0_108_ ( .D(net32[161]), .B(vdd_), .G(vdd_cntl_r[108]),
     .S(vdd_));
pch_hvt  M0_107_ ( .D(net32[162]), .B(vdd_), .G(vdd_cntl_r[107]),
     .S(vdd_));
pch_hvt  M0_106_ ( .D(net32[163]), .B(vdd_), .G(vdd_cntl_r[106]),
     .S(vdd_));
pch_hvt  M0_105_ ( .D(net32[164]), .B(vdd_), .G(vdd_cntl_r[105]),
     .S(vdd_));
pch_hvt  M0_104_ ( .D(net32[165]), .B(vdd_), .G(vdd_cntl_r[104]),
     .S(vdd_));
pch_hvt  M0_103_ ( .D(net32[166]), .B(vdd_), .G(vdd_cntl_r[103]),
     .S(vdd_));
pch_hvt  M0_102_ ( .D(net32[167]), .B(vdd_), .G(vdd_cntl_r[102]),
     .S(vdd_));
pch_hvt  M0_101_ ( .D(net32[168]), .B(vdd_), .G(vdd_cntl_r[101]),
     .S(vdd_));
pch_hvt  M0_100_ ( .D(net32[169]), .B(vdd_), .G(vdd_cntl_r[100]),
     .S(vdd_));
pch_hvt  M0_99_ ( .D(net32[170]), .B(vdd_), .G(vdd_cntl_r[99]),
     .S(vdd_));
pch_hvt  M0_98_ ( .D(net32[171]), .B(vdd_), .G(vdd_cntl_r[98]),
     .S(vdd_));
pch_hvt  M0_97_ ( .D(net32[172]), .B(vdd_), .G(vdd_cntl_r[97]),
     .S(vdd_));
pch_hvt  M0_96_ ( .D(net32[173]), .B(vdd_), .G(vdd_cntl_r[96]),
     .S(vdd_));
pch_hvt  M0_95_ ( .D(net32[174]), .B(vdd_), .G(vdd_cntl_r[95]),
     .S(vdd_));
pch_hvt  M0_94_ ( .D(net32[175]), .B(vdd_), .G(vdd_cntl_r[94]),
     .S(vdd_));
pch_hvt  M0_93_ ( .D(net32[176]), .B(vdd_), .G(vdd_cntl_r[93]),
     .S(vdd_));
pch_hvt  M0_92_ ( .D(net32[177]), .B(vdd_), .G(vdd_cntl_r[92]),
     .S(vdd_));
pch_hvt  M0_91_ ( .D(net32[178]), .B(vdd_), .G(vdd_cntl_r[91]),
     .S(vdd_));
pch_hvt  M0_90_ ( .D(net32[179]), .B(vdd_), .G(vdd_cntl_r[90]),
     .S(vdd_));
pch_hvt  M0_89_ ( .D(net32[180]), .B(vdd_), .G(vdd_cntl_r[89]),
     .S(vdd_));
pch_hvt  M0_88_ ( .D(net32[181]), .B(vdd_), .G(vdd_cntl_r[88]),
     .S(vdd_));
pch_hvt  M0_87_ ( .D(net32[182]), .B(vdd_), .G(vdd_cntl_r[87]),
     .S(vdd_));
pch_hvt  M0_86_ ( .D(net32[183]), .B(vdd_), .G(vdd_cntl_r[86]),
     .S(vdd_));
pch_hvt  M0_85_ ( .D(net32[184]), .B(vdd_), .G(vdd_cntl_r[85]),
     .S(vdd_));
pch_hvt  M0_84_ ( .D(net32[185]), .B(vdd_), .G(vdd_cntl_r[84]),
     .S(vdd_));
pch_hvt  M0_83_ ( .D(net32[186]), .B(vdd_), .G(vdd_cntl_r[83]),
     .S(vdd_));
pch_hvt  M0_82_ ( .D(net32[187]), .B(vdd_), .G(vdd_cntl_r[82]),
     .S(vdd_));
pch_hvt  M0_81_ ( .D(net32[188]), .B(vdd_), .G(vdd_cntl_r[81]),
     .S(vdd_));
pch_hvt  M0_80_ ( .D(net32[189]), .B(vdd_), .G(vdd_cntl_r[80]),
     .S(vdd_));
pch_hvt  M0_79_ ( .D(net32[190]), .B(vdd_), .G(vdd_cntl_r[79]),
     .S(vdd_));
pch_hvt  M0_78_ ( .D(net32[191]), .B(vdd_), .G(vdd_cntl_r[78]),
     .S(vdd_));
pch_hvt  M0_77_ ( .D(net32[192]), .B(vdd_), .G(vdd_cntl_r[77]),
     .S(vdd_));
pch_hvt  M0_76_ ( .D(net32[193]), .B(vdd_), .G(vdd_cntl_r[76]),
     .S(vdd_));
pch_hvt  M0_75_ ( .D(net32[194]), .B(vdd_), .G(vdd_cntl_r[75]),
     .S(vdd_));
pch_hvt  M0_74_ ( .D(net32[195]), .B(vdd_), .G(vdd_cntl_r[74]),
     .S(vdd_));
pch_hvt  M0_73_ ( .D(net32[196]), .B(vdd_), .G(vdd_cntl_r[73]),
     .S(vdd_));
pch_hvt  M0_72_ ( .D(net32[197]), .B(vdd_), .G(vdd_cntl_r[72]),
     .S(vdd_));
pch_hvt  M0_71_ ( .D(net32[198]), .B(vdd_), .G(vdd_cntl_r[71]),
     .S(vdd_));
pch_hvt  M0_70_ ( .D(net32[199]), .B(vdd_), .G(vdd_cntl_r[70]),
     .S(vdd_));
pch_hvt  M0_69_ ( .D(net32[200]), .B(vdd_), .G(vdd_cntl_r[69]),
     .S(vdd_));
pch_hvt  M0_68_ ( .D(net32[201]), .B(vdd_), .G(vdd_cntl_r[68]),
     .S(vdd_));
pch_hvt  M0_67_ ( .D(net32[202]), .B(vdd_), .G(vdd_cntl_r[67]),
     .S(vdd_));
pch_hvt  M0_66_ ( .D(net32[203]), .B(vdd_), .G(vdd_cntl_r[66]),
     .S(vdd_));
pch_hvt  M0_65_ ( .D(net32[204]), .B(vdd_), .G(vdd_cntl_r[65]),
     .S(vdd_));
pch_hvt  M0_64_ ( .D(net32[205]), .B(vdd_), .G(vdd_cntl_r[64]),
     .S(vdd_));
pch_hvt  M0_63_ ( .D(net32[206]), .B(vdd_), .G(vdd_cntl_r[63]),
     .S(vdd_));
pch_hvt  M0_62_ ( .D(net32[207]), .B(vdd_), .G(vdd_cntl_r[62]),
     .S(vdd_));
pch_hvt  M0_61_ ( .D(net32[208]), .B(vdd_), .G(vdd_cntl_r[61]),
     .S(vdd_));
pch_hvt  M0_60_ ( .D(net32[209]), .B(vdd_), .G(vdd_cntl_r[60]),
     .S(vdd_));
pch_hvt  M0_59_ ( .D(net32[210]), .B(vdd_), .G(vdd_cntl_r[59]),
     .S(vdd_));
pch_hvt  M0_58_ ( .D(net32[211]), .B(vdd_), .G(vdd_cntl_r[58]),
     .S(vdd_));
pch_hvt  M0_57_ ( .D(net32[212]), .B(vdd_), .G(vdd_cntl_r[57]),
     .S(vdd_));
pch_hvt  M0_56_ ( .D(net32[213]), .B(vdd_), .G(vdd_cntl_r[56]),
     .S(vdd_));
pch_hvt  M0_55_ ( .D(net32[214]), .B(vdd_), .G(vdd_cntl_r[55]),
     .S(vdd_));
pch_hvt  M0_54_ ( .D(net32[215]), .B(vdd_), .G(vdd_cntl_r[54]),
     .S(vdd_));
pch_hvt  M0_53_ ( .D(net32[216]), .B(vdd_), .G(vdd_cntl_r[53]),
     .S(vdd_));
pch_hvt  M0_52_ ( .D(net32[217]), .B(vdd_), .G(vdd_cntl_r[52]),
     .S(vdd_));
pch_hvt  M0_51_ ( .D(net32[218]), .B(vdd_), .G(vdd_cntl_r[51]),
     .S(vdd_));
pch_hvt  M0_50_ ( .D(net32[219]), .B(vdd_), .G(vdd_cntl_r[50]),
     .S(vdd_));
pch_hvt  M0_49_ ( .D(net32[220]), .B(vdd_), .G(vdd_cntl_r[49]),
     .S(vdd_));
pch_hvt  M0_48_ ( .D(net32[221]), .B(vdd_), .G(vdd_cntl_r[48]),
     .S(vdd_));
pch_hvt  M0_47_ ( .D(net32[222]), .B(vdd_), .G(vdd_cntl_r[47]),
     .S(vdd_));
pch_hvt  M0_46_ ( .D(net32[223]), .B(vdd_), .G(vdd_cntl_r[46]),
     .S(vdd_));
pch_hvt  M0_45_ ( .D(net32[224]), .B(vdd_), .G(vdd_cntl_r[45]),
     .S(vdd_));
pch_hvt  M0_44_ ( .D(net32[225]), .B(vdd_), .G(vdd_cntl_r[44]),
     .S(vdd_));
pch_hvt  M0_43_ ( .D(net32[226]), .B(vdd_), .G(vdd_cntl_r[43]),
     .S(vdd_));
pch_hvt  M0_42_ ( .D(net32[227]), .B(vdd_), .G(vdd_cntl_r[42]),
     .S(vdd_));
pch_hvt  M0_41_ ( .D(net32[228]), .B(vdd_), .G(vdd_cntl_r[41]),
     .S(vdd_));
pch_hvt  M0_40_ ( .D(net32[229]), .B(vdd_), .G(vdd_cntl_r[40]),
     .S(vdd_));
pch_hvt  M0_39_ ( .D(net32[230]), .B(vdd_), .G(vdd_cntl_r[39]),
     .S(vdd_));
pch_hvt  M0_38_ ( .D(net32[231]), .B(vdd_), .G(vdd_cntl_r[38]),
     .S(vdd_));
pch_hvt  M0_37_ ( .D(net32[232]), .B(vdd_), .G(vdd_cntl_r[37]),
     .S(vdd_));
pch_hvt  M0_36_ ( .D(net32[233]), .B(vdd_), .G(vdd_cntl_r[36]),
     .S(vdd_));
pch_hvt  M0_35_ ( .D(net32[234]), .B(vdd_), .G(vdd_cntl_r[35]),
     .S(vdd_));
pch_hvt  M0_34_ ( .D(net32[235]), .B(vdd_), .G(vdd_cntl_r[34]),
     .S(vdd_));
pch_hvt  M0_33_ ( .D(net32[236]), .B(vdd_), .G(vdd_cntl_r[33]),
     .S(vdd_));
pch_hvt  M0_32_ ( .D(net32[237]), .B(vdd_), .G(vdd_cntl_r[32]),
     .S(vdd_));
pch_hvt  M0_31_ ( .D(net32[238]), .B(vdd_), .G(vdd_cntl_r[31]),
     .S(vdd_));
pch_hvt  M0_30_ ( .D(net32[239]), .B(vdd_), .G(vdd_cntl_r[30]),
     .S(vdd_));
pch_hvt  M0_29_ ( .D(net32[240]), .B(vdd_), .G(vdd_cntl_r[29]),
     .S(vdd_));
pch_hvt  M0_28_ ( .D(net32[241]), .B(vdd_), .G(vdd_cntl_r[28]),
     .S(vdd_));
pch_hvt  M0_27_ ( .D(net32[242]), .B(vdd_), .G(vdd_cntl_r[27]),
     .S(vdd_));
pch_hvt  M0_26_ ( .D(net32[243]), .B(vdd_), .G(vdd_cntl_r[26]),
     .S(vdd_));
pch_hvt  M0_25_ ( .D(net32[244]), .B(vdd_), .G(vdd_cntl_r[25]),
     .S(vdd_));
pch_hvt  M0_24_ ( .D(net32[245]), .B(vdd_), .G(vdd_cntl_r[24]),
     .S(vdd_));
pch_hvt  M0_23_ ( .D(net32[246]), .B(vdd_), .G(vdd_cntl_r[23]),
     .S(vdd_));
pch_hvt  M0_22_ ( .D(net32[247]), .B(vdd_), .G(vdd_cntl_r[22]),
     .S(vdd_));
pch_hvt  M0_21_ ( .D(net32[248]), .B(vdd_), .G(vdd_cntl_r[21]),
     .S(vdd_));
pch_hvt  M0_20_ ( .D(net32[249]), .B(vdd_), .G(vdd_cntl_r[20]),
     .S(vdd_));
pch_hvt  M0_19_ ( .D(net32[250]), .B(vdd_), .G(vdd_cntl_r[19]),
     .S(vdd_));
pch_hvt  M0_18_ ( .D(net32[251]), .B(vdd_), .G(vdd_cntl_r[18]),
     .S(vdd_));
pch_hvt  M0_17_ ( .D(net32[252]), .B(vdd_), .G(vdd_cntl_r[17]),
     .S(vdd_));
pch_hvt  M0_16_ ( .D(net32[253]), .B(vdd_), .G(vdd_cntl_r[16]),
     .S(vdd_));
pch_hvt  M0_15_ ( .D(net32[254]), .B(vdd_), .G(vdd_cntl_r[15]),
     .S(vdd_));
pch_hvt  M0_14_ ( .D(net32[255]), .B(vdd_), .G(vdd_cntl_r[14]),
     .S(vdd_));
pch_hvt  M0_13_ ( .D(net32[256]), .B(vdd_), .G(vdd_cntl_r[13]),
     .S(vdd_));
pch_hvt  M0_12_ ( .D(net32[257]), .B(vdd_), .G(vdd_cntl_r[12]),
     .S(vdd_));
pch_hvt  M0_11_ ( .D(net32[258]), .B(vdd_), .G(vdd_cntl_r[11]),
     .S(vdd_));
pch_hvt  M0_10_ ( .D(net32[259]), .B(vdd_), .G(vdd_cntl_r[10]),
     .S(vdd_));
pch_hvt  M0_9_ ( .D(net32[260]), .B(vdd_), .G(vdd_cntl_r[9]),
     .S(vdd_));
pch_hvt  M0_8_ ( .D(net32[261]), .B(vdd_), .G(vdd_cntl_r[8]),
     .S(vdd_));
pch_hvt  M0_7_ ( .D(net32[262]), .B(vdd_), .G(vdd_cntl_r[7]),
     .S(vdd_));
pch_hvt  M0_6_ ( .D(net32[263]), .B(vdd_), .G(vdd_cntl_r[6]),
     .S(vdd_));
pch_hvt  M0_5_ ( .D(net32[264]), .B(vdd_), .G(vdd_cntl_r[5]),
     .S(vdd_));
pch_hvt  M0_4_ ( .D(net32[265]), .B(vdd_), .G(vdd_cntl_r[4]),
     .S(vdd_));
pch_hvt  M0_3_ ( .D(net32[266]), .B(vdd_), .G(vdd_cntl_r[3]),
     .S(vdd_));
pch_hvt  M0_2_ ( .D(net32[267]), .B(vdd_), .G(vdd_cntl_r[2]),
     .S(vdd_));
pch_hvt  M0_1_ ( .D(net32[268]), .B(vdd_), .G(vdd_cntl_r[1]),
     .S(vdd_));
pch_hvt  M0_0_ ( .D(net32[269]), .B(vdd_), .G(vdd_cntl_r[0]),
     .S(vdd_));
pch_hvt  vdd_cntrl_269_ ( .D(net43[0]), .B(vdd_), .G(vdd_cntl_l[269]),
     .S(vdd_));
pch_hvt  vdd_cntrl_268_ ( .D(net43[1]), .B(vdd_), .G(vdd_cntl_l[268]),
     .S(vdd_));
pch_hvt  vdd_cntrl_267_ ( .D(net43[2]), .B(vdd_), .G(vdd_cntl_l[267]),
     .S(vdd_));
pch_hvt  vdd_cntrl_266_ ( .D(net43[3]), .B(vdd_), .G(vdd_cntl_l[266]),
     .S(vdd_));
pch_hvt  vdd_cntrl_265_ ( .D(net43[4]), .B(vdd_), .G(vdd_cntl_l[265]),
     .S(vdd_));
pch_hvt  vdd_cntrl_264_ ( .D(net43[5]), .B(vdd_), .G(vdd_cntl_l[264]),
     .S(vdd_));
pch_hvt  vdd_cntrl_263_ ( .D(net43[6]), .B(vdd_), .G(vdd_cntl_l[263]),
     .S(vdd_));
pch_hvt  vdd_cntrl_262_ ( .D(net43[7]), .B(vdd_), .G(vdd_cntl_l[262]),
     .S(vdd_));
pch_hvt  vdd_cntrl_261_ ( .D(net43[8]), .B(vdd_), .G(vdd_cntl_l[261]),
     .S(vdd_));
pch_hvt  vdd_cntrl_260_ ( .D(net43[9]), .B(vdd_), .G(vdd_cntl_l[260]),
     .S(vdd_));
pch_hvt  vdd_cntrl_259_ ( .D(net43[10]), .B(vdd_), .G(vdd_cntl_l[259]),
     .S(vdd_));
pch_hvt  vdd_cntrl_258_ ( .D(net43[11]), .B(vdd_), .G(vdd_cntl_l[258]),
     .S(vdd_));
pch_hvt  vdd_cntrl_257_ ( .D(net43[12]), .B(vdd_), .G(vdd_cntl_l[257]),
     .S(vdd_));
pch_hvt  vdd_cntrl_256_ ( .D(net43[13]), .B(vdd_), .G(vdd_cntl_l[256]),
     .S(vdd_));
pch_hvt  vdd_cntrl_255_ ( .D(net43[14]), .B(vdd_), .G(vdd_cntl_l[255]),
     .S(vdd_));
pch_hvt  vdd_cntrl_254_ ( .D(net43[15]), .B(vdd_), .G(vdd_cntl_l[254]),
     .S(vdd_));
pch_hvt  vdd_cntrl_253_ ( .D(net43[16]), .B(vdd_), .G(vdd_cntl_l[253]),
     .S(vdd_));
pch_hvt  vdd_cntrl_252_ ( .D(net43[17]), .B(vdd_), .G(vdd_cntl_l[252]),
     .S(vdd_));
pch_hvt  vdd_cntrl_251_ ( .D(net43[18]), .B(vdd_), .G(vdd_cntl_l[251]),
     .S(vdd_));
pch_hvt  vdd_cntrl_250_ ( .D(net43[19]), .B(vdd_), .G(vdd_cntl_l[250]),
     .S(vdd_));
pch_hvt  vdd_cntrl_249_ ( .D(net43[20]), .B(vdd_), .G(vdd_cntl_l[249]),
     .S(vdd_));
pch_hvt  vdd_cntrl_248_ ( .D(net43[21]), .B(vdd_), .G(vdd_cntl_l[248]),
     .S(vdd_));
pch_hvt  vdd_cntrl_247_ ( .D(net43[22]), .B(vdd_), .G(vdd_cntl_l[247]),
     .S(vdd_));
pch_hvt  vdd_cntrl_246_ ( .D(net43[23]), .B(vdd_), .G(vdd_cntl_l[246]),
     .S(vdd_));
pch_hvt  vdd_cntrl_245_ ( .D(net43[24]), .B(vdd_), .G(vdd_cntl_l[245]),
     .S(vdd_));
pch_hvt  vdd_cntrl_244_ ( .D(net43[25]), .B(vdd_), .G(vdd_cntl_l[244]),
     .S(vdd_));
pch_hvt  vdd_cntrl_243_ ( .D(net43[26]), .B(vdd_), .G(vdd_cntl_l[243]),
     .S(vdd_));
pch_hvt  vdd_cntrl_242_ ( .D(net43[27]), .B(vdd_), .G(vdd_cntl_l[242]),
     .S(vdd_));
pch_hvt  vdd_cntrl_241_ ( .D(net43[28]), .B(vdd_), .G(vdd_cntl_l[241]),
     .S(vdd_));
pch_hvt  vdd_cntrl_240_ ( .D(net43[29]), .B(vdd_), .G(vdd_cntl_l[240]),
     .S(vdd_));
pch_hvt  vdd_cntrl_239_ ( .D(net43[30]), .B(vdd_), .G(vdd_cntl_l[239]),
     .S(vdd_));
pch_hvt  vdd_cntrl_238_ ( .D(net43[31]), .B(vdd_), .G(vdd_cntl_l[238]),
     .S(vdd_));
pch_hvt  vdd_cntrl_237_ ( .D(net43[32]), .B(vdd_), .G(vdd_cntl_l[237]),
     .S(vdd_));
pch_hvt  vdd_cntrl_236_ ( .D(net43[33]), .B(vdd_), .G(vdd_cntl_l[236]),
     .S(vdd_));
pch_hvt  vdd_cntrl_235_ ( .D(net43[34]), .B(vdd_), .G(vdd_cntl_l[235]),
     .S(vdd_));
pch_hvt  vdd_cntrl_234_ ( .D(net43[35]), .B(vdd_), .G(vdd_cntl_l[234]),
     .S(vdd_));
pch_hvt  vdd_cntrl_233_ ( .D(net43[36]), .B(vdd_), .G(vdd_cntl_l[233]),
     .S(vdd_));
pch_hvt  vdd_cntrl_232_ ( .D(net43[37]), .B(vdd_), .G(vdd_cntl_l[232]),
     .S(vdd_));
pch_hvt  vdd_cntrl_231_ ( .D(net43[38]), .B(vdd_), .G(vdd_cntl_l[231]),
     .S(vdd_));
pch_hvt  vdd_cntrl_230_ ( .D(net43[39]), .B(vdd_), .G(vdd_cntl_l[230]),
     .S(vdd_));
pch_hvt  vdd_cntrl_229_ ( .D(net43[40]), .B(vdd_), .G(vdd_cntl_l[229]),
     .S(vdd_));
pch_hvt  vdd_cntrl_228_ ( .D(net43[41]), .B(vdd_), .G(vdd_cntl_l[228]),
     .S(vdd_));
pch_hvt  vdd_cntrl_227_ ( .D(net43[42]), .B(vdd_), .G(vdd_cntl_l[227]),
     .S(vdd_));
pch_hvt  vdd_cntrl_226_ ( .D(net43[43]), .B(vdd_), .G(vdd_cntl_l[226]),
     .S(vdd_));
pch_hvt  vdd_cntrl_225_ ( .D(net43[44]), .B(vdd_), .G(vdd_cntl_l[225]),
     .S(vdd_));
pch_hvt  vdd_cntrl_224_ ( .D(net43[45]), .B(vdd_), .G(vdd_cntl_l[224]),
     .S(vdd_));
pch_hvt  vdd_cntrl_223_ ( .D(net43[46]), .B(vdd_), .G(vdd_cntl_l[223]),
     .S(vdd_));
pch_hvt  vdd_cntrl_222_ ( .D(net43[47]), .B(vdd_), .G(vdd_cntl_l[222]),
     .S(vdd_));
pch_hvt  vdd_cntrl_221_ ( .D(net43[48]), .B(vdd_), .G(vdd_cntl_l[221]),
     .S(vdd_));
pch_hvt  vdd_cntrl_220_ ( .D(net43[49]), .B(vdd_), .G(vdd_cntl_l[220]),
     .S(vdd_));
pch_hvt  vdd_cntrl_219_ ( .D(net43[50]), .B(vdd_), .G(vdd_cntl_l[219]),
     .S(vdd_));
pch_hvt  vdd_cntrl_218_ ( .D(net43[51]), .B(vdd_), .G(vdd_cntl_l[218]),
     .S(vdd_));
pch_hvt  vdd_cntrl_217_ ( .D(net43[52]), .B(vdd_), .G(vdd_cntl_l[217]),
     .S(vdd_));
pch_hvt  vdd_cntrl_216_ ( .D(net43[53]), .B(vdd_), .G(vdd_cntl_l[216]),
     .S(vdd_));
pch_hvt  vdd_cntrl_215_ ( .D(net43[54]), .B(vdd_), .G(vdd_cntl_l[215]),
     .S(vdd_));
pch_hvt  vdd_cntrl_214_ ( .D(net43[55]), .B(vdd_), .G(vdd_cntl_l[214]),
     .S(vdd_));
pch_hvt  vdd_cntrl_213_ ( .D(net43[56]), .B(vdd_), .G(vdd_cntl_l[213]),
     .S(vdd_));
pch_hvt  vdd_cntrl_212_ ( .D(net43[57]), .B(vdd_), .G(vdd_cntl_l[212]),
     .S(vdd_));
pch_hvt  vdd_cntrl_211_ ( .D(net43[58]), .B(vdd_), .G(vdd_cntl_l[211]),
     .S(vdd_));
pch_hvt  vdd_cntrl_210_ ( .D(net43[59]), .B(vdd_), .G(vdd_cntl_l[210]),
     .S(vdd_));
pch_hvt  vdd_cntrl_209_ ( .D(net43[60]), .B(vdd_), .G(vdd_cntl_l[209]),
     .S(vdd_));
pch_hvt  vdd_cntrl_208_ ( .D(net43[61]), .B(vdd_), .G(vdd_cntl_l[208]),
     .S(vdd_));
pch_hvt  vdd_cntrl_207_ ( .D(net43[62]), .B(vdd_), .G(vdd_cntl_l[207]),
     .S(vdd_));
pch_hvt  vdd_cntrl_206_ ( .D(net43[63]), .B(vdd_), .G(vdd_cntl_l[206]),
     .S(vdd_));
pch_hvt  vdd_cntrl_205_ ( .D(net43[64]), .B(vdd_), .G(vdd_cntl_l[205]),
     .S(vdd_));
pch_hvt  vdd_cntrl_204_ ( .D(net43[65]), .B(vdd_), .G(vdd_cntl_l[204]),
     .S(vdd_));
pch_hvt  vdd_cntrl_203_ ( .D(net43[66]), .B(vdd_), .G(vdd_cntl_l[203]),
     .S(vdd_));
pch_hvt  vdd_cntrl_202_ ( .D(net43[67]), .B(vdd_), .G(vdd_cntl_l[202]),
     .S(vdd_));
pch_hvt  vdd_cntrl_201_ ( .D(net43[68]), .B(vdd_), .G(vdd_cntl_l[201]),
     .S(vdd_));
pch_hvt  vdd_cntrl_200_ ( .D(net43[69]), .B(vdd_), .G(vdd_cntl_l[200]),
     .S(vdd_));
pch_hvt  vdd_cntrl_199_ ( .D(net43[70]), .B(vdd_), .G(vdd_cntl_l[199]),
     .S(vdd_));
pch_hvt  vdd_cntrl_198_ ( .D(net43[71]), .B(vdd_), .G(vdd_cntl_l[198]),
     .S(vdd_));
pch_hvt  vdd_cntrl_197_ ( .D(net43[72]), .B(vdd_), .G(vdd_cntl_l[197]),
     .S(vdd_));
pch_hvt  vdd_cntrl_196_ ( .D(net43[73]), .B(vdd_), .G(vdd_cntl_l[196]),
     .S(vdd_));
pch_hvt  vdd_cntrl_195_ ( .D(net43[74]), .B(vdd_), .G(vdd_cntl_l[195]),
     .S(vdd_));
pch_hvt  vdd_cntrl_194_ ( .D(net43[75]), .B(vdd_), .G(vdd_cntl_l[194]),
     .S(vdd_));
pch_hvt  vdd_cntrl_193_ ( .D(net43[76]), .B(vdd_), .G(vdd_cntl_l[193]),
     .S(vdd_));
pch_hvt  vdd_cntrl_192_ ( .D(net43[77]), .B(vdd_), .G(vdd_cntl_l[192]),
     .S(vdd_));
pch_hvt  vdd_cntrl_191_ ( .D(net43[78]), .B(vdd_), .G(vdd_cntl_l[191]),
     .S(vdd_));
pch_hvt  vdd_cntrl_190_ ( .D(net43[79]), .B(vdd_), .G(vdd_cntl_l[190]),
     .S(vdd_));
pch_hvt  vdd_cntrl_189_ ( .D(net43[80]), .B(vdd_), .G(vdd_cntl_l[189]),
     .S(vdd_));
pch_hvt  vdd_cntrl_188_ ( .D(net43[81]), .B(vdd_), .G(vdd_cntl_l[188]),
     .S(vdd_));
pch_hvt  vdd_cntrl_187_ ( .D(net43[82]), .B(vdd_), .G(vdd_cntl_l[187]),
     .S(vdd_));
pch_hvt  vdd_cntrl_186_ ( .D(net43[83]), .B(vdd_), .G(vdd_cntl_l[186]),
     .S(vdd_));
pch_hvt  vdd_cntrl_185_ ( .D(net43[84]), .B(vdd_), .G(vdd_cntl_l[185]),
     .S(vdd_));
pch_hvt  vdd_cntrl_184_ ( .D(net43[85]), .B(vdd_), .G(vdd_cntl_l[184]),
     .S(vdd_));
pch_hvt  vdd_cntrl_183_ ( .D(net43[86]), .B(vdd_), .G(vdd_cntl_l[183]),
     .S(vdd_));
pch_hvt  vdd_cntrl_182_ ( .D(net43[87]), .B(vdd_), .G(vdd_cntl_l[182]),
     .S(vdd_));
pch_hvt  vdd_cntrl_181_ ( .D(net43[88]), .B(vdd_), .G(vdd_cntl_l[181]),
     .S(vdd_));
pch_hvt  vdd_cntrl_180_ ( .D(net43[89]), .B(vdd_), .G(vdd_cntl_l[180]),
     .S(vdd_));
pch_hvt  vdd_cntrl_179_ ( .D(net43[90]), .B(vdd_), .G(vdd_cntl_l[179]),
     .S(vdd_));
pch_hvt  vdd_cntrl_178_ ( .D(net43[91]), .B(vdd_), .G(vdd_cntl_l[178]),
     .S(vdd_));
pch_hvt  vdd_cntrl_177_ ( .D(net43[92]), .B(vdd_), .G(vdd_cntl_l[177]),
     .S(vdd_));
pch_hvt  vdd_cntrl_176_ ( .D(net43[93]), .B(vdd_), .G(vdd_cntl_l[176]),
     .S(vdd_));
pch_hvt  vdd_cntrl_175_ ( .D(net43[94]), .B(vdd_), .G(vdd_cntl_l[175]),
     .S(vdd_));
pch_hvt  vdd_cntrl_174_ ( .D(net43[95]), .B(vdd_), .G(vdd_cntl_l[174]),
     .S(vdd_));
pch_hvt  vdd_cntrl_173_ ( .D(net43[96]), .B(vdd_), .G(vdd_cntl_l[173]),
     .S(vdd_));
pch_hvt  vdd_cntrl_172_ ( .D(net43[97]), .B(vdd_), .G(vdd_cntl_l[172]),
     .S(vdd_));
pch_hvt  vdd_cntrl_171_ ( .D(net43[98]), .B(vdd_), .G(vdd_cntl_l[171]),
     .S(vdd_));
pch_hvt  vdd_cntrl_170_ ( .D(net43[99]), .B(vdd_), .G(vdd_cntl_l[170]),
     .S(vdd_));
pch_hvt  vdd_cntrl_169_ ( .D(net43[100]), .B(vdd_),
     .G(vdd_cntl_l[169]), .S(vdd_));
pch_hvt  vdd_cntrl_168_ ( .D(net43[101]), .B(vdd_),
     .G(vdd_cntl_l[168]), .S(vdd_));
pch_hvt  vdd_cntrl_167_ ( .D(net43[102]), .B(vdd_),
     .G(vdd_cntl_l[167]), .S(vdd_));
pch_hvt  vdd_cntrl_166_ ( .D(net43[103]), .B(vdd_),
     .G(vdd_cntl_l[166]), .S(vdd_));
pch_hvt  vdd_cntrl_165_ ( .D(net43[104]), .B(vdd_),
     .G(vdd_cntl_l[165]), .S(vdd_));
pch_hvt  vdd_cntrl_164_ ( .D(net43[105]), .B(vdd_),
     .G(vdd_cntl_l[164]), .S(vdd_));
pch_hvt  vdd_cntrl_163_ ( .D(net43[106]), .B(vdd_),
     .G(vdd_cntl_l[163]), .S(vdd_));
pch_hvt  vdd_cntrl_162_ ( .D(net43[107]), .B(vdd_),
     .G(vdd_cntl_l[162]), .S(vdd_));
pch_hvt  vdd_cntrl_161_ ( .D(net43[108]), .B(vdd_),
     .G(vdd_cntl_l[161]), .S(vdd_));
pch_hvt  vdd_cntrl_160_ ( .D(net43[109]), .B(vdd_),
     .G(vdd_cntl_l[160]), .S(vdd_));
pch_hvt  vdd_cntrl_159_ ( .D(net43[110]), .B(vdd_),
     .G(vdd_cntl_l[159]), .S(vdd_));
pch_hvt  vdd_cntrl_158_ ( .D(net43[111]), .B(vdd_),
     .G(vdd_cntl_l[158]), .S(vdd_));
pch_hvt  vdd_cntrl_157_ ( .D(net43[112]), .B(vdd_),
     .G(vdd_cntl_l[157]), .S(vdd_));
pch_hvt  vdd_cntrl_156_ ( .D(net43[113]), .B(vdd_),
     .G(vdd_cntl_l[156]), .S(vdd_));
pch_hvt  vdd_cntrl_155_ ( .D(net43[114]), .B(vdd_),
     .G(vdd_cntl_l[155]), .S(vdd_));
pch_hvt  vdd_cntrl_154_ ( .D(net43[115]), .B(vdd_),
     .G(vdd_cntl_l[154]), .S(vdd_));
pch_hvt  vdd_cntrl_153_ ( .D(net43[116]), .B(vdd_),
     .G(vdd_cntl_l[153]), .S(vdd_));
pch_hvt  vdd_cntrl_152_ ( .D(net43[117]), .B(vdd_),
     .G(vdd_cntl_l[152]), .S(vdd_));
pch_hvt  vdd_cntrl_151_ ( .D(net43[118]), .B(vdd_),
     .G(vdd_cntl_l[151]), .S(vdd_));
pch_hvt  vdd_cntrl_150_ ( .D(net43[119]), .B(vdd_),
     .G(vdd_cntl_l[150]), .S(vdd_));
pch_hvt  vdd_cntrl_149_ ( .D(net43[120]), .B(vdd_),
     .G(vdd_cntl_l[149]), .S(vdd_));
pch_hvt  vdd_cntrl_148_ ( .D(net43[121]), .B(vdd_),
     .G(vdd_cntl_l[148]), .S(vdd_));
pch_hvt  vdd_cntrl_147_ ( .D(net43[122]), .B(vdd_),
     .G(vdd_cntl_l[147]), .S(vdd_));
pch_hvt  vdd_cntrl_146_ ( .D(net43[123]), .B(vdd_),
     .G(vdd_cntl_l[146]), .S(vdd_));
pch_hvt  vdd_cntrl_145_ ( .D(net43[124]), .B(vdd_),
     .G(vdd_cntl_l[145]), .S(vdd_));
pch_hvt  vdd_cntrl_144_ ( .D(net43[125]), .B(vdd_),
     .G(vdd_cntl_l[144]), .S(vdd_));
pch_hvt  vdd_cntrl_143_ ( .D(net43[126]), .B(vdd_),
     .G(vdd_cntl_l[143]), .S(vdd_));
pch_hvt  vdd_cntrl_142_ ( .D(net43[127]), .B(vdd_),
     .G(vdd_cntl_l[142]), .S(vdd_));
pch_hvt  vdd_cntrl_141_ ( .D(net43[128]), .B(vdd_),
     .G(vdd_cntl_l[141]), .S(vdd_));
pch_hvt  vdd_cntrl_140_ ( .D(net43[129]), .B(vdd_),
     .G(vdd_cntl_l[140]), .S(vdd_));
pch_hvt  vdd_cntrl_139_ ( .D(net43[130]), .B(vdd_),
     .G(vdd_cntl_l[139]), .S(vdd_));
pch_hvt  vdd_cntrl_138_ ( .D(net43[131]), .B(vdd_),
     .G(vdd_cntl_l[138]), .S(vdd_));
pch_hvt  vdd_cntrl_137_ ( .D(net43[132]), .B(vdd_),
     .G(vdd_cntl_l[137]), .S(vdd_));
pch_hvt  vdd_cntrl_136_ ( .D(net43[133]), .B(vdd_),
     .G(vdd_cntl_l[136]), .S(vdd_));
pch_hvt  vdd_cntrl_135_ ( .D(net43[134]), .B(vdd_),
     .G(vdd_cntl_l[135]), .S(vdd_));
pch_hvt  vdd_cntrl_134_ ( .D(net43[135]), .B(vdd_),
     .G(vdd_cntl_l[134]), .S(vdd_));
pch_hvt  vdd_cntrl_133_ ( .D(net43[136]), .B(vdd_),
     .G(vdd_cntl_l[133]), .S(vdd_));
pch_hvt  vdd_cntrl_132_ ( .D(net43[137]), .B(vdd_),
     .G(vdd_cntl_l[132]), .S(vdd_));
pch_hvt  vdd_cntrl_131_ ( .D(net43[138]), .B(vdd_),
     .G(vdd_cntl_l[131]), .S(vdd_));
pch_hvt  vdd_cntrl_130_ ( .D(net43[139]), .B(vdd_),
     .G(vdd_cntl_l[130]), .S(vdd_));
pch_hvt  vdd_cntrl_129_ ( .D(net43[140]), .B(vdd_),
     .G(vdd_cntl_l[129]), .S(vdd_));
pch_hvt  vdd_cntrl_128_ ( .D(net43[141]), .B(vdd_),
     .G(vdd_cntl_l[128]), .S(vdd_));
pch_hvt  vdd_cntrl_127_ ( .D(net43[142]), .B(vdd_),
     .G(vdd_cntl_l[127]), .S(vdd_));
pch_hvt  vdd_cntrl_126_ ( .D(net43[143]), .B(vdd_),
     .G(vdd_cntl_l[126]), .S(vdd_));
pch_hvt  vdd_cntrl_125_ ( .D(net43[144]), .B(vdd_),
     .G(vdd_cntl_l[125]), .S(vdd_));
pch_hvt  vdd_cntrl_124_ ( .D(net43[145]), .B(vdd_),
     .G(vdd_cntl_l[124]), .S(vdd_));
pch_hvt  vdd_cntrl_123_ ( .D(net43[146]), .B(vdd_),
     .G(vdd_cntl_l[123]), .S(vdd_));
pch_hvt  vdd_cntrl_122_ ( .D(net43[147]), .B(vdd_),
     .G(vdd_cntl_l[122]), .S(vdd_));
pch_hvt  vdd_cntrl_121_ ( .D(net43[148]), .B(vdd_),
     .G(vdd_cntl_l[121]), .S(vdd_));
pch_hvt  vdd_cntrl_120_ ( .D(net43[149]), .B(vdd_),
     .G(vdd_cntl_l[120]), .S(vdd_));
pch_hvt  vdd_cntrl_119_ ( .D(net43[150]), .B(vdd_),
     .G(vdd_cntl_l[119]), .S(vdd_));
pch_hvt  vdd_cntrl_118_ ( .D(net43[151]), .B(vdd_),
     .G(vdd_cntl_l[118]), .S(vdd_));
pch_hvt  vdd_cntrl_117_ ( .D(net43[152]), .B(vdd_),
     .G(vdd_cntl_l[117]), .S(vdd_));
pch_hvt  vdd_cntrl_116_ ( .D(net43[153]), .B(vdd_),
     .G(vdd_cntl_l[116]), .S(vdd_));
pch_hvt  vdd_cntrl_115_ ( .D(net43[154]), .B(vdd_),
     .G(vdd_cntl_l[115]), .S(vdd_));
pch_hvt  vdd_cntrl_114_ ( .D(net43[155]), .B(vdd_),
     .G(vdd_cntl_l[114]), .S(vdd_));
pch_hvt  vdd_cntrl_113_ ( .D(net43[156]), .B(vdd_),
     .G(vdd_cntl_l[113]), .S(vdd_));
pch_hvt  vdd_cntrl_112_ ( .D(net43[157]), .B(vdd_),
     .G(vdd_cntl_l[112]), .S(vdd_));
pch_hvt  vdd_cntrl_111_ ( .D(net43[158]), .B(vdd_),
     .G(vdd_cntl_l[111]), .S(vdd_));
pch_hvt  vdd_cntrl_110_ ( .D(net43[159]), .B(vdd_),
     .G(vdd_cntl_l[110]), .S(vdd_));
pch_hvt  vdd_cntrl_109_ ( .D(net43[160]), .B(vdd_),
     .G(vdd_cntl_l[109]), .S(vdd_));
pch_hvt  vdd_cntrl_108_ ( .D(net43[161]), .B(vdd_),
     .G(vdd_cntl_l[108]), .S(vdd_));
pch_hvt  vdd_cntrl_107_ ( .D(net43[162]), .B(vdd_),
     .G(vdd_cntl_l[107]), .S(vdd_));
pch_hvt  vdd_cntrl_106_ ( .D(net43[163]), .B(vdd_),
     .G(vdd_cntl_l[106]), .S(vdd_));
pch_hvt  vdd_cntrl_105_ ( .D(net43[164]), .B(vdd_),
     .G(vdd_cntl_l[105]), .S(vdd_));
pch_hvt  vdd_cntrl_104_ ( .D(net43[165]), .B(vdd_),
     .G(vdd_cntl_l[104]), .S(vdd_));
pch_hvt  vdd_cntrl_103_ ( .D(net43[166]), .B(vdd_),
     .G(vdd_cntl_l[103]), .S(vdd_));
pch_hvt  vdd_cntrl_102_ ( .D(net43[167]), .B(vdd_),
     .G(vdd_cntl_l[102]), .S(vdd_));
pch_hvt  vdd_cntrl_101_ ( .D(net43[168]), .B(vdd_),
     .G(vdd_cntl_l[101]), .S(vdd_));
pch_hvt  vdd_cntrl_100_ ( .D(net43[169]), .B(vdd_),
     .G(vdd_cntl_l[100]), .S(vdd_));
pch_hvt  vdd_cntrl_99_ ( .D(net43[170]), .B(vdd_), .G(vdd_cntl_l[99]),
     .S(vdd_));
pch_hvt  vdd_cntrl_98_ ( .D(net43[171]), .B(vdd_), .G(vdd_cntl_l[98]),
     .S(vdd_));
pch_hvt  vdd_cntrl_97_ ( .D(net43[172]), .B(vdd_), .G(vdd_cntl_l[97]),
     .S(vdd_));
pch_hvt  vdd_cntrl_96_ ( .D(net43[173]), .B(vdd_), .G(vdd_cntl_l[96]),
     .S(vdd_));
pch_hvt  vdd_cntrl_95_ ( .D(net43[174]), .B(vdd_), .G(vdd_cntl_l[95]),
     .S(vdd_));
pch_hvt  vdd_cntrl_94_ ( .D(net43[175]), .B(vdd_), .G(vdd_cntl_l[94]),
     .S(vdd_));
pch_hvt  vdd_cntrl_93_ ( .D(net43[176]), .B(vdd_), .G(vdd_cntl_l[93]),
     .S(vdd_));
pch_hvt  vdd_cntrl_92_ ( .D(net43[177]), .B(vdd_), .G(vdd_cntl_l[92]),
     .S(vdd_));
pch_hvt  vdd_cntrl_91_ ( .D(net43[178]), .B(vdd_), .G(vdd_cntl_l[91]),
     .S(vdd_));
pch_hvt  vdd_cntrl_90_ ( .D(net43[179]), .B(vdd_), .G(vdd_cntl_l[90]),
     .S(vdd_));
pch_hvt  vdd_cntrl_89_ ( .D(net43[180]), .B(vdd_), .G(vdd_cntl_l[89]),
     .S(vdd_));
pch_hvt  vdd_cntrl_88_ ( .D(net43[181]), .B(vdd_), .G(vdd_cntl_l[88]),
     .S(vdd_));
pch_hvt  vdd_cntrl_87_ ( .D(net43[182]), .B(vdd_), .G(vdd_cntl_l[87]),
     .S(vdd_));
pch_hvt  vdd_cntrl_86_ ( .D(net43[183]), .B(vdd_), .G(vdd_cntl_l[86]),
     .S(vdd_));
pch_hvt  vdd_cntrl_85_ ( .D(net43[184]), .B(vdd_), .G(vdd_cntl_l[85]),
     .S(vdd_));
pch_hvt  vdd_cntrl_84_ ( .D(net43[185]), .B(vdd_), .G(vdd_cntl_l[84]),
     .S(vdd_));
pch_hvt  vdd_cntrl_83_ ( .D(net43[186]), .B(vdd_), .G(vdd_cntl_l[83]),
     .S(vdd_));
pch_hvt  vdd_cntrl_82_ ( .D(net43[187]), .B(vdd_), .G(vdd_cntl_l[82]),
     .S(vdd_));
pch_hvt  vdd_cntrl_81_ ( .D(net43[188]), .B(vdd_), .G(vdd_cntl_l[81]),
     .S(vdd_));
pch_hvt  vdd_cntrl_80_ ( .D(net43[189]), .B(vdd_), .G(vdd_cntl_l[80]),
     .S(vdd_));
pch_hvt  vdd_cntrl_79_ ( .D(net43[190]), .B(vdd_), .G(vdd_cntl_l[79]),
     .S(vdd_));
pch_hvt  vdd_cntrl_78_ ( .D(net43[191]), .B(vdd_), .G(vdd_cntl_l[78]),
     .S(vdd_));
pch_hvt  vdd_cntrl_77_ ( .D(net43[192]), .B(vdd_), .G(vdd_cntl_l[77]),
     .S(vdd_));
pch_hvt  vdd_cntrl_76_ ( .D(net43[193]), .B(vdd_), .G(vdd_cntl_l[76]),
     .S(vdd_));
pch_hvt  vdd_cntrl_75_ ( .D(net43[194]), .B(vdd_), .G(vdd_cntl_l[75]),
     .S(vdd_));
pch_hvt  vdd_cntrl_74_ ( .D(net43[195]), .B(vdd_), .G(vdd_cntl_l[74]),
     .S(vdd_));
pch_hvt  vdd_cntrl_73_ ( .D(net43[196]), .B(vdd_), .G(vdd_cntl_l[73]),
     .S(vdd_));
pch_hvt  vdd_cntrl_72_ ( .D(net43[197]), .B(vdd_), .G(vdd_cntl_l[72]),
     .S(vdd_));
pch_hvt  vdd_cntrl_71_ ( .D(net43[198]), .B(vdd_), .G(vdd_cntl_l[71]),
     .S(vdd_));
pch_hvt  vdd_cntrl_70_ ( .D(net43[199]), .B(vdd_), .G(vdd_cntl_l[70]),
     .S(vdd_));
pch_hvt  vdd_cntrl_69_ ( .D(net43[200]), .B(vdd_), .G(vdd_cntl_l[69]),
     .S(vdd_));
pch_hvt  vdd_cntrl_68_ ( .D(net43[201]), .B(vdd_), .G(vdd_cntl_l[68]),
     .S(vdd_));
pch_hvt  vdd_cntrl_67_ ( .D(net43[202]), .B(vdd_), .G(vdd_cntl_l[67]),
     .S(vdd_));
pch_hvt  vdd_cntrl_66_ ( .D(net43[203]), .B(vdd_), .G(vdd_cntl_l[66]),
     .S(vdd_));
pch_hvt  vdd_cntrl_65_ ( .D(net43[204]), .B(vdd_), .G(vdd_cntl_l[65]),
     .S(vdd_));
pch_hvt  vdd_cntrl_64_ ( .D(net43[205]), .B(vdd_), .G(vdd_cntl_l[64]),
     .S(vdd_));
pch_hvt  vdd_cntrl_63_ ( .D(net43[206]), .B(vdd_), .G(vdd_cntl_l[63]),
     .S(vdd_));
pch_hvt  vdd_cntrl_62_ ( .D(net43[207]), .B(vdd_), .G(vdd_cntl_l[62]),
     .S(vdd_));
pch_hvt  vdd_cntrl_61_ ( .D(net43[208]), .B(vdd_), .G(vdd_cntl_l[61]),
     .S(vdd_));
pch_hvt  vdd_cntrl_60_ ( .D(net43[209]), .B(vdd_), .G(vdd_cntl_l[60]),
     .S(vdd_));
pch_hvt  vdd_cntrl_59_ ( .D(net43[210]), .B(vdd_), .G(vdd_cntl_l[59]),
     .S(vdd_));
pch_hvt  vdd_cntrl_58_ ( .D(net43[211]), .B(vdd_), .G(vdd_cntl_l[58]),
     .S(vdd_));
pch_hvt  vdd_cntrl_57_ ( .D(net43[212]), .B(vdd_), .G(vdd_cntl_l[57]),
     .S(vdd_));
pch_hvt  vdd_cntrl_56_ ( .D(net43[213]), .B(vdd_), .G(vdd_cntl_l[56]),
     .S(vdd_));
pch_hvt  vdd_cntrl_55_ ( .D(net43[214]), .B(vdd_), .G(vdd_cntl_l[55]),
     .S(vdd_));
pch_hvt  vdd_cntrl_54_ ( .D(net43[215]), .B(vdd_), .G(vdd_cntl_l[54]),
     .S(vdd_));
pch_hvt  vdd_cntrl_53_ ( .D(net43[216]), .B(vdd_), .G(vdd_cntl_l[53]),
     .S(vdd_));
pch_hvt  vdd_cntrl_52_ ( .D(net43[217]), .B(vdd_), .G(vdd_cntl_l[52]),
     .S(vdd_));
pch_hvt  vdd_cntrl_51_ ( .D(net43[218]), .B(vdd_), .G(vdd_cntl_l[51]),
     .S(vdd_));
pch_hvt  vdd_cntrl_50_ ( .D(net43[219]), .B(vdd_), .G(vdd_cntl_l[50]),
     .S(vdd_));
pch_hvt  vdd_cntrl_49_ ( .D(net43[220]), .B(vdd_), .G(vdd_cntl_l[49]),
     .S(vdd_));
pch_hvt  vdd_cntrl_48_ ( .D(net43[221]), .B(vdd_), .G(vdd_cntl_l[48]),
     .S(vdd_));
pch_hvt  vdd_cntrl_47_ ( .D(net43[222]), .B(vdd_), .G(vdd_cntl_l[47]),
     .S(vdd_));
pch_hvt  vdd_cntrl_46_ ( .D(net43[223]), .B(vdd_), .G(vdd_cntl_l[46]),
     .S(vdd_));
pch_hvt  vdd_cntrl_45_ ( .D(net43[224]), .B(vdd_), .G(vdd_cntl_l[45]),
     .S(vdd_));
pch_hvt  vdd_cntrl_44_ ( .D(net43[225]), .B(vdd_), .G(vdd_cntl_l[44]),
     .S(vdd_));
pch_hvt  vdd_cntrl_43_ ( .D(net43[226]), .B(vdd_), .G(vdd_cntl_l[43]),
     .S(vdd_));
pch_hvt  vdd_cntrl_42_ ( .D(net43[227]), .B(vdd_), .G(vdd_cntl_l[42]),
     .S(vdd_));
pch_hvt  vdd_cntrl_41_ ( .D(net43[228]), .B(vdd_), .G(vdd_cntl_l[41]),
     .S(vdd_));
pch_hvt  vdd_cntrl_40_ ( .D(net43[229]), .B(vdd_), .G(vdd_cntl_l[40]),
     .S(vdd_));
pch_hvt  vdd_cntrl_39_ ( .D(net43[230]), .B(vdd_), .G(vdd_cntl_l[39]),
     .S(vdd_));
pch_hvt  vdd_cntrl_38_ ( .D(net43[231]), .B(vdd_), .G(vdd_cntl_l[38]),
     .S(vdd_));
pch_hvt  vdd_cntrl_37_ ( .D(net43[232]), .B(vdd_), .G(vdd_cntl_l[37]),
     .S(vdd_));
pch_hvt  vdd_cntrl_36_ ( .D(net43[233]), .B(vdd_), .G(vdd_cntl_l[36]),
     .S(vdd_));
pch_hvt  vdd_cntrl_35_ ( .D(net43[234]), .B(vdd_), .G(vdd_cntl_l[35]),
     .S(vdd_));
pch_hvt  vdd_cntrl_34_ ( .D(net43[235]), .B(vdd_), .G(vdd_cntl_l[34]),
     .S(vdd_));
pch_hvt  vdd_cntrl_33_ ( .D(net43[236]), .B(vdd_), .G(vdd_cntl_l[33]),
     .S(vdd_));
pch_hvt  vdd_cntrl_32_ ( .D(net43[237]), .B(vdd_), .G(vdd_cntl_l[32]),
     .S(vdd_));
pch_hvt  vdd_cntrl_31_ ( .D(net43[238]), .B(vdd_), .G(vdd_cntl_l[31]),
     .S(vdd_));
pch_hvt  vdd_cntrl_30_ ( .D(net43[239]), .B(vdd_), .G(vdd_cntl_l[30]),
     .S(vdd_));
pch_hvt  vdd_cntrl_29_ ( .D(net43[240]), .B(vdd_), .G(vdd_cntl_l[29]),
     .S(vdd_));
pch_hvt  vdd_cntrl_28_ ( .D(net43[241]), .B(vdd_), .G(vdd_cntl_l[28]),
     .S(vdd_));
pch_hvt  vdd_cntrl_27_ ( .D(net43[242]), .B(vdd_), .G(vdd_cntl_l[27]),
     .S(vdd_));
pch_hvt  vdd_cntrl_26_ ( .D(net43[243]), .B(vdd_), .G(vdd_cntl_l[26]),
     .S(vdd_));
pch_hvt  vdd_cntrl_25_ ( .D(net43[244]), .B(vdd_), .G(vdd_cntl_l[25]),
     .S(vdd_));
pch_hvt  vdd_cntrl_24_ ( .D(net43[245]), .B(vdd_), .G(vdd_cntl_l[24]),
     .S(vdd_));
pch_hvt  vdd_cntrl_23_ ( .D(net43[246]), .B(vdd_), .G(vdd_cntl_l[23]),
     .S(vdd_));
pch_hvt  vdd_cntrl_22_ ( .D(net43[247]), .B(vdd_), .G(vdd_cntl_l[22]),
     .S(vdd_));
pch_hvt  vdd_cntrl_21_ ( .D(net43[248]), .B(vdd_), .G(vdd_cntl_l[21]),
     .S(vdd_));
pch_hvt  vdd_cntrl_20_ ( .D(net43[249]), .B(vdd_), .G(vdd_cntl_l[20]),
     .S(vdd_));
pch_hvt  vdd_cntrl_19_ ( .D(net43[250]), .B(vdd_), .G(vdd_cntl_l[19]),
     .S(vdd_));
pch_hvt  vdd_cntrl_18_ ( .D(net43[251]), .B(vdd_), .G(vdd_cntl_l[18]),
     .S(vdd_));
pch_hvt  vdd_cntrl_17_ ( .D(net43[252]), .B(vdd_), .G(vdd_cntl_l[17]),
     .S(vdd_));
pch_hvt  vdd_cntrl_16_ ( .D(net43[253]), .B(vdd_), .G(vdd_cntl_l[16]),
     .S(vdd_));
pch_hvt  vdd_cntrl_15_ ( .D(net43[254]), .B(vdd_), .G(vdd_cntl_l[15]),
     .S(vdd_));
pch_hvt  vdd_cntrl_14_ ( .D(net43[255]), .B(vdd_), .G(vdd_cntl_l[14]),
     .S(vdd_));
pch_hvt  vdd_cntrl_13_ ( .D(net43[256]), .B(vdd_), .G(vdd_cntl_l[13]),
     .S(vdd_));
pch_hvt  vdd_cntrl_12_ ( .D(net43[257]), .B(vdd_), .G(vdd_cntl_l[12]),
     .S(vdd_));
pch_hvt  vdd_cntrl_11_ ( .D(net43[258]), .B(vdd_), .G(vdd_cntl_l[11]),
     .S(vdd_));
pch_hvt  vdd_cntrl_10_ ( .D(net43[259]), .B(vdd_), .G(vdd_cntl_l[10]),
     .S(vdd_));
pch_hvt  vdd_cntrl_9_ ( .D(net43[260]), .B(vdd_), .G(vdd_cntl_l[9]),
     .S(vdd_));
pch_hvt  vdd_cntrl_8_ ( .D(net43[261]), .B(vdd_), .G(vdd_cntl_l[8]),
     .S(vdd_));
pch_hvt  vdd_cntrl_7_ ( .D(net43[262]), .B(vdd_), .G(vdd_cntl_l[7]),
     .S(vdd_));
pch_hvt  vdd_cntrl_6_ ( .D(net43[263]), .B(vdd_), .G(vdd_cntl_l[6]),
     .S(vdd_));
pch_hvt  vdd_cntrl_5_ ( .D(net43[264]), .B(vdd_), .G(vdd_cntl_l[5]),
     .S(vdd_));
pch_hvt  vdd_cntrl_4_ ( .D(net43[265]), .B(vdd_), .G(vdd_cntl_l[4]),
     .S(vdd_));
pch_hvt  vdd_cntrl_3_ ( .D(net43[266]), .B(vdd_), .G(vdd_cntl_l[3]),
     .S(vdd_));
pch_hvt  vdd_cntrl_2_ ( .D(net43[267]), .B(vdd_), .G(vdd_cntl_l[2]),
     .S(vdd_));
pch_hvt  vdd_cntrl_1_ ( .D(net43[268]), .B(vdd_), .G(vdd_cntl_l[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(net43[269]), .B(vdd_), .G(vdd_cntl_l[0]),
     .S(vdd_));

endmodule
// Library - leafcell, Cell - lowla_modified, View - schematic
// LAST TIME SAVED: Sep 15 13:19:27 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module lowla_modified ( lao, clk, min );
output  lao;

input  clk, min;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I289 ( .A(net29), .Y(lao));
inv_hvt I290 ( .A(st2), .Y(net29));
inv_hvt I_inv ( .A(clk), .Y(cbitb));
inv_hvt I_inv3 ( .A(cbitb), .Y(clkd));
txgate_hvt I249 ( .in(lao), .out(st2), .pp(cbitb), .nn(clkd));
txgate_hvt I248 ( .in(min), .out(st2), .pp(clkd), .nn(cbitb));

endmodule
// Library - leafcell, Cell - bram_bufferx4x6, View - schematic
// LAST TIME SAVED: Sep 15 13:53:57 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module bram_bufferx4x6 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx4 I4 ( .in(d1), .out(d2));
bram_bufferx4 I5 ( .in(d2), .out(d3));
bram_bufferx4 I6 ( .in(d3), .out(d4));
bram_bufferx4 I7 ( .in(d4), .out(out));
bram_bufferx4 I3 ( .in(d0), .out(d1));
bram_bufferx4 I0 ( .in(in), .out(d0));

endmodule
// Library - leafcell, Cell - tckbufx16, View - schematic
// LAST TIME SAVED: Jan 31 14:34:05 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module tckbufx16 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - clk_colbuf8k, View - schematic
// LAST TIME SAVED: Jan 15 15:48:29 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module clk_colbuf8k ( clko, clki );
output  clko;

input  clki;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I19 ( .A(clkb), .Y(clko));
inv_hvt I22 ( .A(clki), .Y(clkb));

endmodule
// Library - leafcell, Cell - clk_colbuf8kx8, View - schematic
// LAST TIME SAVED: Jan 23 09:43:03 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module clk_colbuf8kx8 ( clko, clki );


output [7:0]  clko;

input [7:0]  clki;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



clk_colbuf8k iclk_colbuf_7_ ( .clki(clki[7]), .clko(clko[7]));
clk_colbuf8k iclk_colbuf_6_ ( .clki(clki[6]), .clko(clko[6]));
clk_colbuf8k iclk_colbuf_5_ ( .clki(clki[5]), .clko(clko[5]));
clk_colbuf8k iclk_colbuf_4_ ( .clki(clki[4]), .clko(clko[4]));
clk_colbuf8k iclk_colbuf_3_ ( .clki(clki[3]), .clko(clko[3]));
clk_colbuf8k iclk_colbuf_2_ ( .clki(clki[2]), .clko(clko[2]));
clk_colbuf8k iclk_colbuf_1_ ( .clki(clki[1]), .clko(clko[1]));
clk_colbuf8k iclk_colbuf_0_ ( .clki(clki[0]), .clko(clko[0]));

endmodule
// Library - leafcell, Cell - fabric_buf8k, View - schematic
// LAST TIME SAVED: Jan 15 15:42:13 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module fabric_buf8k ( f_out, f_in );
output  f_out;

input  f_in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I252 ( .A(net6), .Y(f_out));
inv_hvt I248 ( .A(f_in), .Y(net6));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev0, View - schematic
// LAST TIME SAVED: Jun  2 13:19:45 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module clkmandcmuxrev0 ( clk, clkb, glb2local, s_r, cbit, cbitb,
     glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, min0, min1,
     min2, min3, prog );
output  clk, clkb, s_r;

input  prog;

output [3:0]  glb2local;

input [7:0]  min3;
input [7:0]  min1;
input [7:0]  min0;
input [7:0]  min2;
input [31:0]  cbitb;
input [7:0]  glb_netwk;
input [5:0]  lc_trk_g0;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g3;
input [31:0]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sr_clkm8to1 I296 ( .mout(s_r), .cbitb(cbitb[12:9]), .min({lc_trk_g3[5],
     lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4], glb_netwk[6],
     glb_netwk[4], glb_netwk[2], glb_netwk[0]}), .cbit(cbit[12:9]),
     .prog(prog));
ce_clkm8to1 I283 ( .moutb(ceb), .cbitb(cbitb[8:5]), .cbit(cbit[8:5]),
     .prog(prog), .min({lc_trk_g3[3], lc_trk_g2[2], lc_trk_g1[3],
     lc_trk_g0[2], glb_netwk[7], glb_netwk[5], glb_netwk[3],
     glb_netwk[1]}));
clk_mux12to1 I298 ( .cbitb({cbitb[31], cbitb[4], cbitb[3], cbitb[2],
     cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3], cbit[2],
     cbit[1], cbit[0]}), .prog(prog), .min({lc_trk_g3[1], lc_trk_g2[0],
     lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}), .clk(clk),
     .clkb(clkb), .cenb(ceb));
clk_mux8to1 I285 ( .min(min3[7:0]), .prog(prog), .inmuxo(glb2local[0]),
     .cbit(cbit[16:13]), .cbitb(cbitb[16:13]));
clk_mux8to1 I293 ( .prog(prog), .inmuxo(glb2local[1]), .min(min2[7:0]),
     .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I294 ( .prog(prog), .inmuxo(glb2local[2]), .min(min1[7:0]),
     .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
clk_mux8to1 I295 ( .prog(prog), .inmuxo(glb2local[3]), .min(min0[7:0]),
     .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));

endmodule
// Library - leafcell, Cell - sbox1, View - schematic
// LAST TIME SAVED: Jun  8 15:19:03 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox1 ( b, l, r, t, c, cb, prog );
inout  b, l, r, t;

input  prog;

input [7:0]  cb;
input [7:0]  c;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sbox1m3to1 I232 ( .in2(r), .cb(cb[7:6]), .op(t), .in0(l), .in1(b),
     .c(c[7:6]), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb(cb[3:2]), .op(l), .in0(b), .in1(t),
     .c(c[3:2]), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb(cb[1:0]), .op(b), .in0(l), .in1(t),
     .c(c[1:0]), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb(cb[5:4]), .op(r), .in0(l), .in1(t),
     .c(c[5:4]), .prog(prog));

endmodule
// Library - xpmem, Cell - cram16x4, View - schematic
// LAST TIME SAVED: Jul 28 08:31:30 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module cram16x4 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [63:0]  q_b;
output [63:0]  q;

inout [3:0]  bl;

input [15:0]  pgate;
input [15:0]  r_gnd;
input [15:0]  wl;
input [15:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 I16_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[1:0]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[15:14]));
cram2x2 I16_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[1:0]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[13:12]));
cram2x2 I16_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[1:0]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[11:10]));
cram2x2 I16_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[1:0]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[9:8]));
cram2x2 I16_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[1:0]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[7:6]));
cram2x2 I16_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[1:0]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[5:4]));
cram2x2 I16_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[1:0]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[3:2]));
cram2x2 I16_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset_b[15:14]), .r_vdd(r_gnd[15:14]),
     .pgate(pgate[15:14]), .bl(bl[3:2]), .q_b(q_b[63:60]),
     .q(q[63:60]), .wl(wl[15:14]));
cram2x2 Imstake_6_ ( .reset(reset_b[13:12]), .r_vdd(r_gnd[13:12]),
     .pgate(pgate[13:12]), .bl(bl[3:2]), .q_b(q_b[59:56]),
     .q(q[59:56]), .wl(wl[13:12]));
cram2x2 Imstake_5_ ( .reset(reset_b[11:10]), .r_vdd(r_gnd[11:10]),
     .pgate(pgate[11:10]), .bl(bl[3:2]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[11:10]));
cram2x2 Imstake_4_ ( .reset(reset_b[9:8]), .r_vdd(r_gnd[9:8]),
     .pgate(pgate[9:8]), .bl(bl[3:2]), .q_b(q_b[51:48]), .q(q[51:48]),
     .wl(wl[9:8]));
cram2x2 Imstake_3_ ( .reset(reset_b[7:6]), .r_vdd(r_gnd[7:6]),
     .pgate(pgate[7:6]), .bl(bl[3:2]), .q_b(q_b[47:44]), .q(q[47:44]),
     .wl(wl[7:6]));
cram2x2 Imstake_2_ ( .reset(reset_b[5:4]), .r_vdd(r_gnd[5:4]),
     .pgate(pgate[5:4]), .bl(bl[3:2]), .q_b(q_b[43:40]), .q(q[43:40]),
     .wl(wl[5:4]));
cram2x2 Imstake_1_ ( .reset(reset_b[3:2]), .r_vdd(r_gnd[3:2]),
     .pgate(pgate[3:2]), .bl(bl[3:2]), .q_b(q_b[39:36]), .q(q[39:36]),
     .wl(wl[3:2]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[35:32]), .q(q[35:32]),
     .wl(wl[1:0]));

endmodule
// Library - xpmem, Cell - ml_rowdrv2, View - schematic
// LAST TIME SAVED: Aug 23 15:16:05 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_rowdrv2 ( pgate, reset, smc_rsr_out, vddctrl, wl, wl_rd_sup,
     wl_rden_b, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     por_rst, rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write );
output  pgate, reset, smc_rsr_out, vddctrl, wl;

inout  wl_rd_sup, wl_rden_b;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I163 ( .A(smc_rsr_out), .B(cram_rst), .Y(net056),
     .C(por_rst));
pch  MP0 ( .D(wl), .B(vdd_), .G(act_rd_b), .S(wl_rd_sup));
nch  M1 ( .D(wl), .B(gnd_), .G(act_rd), .S(wl_rd_sup));
nand2_hvt I182 ( .A(cram_wl_en), .Y(net057), .B(smc_rsr_out));
nand2_hvt I184 ( .A(smc_write), .Y(act_wrt_b), .B(net075));
nand2_hvt I171 ( .A(act_rd_b), .Y(off_b), .B(act_wrt_b));
nand2_hvt I159 ( .A(smc_rsr_out), .Y(net054), .B(cram_vddoff));
nand2_hvt I185 ( .A(net075), .Y(act_rd_b), .B(net073));
nand2_hvt I215 ( .A(smc_rsr_out), .Y(net0165), .B(cram_pgateoff));
inv_hvt I186 ( .A(net83), .Y(smc_rsr_out));
inv_hvt I167 ( .A(net054), .Y(vddctrl));
inv_hvt I165 ( .A(net056), .Y(reset));
inv_hvt I183 ( .A(off_b), .Y(off));
inv_hvt I170 ( .A(act_rd_b), .Y(act_rd));
inv_hvt I178 ( .A(smc_write), .Y(net073));
inv_hvt I180 ( .A(net057), .Y(net075));
inv_hvt I216 ( .A(net0165), .Y(pgate));
ml_dff_schematic I146 ( .R(rsr_rst), .D(smc_rsr_in), .CLK(smc_rsr_inc),
     .QN(net83), .Q(net0197));
nch_hvt  MN16 ( .D(wl_rden_b), .B(gnd_), .G(act_rd), .S(gnd_));
nch_hvt  MN10 ( .D(wl), .B(gnd_), .G(off), .S(gnd_));
pch_hvt  MP13 ( .D(wl), .B(vdd_), .G(act_wrt_b), .S(vdd_));

endmodule
// Library - leafcell, Cell - misc_module4rev0, View - schematic
// LAST TIME SAVED: Jun  2 13:24:00 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module misc_module4rev0 ( S_R, clk, clkb, glb2local, sp4, bl, b,
     glb_netwk, l, lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, m, min0,
     min1, min2, min3, pgate, prog, r, reset_b, sp12, vdd_cntl, wl );
output  S_R, clk, clkb;


input  prog;

output [3:0]  glb2local;
output [7:0]  sp4;

inout [3:0]  bl;

input [15:0]  wl;
input [1:0]  b;
input [1:0]  r;
input [7:0]  sp12;
input [7:0]  min3;
input [5:0]  lc_trk_g0;
input [15:0]  vdd_cntl;
input [5:0]  lc_trk_g2;
input [7:0]  min2;
input [7:0]  min1;
input [15:0]  pgate;
input [7:0]  min0;
input [5:0]  lc_trk_g3;
input [1:0]  l;
input [1:0]  m;
input [15:0]  reset_b;
input [5:0]  lc_trk_g1;
input [7:0]  glb_netwk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  r_vdd;

wire  [63:0]  cbit;

wire  [63:0]  cbitb;



clkmandcmuxrev0 Itclkm ( .min2(min2[7:0]), .min1(min1[7:0]),
     .min0(min0[7:0]), .min3(min3[7:0]), .cbit({cbit[2], cbit[1],
     cbit[0], cbit[27], cbit[25], cbit[26], cbit[24], cbit[23],
     cbit[21], cbit[22], cbit[20], cbit[19], cbit[17], cbit[18],
     cbit[16], cbit[15], cbit[13], cbit[14], cbit[12], cbit[31],
     cbit[29], cbit[30], cbit[28], cbit[11], cbit[9], cbit[10],
     cbit[8], cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}), .glb2local(glb2local[3:0]),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .glb_netwk(glb_netwk[7:0]), .prog(prog), .clk(clk), .clkb(clkb),
     .s_r(S_R));
pch_hvt  vdd_cntrl_15_ ( .D(r_vdd[15]), .B(vdd_), .G(vdd_cntl[15]),
     .S(vdd_));
pch_hvt  vdd_cntrl_14_ ( .D(r_vdd[14]), .B(vdd_), .G(vdd_cntl[14]),
     .S(vdd_));
pch_hvt  vdd_cntrl_13_ ( .D(r_vdd[13]), .B(vdd_), .G(vdd_cntl[13]),
     .S(vdd_));
pch_hvt  vdd_cntrl_12_ ( .D(r_vdd[12]), .B(vdd_), .G(vdd_cntl[12]),
     .S(vdd_));
pch_hvt  vdd_cntrl_11_ ( .D(r_vdd[11]), .B(vdd_), .G(vdd_cntl[11]),
     .S(vdd_));
pch_hvt  vdd_cntrl_10_ ( .D(r_vdd[10]), .B(vdd_), .G(vdd_cntl[10]),
     .S(vdd_));
pch_hvt  vdd_cntrl_9_ ( .D(r_vdd[9]), .B(vdd_), .G(vdd_cntl[9]),
     .S(vdd_));
pch_hvt  vdd_cntrl_8_ ( .D(r_vdd[8]), .B(vdd_), .G(vdd_cntl[8]),
     .S(vdd_));
pch_hvt  vdd_cntrl_7_ ( .D(r_vdd[7]), .B(vdd_), .G(vdd_cntl[7]),
     .S(vdd_));
pch_hvt  vdd_cntrl_6_ ( .D(r_vdd[6]), .B(vdd_), .G(vdd_cntl[6]),
     .S(vdd_));
pch_hvt  vdd_cntrl_5_ ( .D(r_vdd[5]), .B(vdd_), .G(vdd_cntl[5]),
     .S(vdd_));
pch_hvt  vdd_cntrl_4_ ( .D(r_vdd[4]), .B(vdd_), .G(vdd_cntl[4]),
     .S(vdd_));
pch_hvt  vdd_cntrl_3_ ( .D(r_vdd[3]), .B(vdd_), .G(vdd_cntl[3]),
     .S(vdd_));
pch_hvt  vdd_cntrl_2_ ( .D(r_vdd[2]), .B(vdd_), .G(vdd_cntl[2]),
     .S(vdd_));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sp12to4 Isp12to4_7_ ( .triout(sp4[7]), .cbitb(cbitb[62]),
     .drv(sp12[7]), .prog(net109));
sp12to4 Isp12to4_6_ ( .triout(sp4[6]), .cbitb(cbitb[58]),
     .drv(sp12[6]), .prog(net109));
sp12to4 Isp12to4_5_ ( .triout(sp4[5]), .cbitb(cbitb[54]),
     .drv(sp12[5]), .prog(net109));
sp12to4 Isp12to4_4_ ( .triout(sp4[4]), .cbitb(cbitb[50]),
     .drv(sp12[4]), .prog(net109));
sp12to4 Isp12to4_3_ ( .triout(sp4[3]), .cbitb(cbitb[46]),
     .drv(sp12[3]), .prog(net109));
sp12to4 Isp12to4_2_ ( .triout(sp4[2]), .cbitb(cbitb[42]),
     .drv(sp12[2]), .prog(net109));
sp12to4 Isp12to4_1_ ( .triout(sp4[1]), .cbitb(cbitb[5]), .drv(sp12[1]),
     .prog(net109));
sp12to4 Isp12to4_0_ ( .triout(sp4[0]), .cbitb(cbitb[34]),
     .drv(sp12[0]), .prog(net109));
sbox1 Isp12_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(prog));
sbox1 Isp12_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(prog));
cram16x4 Ic64 ( .r_gnd(r_vdd[15:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .q(cbit[63:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net109));

endmodule
// Library - leafcell, Cell - logic_cell, View - schematic
// LAST TIME SAVED: Aug 28 17:23:08 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module logic_cell ( carry_out, out, carry_in, cbit, clk, clkb, in0,
     in1, in2, in3, prog, purst, s_r );
output  carry_out, out;

input  carry_in, clk, clkb, in0, in1, in2, in3, prog, purst, s_r;

input [20:0]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



coredffr REG ( .purst(purst), .d(LUT4_outd), .q(rego),
     .cbit(cbit[17:16]), .clkb(clkb), .clk(clk), .S_R(s_r));
carry_logic ICARRY_LOGIC ( .b_bar(in1b1), .carry_in(carry_in), .b(in1),
     .cout(carry_out), .a(in2), .a_bar(in2b1), .vg_en(cbit[20]));
o_mux Iomux ( .in1(rego), .out(out), .cbit(cbit[19]), .prog(prog),
     .in0(LUT4_outd));
clut4 iclut4 ( .in0b(in0b1), .in3b(in3b1), .in2b(in2b1),
     .lut4(LUT4_outd), .in1b(in1b1), .in2(in2), .in1(in1), .in0(in0),
     .in3(in3), .cbit(cbit[15:0]));
inv_hvt I163 ( .A(in3), .Y(in3b1));
inv_hvt I164 ( .A(in1), .Y(in1b1));
inv_hvt I162 ( .A(in2), .Y(in2b1));
inv_hvt I161 ( .A(in0), .Y(in0b1));

endmodule
// Library - leafcell, Cell - odrv12_30, View - schematic
// LAST TIME SAVED: Jun  5 15:34:53 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module odrv12_30 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_h_r;

input  prog, slfop;

output [2:0]  sp4_h_r;
output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_r_v_b;

input [11:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



odrv12 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b[1]));
odrv12 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp12(sp12_v_b[0]));
odrv12 I70 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r));
odrv4 I69_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I71_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[2]));
odrv4 I71_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[1]));
odrv4 I71_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp4(sp4_v_b[0]));
odrv4 I73_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I73_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I73_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - xpmem, Cell - cram_2x28, View - schematic
// LAST TIME SAVED: Jul 28 08:32:33 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module cram_2x28 ( q, q_b, bl, pgate, r_vdd, reset, wl );



output [55:0]  q;
output [55:0]  q_b;

inout [27:0]  bl;

input [1:0]  wl;
input [1:0]  reset;
input [1:0]  r_vdd;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_13_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[27:26]), .q_b(q_b[55:52]),
     .q(q[55:52]), .wl(wl[1:0]));
cram2x2 Imstake_12_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[25:24]), .q_b(q_b[51:48]),
     .q(q[51:48]), .wl(wl[1:0]));
cram2x2 Imstake_11_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[23:22]), .q_b(q_b[47:44]),
     .q(q[47:44]), .wl(wl[1:0]));
cram2x2 Imstake_10_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[21:20]), .q_b(q_b[43:40]),
     .q(q[43:40]), .wl(wl[1:0]));
cram2x2 Imstake_9_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[19:18]), .q_b(q_b[39:36]),
     .q(q[39:36]), .wl(wl[1:0]));
cram2x2 Imstake_8_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[17:16]), .q_b(q_b[35:32]),
     .q(q[35:32]), .wl(wl[1:0]));
cram2x2 Imstake_7_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[15:14]), .q_b(q_b[31:28]),
     .q(q[31:28]), .wl(wl[1:0]));
cram2x2 Imstake_6_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[13:12]), .q_b(q_b[27:24]),
     .q(q[27:24]), .wl(wl[1:0]));
cram2x2 Imstake_5_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - lcmuxod3_0rev, View - schematic
// LAST TIME SAVED: Jun  2 13:13:15 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module lcmuxod3_0rev ( carry_out, cbit, cbitb, op, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1,
     min2, min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_h_r;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_v_b;
output [1:0]  sp12_v_b;
output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [55:0]  cbit;
output [55:0]  cbitb;

input [15:0]  min3;
input [27:0]  bl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [15:0]  min2;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  wl;
input [15:0]  min1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
odrv12_30 Iodrv30 ( .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - lcmuxod3_0, View - schematic
// LAST TIME SAVED: Aug 21 17:57:09 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module lcmuxod3_0 ( carry_out, op, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_h_r;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min2;
input [1:0]  wl;
input [15:0]  min3;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [27:0]  bl;
input [1:0]  pgate;
input [15:0]  min1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
odrv12_30 Iodrv30 ( .sp4_r_v_b(sp4_r_v_b[2:0]), .cbitb({cbitb[53],
     cbitb[55], cbitb[52], cbitb[54], cbitb[51], cbitb[49], cbitb[44],
     cbitb[46], cbitb[43], cbitb[41], cbitb[42], cbitb[40]}),
     .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - odrv12_74, View - schematic
// LAST TIME SAVED: Jun  5 15:30:49 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module odrv12_74 ( sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b,
     cbitb, prog, slfop );
output  sp12_v_b;

input  prog, slfop;

output [2:0]  sp4_v_b;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_h_r;

input [11:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



odrv12 I69_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[4]),
     .sp12(sp12_h_r[1]));
odrv12 I69_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[3]),
     .sp12(sp12_h_r[0]));
odrv12 I71 ( .slfop(slfop), .prog(prog), .cbitb(cbitb[8]),
     .sp12(sp12_v_b));
odrv4 I68_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[2]),
     .sp4(sp4_h_r[2]));
odrv4 I68_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[1]),
     .sp4(sp4_h_r[1]));
odrv4 I68_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[0]),
     .sp4(sp4_h_r[0]));
odrv4 I70_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[7]),
     .sp4(sp4_v_b[2]));
odrv4 I70_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[6]),
     .sp4(sp4_v_b[1]));
odrv4 I70_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[5]),
     .sp4(sp4_v_b[0]));
odrv4 I72_2_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[11]),
     .sp4(sp4_r_v_b[2]));
odrv4 I72_1_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[10]),
     .sp4(sp4_r_v_b[1]));
odrv4 I72_0_ ( .slfop(slfop), .prog(prog), .cbitb(cbitb[9]),
     .sp4(sp4_r_v_b[0]));

endmodule
// Library - leafcell, Cell - lcmuxod7_4, View - schematic
// LAST TIME SAVED: Aug 21 17:56:42 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module lcmuxod7_4 ( carry_out, op, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bl, carry_in, clk, clkb, min0, min1, min2,
     min3, pgate, prog, purst, reset_b, s_r, vdd_cntl, wl );
output  carry_out, op, sp12_v_b;

input  carry_in, clk, clkb, prog, purst, s_r;

output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [1:0]  sp12_h_r;
output [2:0]  sp4_v_b;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [15:0]  min2;
input [1:0]  reset_b;
input [15:0]  min3;
input [15:0]  min0;
input [27:0]  bl;
input [15:0]  min1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
in_mux in1mux ( .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}),
     .min(min1[15:0]), .prog(prog), .inmuxo(in1));
in_mux in0mux ( .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}),
     .min(min0[15:0]), .prog(prog), .inmuxo(in0));
in_mux in2mux ( .cbit({cbit[12], cbit[13], cbit[16], cbit[19],
     cbit[17]}), .cbitb({cbitb[12], cbitb[13], cbitb[16], cbitb[19],
     cbitb[17]}), .min(min2[15:0]), .prog(prog), .inmuxo(in2));
in_mux in3mux ( .min(min3[15:0]), .cbit({cbit[14], cbit[15], cbit[18],
     cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15], cbitb[18],
     cbitb[11], cbitb[9]}), .prog(prog), .inmuxo(in3));
logic_cell ILC ( .purst(purst), .in1(in1), .in3(in3), .in2(in2),
     .in0(in0), .s_r(s_r), .cbit({cbit[38], cbit[39], cbit[39],
     cbit[37], cbit[36], cbit[22], cbit[20], cbit[21], cbit[23],
     cbit[26], cbit[24], cbit[25], cbit[27], cbit[35], cbit[33],
     cbit[32], cbit[34], cbit[31], cbit[29], cbit[28], cbit[30]}),
     .prog(prog), .clkb(clkb), .carry_in(carry_in),
     .carry_out(carry_out), .clk(clk), .out(op));
odrv12_74 Iodrv74 ( .cbitb({cbitb[53], cbitb[55], cbitb[52], cbitb[54],
     cbitb[51], cbitb[49], cbitb[44], cbitb[46], cbitb[43], cbitb[41],
     cbitb[42], cbitb[40]}), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_h_r(sp4_h_r[2:0]),
     .sp12_v_b(sp12_v_b), .sp12_h_r(sp12_h_r[1:0]), .slfop(op),
     .prog(prog));
cram_2x28 I41 ( .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]), .q(cbit[55:0]), .wl(wl[1:0]), .bl(bl[27:0]),
     .q_b(cbitb[55:0]));

endmodule
// Library - leafcell, Cell - lccol_rev0, View - schematic
// LAST TIME SAVED: Jun 13 13:29:57 2008
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module lccol_rev0 ( carry_out, slf_op, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, cin2local, clk, clkb, lc_trk_g0, lc_trk_g1,
     lc_trk_g2, lc_trk_g3, pgate, prog, purst, reset_b, s_r, vdd_cntl,
     wl );
output  carry_out;


input  cin2local, clk, clkb, prog, purst, s_r;

output [7:0]  slf_op;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [27:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_r_v_b;

input [15:0]  wl;
input [15:0]  pgate;
input [15:0]  reset_b;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g1;
input [7:0]  lc_trk_g2;
input [7:0]  lc_trk_g3;
input [15:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [55:0]  cbit;

wire  [55:0]  cbitb;



lcmuxod3_0rev ILC_00 ( .cbitb(cbitb[55:0]), .cbit(cbit[55:0]),
     .vdd_cntl(vdd_cntl[1:0]), .purst(purst), .pgate(pgate[1:0]),
     .sp4_r_v_b({sp4_r_v_b[33], sp4_r_v_b[17], sp4_r_v_b[1]}),
     .sp12_h_r(sp12_h_r[8]), .sp12_v_b({sp12_v_b[16], sp12_v_b[0]}),
     .sp4_h_r({sp4_h_r[32], sp4_h_r[16], sp4_h_r[0]}),
     .sp4_v_b({sp4_v_b[32], sp4_v_b[16], sp4_v_b[0]}), .clk(clk),
     .carry_in(cin), .op(slf_op[0]), .carry_out(c_01), .s_r(s_r),
     .reset_b(reset_b[1:0]), .bl(bl[27:0]), .wl(wl[1:0]),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], cin}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}));
mux_4carry Icarry_cnt ( .cin(cin2local), .lcl_cin(cin),
     .cbitb({cbitb[45], cbitb[48]}), .prog(prog), .cbit({cbit[45],
     cbit[48]}));
lcmuxod3_0 ILC_02 ( .vdd_cntl(vdd_cntl[5:4]), .purst(purst),
     .pgate(pgate[5:4]), .sp4_r_v_b({sp4_r_v_b[37], sp4_r_v_b[21],
     sp4_r_v_b[5]}), .sp12_h_r(sp12_h_r[12]), .sp12_v_b({sp12_v_b[20],
     sp12_v_b[4]}), .sp4_h_r({sp4_h_r[36], sp4_h_r[20], sp4_h_r[4]}),
     .sp4_v_b({sp4_v_b[36], sp4_v_b[20], sp4_v_b[4]}), .clk(clk),
     .carry_in(c_12), .op(slf_op[2]), .carry_out(c_23), .s_r(s_r),
     .reset_b(reset_b[5:4]), .bl(bl[27:0]), .wl(wl[5:4]),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_12}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}));
lcmuxod3_0 ILC_03 ( .vdd_cntl(vdd_cntl[7:6]), .purst(purst),
     .pgate(pgate[7:6]), .sp4_r_v_b({sp4_r_v_b[39], sp4_r_v_b[23],
     sp4_r_v_b[7]}), .sp12_h_r(sp12_h_r[14]), .sp12_v_b({sp12_v_b[22],
     sp12_v_b[6]}), .sp4_h_r({sp4_h_r[38], sp4_h_r[22], sp4_h_r[6]}),
     .sp4_v_b({sp4_v_b[38], sp4_v_b[22], sp4_v_b[6]}), .clk(clk),
     .carry_in(c_23), .op(slf_op[3]), .carry_out(c_34), .s_r(s_r),
     .reset_b(reset_b[7:6]), .bl(bl[27:0]), .wl(wl[7:6]),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_23}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}));
lcmuxod3_0 ILC_01 ( .vdd_cntl(vdd_cntl[3:2]), .purst(purst),
     .pgate(pgate[3:2]), .sp4_r_v_b({sp4_r_v_b[35], sp4_r_v_b[19],
     sp4_r_v_b[3]}), .sp12_h_r(sp12_h_r[10]), .sp12_v_b({sp12_v_b[18],
     sp12_v_b[2]}), .sp4_h_r({sp4_h_r[34], sp4_h_r[18], sp4_h_r[2]}),
     .sp4_v_b({sp4_v_b[34], sp4_v_b[18], sp4_v_b[2]}), .clk(clk),
     .carry_in(c_01), .op(slf_op[1]), .carry_out(c_12), .s_r(s_r),
     .reset_b(reset_b[3:2]), .bl(bl[27:0]), .wl(wl[3:2]),
     .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_01}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}));
lcmuxod7_4 ILC_07 ( .vdd_cntl(vdd_cntl[15:14]), .purst(purst),
     .pgate(pgate[15:14]), .sp4_r_v_b({sp4_r_v_b[47], sp4_r_v_b[31],
     sp4_r_v_b[15]}), .sp12_h_r({sp12_h_r[22], sp12_h_r[6]}),
     .sp12_v_b(sp12_v_b[14]), .sp4_h_r({sp4_h_r[46], sp4_h_r[30],
     sp4_h_r[14]}), .sp4_v_b({sp4_v_b[46], sp4_v_b[30], sp4_v_b[14]}),
     .clk(clk), .carry_in(c_67), .op(slf_op[7]), .carry_out(carry_out),
     .s_r(s_r), .reset_b(reset_b[15:14]), .bl(bl[27:0]),
     .wl(wl[15:14]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_67}),
     .prog(prog), .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}));
lcmuxod7_4 ILC_06 ( .vdd_cntl(vdd_cntl[13:12]), .purst(purst),
     .pgate(pgate[13:12]), .sp4_r_v_b({sp4_r_v_b[45], sp4_r_v_b[29],
     sp4_r_v_b[13]}), .sp12_h_r({sp12_h_r[20], sp12_h_r[4]}),
     .sp12_v_b(sp12_v_b[12]), .sp4_h_r({sp4_h_r[44], sp4_h_r[28],
     sp4_h_r[12]}), .sp4_v_b({sp4_v_b[44], sp4_v_b[28], sp4_v_b[12]}),
     .clk(clk), .carry_in(c_56), .op(slf_op[6]), .carry_out(c_67),
     .s_r(s_r), .reset_b(reset_b[13:12]), .bl(bl[27:0]),
     .wl(wl[13:12]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_56}),
     .prog(prog), .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}));
lcmuxod7_4 ILC_04 ( .vdd_cntl(vdd_cntl[9:8]), .purst(purst),
     .pgate(pgate[9:8]), .sp4_r_v_b({sp4_r_v_b[41], sp4_r_v_b[25],
     sp4_r_v_b[9]}), .sp12_h_r({sp12_h_r[16], sp12_h_r[0]}),
     .sp12_v_b(sp12_v_b[8]), .sp4_h_r({sp4_h_r[40], sp4_h_r[24],
     sp4_h_r[8]}), .sp4_v_b({sp4_v_b[40], sp4_v_b[24], sp4_v_b[8]}),
     .clk(clk), .carry_in(c_34), .op(slf_op[4]), .carry_out(c_45),
     .s_r(s_r), .reset_b(reset_b[9:8]), .bl(bl[27:0]), .wl(wl[9:8]),
     .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], c_34}), .prog(prog),
     .clkb(clkb), .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3],
     lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2],
     lc_trk_g0[0]}));
lcmuxod7_4 ILC_05 ( .vdd_cntl(vdd_cntl[11:10]), .purst(purst),
     .pgate(pgate[11:10]), .sp4_r_v_b({sp4_r_v_b[43], sp4_r_v_b[27],
     sp4_r_v_b[11]}), .sp12_h_r({sp12_h_r[18], sp12_h_r[2]}),
     .sp12_v_b(sp12_v_b[10]), .sp4_h_r({sp4_h_r[42], sp4_h_r[26],
     sp4_h_r[10]}), .sp4_v_b({sp4_v_b[42], sp4_v_b[26], sp4_v_b[10]}),
     .clk(clk), .carry_in(c_45), .op(slf_op[5]), .carry_out(c_56),
     .s_r(s_r), .reset_b(reset_b[11:10]), .bl(bl[27:0]),
     .wl(wl[11:10]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], c_45}),
     .prog(prog), .clkb(clkb), .min2({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}));

endmodule
// Library - xpmem, Cell - cram2x2x5, View - schematic
// LAST TIME SAVED: Jul 28 08:25:47 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module cram2x2x5 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [19:0]  q_b;
output [19:0]  q;

inout [9:0]  bl;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  r_gnd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile_last, View - schematic
// LAST TIME SAVED: Aug  9 15:08:40 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_rowdrv_tile_last ( pgate, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  wl;
output [15:0]  reset;
output [15:0]  pgate;
output [15:0]  vddctrl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  smc_rsr_out;



nor2_hvt I211 ( .A(smc_rsr_out[15]), .Y(net049), .B(smc_rsr_inc_out));
ml_rowdrv2_last Iml_rowdrv2_last ( .smc_rsr_inc(smc_rsr_inc_last),
     .smc_rsr_in(smc_rsr_out[14]), .rsr_rst(rsr_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_rst(cram_rst_buf),
     .smc_rsr_out(smc_rsr_out[15]), .reset(reset[15]), .wl(wl[15]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]));
inv_hvt I391 ( .A(net049), .Y(smc_rsr_inc_last));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I194 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I195 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I198 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I207 ( .A(net041), .Y(por_rst_buf));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net079));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I200 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I206 ( .A(net047), .Y(rsr_rst_buf));
inv_hvt I190 ( .A(net079), .Y(smc_rsr_1st_out));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_buf), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - leafcell, Cell - sbox11to9_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:54:03 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox11to9_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[4]), .in5(t[10]), .in4(r[2]), .in3(r[10]),
     .in2(r[7]), .in1(b[10]), .in0(b[5]), .out(l[10]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[5]), .in5(t[11]), .in4(r[3]), .in3(r[11]),
     .in2(r[8]), .in1(b[11]), .in0(b[6]), .out(l[11]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[3]), .in5(t[9]), .in4(r[1]), .in3(r[9]),
     .in2(r[6]), .in1(b[9]), .in0(b[4]), .out(l[9]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[3]), .in5(r[9]), .in4(b[1]), .in3(b[9]),
     .in2(b[6]), .in1(l[9]), .in0(l[4]), .out(t[9]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[5]), .in5(r[11]), .in4(b[3]), .in3(b[11]),
     .in2(b[8]), .in1(l[11]), .in0(l[6]), .out(t[11]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[4]), .in5(r[10]), .in4(b[2]), .in3(b[10]),
     .in2(b[7]), .in1(l[10]), .in0(l[5]), .out(t[10]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox11to9_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:53:32 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox11to9_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  b;

input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[4]), .in5(b[10]), .in4(l[2]), .in3(l[10]),
     .in2(l[7]), .in1(t[10]), .in0(t[5]), .out(r[10]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[5]), .in5(b[11]), .in4(l[3]), .in3(l[11]),
     .in2(l[8]), .in1(t[11]), .in0(t[6]), .out(r[11]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[3]), .in5(b[9]), .in4(l[1]), .in3(l[9]),
     .in2(l[6]), .in1(t[9]), .in0(t[4]), .out(r[9]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[4]), .in5(l[10]), .in4(t[2]), .in3(t[10]),
     .in2(t[7]), .in1(r[10]), .in0(r[5]), .out(b[10]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[5]), .in5(l[11]), .in4(t[3]), .in3(t[11]),
     .in2(t[8]), .in1(r[11]), .in0(r[6]), .out(b[11]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[3]), .in5(l[9]), .in4(t[1]), .in3(t[9]),
     .in2(t[6]), .in1(r[9]), .in0(r[4]), .out(b[9]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox8to6_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:52:49 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox8to6_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  t;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;

input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[1]), .in5(t[7]), .in4(r[11]), .in3(r[7]),
     .in2(r[4]), .in1(b[7]), .in0(b[2]), .out(l[7]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[2]), .in5(t[8]), .in4(r[0]), .in3(r[8]),
     .in2(r[5]), .in1(b[8]), .in0(b[3]), .out(l[8]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[0]), .in5(t[6]), .in4(r[10]), .in3(r[6]),
     .in2(r[3]), .in1(b[6]), .in0(b[1]), .out(l[6]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[0]), .in5(r[6]), .in4(b[10]), .in3(b[6]),
     .in2(b[3]), .in1(l[6]), .in0(l[1]), .out(t[6]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[2]), .in5(r[8]), .in4(b[0]), .in3(b[8]),
     .in2(b[5]), .in1(l[8]), .in0(l[3]), .out(t[8]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[1]), .in5(r[7]), .in4(b[11]), .in3(b[7]),
     .in2(b[4]), .in1(l[7]), .in0(l[2]), .out(t[7]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox8to6_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:36:51 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox8to6_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  cbit;

wire  [19:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[1]), .in5(b[7]), .in4(l[11]), .in3(l[7]),
     .in2(l[4]), .in1(t[7]), .in0(t[2]), .out(r[7]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[2]), .in5(b[8]), .in4(l[0]), .in3(l[8]),
     .in2(l[5]), .in1(t[8]), .in0(t[3]), .out(r[8]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[0]), .in5(b[6]), .in4(l[10]), .in3(l[6]),
     .in2(l[3]), .in1(t[6]), .in0(t[1]), .out(r[6]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[1]), .in5(l[7]), .in4(t[11]), .in3(t[7]),
     .in2(t[4]), .in1(r[7]), .in0(r[2]), .out(b[7]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[2]), .in5(l[8]), .in4(t[0]), .in3(t[8]),
     .in2(t[5]), .in1(r[8]), .in0(r[3]), .out(b[8]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[0]), .in5(l[6]), .in4(t[10]), .in3(t[6]),
     .in2(t[3]), .in1(r[6]), .in0(r[1]), .out(b[6]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox5to3_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:36:06 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox5to3_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  l;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  t;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[10]), .in5(t[4]), .in4(r[8]), .in3(r[4]),
     .in2(r[1]), .in1(b[4]), .in0(b[11]), .out(l[4]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[11]), .in5(t[5]), .in4(r[9]), .in3(r[5]),
     .in2(r[2]), .in1(b[5]), .in0(b[0]), .out(l[5]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[9]), .in5(t[3]), .in4(r[7]), .in3(r[3]),
     .in2(r[0]), .in1(b[3]), .in0(b[10]), .out(l[3]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[9]), .in5(r[3]), .in4(b[7]), .in3(b[3]),
     .in2(b[0]), .in1(l[3]), .in0(l[10]), .out(t[3]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[11]), .in5(r[5]), .in4(b[9]), .in3(b[5]),
     .in2(b[2]), .in1(l[5]), .in0(l[0]), .out(t[5]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[10]), .in5(r[4]), .in4(b[8]), .in3(b[4]),
     .in2(b[1]), .in1(l[4]), .in0(l[11]), .out(t[4]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 I534 ( .q(cbit[19:0]), .r_gnd(r_vdd[1:0]),
     .reset_b(reset_b[1:0]), .wl(wl[1:0]), .bl(bl[9:0]),
     .q_b(cbitb[19:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - sbox5to3_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:35:35 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox5to3_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;

input [1:0]  wl;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbitb;

wire  [19:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[10]), .in5(b[4]), .in4(l[8]), .in3(l[4]),
     .in2(l[1]), .in1(t[4]), .in0(t[11]), .out(r[4]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[11]), .in5(b[5]), .in4(l[9]), .in3(l[5]),
     .in2(l[2]), .in1(t[5]), .in0(t[0]), .out(r[5]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[9]), .in5(b[3]), .in4(l[7]), .in3(l[3]),
     .in2(l[0]), .in1(t[3]), .in0(t[10]), .out(r[3]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[10]), .in5(l[4]), .in4(t[8]), .in3(t[4]),
     .in2(t[1]), .in1(r[4]), .in0(r[11]), .out(b[4]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[11]), .in5(l[5]), .in4(t[9]), .in3(t[5]),
     .in2(t[2]), .in1(r[5]), .in0(r[0]), .out(b[5]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[9]), .in5(l[3]), .in4(t[7]), .in3(t[3]),
     .in2(t[0]), .in1(r[3]), .in0(r[10]), .out(b[3]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox2to0_220_p2, View - schematic
// LAST TIME SAVED: Aug 21 17:35:04 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox2to0_220_p2 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  l;
inout [11:0]  b;
inout [11:0]  t;
inout [11:0]  r;

input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [19:0]  cbit;

wire  [19:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I525 ( .in6(t[7]), .in5(t[1]), .in4(r[5]), .in3(r[1]),
     .in2(r[10]), .in1(b[1]), .in0(b[8]), .out(l[1]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I526 ( .in6(t[8]), .in5(t[2]), .in4(r[6]), .in3(r[2]),
     .in2(r[11]), .in1(b[2]), .in0(b[9]), .out(l[2]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I527 ( .in6(t[6]), .in5(t[0]), .in4(r[4]), .in3(r[0]),
     .in2(r[9]), .in1(b[0]), .in0(b[7]), .out(l[0]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I528 ( .in6(r[6]), .in5(r[0]), .in4(b[4]), .in3(b[0]),
     .in2(b[9]), .in1(l[0]), .in0(l[7]), .out(t[0]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
sbox7to1_220 I529 ( .in6(r[8]), .in5(r[2]), .in4(b[6]), .in3(b[2]),
     .in2(b[11]), .in1(l[2]), .in0(l[9]), .out(t[2]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I530 ( .in6(r[7]), .in5(r[1]), .in4(b[5]), .in3(b[1]),
     .in2(b[10]), .in1(l[1]), .in0(l[8]), .out(t[1]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - sbox2to0_220_p1, View - schematic
// LAST TIME SAVED: Aug 21 17:34:25 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module sbox2to0_220_p1 ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [11:0]  r;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;
inout [9:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [19:0]  cbit;

wire  [19:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox7to1_220 I509 ( .in6(b[7]), .in5(b[1]), .in4(l[5]), .in3(l[1]),
     .in2(l[10]), .in1(t[1]), .in0(t[8]), .out(r[1]), .c({cbit[10],
     cbit[11], cbit[14]}), .cb({cbitb[10], cbitb[11], cbitb[14]}),
     .prog(prog));
sbox7to1_220 I510 ( .in6(b[8]), .in5(b[2]), .in4(l[6]), .in3(l[2]),
     .in2(l[11]), .in1(t[2]), .in0(t[9]), .out(r[2]), .c({cbit[13],
     cbit[18], cbit[17]}), .cb({cbitb[13], cbitb[18], cbitb[17]}),
     .prog(prog));
sbox7to1_220 I508 ( .in6(b[6]), .in5(b[0]), .in4(l[4]), .in3(l[0]),
     .in2(l[9]), .in1(t[0]), .in0(t[7]), .out(r[0]), .c({cbit[4],
     cbit[3], cbit[0]}), .cb({cbitb[4], cbitb[3], cbitb[0]}),
     .prog(prog));
sbox7to1_220 I523 ( .in6(l[7]), .in5(l[1]), .in4(t[5]), .in3(t[1]),
     .in2(t[10]), .in1(r[1]), .in0(r[8]), .out(b[1]), .c({cbit[9],
     cbit[8], cbit[12]}), .cb({cbitb[9], cbitb[8], cbitb[12]}),
     .prog(prog));
sbox7to1_220 I522 ( .in6(l[8]), .in5(l[2]), .in4(t[6]), .in3(t[2]),
     .in2(t[11]), .in1(r[2]), .in0(r[9]), .out(b[2]), .c({cbit[19],
     cbit[16], cbit[15]}), .cb({cbitb[19], cbitb[16], cbitb[15]}),
     .prog(prog));
sbox7to1_220 I524 ( .in6(l[6]), .in5(l[0]), .in4(t[4]), .in3(t[0]),
     .in2(t[9]), .in1(r[0]), .in0(r[7]), .out(b[0]), .c({cbit[2],
     cbit[1], cbit[6]}), .cb({cbitb[2], cbitb[1], cbitb[6]}),
     .prog(prog));
cram2x2x5 Imem20 ( .pgate(pgate[1:0]), .q(cbit[19:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[9:0]), .q_b(cbitb[19:0]));

endmodule
// Library - leafcell, Cell - span4_switchandmem, View - schematic
// LAST TIME SAVED: Jul 24 12:49:53 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module span4_switchandmem ( b, bl, l, r, t, pgate, prog, reset_b,
     vdd_cntl, wl );

input  prog;

inout [9:0]  bl;
inout [11:0]  b;
inout [11:0]  l;
inout [11:0]  t;
inout [11:0]  r;

input [15:0]  wl;
input [15:0]  reset_b;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sbox11to9_220_p2 I73 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .l(l[11:0]), .r(r[11:0]), .t(t[11:0]),
     .b(b[11:0]), .prog(prog), .wl(wl[15:14]), .bl(bl[9:0]),
     .reset_b(reset_b[15:14]));
sbox11to9_220_p1 I75 ( .vdd_cntl(vdd_cntl[13:12]),
     .pgate(pgate[13:12]), .l(l[11:0]), .r(r[11:0]), .t(t[11:0]),
     .b(b[11:0]), .prog(prog), .wl(wl[13:12]), .bl(bl[9:0]),
     .reset_b(reset_b[13:12]));
sbox8to6_220_p2 I74 ( .vdd_cntl(vdd_cntl[11:10]), .pgate(pgate[11:10]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[11:10]), .bl(bl[9:0]), .reset_b(reset_b[11:10]));
sbox8to6_220_p1 I76 ( .vdd_cntl(vdd_cntl[9:8]), .pgate(pgate[9:8]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[9:8]), .bl(bl[9:0]), .reset_b(reset_b[9:8]));
sbox5to3_220_p2 I71 ( .vdd_cntl(vdd_cntl[7:6]), .pgate(pgate[7:6]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[7:6]), .bl(bl[9:0]), .reset_b(reset_b[7:6]));
sbox5to3_220_p1 I72 ( .vdd_cntl(vdd_cntl[5:4]), .pgate(pgate[5:4]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[5:4]), .bl(bl[9:0]), .reset_b(reset_b[5:4]));
sbox2to0_220_p2 I70 ( .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[3:2]), .bl(bl[9:0]), .reset_b(reset_b[3:2]));
sbox2to0_220_p1 I69 ( .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]),
     .l(l[11:0]), .r(r[11:0]), .t(t[11:0]), .b(b[11:0]), .prog(prog),
     .wl(wl[1:0]), .bl(bl[9:0]), .reset_b(reset_b[1:0]));

endmodule
// Library - leafcell, Cell - span4, View - schematic
// LAST TIME SAVED: Sep  5 23:05:28 2007
// NETLIST TIME: Nov 14 16:17:14 2008
`timescale 1ns / 1ns 

module span4 ( bl, sp4_h_l, sp4_h_r, sp4_v_b, sp4_v_t, pgate, prog,
     reset_b, vdd_cntl, wl );

input  prog;

inout [47:0]  sp4_v_b;
inout [9:0]  bl;
inout [47:0]  sp4_h_l;
inout [47:0]  sp4_v_t;
inout [47:0]  sp4_h_r;

input [15:0]  vdd_cntl;
input [15:0]  reset_b;
input [15:0]  wl;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  sp4_h_r_mid;

wire  [11:0]  sp4_v_b_mid;



rm7  R1_27_ ( .MINUS(sp4_h_r[47]), .PLUS(sp4_h_l[34]));
rm7  R1_26_ ( .MINUS(sp4_h_r[46]), .PLUS(sp4_h_l[35]));
rm7  R1_25_ ( .MINUS(sp4_h_r[45]), .PLUS(sp4_h_l[32]));
rm7  R1_24_ ( .MINUS(sp4_h_r[44]), .PLUS(sp4_h_l[33]));
rm7  R1_23_ ( .MINUS(sp4_h_r[43]), .PLUS(sp4_h_l[30]));
rm7  R1_22_ ( .MINUS(sp4_h_r[42]), .PLUS(sp4_h_l[31]));
rm7  R1_21_ ( .MINUS(sp4_h_r[41]), .PLUS(sp4_h_l[28]));
rm7  R1_20_ ( .MINUS(sp4_h_r[40]), .PLUS(sp4_h_l[29]));
rm7  R1_19_ ( .MINUS(sp4_h_r[39]), .PLUS(sp4_h_l[26]));
rm7  R1_18_ ( .MINUS(sp4_h_r[38]), .PLUS(sp4_h_l[27]));
rm7  R1_17_ ( .MINUS(sp4_h_r[37]), .PLUS(sp4_h_l[24]));
rm7  R1_16_ ( .MINUS(sp4_h_r[36]), .PLUS(sp4_h_l[25]));
rm7  R1_15_ ( .MINUS(sp4_h_r[35]), .PLUS(sp4_h_l[22]));
rm7  R1_14_ ( .MINUS(sp4_h_r[34]), .PLUS(sp4_h_l[23]));
rm7  R1_13_ ( .MINUS(sp4_h_r[23]), .PLUS(sp4_h_l[10]));
rm7  R1_12_ ( .MINUS(sp4_h_r[22]), .PLUS(sp4_h_l[11]));
rm7  R1_11_ ( .MINUS(sp4_h_r_mid[11]), .PLUS(sp4_h_l[46]));
rm7  R1_10_ ( .MINUS(sp4_h_r_mid[10]), .PLUS(sp4_h_l[47]));
rm7  R1_9_ ( .MINUS(sp4_h_r_mid[9]), .PLUS(sp4_h_l[44]));
rm7  R1_8_ ( .MINUS(sp4_h_r_mid[8]), .PLUS(sp4_h_l[45]));
rm7  R1_7_ ( .MINUS(sp4_h_r_mid[7]), .PLUS(sp4_h_l[42]));
rm7  R1_6_ ( .MINUS(sp4_h_r_mid[6]), .PLUS(sp4_h_l[43]));
rm7  R1_5_ ( .MINUS(sp4_h_r_mid[5]), .PLUS(sp4_h_l[40]));
rm7  R1_4_ ( .MINUS(sp4_h_r_mid[4]), .PLUS(sp4_h_l[41]));
rm7  R1_3_ ( .MINUS(sp4_h_r_mid[3]), .PLUS(sp4_h_l[38]));
rm7  R1_2_ ( .MINUS(sp4_h_r_mid[2]), .PLUS(sp4_h_l[39]));
rm7  R1_1_ ( .MINUS(sp4_h_r_mid[1]), .PLUS(sp4_h_l[36]));
rm7  R1_0_ ( .MINUS(sp4_h_r_mid[0]), .PLUS(sp4_h_l[37]));
rm5  R2_19_ ( .MINUS(sp4_h_r[33]), .PLUS(sp4_h_l[20]));
rm5  R2_18_ ( .MINUS(sp4_h_r[32]), .PLUS(sp4_h_l[21]));
rm5  R2_17_ ( .MINUS(sp4_h_r[31]), .PLUS(sp4_h_l[18]));
rm5  R2_16_ ( .MINUS(sp4_h_r[30]), .PLUS(sp4_h_l[19]));
rm5  R2_15_ ( .MINUS(sp4_h_r[29]), .PLUS(sp4_h_l[16]));
rm5  R2_14_ ( .MINUS(sp4_h_r[28]), .PLUS(sp4_h_l[17]));
rm5  R2_13_ ( .MINUS(sp4_h_r[27]), .PLUS(sp4_h_l[14]));
rm5  R2_12_ ( .MINUS(sp4_h_r[26]), .PLUS(sp4_h_l[15]));
rm5  R2_11_ ( .MINUS(sp4_h_r[25]), .PLUS(sp4_h_l[12]));
rm5  R2_10_ ( .MINUS(sp4_h_r[24]), .PLUS(sp4_h_l[13]));
rm5  R2_9_ ( .MINUS(sp4_h_r[21]), .PLUS(sp4_h_l[8]));
rm5  R2_8_ ( .MINUS(sp4_h_r[20]), .PLUS(sp4_h_l[9]));
rm5  R2_7_ ( .MINUS(sp4_h_r[19]), .PLUS(sp4_h_l[6]));
rm5  R2_6_ ( .MINUS(sp4_h_r[18]), .PLUS(sp4_h_l[7]));
rm5  R2_5_ ( .MINUS(sp4_h_r[17]), .PLUS(sp4_h_l[4]));
rm5  R2_4_ ( .MINUS(sp4_h_r[16]), .PLUS(sp4_h_l[5]));
rm5  R2_3_ ( .MINUS(sp4_h_r[15]), .PLUS(sp4_h_l[2]));
rm5  R2_2_ ( .MINUS(sp4_h_r[14]), .PLUS(sp4_h_l[3]));
rm5  R2_1_ ( .MINUS(sp4_h_r[13]), .PLUS(sp4_h_l[0]));
rm5  R2_0_ ( .MINUS(sp4_h_r[12]), .PLUS(sp4_h_l[1]));
rm6  R0_47_ ( .MINUS(sp4_v_b[47]), .PLUS(sp4_v_t[34]));
rm6  R0_46_ ( .MINUS(sp4_v_b[46]), .PLUS(sp4_v_t[35]));
rm6  R0_45_ ( .MINUS(sp4_v_b[45]), .PLUS(sp4_v_t[32]));
rm6  R0_44_ ( .MINUS(sp4_v_b[44]), .PLUS(sp4_v_t[33]));
rm6  R0_43_ ( .MINUS(sp4_v_b[43]), .PLUS(sp4_v_t[30]));
rm6  R0_42_ ( .MINUS(sp4_v_b[42]), .PLUS(sp4_v_t[31]));
rm6  R0_41_ ( .MINUS(sp4_v_b[41]), .PLUS(sp4_v_t[28]));
rm6  R0_40_ ( .MINUS(sp4_v_b[40]), .PLUS(sp4_v_t[29]));
rm6  R0_39_ ( .MINUS(sp4_v_b[39]), .PLUS(sp4_v_t[26]));
rm6  R0_38_ ( .MINUS(sp4_v_b[38]), .PLUS(sp4_v_t[27]));
rm6  R0_37_ ( .MINUS(sp4_v_b[37]), .PLUS(sp4_v_t[24]));
rm6  R0_36_ ( .MINUS(sp4_v_b[36]), .PLUS(sp4_v_t[25]));
rm6  R0_35_ ( .MINUS(sp4_v_b[35]), .PLUS(sp4_v_t[22]));
rm6  R0_34_ ( .MINUS(sp4_v_b[34]), .PLUS(sp4_v_t[23]));
rm6  R0_33_ ( .MINUS(sp4_v_b[33]), .PLUS(sp4_v_t[20]));
rm6  R0_32_ ( .MINUS(sp4_v_b[32]), .PLUS(sp4_v_t[21]));
rm6  R0_31_ ( .MINUS(sp4_v_b[31]), .PLUS(sp4_v_t[18]));
rm6  R0_30_ ( .MINUS(sp4_v_b[30]), .PLUS(sp4_v_t[19]));
rm6  R0_29_ ( .MINUS(sp4_v_b[29]), .PLUS(sp4_v_t[16]));
rm6  R0_28_ ( .MINUS(sp4_v_b[28]), .PLUS(sp4_v_t[17]));
rm6  R0_27_ ( .MINUS(sp4_v_b[27]), .PLUS(sp4_v_t[14]));
rm6  R0_26_ ( .MINUS(sp4_v_b[26]), .PLUS(sp4_v_t[15]));
rm6  R0_25_ ( .MINUS(sp4_v_b[25]), .PLUS(sp4_v_t[12]));
rm6  R0_24_ ( .MINUS(sp4_v_b[24]), .PLUS(sp4_v_t[13]));
rm6  R0_23_ ( .MINUS(sp4_v_b[23]), .PLUS(sp4_v_t[10]));
rm6  R0_22_ ( .MINUS(sp4_v_b[22]), .PLUS(sp4_v_t[11]));
rm6  R0_21_ ( .MINUS(sp4_v_b[21]), .PLUS(sp4_v_t[8]));
rm6  R0_20_ ( .MINUS(sp4_v_b[20]), .PLUS(sp4_v_t[9]));
rm6  R0_19_ ( .MINUS(sp4_v_b[19]), .PLUS(sp4_v_t[6]));
rm6  R0_18_ ( .MINUS(sp4_v_b[18]), .PLUS(sp4_v_t[7]));
rm6  R0_17_ ( .MINUS(sp4_v_b[17]), .PLUS(sp4_v_t[4]));
rm6  R0_16_ ( .MINUS(sp4_v_b[16]), .PLUS(sp4_v_t[5]));
rm6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[2]));
rm6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[3]));
rm6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[0]));
rm6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[1]));
rm6  R0_11_ ( .MINUS(sp4_v_b_mid[11]), .PLUS(sp4_v_t[46]));
rm6  R0_10_ ( .MINUS(sp4_v_b_mid[10]), .PLUS(sp4_v_t[47]));
rm6  R0_9_ ( .MINUS(sp4_v_b_mid[9]), .PLUS(sp4_v_t[44]));
rm6  R0_8_ ( .MINUS(sp4_v_b_mid[8]), .PLUS(sp4_v_t[45]));
rm6  R0_7_ ( .MINUS(sp4_v_b_mid[7]), .PLUS(sp4_v_t[42]));
rm6  R0_6_ ( .MINUS(sp4_v_b_mid[6]), .PLUS(sp4_v_t[43]));
rm6  R0_5_ ( .MINUS(sp4_v_b_mid[5]), .PLUS(sp4_v_t[40]));
rm6  R0_4_ ( .MINUS(sp4_v_b_mid[4]), .PLUS(sp4_v_t[41]));
rm6  R0_3_ ( .MINUS(sp4_v_b_mid[3]), .PLUS(sp4_v_t[38]));
rm6  R0_2_ ( .MINUS(sp4_v_b_mid[2]), .PLUS(sp4_v_t[39]));
rm6  R0_1_ ( .MINUS(sp4_v_b_mid[1]), .PLUS(sp4_v_t[36]));
rm6  R0_0_ ( .MINUS(sp4_v_b_mid[0]), .PLUS(sp4_v_t[37]));
span4_switchandmem ISPAN4_SW ( .vdd_cntl(vdd_cntl[15:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]), .b(sp4_v_b[11:0]),
     .r(sp4_h_r[11:0]), .l(sp4_h_r_mid[11:0]), .prog(prog),
     .wl(wl[15:0]), .t(sp4_v_b_mid[11:0]), .bl(bl[9:0]));

endmodule
// Library - xpmem, Cell - ml_rowdrv_tile, View - schematic
// LAST TIME SAVED: Aug 15 11:21:19 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_rowdrv_tile ( pgate, por_rst_out, reset, smc_rsr_1st_out,
     smc_rsr_inc_out, smcc_rsr_out, vddctrl, wl, cram_pgateoff,
     cram_rst, cram_vddoff, cram_wl_en, por_rst, rsr_rst, smc_rsr_in,
     smc_rsr_inc, smc_write );
output  por_rst_out, smc_rsr_1st_out, smc_rsr_inc_out, smcc_rsr_out;

input  cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en, por_rst,
     rsr_rst, smc_rsr_in, smc_rsr_inc, smc_write;

output [15:0]  vddctrl;
output [15:0]  reset;
output [15:0]  pgate;
output [15:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  smc_rsr_out;



inv_hvt I207 ( .A(net041), .Y(por_rst_out));
inv_hvt I192 ( .A(smc_write), .Y(net069));
inv_hvt I293 ( .A(net069), .Y(smc_write_buf));
inv_hvt I193 ( .A(cram_pgateoff), .Y(net067));
inv_hvt I194 ( .A(net067), .Y(cram_pateoff_buf));
inv_hvt I286 ( .A(smc_rsr_out[15]), .Y(net62));
inv_hvt I195 ( .A(net061), .Y(cram_vddoff_buf));
inv_hvt I196 ( .A(cram_vddoff), .Y(net061));
inv_hvt I197 ( .A(cram_rst), .Y(net057));
inv_hvt I198 ( .A(net057), .Y(cram_rst_buf));
inv_hvt I199 ( .A(cram_wl_en), .Y(net055));
inv_hvt I190 ( .A(net037), .Y(smc_rsr_1st_out));
inv_hvt I203 ( .A(smc_rsr_inc), .Y(net051));
inv_hvt I204 ( .A(net051), .Y(smc_rsr_inc_out));
inv_hvt I191 ( .A(smc_rsr_out[0]), .Y(net037));
inv_hvt I205 ( .A(rsr_rst), .Y(net047));
inv_hvt I208 ( .A(por_rst), .Y(net041));
inv_hvt I200 ( .A(net055), .Y(cram_wl_en_buf));
inv_hvt I281 ( .A(net62), .Y(smcc_rsr_out));
inv_hvt I206 ( .A(net047), .Y(rsr_rst_buf));
ml_rowdrvsup2 Iml_rowdrvsup2 ( .wl_rden_b(wl_rden_b),
     .wl_rd_sup(wl_rd_sup));
ml_rowdrv2 Iml_rowdrv2_15_ ( .reset(reset[15]), .wl(wl[15]),
     .vddctrl(vddctrl[15]), .pgate(pgate[15]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[14]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[15]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_14_ ( .reset(reset[14]), .wl(wl[14]),
     .vddctrl(vddctrl[14]), .pgate(pgate[14]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[14]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_13_ ( .reset(reset[13]), .wl(wl[13]),
     .vddctrl(vddctrl[13]), .pgate(pgate[13]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[13]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_12_ ( .reset(reset[12]), .wl(wl[12]),
     .vddctrl(vddctrl[12]), .pgate(pgate[12]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[12]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_11_ ( .reset(reset[11]), .wl(wl[11]),
     .vddctrl(vddctrl[11]), .pgate(pgate[11]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[11]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_10_ ( .reset(reset[10]), .wl(wl[10]),
     .vddctrl(vddctrl[10]), .pgate(pgate[10]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[10]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_9_ ( .reset(reset[9]), .wl(wl[9]),
     .vddctrl(vddctrl[9]), .pgate(pgate[9]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[9]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_8_ ( .reset(reset[8]), .wl(wl[8]),
     .vddctrl(vddctrl[8]), .pgate(pgate[8]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[8]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_7_ ( .reset(reset[7]), .wl(wl[7]),
     .vddctrl(vddctrl[7]), .pgate(pgate[7]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[7]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_6_ ( .reset(reset[6]), .wl(wl[6]),
     .vddctrl(vddctrl[6]), .pgate(pgate[6]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[6]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_5_ ( .reset(reset[5]), .wl(wl[5]),
     .vddctrl(vddctrl[5]), .pgate(pgate[5]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[5]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_4_ ( .reset(reset[4]), .wl(wl[4]),
     .vddctrl(vddctrl[4]), .pgate(pgate[4]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[4]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_3_ ( .reset(reset[3]), .wl(wl[3]),
     .vddctrl(vddctrl[3]), .pgate(pgate[3]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[3]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_2_ ( .reset(reset[2]), .wl(wl[2]),
     .vddctrl(vddctrl[2]), .pgate(pgate[2]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[2]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_1_ ( .reset(reset[1]), .wl(wl[1]),
     .vddctrl(vddctrl[1]), .pgate(pgate[1]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[1]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));
ml_rowdrv2 Iml_rowdrv2_0_ ( .reset(reset[0]), .wl(wl[0]),
     .vddctrl(vddctrl[0]), .pgate(pgate[0]),
     .smc_rsr_inc(smc_rsr_inc_out), .smc_rsr_in(smc_rsr_in),
     .rsr_rst(rsr_rst_buf), .cram_wl_en(cram_wl_en_buf),
     .cram_rst(cram_rst_buf), .smc_rsr_out(smc_rsr_out[0]),
     .por_rst(por_rst_out), .smc_write(smc_write_buf),
     .cram_vddoff(cram_vddoff_buf), .wl_rd_sup(wl_rd_sup),
     .wl_rden_b(wl_rden_b), .cram_pgateoff(cram_pateoff_buf));

endmodule
// Library - xpmem, Cell - cram2x2x6, View - schematic
// LAST TIME SAVED: Jul 28 08:29:06 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module cram2x2x6 ( q, q_b, bl, pgate, r_gnd, reset_b, wl );



output [23:0]  q;
output [23:0]  q_b;

inout [11:0]  bl;

input [1:0]  reset_b;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  r_gnd;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cram2x2 Imstake_5_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[11:10]), .q_b(q_b[23:20]),
     .q(q[23:20]), .wl(wl[1:0]));
cram2x2 Imstake_4_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[9:8]), .q_b(q_b[19:16]), .q(q[19:16]),
     .wl(wl[1:0]));
cram2x2 Imstake_3_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[7:6]), .q_b(q_b[15:12]), .q(q[15:12]),
     .wl(wl[1:0]));
cram2x2 Imstake_2_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[5:4]), .q_b(q_b[11:8]), .q(q[11:8]),
     .wl(wl[1:0]));
cram2x2 Imstake_1_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[3:2]), .q_b(q_b[7:4]), .q(q[7:4]),
     .wl(wl[1:0]));
cram2x2 Imstake_0_ ( .reset(reset_b[1:0]), .r_vdd(r_gnd[1:0]),
     .pgate(pgate[1:0]), .bl(bl[1:0]), .q_b(q_b[3:0]), .q(q[3:0]),
     .wl(wl[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_base, View - schematic
// LAST TIME SAVED: Sep 13 06:51:33 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_base ( lc_trk_out, sp4_out, bl, min0, min1, min2,
     min3, pgate, prog, reset_b, sp12_in, vdd_cntl, wl );


input  prog;

output [1:0]  sp4_out;
output [3:0]  lc_trk_out;

inout [11:0]  bl;

input [1:0]  wl;
input [1:0]  sp12_in;
input [15:0]  min1;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [15:0]  min3;
input [1:0]  pgate;
input [15:0]  min0;
input [15:0]  min2;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [23:0]  cbitb;

wire  [23:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
g_mux Imux2 ( .min(min2[15:0]), .prog(net60), .inmuxo(lc_trk_out[2]),
     .cbit({cbit[16], cbit[17], cbit[20], cbit[23], cbit[21]}),
     .cbitb({cbitb[16], cbitb[17], cbitb[20], cbitb[23], cbitb[21]}));
g_mux Imux3 ( .min(min3[15:0]), .prog(net60), .inmuxo(lc_trk_out[3]),
     .cbit({cbit[18], cbit[19], cbit[22], cbit[15], cbit[13]}),
     .cbitb({cbitb[18], cbitb[19], cbitb[22], cbitb[15], cbitb[13]}));
g_mux Imux1 ( .min(min1[15:0]), .prog(net60), .inmuxo(lc_trk_out[1]),
     .cbit({cbit[7], cbit[6], cbit[3], cbit[10], cbit[8]}),
     .cbitb({cbitb[7], cbitb[6], cbitb[3], cbitb[10], cbitb[8]}));
g_mux Imux0 ( .min(min0[15:0]), .prog(net60), .inmuxo(lc_trk_out[0]),
     .cbit({cbit[5], cbit[4], cbit[1], cbit[2], cbit[0]}),
     .cbitb({cbitb[5], cbitb[4], cbitb[1], cbitb[2], cbitb[0]}));
cram2x2x6 Imem2x2x6 ( .pgate(pgate[1:0]), .q(cbit[23:0]),
     .r_gnd(r_vdd[1:0]), .reset_b(reset_b[1:0]), .wl(wl[1:0]),
     .bl(bl[11:0]), .q_b(cbitb[23:0]));
sp12to4 Isp12to4_1_ ( .triout(sp4_out[1]), .cbitb(cbitb[11]),
     .drv(sp12_in[1]), .prog(net60));
sp12to4 Isp12to4_0_ ( .triout(sp4_out[0]), .cbitb(cbitb[9]),
     .drv(sp12_in[0]), .prog(net60));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net60));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0a, View - schematic
// LAST TIME SAVED: Jul 24 13:27:07 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g0a ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g0;

inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;

input [7:0]  tnl_op;
input [1:0]  vdd_cntl;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[34], sp4_r_v_b[25]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[33], sp4_r_v_b[26]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[35], sp4_r_v_b[24]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[32], sp4_r_v_b[27]}),
     .sp4_out(sp4_v_b[13:12]), .sp12_in({sp12_v_b[3], sp12_v_b[1]}),
     .lc_trk_out(lc_trk_g0[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g0b, View - schematic
// LAST TIME SAVED: Jul 24 13:26:14 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g0b ( lc_trk_g0, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, glb2local, lft_op,
     pgate, prog, reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op,
     vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g0;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [1:0]  pgate;
input [1:0]  wl;
input [3:0]  glb2local;
input [7:0]  bnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  top_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g0b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], glb2local[1]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], glb2local[2]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], glb2local[0]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], glb2local[3]}),
     .sp4_out(sp4_v_b[15:14]), .sp12_in({sp12_v_b[7], sp12_v_b[5]}),
     .lc_trk_out(lc_trk_g0[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1a, View - schematic
// LAST TIME SAVED: Jul 24 13:25:29 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g1a ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_v_b;

input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [1:0]  wl;
input [7:0]  bnl_op;
input [7:0]  bnr_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[17], sp4_h_r[9], sp4_h_r[1], sp4_v_b[17],
     sp4_v_b[9], sp4_v_b[1], sp12_h_r[17], sp12_h_r[9], sp12_h_r[1],
     lft_op[1], top_op[1], bot_op[1], bnr_op[1], slf_op[1],
     sp4_r_v_b[25], sp4_r_v_b[1]}), .min2({sp4_h_r[18], sp4_h_r[10],
     sp4_h_r[2], sp4_v_b[18], sp4_v_b[10], sp4_v_b[2], sp12_h_r[18],
     sp12_h_r[10], sp12_h_r[2], lft_op[2], top_op[2], bot_op[2],
     bnr_op[2], slf_op[2], sp4_r_v_b[26], sp4_r_v_b[2]}),
     .min0({sp4_h_r[16], sp4_h_r[8], sp4_h_r[0], sp4_v_b[16],
     sp4_v_b[8], sp4_v_b[0], sp12_h_r[16], sp12_h_r[8], sp12_h_r[0],
     lft_op[0], top_op[0], bot_op[0], bnr_op[0], slf_op[0],
     sp4_r_v_b[24], sp4_r_v_b[0]}), .min3({sp4_h_r[19], sp4_h_r[11],
     sp4_h_r[3], sp4_v_b[19], sp4_v_b[11], sp4_v_b[3], sp12_h_r[19],
     sp12_h_r[11], sp12_h_r[3], lft_op[3], top_op[3], bot_op[3],
     bnr_op[3], slf_op[3], sp4_r_v_b[27], sp4_r_v_b[3]}),
     .sp4_out(sp4_v_b[17:16]), .sp12_in({sp12_v_b[11], sp12_v_b[9]}),
     .lc_trk_out(lc_trk_g1[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g1b, View - schematic
// LAST TIME SAVED: Jul 24 13:24:39 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g1b ( lc_trk_g1, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g1;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [7:0]  tnl_op;
input [1:0]  reset_b;
input [7:0]  bnr_op;
input [7:0]  top_op;
input [7:0]  lft_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g1b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[21], sp4_h_r[13], sp4_h_r[5], sp4_v_b[21],
     sp4_v_b[13], sp4_v_b[5], sp12_h_r[21], sp12_h_r[13], sp12_h_r[5],
     lft_op[5], top_op[5], bot_op[5], bnr_op[5], slf_op[5],
     sp4_r_v_b[29], sp4_r_v_b[5]}), .min2({sp4_h_r[22], sp4_h_r[14],
     sp4_h_r[6], sp4_v_b[22], sp4_v_b[14], sp4_v_b[6], sp12_h_r[22],
     sp12_h_r[14], sp12_h_r[6], lft_op[6], top_op[6], bot_op[6],
     bnr_op[6], slf_op[6], sp4_r_v_b[30], sp4_r_v_b[6]}),
     .min0({sp4_h_r[20], sp4_h_r[12], sp4_h_r[4], sp4_v_b[20],
     sp4_v_b[12], sp4_v_b[4], sp12_h_r[20], sp12_h_r[12], sp12_h_r[4],
     lft_op[4], top_op[4], bot_op[4], bnr_op[4], slf_op[4],
     sp4_r_v_b[28], sp4_r_v_b[4]}), .min3({sp4_h_r[23], sp4_h_r[15],
     sp4_h_r[7], sp4_v_b[23], sp4_v_b[15], sp4_v_b[7], sp12_h_r[23],
     sp12_h_r[15], sp12_h_r[7], lft_op[7], top_op[7], bot_op[7],
     bnr_op[7], slf_op[7], sp4_r_v_b[31], sp4_r_v_b[7]}),
     .sp4_out(sp4_v_b[19:18]), .sp12_in({sp12_v_b[15], sp12_v_b[13]}),
     .lc_trk_out(lc_trk_g1[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2a, View - schematic
// LAST TIME SAVED: Jul 24 13:23:46 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g2a ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g2;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;

input [7:0]  lft_op;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  tnl_op;
input [7:0]  slf_op;
input [1:0]  vdd_cntl;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
input [7:0]  bnr_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[33], sp4_r_v_b[9]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[34], sp4_r_v_b[10]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[32], sp4_r_v_b[8]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[35], sp4_r_v_b[11]}),
     .sp4_out(sp4_v_b[21:20]), .sp12_in({sp12_v_b[19], sp12_v_b[17]}),
     .lc_trk_out(lc_trk_g2[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g2b, View - schematic
// LAST TIME SAVED: Jul 24 13:22:58 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g2b ( lc_trk_g2, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g2;

inout [47:0]  sp4_r_v_b;
inout [23:0]  sp12_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [7:0]  bnr_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  slf_op;
input [7:0]  bnl_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g2b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[37], sp4_r_v_b[13]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[38], sp4_r_v_b[14]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[36], sp4_r_v_b[12]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[39], sp4_r_v_b[15]}),
     .sp4_out(sp4_v_b[23:22]), .sp12_in({sp12_v_b[23], sp12_v_b[21]}),
     .lc_trk_out(lc_trk_g2[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3a, View - schematic
// LAST TIME SAVED: Jul 24 13:22:20 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g3a ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [3:0]  lc_trk_g3;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [47:0]  sp4_h_r;

input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  reset_b;
input [7:0]  top_op;
input [1:0]  vdd_cntl;
input [7:0]  bnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [7:0]  bnl_op;
input [7:0]  tnr_op;
input [7:0]  bot_op;
input [1:0]  wl;
input [7:0]  slf_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3a ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[41], sp4_h_r[33], sp4_h_r[25], sp4_v_b[41],
     sp4_v_b[33], sp4_v_b[25], sp12_v_b[17], sp12_v_b[9], sp12_v_b[1],
     rgt_op[1], tnl_op[1], tnr_op[1], bnl_op[1], slf_op[1],
     sp4_r_v_b[41], sp4_r_v_b[17]}), .min2({sp4_h_r[42], sp4_h_r[34],
     sp4_h_r[26], sp4_v_b[42], sp4_v_b[34], sp4_v_b[26], sp12_v_b[18],
     sp12_v_b[10], sp12_v_b[2], rgt_op[2], tnl_op[2], tnr_op[2],
     bnl_op[2], slf_op[2], sp4_r_v_b[42], sp4_r_v_b[18]}),
     .min0({sp4_h_r[40], sp4_h_r[32], sp4_h_r[24], sp4_v_b[40],
     sp4_v_b[32], sp4_v_b[24], sp12_v_b[16], sp12_v_b[8], sp12_v_b[0],
     rgt_op[0], tnl_op[0], tnr_op[0], bnl_op[0], slf_op[0],
     sp4_r_v_b[40], sp4_r_v_b[16]}), .min3({sp4_h_r[43], sp4_h_r[35],
     sp4_h_r[27], sp4_v_b[43], sp4_v_b[35], sp4_v_b[27], sp12_v_b[19],
     sp12_v_b[11], sp12_v_b[3], rgt_op[3], tnl_op[3], tnr_op[3],
     bnl_op[3], slf_op[3], sp4_r_v_b[43], sp4_r_v_b[19]}),
     .sp4_out(sp4_h_r[13:12]), .sp12_in({sp12_h_r[2], sp12_h_r[0]}),
     .lc_trk_out(lc_trk_g3[3:0]), .pgate(pgate[1:0]));

endmodule
// Library - leafcell, Cell - gmux_sp12to4_g3b, View - schematic
// LAST TIME SAVED: Jul 24 13:21:26 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4_g3b ( lc_trk_g3, bl, sp4_h_r, sp4_r_v_b, sp4_v_b,
     sp12_h_r, sp12_v_b, bnl_op, bnr_op, bot_op, lft_op, pgate, prog,
     reset_b, rgt_op, slf_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:4]  lc_trk_g3;

inout [23:0]  sp12_v_b;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [23:0]  sp12_h_r;
inout [11:0]  bl;

input [7:0]  top_op;
input [7:0]  bnr_op;
input [1:0]  reset_b;
input [7:0]  lft_op;
input [1:0]  pgate;
input [1:0]  wl;
input [7:0]  tnr_op;
input [7:0]  tnl_op;
input [7:0]  rgt_op;
input [1:0]  vdd_cntl;
input [7:0]  bnl_op;
input [7:0]  slf_op;
input [7:0]  bot_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_base Igmux_12to4_g3b ( .vdd_cntl(vdd_cntl[1:0]),
     .wl(wl[1:0]), .bl(bl[11:0]), .prog(prog), .reset_b(reset_b[1:0]),
     .min1({sp4_h_r[45], sp4_h_r[37], sp4_h_r[29], sp4_v_b[45],
     sp4_v_b[37], sp4_v_b[29], sp12_v_b[21], sp12_v_b[13], sp12_v_b[5],
     rgt_op[5], tnl_op[5], tnr_op[5], bnl_op[5], slf_op[5],
     sp4_r_v_b[45], sp4_r_v_b[21]}), .min2({sp4_h_r[46], sp4_h_r[38],
     sp4_h_r[30], sp4_v_b[46], sp4_v_b[38], sp4_v_b[30], sp12_v_b[22],
     sp12_v_b[14], sp12_v_b[6], rgt_op[6], tnl_op[6], tnr_op[6],
     bnl_op[6], slf_op[6], sp4_r_v_b[46], sp4_r_v_b[22]}),
     .min0({sp4_h_r[44], sp4_h_r[36], sp4_h_r[28], sp4_v_b[44],
     sp4_v_b[36], sp4_v_b[28], sp12_v_b[20], sp12_v_b[12], sp12_v_b[4],
     rgt_op[4], tnl_op[4], tnr_op[4], bnl_op[4], slf_op[4],
     sp4_r_v_b[44], sp4_r_v_b[20]}), .min3({sp4_h_r[47], sp4_h_r[39],
     sp4_h_r[31], sp4_v_b[47], sp4_v_b[39], sp4_v_b[31], sp12_v_b[23],
     sp12_v_b[15], sp12_v_b[7], rgt_op[7], tnl_op[7], tnr_op[7],
     bnl_op[7], slf_op[7], sp4_r_v_b[47], sp4_r_v_b[23]}),
     .sp4_out(sp4_h_r[15:14]), .sp12_in({sp12_h_r[6], sp12_h_r[4]}),
     .lc_trk_out(lc_trk_g3[7:4]), .pgate(pgate[1:0]));

endmodule
// Library - xpmem, Cell - ml_rowdrv_bank10k, View - schematic
// LAST TIME SAVED: Oct  6 14:43:11 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module ml_rowdrv_bank10k ( jtag_rowtest_mode_b, last_rsr, pgate, reset,
     vddctrl, wl, banksel, cram_pgateoff, cram_rst, cram_vddoff,
     cram_wl_en, jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst,
     smc_rsr_inc, smc_write, trst_b );
output  jtag_rowtest_mode_b, last_rsr;

input  banksel, cram_pgateoff, cram_rst, cram_vddoff, cram_wl_en,
     jtag_clk, jtag_rowtest_rst, por_rst, rsr_rst, smc_rsr_inc,
     smc_write, trst_b;

output [271:0]  pgate;
output [271:0]  vddctrl;
output [271:0]  reset;
output [271:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:0]  smc_rsr_1st_out_buf;

wire  [16:0]  smc_rsr_out;

wire  [0:16]  smc_rsr_1st_out;

wire  [15:0]  smc_rsr_inc_out;

wire  [15:0]  por_rst_out;



tielo I252 ( .tielo(net0130));
tiehi I269 ( .tiehi(net162));
tiehi I249 ( .tiehi(net131));
tiehi I250 ( .tiehi(net132));
ml_buf_ice5_2 I227 ( .in(net131), .o(net134), .sel(net131));
ml_buf_ice5_2 I216 ( .in(net131), .o(net137), .sel(net131));
ml_buf_ice5_2 I198 ( .sel(banksel), .in(cram_wl_en),
     .o(cram_wl_en_buf));
ml_buf_ice5_2 I196 ( .sel(banksel), .in(cram_rst), .o(cram_rst_buf));
ml_buf_ice5_2 I199 ( .sel(net132), .in(por_rst), .o(por_rst_buf));
ml_buf_ice5_2 I197 ( .sel(banksel), .in(cram_vddoff),
     .o(cram_vddoff_buf));
ml_buf_ice5_2 I195 ( .sel(banksel), .in(cram_pgateoff),
     .o(cram_pgateoff_buf));
ml_buf_ice5_2 I201 ( .sel(banksel), .in(smc_write), .o(smc_write_buf));
ml_buf_ice5_2 I203 ( .sel(net184), .in(net184), .o(smc_rsr_inc_buf));
ml_buf_ice5_2 I213 ( .in(net162), .o(net161), .sel(net162));
ml_rowdrv_tile_last Iml_rowdrv_tile_last (
     .smc_rsr_inc_out(smc_rsr_inc_out_last), .pgate(pgate[271:256]),
     .wl(wl[271:256]), .vddctrl(vddctrl[271:256]),
     .reset(reset[271:256]), .smc_rsr_1st_out(smc_rsr_1st_out[16]),
     .smcc_rsr_out(smc_rsr_out[16]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_buf), .smc_rsr_in(smc_rsr_out[15]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[15]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf));
nand2_hvt I233 ( .A(smc_rsr_inc), .B(banksel), .Y(net181));
mux2_hvt I161 ( .in1(jtag_clk), .in0(net263), .out(net184),
     .sel(net256));
nand3_hvt I231 ( .Y(net186), .B(net190), .C(net190), .A(net190));
nand3_hvt I230 ( .Y(net190), .B(net195), .C(net195), .A(net195));
nand3_hvt I224 ( .B(net131), .Y(net195), .A(net131), .C(net131));
nor3_hvt I238 ( .B(por_rst), .Y(net248), .A(net208), .C(trst));
nor3_hvt I232 ( .C(rsr_rst), .A(jtag_rowtest_rst), .B(net0130),
     .Y(net213));
nor3_hvt I218 ( .B(net225), .Y(net215), .A(net225), .C(net225));
nor3_hvt I220 ( .B(net215), .Y(net219), .A(net215), .C(net215));
nor3_hvt I217 ( .C(net131), .A(net131), .B(net131), .Y(net225));
nor3_hvt I244 ( .B(por_rst), .Y(net227), .A(net276),
     .C(smc_rsr_1st_out_buf[0]));
ml_rowdrv_tile Iml_rowdrv_tile_15_ ( .por_rst_out(por_rst_out[15]),
     .smc_rsr_inc_out(smc_rsr_inc_out[15]),
     .smcc_rsr_out(smc_rsr_out[15]),
     .smc_rsr_1st_out(smc_rsr_1st_out[15]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out_last), .smc_rsr_in(smc_rsr_out[14]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[14]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[255:240]), .vddctrl(vddctrl[255:240]),
     .reset(reset[255:240]), .pgate(pgate[255:240]));
ml_rowdrv_tile Iml_rowdrv_tile_14_ ( .por_rst_out(por_rst_out[14]),
     .smc_rsr_inc_out(smc_rsr_inc_out[14]),
     .smcc_rsr_out(smc_rsr_out[14]),
     .smc_rsr_1st_out(smc_rsr_1st_out[14]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[15]), .smc_rsr_in(smc_rsr_out[13]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[13]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[239:224]), .vddctrl(vddctrl[239:224]),
     .reset(reset[239:224]), .pgate(pgate[239:224]));
ml_rowdrv_tile Iml_rowdrv_tile_13_ ( .por_rst_out(por_rst_out[13]),
     .smc_rsr_inc_out(smc_rsr_inc_out[13]),
     .smcc_rsr_out(smc_rsr_out[13]),
     .smc_rsr_1st_out(smc_rsr_1st_out[13]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[14]), .smc_rsr_in(smc_rsr_out[12]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[12]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[223:208]), .vddctrl(vddctrl[223:208]),
     .reset(reset[223:208]), .pgate(pgate[223:208]));
ml_rowdrv_tile Iml_rowdrv_tile_12_ ( .por_rst_out(por_rst_out[12]),
     .smc_rsr_inc_out(smc_rsr_inc_out[12]),
     .smcc_rsr_out(smc_rsr_out[12]),
     .smc_rsr_1st_out(smc_rsr_1st_out[12]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[13]), .smc_rsr_in(smc_rsr_out[11]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[11]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[207:192]), .vddctrl(vddctrl[207:192]),
     .reset(reset[207:192]), .pgate(pgate[207:192]));
ml_rowdrv_tile Iml_rowdrv_tile_11_ ( .por_rst_out(por_rst_out[11]),
     .smc_rsr_inc_out(smc_rsr_inc_out[11]),
     .smcc_rsr_out(smc_rsr_out[11]),
     .smc_rsr_1st_out(smc_rsr_1st_out[11]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[12]), .smc_rsr_in(smc_rsr_out[10]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[10]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[191:176]), .vddctrl(vddctrl[191:176]),
     .reset(reset[191:176]), .pgate(pgate[191:176]));
ml_rowdrv_tile Iml_rowdrv_tile_10_ ( .por_rst_out(por_rst_out[10]),
     .smc_rsr_inc_out(smc_rsr_inc_out[10]),
     .smcc_rsr_out(smc_rsr_out[10]),
     .smc_rsr_1st_out(smc_rsr_1st_out[10]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[11]), .smc_rsr_in(smc_rsr_out[9]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[9]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[175:160]), .vddctrl(vddctrl[175:160]),
     .reset(reset[175:160]), .pgate(pgate[175:160]));
ml_rowdrv_tile Iml_rowdrv_tile_9_ ( .por_rst_out(por_rst_out[9]),
     .smc_rsr_inc_out(smc_rsr_inc_out[9]),
     .smcc_rsr_out(smc_rsr_out[9]),
     .smc_rsr_1st_out(smc_rsr_1st_out[9]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[10]), .smc_rsr_in(smc_rsr_out[8]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[8]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[159:144]), .vddctrl(vddctrl[159:144]),
     .reset(reset[159:144]), .pgate(pgate[159:144]));
ml_rowdrv_tile Iml_rowdrv_tile_8_ ( .por_rst_out(por_rst_out[8]),
     .smc_rsr_inc_out(smc_rsr_inc_out[8]),
     .smcc_rsr_out(smc_rsr_out[8]),
     .smc_rsr_1st_out(smc_rsr_1st_out[8]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[9]), .smc_rsr_in(smc_rsr_out[7]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[7]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[143:128]), .vddctrl(vddctrl[143:128]),
     .reset(reset[143:128]), .pgate(pgate[143:128]));
ml_rowdrv_tile Iml_rowdrv_tile_7_ ( .por_rst_out(por_rst_out[7]),
     .smc_rsr_inc_out(smc_rsr_inc_out[7]),
     .smcc_rsr_out(smc_rsr_out[7]),
     .smc_rsr_1st_out(smc_rsr_1st_out[7]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[8]), .smc_rsr_in(smc_rsr_out[6]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[6]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[127:112]), .vddctrl(vddctrl[127:112]),
     .reset(reset[127:112]), .pgate(pgate[127:112]));
ml_rowdrv_tile Iml_rowdrv_tile_6_ ( .por_rst_out(por_rst_out[6]),
     .smc_rsr_inc_out(smc_rsr_inc_out[6]),
     .smcc_rsr_out(smc_rsr_out[6]),
     .smc_rsr_1st_out(smc_rsr_1st_out[6]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[7]), .smc_rsr_in(smc_rsr_out[5]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[5]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[111:96]), .vddctrl(vddctrl[111:96]), .reset(reset[111:96]),
     .pgate(pgate[111:96]));
ml_rowdrv_tile Iml_rowdrv_tile_5_ ( .por_rst_out(por_rst_out[5]),
     .smc_rsr_inc_out(smc_rsr_inc_out[5]),
     .smcc_rsr_out(smc_rsr_out[5]),
     .smc_rsr_1st_out(smc_rsr_1st_out[5]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[6]), .smc_rsr_in(smc_rsr_out[4]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[4]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[95:80]), .vddctrl(vddctrl[95:80]), .reset(reset[95:80]),
     .pgate(pgate[95:80]));
ml_rowdrv_tile Iml_rowdrv_tile_4_ ( .por_rst_out(por_rst_out[4]),
     .smc_rsr_inc_out(smc_rsr_inc_out[4]),
     .smcc_rsr_out(smc_rsr_out[4]),
     .smc_rsr_1st_out(smc_rsr_1st_out[4]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[5]), .smc_rsr_in(smc_rsr_out[3]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[3]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[79:64]), .vddctrl(vddctrl[79:64]), .reset(reset[79:64]),
     .pgate(pgate[79:64]));
ml_rowdrv_tile Iml_rowdrv_tile_3_ ( .por_rst_out(por_rst_out[3]),
     .smc_rsr_inc_out(smc_rsr_inc_out[3]),
     .smcc_rsr_out(smc_rsr_out[3]),
     .smc_rsr_1st_out(smc_rsr_1st_out[3]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[4]), .smc_rsr_in(smc_rsr_out[2]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[2]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[63:48]), .vddctrl(vddctrl[63:48]), .reset(reset[63:48]),
     .pgate(pgate[63:48]));
ml_rowdrv_tile Iml_rowdrv_tile_2_ ( .por_rst_out(por_rst_out[2]),
     .smc_rsr_inc_out(smc_rsr_inc_out[2]),
     .smcc_rsr_out(smc_rsr_out[2]),
     .smc_rsr_1st_out(smc_rsr_1st_out[2]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[3]), .smc_rsr_in(smc_rsr_out[1]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[1]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[47:32]), .vddctrl(vddctrl[47:32]), .reset(reset[47:32]),
     .pgate(pgate[47:32]));
ml_rowdrv_tile Iml_rowdrv_tile_1_ ( .por_rst_out(por_rst_out[1]),
     .smc_rsr_inc_out(smc_rsr_inc_out[1]),
     .smcc_rsr_out(smc_rsr_out[1]),
     .smc_rsr_1st_out(smc_rsr_1st_out[1]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[2]), .smc_rsr_in(smc_rsr_out[0]),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_out[0]),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[31:16]), .vddctrl(vddctrl[31:16]), .reset(reset[31:16]),
     .pgate(pgate[31:16]));
ml_rowdrv_tile Iml_rowdrv_tile_0_ ( .por_rst_out(por_rst_out[0]),
     .smc_rsr_inc_out(smc_rsr_inc_out[0]),
     .smcc_rsr_out(smc_rsr_out[0]),
     .smc_rsr_1st_out(smc_rsr_1st_out[0]), .smc_write(smc_write_buf),
     .smc_rsr_inc(smc_rsr_inc_out[1]), .smc_rsr_in(smc_rsr_in_1st),
     .rsr_rst(rst_row_reg), .por_rst(por_rst_buf),
     .cram_wl_en(cram_wl_en_buf), .cram_vddoff(cram_vddoff_buf),
     .cram_rst(cram_rst_buf), .cram_pgateoff(cram_pgateoff_buf),
     .wl(wl[15:0]), .vddctrl(vddctrl[15:0]), .reset(reset[15:0]),
     .pgate(pgate[15:0]));
nor2_hvt I239 ( .A(jtag_rowtest_rst), .B(net248), .Y(net208));
nor2_hvt I193 ( .A(por_rst), .B(rsr_set_1st), .Y(net252));
nor2_hvt I245 ( .A(rsr_set_1st), .B(net227), .Y(net276));
inv_hvt I247 ( .A(net256), .Y(jtag_rowtest_mode_b));
inv_hvt I241 ( .A(net208), .Y(net256));
inv_hvt I192 ( .A(net213), .Y(rsr_set_1st));
inv_hvt I234 ( .A(net181), .Y(net263));
inv_hvt I35 ( .A(net264), .Y(smc_rsr_1st_out_buf[0]));
inv_hvt I240 ( .A(trst_b), .Y(trst));
inv_hvt I210 ( .A(net268), .Y(last_rsr));
inv_hvt I391 ( .A(net252), .Y(rst_row_reg));
inv_hvt I36 ( .A(smc_rsr_1st_out[0]), .Y(net264));
inv_hvt I209 ( .A(smc_rsr_out[16]), .Y(net268));
inv_hvt I205 ( .A(net276), .Y(smc_rsr_in_1st));

endmodule
// Library - leafcell, Cell - gmux_sp12to4, View - schematic
// LAST TIME SAVED: Jul 25 23:13:29 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module gmux_sp12to4 ( lc_trk_g0, lc_trk_g1, lc_trk_g2, lc_trk_g3, bl,
     sp4_h_r, sp4_r_v_b, sp4_v_b, sp12_h_r, sp12_v_b, bnl_op, bnr_op,
     bot_op, glb2local, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g3;

inout [23:0]  sp12_h_r;
inout [47:0]  sp4_h_r;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_r_v_b;
inout [11:0]  bl;
inout [23:0]  sp12_v_b;

input [7:0]  slf_op;
input [7:0]  top_op;
input [7:0]  tnr_op;
input [7:0]  rgt_op;
input [7:0]  bot_op;
input [7:0]  lft_op;
input [7:0]  tnl_op;
input [7:0]  bnr_op;
input [3:0]  glb2local;
input [15:0]  vdd_cntl;
input [15:0]  pgate;
input [15:0]  reset_b;
input [7:0]  bnl_op;
input [15:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



gmux_sp12to4_g0a Ig0_30 ( .vdd_cntl(vdd_cntl[1:0]), .pgate(pgate[1:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp12_v_b(sp12_v_b[23:0]),
     .lc_trk_g0(lc_trk_g0[3:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[1:0]), .reset_b(reset_b[1:0]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g0b Ig0_74 ( .vdd_cntl(vdd_cntl[3:2]), .pgate(pgate[3:2]),
     .glb2local(glb2local[3:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .lc_trk_g0(lc_trk_g0[7:4]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g1a Ig1_30 ( .vdd_cntl(vdd_cntl[5:4]), .pgate(pgate[5:4]),
     .bl(bl[11:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .bot_op(bot_op[7:0]), .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]),
     .lft_op(lft_op[7:0]), .prog(prog), .rgt_op(rgt_op[7:0]),
     .reset_b(reset_b[5:4]), .slf_op(slf_op[7:0]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .wl(wl[5:4]), .lc_trk_g1(lc_trk_g1[3:0]));
gmux_sp12to4_g1b Ig1_74 ( .vdd_cntl(vdd_cntl[7:6]), .pgate(pgate[7:6]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .lc_trk_g1(lc_trk_g1[7:4]),
     .top_op(top_op[7:0]), .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]),
     .wl(wl[7:6]), .reset_b(reset_b[7:6]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g2a Ig2_30 ( .vdd_cntl(vdd_cntl[9:8]), .wl(wl[9:8]),
     .reset_b(reset_b[9:8]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[3:0]), .pgate(pgate[9:8]));
gmux_sp12to4_g2b Ig2_74 ( .vdd_cntl(vdd_cntl[11:10]),
     .pgate(pgate[11:10]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g2(lc_trk_g2[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .wl(wl[11:10]),
     .reset_b(reset_b[11:10]), .prog(prog), .bl(bl[11:0]));
gmux_sp12to4_g3a Ig3_30 ( .vdd_cntl(vdd_cntl[13:12]), .wl(wl[13:12]),
     .reset_b(reset_b[13:12]), .prog(prog), .bl(bl[11:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]),
     .bnl_op(bnl_op[7:0]), .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]),
     .rgt_op(rgt_op[7:0]), .slf_op(slf_op[7:0]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .pgate(pgate[13:12]), .lc_trk_g3(lc_trk_g3[3:0]));
gmux_sp12to4_g3b Ig3_74 ( .vdd_cntl(vdd_cntl[15:14]),
     .pgate(pgate[15:14]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp12_h_r(sp12_h_r[23:0]), .sp12_v_b(sp12_v_b[23:0]),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .lc_trk_g3(lc_trk_g3[7:4]), .top_op(top_op[7:0]),
     .tnl_op(tnl_op[7:0]), .tnr_op(tnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bnr_op(bnr_op[7:0]), .lft_op(lft_op[7:0]), .rgt_op(rgt_op[7:0]),
     .slf_op(slf_op[7:0]), .bot_op(bot_op[7:0]), .prog(prog),
     .bl(bl[11:0]), .reset_b(reset_b[15:14]), .wl(wl[15:14]));

endmodule
// Library - leafcell, Cell - ltile4rev0, View - schematic
// LAST TIME SAVED: Jun  2 13:31:12 2008
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module ltile4rev0 ( carry_out, slf_op, bl, sp4_h_l, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp4_v_t, sp12_h_l, sp12_h_r, sp12_v_b, sp12_v_t, bnl_op,
     bnr_op, bot_op, carry_in, glb_netwk, lft_op, pgate, prog, purst,
     reset_b, rgt_op, tnl_op, tnr_op, top_op, vdd_cntl, wl );
output  carry_out;


input  carry_in, prog, purst;

output [7:0]  slf_op;

inout [23:0]  sp12_v_t;
inout [47:0]  sp4_h_l;
inout [23:0]  sp12_h_l;
inout [23:0]  sp12_v_b;
inout [47:0]  sp4_v_t;
inout [53:0]  bl;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_h_r;
inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;

input [15:0]  pgate;
input [7:0]  tnl_op;
input [7:0]  bot_op;
input [7:0]  top_op;
input [7:0]  glb_netwk;
input [7:0]  lft_op;
input [15:0]  reset_b;
input [7:0]  rgt_op;
input [7:0]  tnr_op;
input [15:0]  vdd_cntl;
input [7:0]  bnr_op;
input [15:0]  wl;
input [7:0]  bnl_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net_glb2local;

wire  [7:0]  lc_trk_g3;

wire  [1:0]  sp12_h_r_mid;

wire  [7:0]  lc_trk_g2;

wire  [1:0]  sp12_v_b_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



misc_module4rev0 Ickmux_sp12to4_sp12sw ( .vdd_cntl({vdd_cntl[14],
     vdd_cntl[15], vdd_cntl[12], vdd_cntl[13], vdd_cntl[10],
     vdd_cntl[11], vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7],
     vdd_cntl[4], vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0],
     vdd_cntl[1]}), .glb_netwk(glb_netwk[7:0]), .l(sp12_h_r_mid[1:0]),
     .m(sp12_v_b_mid[1:0]), .r(sp12_h_r[1:0]), .b(sp12_v_b[1:0]),
     .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18], sp12_h_r[16],
     sp12_h_r[14], sp12_h_r[12], sp12_h_r[10], sp12_h_r[8]}),
     .sp4(sp4_h_r[23:16]), .min3(glb_netwk[7:0]),
     .min0(glb_netwk[7:0]), .min1(glb_netwk[7:0]),
     .min2(glb_netwk[7:0]), .prog(progd), .lc_trk_g0(lc_trk_g0[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .lc_trk_g1(lc_trk_g1[5:0]), .wl({wl[14], wl[15], wl[12], wl[13],
     wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2],
     wl[3], wl[0], wl[1]}), .S_R(s_r), .clkb(clkb), .bl(bl[3:0]),
     .clk(clk), .reset_b({reset_b[14], reset_b[15], reset_b[12],
     reset_b[13], reset_b[10], reset_b[11], reset_b[8], reset_b[9],
     reset_b[6], reset_b[7], reset_b[4], reset_b[5], reset_b[2],
     reset_b[3], reset_b[0], reset_b[1]}), .pgate({pgate[14],
     pgate[15], pgate[12], pgate[13], pgate[10], pgate[11], pgate[8],
     pgate[9], pgate[6], pgate[7], pgate[4], pgate[5], pgate[2],
     pgate[3], pgate[0], pgate[1]}), .glb2local(net_glb2local[3:0]));
lccol_rev0 I_lcx8 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .s_r(s_r), .reset_b({reset_b[14], reset_b[15], reset_b[12],
     reset_b[13], reset_b[10], reset_b[11], reset_b[8], reset_b[9],
     reset_b[6], reset_b[7], reset_b[4], reset_b[5], reset_b[2],
     reset_b[3], reset_b[0], reset_b[1]}), .purst(purst), .prog(progd),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .lc_trk_g3(lc_trk_g3[7:0]), .lc_trk_g2(lc_trk_g2[7:0]),
     .lc_trk_g1(lc_trk_g1[7:0]), .lc_trk_g0(lc_trk_g0[7:0]),
     .clkb(clkb), .clk(clk), .cin2local(carry_in),
     .slf_op(slf_op[7:0]), .carry_out(carry_out),
     .sp12_v_b(sp12_v_b[23:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_r_v_b(sp4_r_v_b[47:0]),
     .sp4_h_r(sp4_h_r[47:0]), .bl(bl[53:26]));
rm6  R3_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm6  R3_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm6  R3_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm6  R3_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm6  R3_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm6  R3_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm6  R3_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm6  R3_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm6  R3_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm6  R3_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm6  R3_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm6  R3_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm6  R3_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm6  R3_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm6  R3_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm6  R3_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm6  R3_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm6  R3_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm6  R3_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm6  R3_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm6  R3_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm6  R3_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm6  R3_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm6  R3_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
rm7  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
span4 Isp4_sw ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15], vdd_cntl[12],
     vdd_cntl[13], vdd_cntl[10], vdd_cntl[11], vdd_cntl[8],
     vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4], vdd_cntl[5],
     vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .sp4_h_r(sp4_h_r[47:0]), .sp4_v_b(sp4_v_b[47:0]),
     .sp4_h_l(sp4_h_l[47:0]), .sp4_v_t(sp4_v_t[47:0]),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(progd), .wl({wl[14], wl[15], wl[12], wl[13],
     wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5], wl[2],
     wl[3], wl[0], wl[1]}), .bl(bl[13:4]));
gmux_sp12to4 Igmux_sp12to4 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .reset_b({reset_b[14], reset_b[15], reset_b[12], reset_b[13],
     reset_b[10], reset_b[11], reset_b[8], reset_b[9], reset_b[6],
     reset_b[7], reset_b[4], reset_b[5], reset_b[2], reset_b[3],
     reset_b[0], reset_b[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .glb2local(net_glb2local[3:0]),
     .sp12_v_b(sp12_v_b[23:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_r(sp4_h_r[47:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g3(lc_trk_g3[7:0]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .bot_op(bot_op[7:0]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .prog(progd),
     .lft_op(lft_op[7:0]), .bnr_op(bnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .bl(bl[25:14]));
inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(progd));

endmodule
// Library - leafcell, Cell - array_LT1x16, View - schematic
// LAST TIME SAVED: Jun 12 09:45:55 2008
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module array_LT1x16 ( carry_out, glb_netwk, slf_op_01, slf_op_02,
     slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07, slf_op_08,
     slf_op_09, slf_op_10, slf_op_11, slf_op_12, slf_op_13, slf_op_14,
     slf_op_15, slf_op_16, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02,
     sp4_h_l_03, sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07,
     sp4_h_l_08, sp4_h_l_09, sp4_h_l_10, sp4_h_l_11, sp4_h_l_12,
     sp4_h_l_13, sp4_h_l_14, sp4_h_l_15, sp4_h_l_16, sp4_h_r_01,
     sp4_h_r_02, sp4_h_r_03, sp4_h_r_04, sp4_h_r_05, sp4_h_r_06,
     sp4_h_r_07, sp4_h_r_08, sp4_h_r_09, sp4_h_r_10, sp4_h_r_11,
     sp4_h_r_12, sp4_h_r_13, sp4_h_r_14, sp4_h_r_15, sp4_h_r_16,
     sp4_r_v_b_01, sp4_r_v_b_02, sp4_r_v_b_03, sp4_r_v_b_04,
     sp4_r_v_b_05, sp4_r_v_b_06, sp4_r_v_b_07, sp4_r_v_b_08,
     sp4_r_v_b_09, sp4_r_v_b_10, sp4_r_v_b_11, sp4_r_v_b_12,
     sp4_r_v_b_13, sp4_r_v_b_14, sp4_r_v_b_15, sp4_r_v_b_16,
     sp4_v_b_01, sp4_v_b_02, sp4_v_b_03, sp4_v_b_04, sp4_v_b_05,
     sp4_v_b_06, sp4_v_b_07, sp4_v_b_08, sp4_v_b_09, sp4_v_b_10,
     sp4_v_b_11, sp4_v_b_12, sp4_v_b_13, sp4_v_b_14, sp4_v_b_15,
     sp4_v_b_16, sp4_v_t_16, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03,
     sp12_h_l_04, sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08,
     sp12_h_l_09, sp12_h_l_10, sp12_h_l_11, sp12_h_l_12, sp12_h_l_13,
     sp12_h_l_14, sp12_h_l_15, sp12_h_l_16, sp12_h_r_01, sp12_h_r_02,
     sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06, sp12_h_r_07,
     sp12_h_r_08, sp12_h_r_09, sp12_h_r_10, sp12_h_r_11, sp12_h_r_12,
     sp12_h_r_13, sp12_h_r_14, sp12_h_r_15, sp12_h_r_16, sp12_v_b_01,
     sp12_v_t_16, vdd_cntl, wl, bnl_op_01, bnr_op_01, bot_op_01,
     carry_in, glb_netwk_col, lft_op_01, lft_op_02, lft_op_03,
     lft_op_04, lft_op_05, lft_op_06, lft_op_07, lft_op_08, lft_op_09,
     lft_op_10, lft_op_11, lft_op_12, lft_op_13, lft_op_14, lft_op_15,
     lft_op_16, prog, purst, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, rgt_op_09,
     rgt_op_10, rgt_op_11, rgt_op_12, rgt_op_13, rgt_op_14, rgt_op_15,
     rgt_op_16, tnl_op_16, tnr_op_16, top_op_16 );
output  carry_out;


input  carry_in, prog, purst;

output [7:0]  slf_op_01;
output [7:0]  slf_op_10;
output [7:0]  slf_op_08;
output [7:0]  slf_op_16;
output [7:0]  slf_op_02;
output [7:0]  slf_op_12;
output [7:0]  glb_netwk;
output [7:0]  slf_op_06;
output [7:0]  slf_op_03;
output [7:0]  slf_op_11;
output [7:0]  slf_op_09;
output [7:0]  slf_op_13;
output [7:0]  slf_op_15;
output [7:0]  slf_op_04;
output [7:0]  slf_op_05;
output [7:0]  slf_op_14;
output [7:0]  slf_op_07;

inout [47:0]  sp4_v_b_03;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_h_r_09;
inout [47:0]  sp4_h_r_16;
inout [23:0]  sp12_h_l_04;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_v_b_05;
inout [47:0]  sp4_v_b_16;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_r_v_b_12;
inout [23:0]  sp12_h_r_13;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_v_b_15;
inout [47:0]  sp4_r_v_b_05;
inout [47:0]  sp4_v_b_13;
inout [23:0]  sp12_h_r_15;
inout [47:0]  sp4_h_l_10;
inout [47:0]  sp4_h_l_16;
inout [47:0]  sp4_h_r_13;
inout [47:0]  sp4_v_b_09;
inout [23:0]  sp12_h_r_11;
inout [47:0]  sp4_v_b_14;
inout [47:0]  sp4_h_r_11;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_h_r_08;
inout [23:0]  sp12_h_l_11;
inout [23:0]  sp12_h_r_14;
inout [23:0]  sp12_h_l_12;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_r_v_b_03;
inout [23:0]  sp12_h_l_05;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_r_v_b_14;
inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_h_l_13;
inout [47:0]  sp4_h_l_11;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_h_l_06;
inout [255:0]  wl;
inout [255:0]  reset_b;
inout [47:0]  sp4_h_l_14;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_v_t_16;
inout [47:0]  sp4_h_l_13;
inout [23:0]  sp12_h_l_16;
inout [23:0]  sp12_h_r_08;
inout [47:0]  sp4_h_r_01;
inout [23:0]  sp12_h_l_09;
inout [23:0]  sp12_h_r_10;
inout [47:0]  sp4_h_r_05;
inout [23:0]  sp12_h_r_01;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_h_r_12;
inout [23:0]  sp12_h_r_12;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_v_b_10;
inout [23:0]  sp12_h_r_16;
inout [47:0]  sp4_h_r_02;
inout [23:0]  sp12_h_l_08;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_h_l_01;
inout [255:0]  vdd_cntl;
inout [23:0]  sp12_v_t_16;
inout [47:0]  sp4_r_v_b_16;
inout [47:0]  sp4_h_r_04;
inout [23:0]  sp12_h_l_10;
inout [47:0]  sp4_h_l_15;
inout [47:0]  sp4_v_b_06;
inout [47:0]  sp4_v_b_01;
inout [23:0]  sp12_h_l_15;
inout [23:0]  sp12_h_r_03;
inout [23:0]  sp12_h_r_09;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_h_l_09;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_v_b_12;
inout [47:0]  sp4_r_v_b_10;
inout [23:0]  sp12_h_r_07;
inout [255:0]  pgate;
inout [23:0]  sp12_h_r_04;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_r_v_b_13;
inout [47:0]  sp4_h_l_12;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_r_v_b_15;
inout [47:0]  sp4_r_v_b_09;
inout [53:0]  bl;
inout [47:0]  sp4_h_r_10;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_h_r_15;
inout [47:0]  sp4_v_b_11;
inout [23:0]  sp12_v_b_01;
inout [47:0]  sp4_h_l_03;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_r_v_b_11;
inout [47:0]  sp4_h_r_14;
inout [23:0]  sp12_h_l_14;
inout [47:0]  sp4_h_l_04;

input [7:0]  lft_op_11;
input [7:0]  rgt_op_15;
input [7:0]  rgt_op_02;
input [7:0]  lft_op_03;
input [7:0]  glb_netwk_col;
input [7:0]  lft_op_08;
input [7:0]  lft_op_04;
input [7:0]  rgt_op_06;
input [7:0]  tnr_op_16;
input [7:0]  lft_op_06;
input [7:0]  lft_op_15;
input [7:0]  rgt_op_10;
input [7:0]  tnl_op_16;
input [7:0]  rgt_op_12;
input [7:0]  bnl_op_01;
input [7:0]  bot_op_01;
input [7:0]  lft_op_05;
input [7:0]  bnr_op_01;
input [7:0]  lft_op_16;
input [7:0]  rgt_op_04;
input [7:0]  rgt_op_14;
input [7:0]  rgt_op_16;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_09;
input [7:0]  rgt_op_13;
input [7:0]  lft_op_07;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_10;
input [7:0]  lft_op_12;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_11;
input [7:0]  lft_op_02;
input [7:0]  lft_op_09;
input [7:0]  lft_op_14;
input [7:0]  top_op_16;
input [7:0]  lft_op_13;
input [7:0]  rgt_op_08;
input [7:0]  lft_op_01;
input [7:0]  rgt_op_01;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:23]  net840;

wire  [0:23]  net644;

wire  [0:23]  net896;

wire  [0:23]  net756;

wire  [0:23]  net700;

wire  [0:23]  net980;

wire  [0:23]  net672;

wire  [0:23]  net1036;

wire  [0:23]  net1008;

wire  [0:23]  net924;

wire  [0:23]  net812;

wire  [0:23]  net728;

wire  [0:23]  net616;

wire  [0:23]  net868;

wire  [0:23]  net952;



ltile4rev0 I_LT06 ( .prog(prog), .carry_out(net608),
     .lft_op(lft_op_06[7:0]), .sp12_h_l(sp12_h_l_06[23:0]),
     .sp4_h_l(sp4_h_l_06[47:0]), .sp4_v_b(sp4_v_b_06[47:0]),
     .sp12_v_b(net700[0:23]), .sp12_h_r(sp12_h_r_06[23:0]),
     .sp4_h_r(sp4_h_r_06[47:0]), .sp12_v_t(net616[0:23]),
     .sp4_v_t(sp4_v_b_07[47:0]), .sp4_r_v_b(sp4_r_v_b_06[47:0]),
     .wl(wl[95:80]), .top_op(slf_op_07[7:0]), .rgt_op(rgt_op_06[7:0]),
     .bot_op(slf_op_05[7:0]), .bl(bl[53:0]), .reset_b(reset_b[95:80]),
     .vdd_cntl(vdd_cntl[95:80]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net692), .purst(purst), .slf_op(slf_op_06[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_05[7:0]),
     .bnl_op(lft_op_05[7:0]), .tnr_op(rgt_op_07[7:0]),
     .tnl_op(lft_op_07[7:0]));
ltile4rev0 I_LT03 ( .prog(prog), .carry_out(net636),
     .lft_op(lft_op_03[7:0]), .sp12_h_l(sp12_h_l_03[23:0]),
     .sp4_h_l(sp4_h_l_03[47:0]), .sp4_v_b(sp4_v_b_03[47:0]),
     .sp12_v_b(net924[0:23]), .sp12_h_r(sp12_h_r_03[23:0]),
     .sp4_h_r(sp4_h_r_03[47:0]), .sp12_v_t(net644[0:23]),
     .sp4_v_t(sp4_v_b_04[47:0]), .sp4_r_v_b(sp4_r_v_b_03[47:0]),
     .wl(wl[47:32]), .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net916), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4rev0 I_LT04 ( .prog(prog), .carry_out(net664),
     .lft_op(lft_op_04[7:0]), .sp12_h_l(sp12_h_l_04[23:0]),
     .sp4_h_l(sp4_h_l_04[47:0]), .sp4_v_b(sp4_v_b_04[47:0]),
     .sp12_v_b(net644[0:23]), .sp12_h_r(sp12_h_r_04[23:0]),
     .sp4_h_r(sp4_h_r_04[47:0]), .sp12_v_t(net672[0:23]),
     .sp4_v_t(sp4_v_b_05[47:0]), .sp4_r_v_b(sp4_r_v_b_04[47:0]),
     .wl(wl[63:48]), .top_op(slf_op_05[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net636), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(rgt_op_05[7:0]),
     .tnl_op(lft_op_05[7:0]));
ltile4rev0 I_LT05 ( .prog(prog), .carry_out(net692),
     .lft_op(lft_op_05[7:0]), .sp12_h_l(sp12_h_l_05[23:0]),
     .sp4_h_l(sp4_h_l_05[47:0]), .sp4_v_b(sp4_v_b_05[47:0]),
     .sp12_v_b(net672[0:23]), .sp12_h_r(sp12_h_r_05[23:0]),
     .sp4_h_r(sp4_h_r_05[47:0]), .sp12_v_t(net700[0:23]),
     .sp4_v_t(sp4_v_b_06[47:0]), .sp4_r_v_b(sp4_r_v_b_05[47:0]),
     .wl(wl[79:64]), .top_op(slf_op_06[7:0]), .rgt_op(rgt_op_05[7:0]),
     .bot_op(slf_op_04[7:0]), .bl(bl[53:0]), .reset_b(reset_b[79:64]),
     .vdd_cntl(vdd_cntl[79:64]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net664), .purst(purst), .slf_op(slf_op_05[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_04[7:0]),
     .bnl_op(lft_op_04[7:0]), .tnr_op(rgt_op_06[7:0]),
     .tnl_op(lft_op_06[7:0]));
ltile4rev0 I_LT12 ( .prog(prog), .carry_out(net720),
     .lft_op(lft_op_12[7:0]), .sp12_h_l(sp12_h_l_12[23:0]),
     .sp4_h_l(sp4_h_l_12[47:0]), .sp4_v_b(sp4_v_b_12[47:0]),
     .sp12_v_b(net756[0:23]), .sp12_h_r(sp12_h_r_12[23:0]),
     .sp4_h_r(sp4_h_r_12[47:0]), .sp12_v_t(net728[0:23]),
     .sp4_v_t(sp4_v_b_13[47:0]), .sp4_r_v_b(sp4_r_v_b_12[47:0]),
     .wl(wl[191:176]), .top_op(slf_op_13[7:0]),
     .rgt_op(rgt_op_12[7:0]), .bot_op(slf_op_11[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[191:176]), .vdd_cntl(vdd_cntl[191:176]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net748), .purst(purst),
     .slf_op(slf_op_12[7:0]), .pgate(pgate[191:176]),
     .bnr_op(rgt_op_11[7:0]), .bnl_op(lft_op_11[7:0]),
     .tnr_op(rgt_op_13[7:0]), .tnl_op(lft_op_13[7:0]));
ltile4rev0 I_LT11 ( .prog(prog), .carry_out(net748),
     .lft_op(lft_op_11[7:0]), .sp12_h_l(sp12_h_l_11[23:0]),
     .sp4_h_l(sp4_h_l_11[47:0]), .sp4_v_b(sp4_v_b_11[47:0]),
     .sp12_v_b(net952[0:23]), .sp12_h_r(sp12_h_r_11[23:0]),
     .sp4_h_r(sp4_h_r_11[47:0]), .sp12_v_t(net756[0:23]),
     .sp4_v_t(sp4_v_b_12[47:0]), .sp4_r_v_b(sp4_r_v_b_11[47:0]),
     .wl(wl[175:160]), .top_op(slf_op_12[7:0]),
     .rgt_op(rgt_op_11[7:0]), .bot_op(slf_op_10[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[175:160]), .vdd_cntl(vdd_cntl[175:160]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net944), .purst(purst),
     .slf_op(slf_op_11[7:0]), .pgate(pgate[175:160]),
     .bnr_op(rgt_op_10[7:0]), .bnl_op(lft_op_10[7:0]),
     .tnr_op(rgt_op_12[7:0]), .tnl_op(lft_op_12[7:0]));
ltile4rev0 I_LT16 ( .prog(prog), .carry_out(carry_out),
     .lft_op(lft_op_16[7:0]), .sp12_h_l(sp12_h_l_16[23:0]),
     .sp4_h_l(sp4_h_l_16[47:0]), .sp4_v_b(sp4_v_b_16[47:0]),
     .sp12_v_b(net868[0:23]), .sp12_h_r(sp12_h_r_16[23:0]),
     .sp4_h_r(sp4_h_r_16[47:0]), .sp12_v_t(sp12_v_t_16[23:0]),
     .sp4_v_t(sp4_v_t_16[47:0]), .sp4_r_v_b(sp4_r_v_b_16[47:0]),
     .wl(wl[255:240]), .top_op(top_op_16[7:0]),
     .rgt_op(rgt_op_16[7:0]), .bot_op(slf_op_15[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[255:240]), .vdd_cntl(vdd_cntl[255:240]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net860), .purst(purst),
     .slf_op(slf_op_16[7:0]), .pgate(pgate[255:240]),
     .bnr_op(rgt_op_15[7:0]), .bnl_op(lft_op_15[7:0]),
     .tnr_op(tnr_op_16[7:0]), .tnl_op(tnl_op_16[7:0]));
ltile4rev0 I_LT14 ( .prog(prog), .carry_out(net804),
     .lft_op(lft_op_14[7:0]), .sp12_h_l(sp12_h_l_14[23:0]),
     .sp4_h_l(sp4_h_l_14[47:0]), .sp4_v_b(sp4_v_b_14[47:0]),
     .sp12_v_b(net840[0:23]), .sp12_h_r(sp12_h_r_14[23:0]),
     .sp4_h_r(sp4_h_r_14[47:0]), .sp12_v_t(net812[0:23]),
     .sp4_v_t(sp4_v_b_15[47:0]), .sp4_r_v_b(sp4_r_v_b_14[47:0]),
     .wl(wl[223:208]), .top_op(slf_op_15[7:0]),
     .rgt_op(rgt_op_14[7:0]), .bot_op(slf_op_13[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[223:208]), .vdd_cntl(vdd_cntl[223:208]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net832), .purst(purst),
     .slf_op(slf_op_14[7:0]), .pgate(pgate[223:208]),
     .bnr_op(rgt_op_13[7:0]), .bnl_op(lft_op_13[7:0]),
     .tnr_op(rgt_op_15[7:0]), .tnl_op(lft_op_15[7:0]));
ltile4rev0 I_LT13 ( .prog(prog), .carry_out(net832),
     .lft_op(lft_op_13[7:0]), .sp12_h_l(sp12_h_l_13[23:0]),
     .sp4_h_l(sp4_h_l_13[47:0]), .sp4_v_b(sp4_v_b_13[47:0]),
     .sp12_v_b(net728[0:23]), .sp12_h_r(sp12_h_r_13[23:0]),
     .sp4_h_r(sp4_h_r_13[47:0]), .sp12_v_t(net840[0:23]),
     .sp4_v_t(sp4_v_b_14[47:0]), .sp4_r_v_b(sp4_r_v_b_13[47:0]),
     .wl(wl[207:192]), .top_op(slf_op_14[7:0]),
     .rgt_op(rgt_op_13[7:0]), .bot_op(slf_op_12[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[207:192]), .vdd_cntl(vdd_cntl[207:192]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net720), .purst(purst),
     .slf_op(slf_op_13[7:0]), .pgate(pgate[207:192]),
     .bnr_op(rgt_op_12[7:0]), .bnl_op(lft_op_12[7:0]),
     .tnr_op(rgt_op_14[7:0]), .tnl_op(lft_op_14[7:0]));
ltile4rev0 I_LT15 ( .prog(prog), .carry_out(net860),
     .lft_op(lft_op_15[7:0]), .sp12_h_l(sp12_h_l_15[23:0]),
     .sp4_h_l(sp4_h_l_15[47:0]), .sp4_v_b(sp4_v_b_15[47:0]),
     .sp12_v_b(net812[0:23]), .sp12_h_r(sp12_h_r_15[23:0]),
     .sp4_h_r(sp4_h_r_15[47:0]), .sp12_v_t(net868[0:23]),
     .sp4_v_t(sp4_v_b_16[47:0]), .sp4_r_v_b(sp4_r_v_b_15[47:0]),
     .wl(wl[239:224]), .top_op(slf_op_16[7:0]),
     .rgt_op(rgt_op_15[7:0]), .bot_op(slf_op_14[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[239:224]), .vdd_cntl(vdd_cntl[239:224]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net804), .purst(purst),
     .slf_op(slf_op_15[7:0]), .pgate(pgate[239:224]),
     .bnr_op(rgt_op_14[7:0]), .bnl_op(lft_op_14[7:0]),
     .tnr_op(rgt_op_16[7:0]), .tnl_op(lft_op_16[7:0]));
ltile4rev0 I_LT01 ( .prog(prog), .carry_out(net888),
     .lft_op(lft_op_01[7:0]), .sp12_h_l(sp12_h_l_01[23:0]),
     .sp4_h_l(sp4_h_l_01[47:0]), .sp4_v_b(sp4_v_b_01[47:0]),
     .sp12_v_b(sp12_v_b_01[23:0]), .sp12_h_r(sp12_h_r_01[23:0]),
     .sp4_h_r(sp4_h_r_01[47:0]), .sp12_v_t(net896[0:23]),
     .sp4_v_t(sp4_v_b_02[47:0]), .sp4_r_v_b(sp4_r_v_b_01[47:0]),
     .wl(wl[15:0]), .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4rev0 I_LT02 ( .prog(prog), .carry_out(net916),
     .lft_op(lft_op_02[7:0]), .sp12_h_l(sp12_h_l_02[23:0]),
     .sp4_h_l(sp4_h_l_02[47:0]), .sp4_v_b(sp4_v_b_02[47:0]),
     .sp12_v_b(net896[0:23]), .sp12_h_r(sp12_h_r_02[23:0]),
     .sp4_h_r(sp4_h_r_02[47:0]), .sp12_v_t(net924[0:23]),
     .sp4_v_t(sp4_v_b_03[47:0]), .sp4_r_v_b(sp4_r_v_b_02[47:0]),
     .wl(wl[31:16]), .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net888), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));
ltile4rev0 I_LT10 ( .prog(prog), .carry_out(net944),
     .lft_op(lft_op_10[7:0]), .sp12_h_l(sp12_h_l_10[23:0]),
     .sp4_h_l(sp4_h_l_10[47:0]), .sp4_v_b(sp4_v_b_10[47:0]),
     .sp12_v_b(net1036[0:23]), .sp12_h_r(sp12_h_r_10[23:0]),
     .sp4_h_r(sp4_h_r_10[47:0]), .sp12_v_t(net952[0:23]),
     .sp4_v_t(sp4_v_b_11[47:0]), .sp4_r_v_b(sp4_r_v_b_10[47:0]),
     .wl(wl[159:144]), .top_op(slf_op_11[7:0]),
     .rgt_op(rgt_op_10[7:0]), .bot_op(slf_op_09[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[159:144]), .vdd_cntl(vdd_cntl[159:144]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net1028), .purst(purst),
     .slf_op(slf_op_10[7:0]), .pgate(pgate[159:144]),
     .bnr_op(rgt_op_09[7:0]), .bnl_op(lft_op_09[7:0]),
     .tnr_op(rgt_op_11[7:0]), .tnl_op(lft_op_11[7:0]));
ltile4rev0 I_LT08 ( .prog(prog), .carry_out(net972),
     .lft_op(lft_op_08[7:0]), .sp12_h_l(sp12_h_l_08[23:0]),
     .sp4_h_l(sp4_h_l_08[47:0]), .sp4_v_b(sp4_v_b_08[47:0]),
     .sp12_v_b(net1008[0:23]), .sp12_h_r(sp12_h_r_08[23:0]),
     .sp4_h_r(sp4_h_r_08[47:0]), .sp12_v_t(net980[0:23]),
     .sp4_v_t(sp4_v_b_09[47:0]), .sp4_r_v_b(sp4_r_v_b_08[47:0]),
     .wl(wl[127:112]), .top_op(slf_op_09[7:0]),
     .rgt_op(rgt_op_08[7:0]), .bot_op(slf_op_07[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[127:112]), .vdd_cntl(vdd_cntl[127:112]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net1000), .purst(purst),
     .slf_op(slf_op_08[7:0]), .pgate(pgate[127:112]),
     .bnr_op(rgt_op_07[7:0]), .bnl_op(lft_op_07[7:0]),
     .tnr_op(rgt_op_09[7:0]), .tnl_op(lft_op_09[7:0]));
ltile4rev0 I_LT07 ( .prog(prog), .carry_out(net1000),
     .lft_op(lft_op_07[7:0]), .sp12_h_l(sp12_h_l_07[23:0]),
     .sp4_h_l(sp4_h_l_07[47:0]), .sp4_v_b(sp4_v_b_07[47:0]),
     .sp12_v_b(net616[0:23]), .sp12_h_r(sp12_h_r_07[23:0]),
     .sp4_h_r(sp4_h_r_07[47:0]), .sp12_v_t(net1008[0:23]),
     .sp4_v_t(sp4_v_b_08[47:0]), .sp4_r_v_b(sp4_r_v_b_07[47:0]),
     .wl(wl[111:96]), .top_op(slf_op_08[7:0]), .rgt_op(rgt_op_07[7:0]),
     .bot_op(slf_op_06[7:0]), .bl(bl[53:0]), .reset_b(reset_b[111:96]),
     .vdd_cntl(vdd_cntl[111:96]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net608), .purst(purst), .slf_op(slf_op_07[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_06[7:0]),
     .bnl_op(lft_op_06[7:0]), .tnr_op(rgt_op_08[7:0]),
     .tnl_op(lft_op_08[7:0]));
ltile4rev0 I_LT09 ( .prog(prog), .carry_out(net1028),
     .lft_op(lft_op_09[7:0]), .sp12_h_l(sp12_h_l_09[23:0]),
     .sp4_h_l(sp4_h_l_09[47:0]), .sp4_v_b(sp4_v_b_09[47:0]),
     .sp12_v_b(net980[0:23]), .sp12_h_r(sp12_h_r_09[23:0]),
     .sp4_h_r(sp4_h_r_09[47:0]), .sp12_v_t(net1036[0:23]),
     .sp4_v_t(sp4_v_b_10[47:0]), .sp4_r_v_b(sp4_r_v_b_09[47:0]),
     .wl(wl[143:128]), .top_op(slf_op_10[7:0]),
     .rgt_op(rgt_op_09[7:0]), .bot_op(slf_op_08[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[143:128]), .vdd_cntl(vdd_cntl[143:128]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net972), .purst(purst),
     .slf_op(slf_op_09[7:0]), .pgate(pgate[143:128]),
     .bnr_op(rgt_op_08[7:0]), .bnl_op(lft_op_08[7:0]),
     .tnr_op(rgt_op_10[7:0]), .tnl_op(lft_op_10[7:0]));
clk_colbuf8kx8 I78 ( .clko(glb_netwk[7:0]), .clki(glb_netwk_col[7:0]));

endmodule
// Library - leafcell, Cell - clkmandcmuxrev, View - schematic
// LAST TIME SAVED: Jul 24 09:36:22 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module clkmandcmuxrev ( cin2lcl, clk, clkb, glb2local, s_r, carry_in,
     cbit, cbitb, glb_netwk, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, min0, min1, min2, min3, prog );
output  cin2lcl, clk, clkb, s_r;

input  carry_in, prog;

output [3:0]  glb2local;

input [7:0]  min0;
input [7:0]  min3;
input [7:0]  glb_netwk;
input [31:0]  cbit;
input [31:0]  cbitb;
input [5:0]  lc_trk_g1;
input [5:0]  lc_trk_g0;
input [7:0]  min2;
input [7:0]  min1;
input [5:0]  lc_trk_g2;
input [5:0]  lc_trk_g3;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



sr_clkm8to1 I296 ( .mout(s_r), .cbitb(cbitb[12:9]), .min({lc_trk_g3[5],
     lc_trk_g2[4], lc_trk_g1[5], lc_trk_g0[4], glb_netwk[6],
     glb_netwk[4], glb_netwk[2], glb_netwk[0]}), .cbit(cbit[12:9]),
     .prog(prog));
ce_clkm8to1 I283 ( .moutb(ceb), .cbitb(cbitb[8:5]), .cbit(cbit[8:5]),
     .prog(prog), .min({lc_trk_g3[3], lc_trk_g2[2], lc_trk_g1[3],
     lc_trk_g0[2], glb_netwk[7], glb_netwk[5], glb_netwk[3],
     glb_netwk[1]}));
clk_mux12to1 I298 ( .cbitb({cbitb[31], cbitb[4], cbitb[3], cbitb[2],
     cbitb[1], cbitb[0]}), .cbit({cbit[31], cbit[4], cbit[3], cbit[2],
     cbit[1], cbit[0]}), .prog(prog), .min({lc_trk_g3[1], lc_trk_g2[0],
     lc_trk_g1[1], lc_trk_g0[0], glb_netwk[7:0]}), .clk(clk),
     .clkb(clkb), .cenb(ceb));
clk_mux8to1 I285 ( .min(min3[7:0]), .prog(prog), .inmuxo(glb2local[0]),
     .cbit(cbit[16:13]), .cbitb(cbitb[16:13]));
clk_mux8to1 I293 ( .prog(prog), .inmuxo(glb2local[1]), .min(min2[7:0]),
     .cbit(cbit[20:17]), .cbitb(cbitb[20:17]));
clk_mux8to1 I294 ( .prog(prog), .inmuxo(glb2local[2]), .min(min1[7:0]),
     .cbit(cbit[24:21]), .cbitb(cbitb[24:21]));
clk_mux8to1 I295 ( .prog(prog), .inmuxo(glb2local[3]), .min(min0[7:0]),
     .cbit(cbit[28:25]), .cbitb(cbitb[28:25]));
mux_4carry Icarry_cnt ( .cin(carry_in), .lcl_cin(cin2lcl),
     .cbitb(cbitb[30:29]), .prog(prog), .cbit(cbit[30:29]));

endmodule
// Library - leafcell, Cell - misc_module4rev, View - schematic
// LAST TIME SAVED: Aug 21 17:26:57 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module misc_module4rev ( S_R, cin2lcl, clk, clkb, glb2local, sp4, bl,
     b, carry_in, glb_netwk, l, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, m, min0, min1, min2, min3, pgate, prog, r, reset_b,
     sp12, vdd_cntl, wl );
output  S_R, cin2lcl, clk, clkb;


input  carry_in, prog;

output [7:0]  sp4;
output [3:0]  glb2local;

inout [3:0]  bl;

input [15:0]  reset_b;
input [15:0]  pgate;
input [7:0]  sp12;
input [1:0]  m;
input [7:0]  min0;
input [15:0]  vdd_cntl;
input [5:0]  lc_trk_g0;
input [1:0]  l;
input [5:0]  lc_trk_g2;
input [15:0]  wl;
input [1:0]  b;
input [7:0]  min3;
input [7:0]  glb_netwk;
input [7:0]  min1;
input [5:0]  lc_trk_g3;
input [5:0]  lc_trk_g1;
input [7:0]  min2;
input [1:0]  r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [63:0]  cbitb;

wire  [15:0]  r_vdd;

wire  [63:0]  cbit;



pch_hvt  vdd_cntrl_15_ ( .D(r_vdd[15]), .B(vdd_), .G(vdd_cntl[15]),
     .S(vdd_));
pch_hvt  vdd_cntrl_14_ ( .D(r_vdd[14]), .B(vdd_), .G(vdd_cntl[14]),
     .S(vdd_));
pch_hvt  vdd_cntrl_13_ ( .D(r_vdd[13]), .B(vdd_), .G(vdd_cntl[13]),
     .S(vdd_));
pch_hvt  vdd_cntrl_12_ ( .D(r_vdd[12]), .B(vdd_), .G(vdd_cntl[12]),
     .S(vdd_));
pch_hvt  vdd_cntrl_11_ ( .D(r_vdd[11]), .B(vdd_), .G(vdd_cntl[11]),
     .S(vdd_));
pch_hvt  vdd_cntrl_10_ ( .D(r_vdd[10]), .B(vdd_), .G(vdd_cntl[10]),
     .S(vdd_));
pch_hvt  vdd_cntrl_9_ ( .D(r_vdd[9]), .B(vdd_), .G(vdd_cntl[9]),
     .S(vdd_));
pch_hvt  vdd_cntrl_8_ ( .D(r_vdd[8]), .B(vdd_), .G(vdd_cntl[8]),
     .S(vdd_));
pch_hvt  vdd_cntrl_7_ ( .D(r_vdd[7]), .B(vdd_), .G(vdd_cntl[7]),
     .S(vdd_));
pch_hvt  vdd_cntrl_6_ ( .D(r_vdd[6]), .B(vdd_), .G(vdd_cntl[6]),
     .S(vdd_));
pch_hvt  vdd_cntrl_5_ ( .D(r_vdd[5]), .B(vdd_), .G(vdd_cntl[5]),
     .S(vdd_));
pch_hvt  vdd_cntrl_4_ ( .D(r_vdd[4]), .B(vdd_), .G(vdd_cntl[4]),
     .S(vdd_));
pch_hvt  vdd_cntrl_3_ ( .D(r_vdd[3]), .B(vdd_), .G(vdd_cntl[3]),
     .S(vdd_));
pch_hvt  vdd_cntrl_2_ ( .D(r_vdd[2]), .B(vdd_), .G(vdd_cntl[2]),
     .S(vdd_));
pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clkmandcmuxrev Itclkm ( .min2(min2[7:0]), .min1(min1[7:0]),
     .min0(min0[7:0]), .min3(min3[7:0]), .cbit({cbit[2], cbit[1],
     cbit[0], cbit[27], cbit[25], cbit[26], cbit[24], cbit[23],
     cbit[21], cbit[22], cbit[20], cbit[19], cbit[17], cbit[18],
     cbit[16], cbit[15], cbit[13], cbit[14], cbit[12], cbit[31],
     cbit[29], cbit[30], cbit[28], cbit[11], cbit[9], cbit[10],
     cbit[8], cbit[38], cbit[36], cbit[7], cbit[6], cbit[4]}),
     .cbitb({cbitb[2], cbitb[1], cbitb[0], cbitb[27], cbitb[25],
     cbitb[26], cbitb[24], cbitb[23], cbitb[21], cbitb[22], cbitb[20],
     cbitb[19], cbitb[17], cbitb[18], cbitb[16], cbitb[15], cbitb[13],
     cbitb[14], cbitb[12], cbitb[31], cbitb[29], cbitb[30], cbitb[28],
     cbitb[11], cbitb[9], cbitb[10], cbitb[8], cbitb[38], cbitb[36],
     cbitb[7], cbitb[6], cbitb[4]}), .glb2local(glb2local[3:0]),
     .lc_trk_g0(lc_trk_g0[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .lc_trk_g2(lc_trk_g2[5:0]), .lc_trk_g3(lc_trk_g3[5:0]),
     .glb_netwk(glb_netwk[7:0]), .prog(prog), .cin2lcl(cin2lcl),
     .clk(clk), .clkb(clkb), .s_r(S_R), .carry_in(carry_in));
sp12to4 Isp12to4_7_ ( .triout(sp4[7]), .cbitb(cbitb[62]),
     .drv(sp12[7]), .prog(net109));
sp12to4 Isp12to4_6_ ( .triout(sp4[6]), .cbitb(cbitb[58]),
     .drv(sp12[6]), .prog(net109));
sp12to4 Isp12to4_5_ ( .triout(sp4[5]), .cbitb(cbitb[54]),
     .drv(sp12[5]), .prog(net109));
sp12to4 Isp12to4_4_ ( .triout(sp4[4]), .cbitb(cbitb[50]),
     .drv(sp12[4]), .prog(net109));
sp12to4 Isp12to4_3_ ( .triout(sp4[3]), .cbitb(cbitb[46]),
     .drv(sp12[3]), .prog(net109));
sp12to4 Isp12to4_2_ ( .triout(sp4[2]), .cbitb(cbitb[42]),
     .drv(sp12[2]), .prog(net109));
sp12to4 Isp12to4_1_ ( .triout(sp4[1]), .cbitb(cbitb[5]), .drv(sp12[1]),
     .prog(net109));
sp12to4 Isp12to4_0_ ( .triout(sp4[0]), .cbitb(cbitb[34]),
     .drv(sp12[0]), .prog(net109));
sbox1 Isp12_1_ ( .l(l[1]), .cb({cbitb[63], cbitb[61], cbitb[59],
     cbitb[57], cbitb[55], cbitb[53], cbitb[51], cbitb[49]}), .r(r[1]),
     .t(m[1]), .b(b[1]), .c({cbit[63], cbit[61], cbit[59], cbit[57],
     cbit[55], cbit[53], cbit[51], cbit[49]}), .prog(prog));
sbox1 Isp12_0_ ( .l(l[0]), .cb({cbitb[47], cbitb[45], cbitb[43],
     cbitb[41], cbitb[39], cbitb[37], cbitb[35], cbitb[33]}), .r(r[0]),
     .t(m[0]), .b(b[0]), .c({cbit[47], cbit[45], cbit[43], cbit[41],
     cbit[39], cbit[37], cbit[35], cbit[33]}), .prog(prog));
cram16x4 Ic64 ( .r_gnd(r_vdd[15:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .q(cbit[63:0]), .wl(wl[15:0]),
     .q_b(cbitb[63:0]), .bl(bl[3:0]));
inv_hvt I61 ( .A(prog), .Y(progb));
inv_hvt I62 ( .A(progb), .Y(net109));

endmodule
// Library - leafcell, Cell - bram_routing_tracks4rev, View - schematic
// LAST TIME SAVED: Nov  2 15:55:57 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_routing_tracks4rev ( clk, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, s_r, bl, sp4_h_l, sp4_h_r, sp4_r_v_b, sp4_v_b, sp4_v_t,
     sp12_h_l, sp12_h_r, sp12_v_b, sp12_v_t, bnl_op, bnr_op, bot_op,
     carry_in, glb_netwk, lft_op, pgate, prog, reset_b, rgt_op, slf_op,
     tnl_op, tnr_op, top_op, vdd_cntl, wl );
output  clk, s_r;


input  carry_in, prog;

output [7:0]  lc_trk_g2;
output [7:0]  lc_trk_g0;
output [7:0]  lc_trk_g3;
output [7:0]  lc_trk_g1;

inout [47:0]  sp4_r_v_b;
inout [47:0]  sp4_v_b;
inout [47:0]  sp4_h_l;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_v_t;
inout [23:0]  sp12_h_r;
inout [23:0]  sp12_v_b;
inout [25:0]  bl;
inout [47:0]  sp4_h_r;
inout [23:0]  sp12_v_t;

input [15:0]  reset_b;
input [7:0]  bnl_op;
input [7:0]  lft_op;
input [7:0]  bot_op;
input [15:0]  pgate;
input [7:0]  top_op;
input [7:0]  rgt_op;
input [7:0]  bnr_op;
input [7:0]  tnl_op;
input [7:0]  tnr_op;
input [15:0]  wl;
input [7:0]  glb_netwk;
input [7:0]  slf_op;
input [15:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  net_glb2local;

wire  [1:0]  sp12_v_b_mid;

wire  [1:0]  sp12_h_r_mid;



rm6  R0_23_ ( .MINUS(sp12_h_r[23]), .PLUS(sp12_h_l[20]));
rm6  R0_22_ ( .MINUS(sp12_h_r[22]), .PLUS(sp12_h_l[21]));
rm6  R0_21_ ( .MINUS(sp12_h_r[21]), .PLUS(sp12_h_l[18]));
rm6  R0_20_ ( .MINUS(sp12_h_r[20]), .PLUS(sp12_h_l[19]));
rm6  R0_19_ ( .MINUS(sp12_h_r[19]), .PLUS(sp12_h_l[16]));
rm6  R0_18_ ( .MINUS(sp12_h_r[18]), .PLUS(sp12_h_l[17]));
rm6  R0_17_ ( .MINUS(sp12_h_r[17]), .PLUS(sp12_h_l[14]));
rm6  R0_16_ ( .MINUS(sp12_h_r[16]), .PLUS(sp12_h_l[15]));
rm6  R0_15_ ( .MINUS(sp12_h_r[15]), .PLUS(sp12_h_l[12]));
rm6  R0_14_ ( .MINUS(sp12_h_r[14]), .PLUS(sp12_h_l[13]));
rm6  R0_13_ ( .MINUS(sp12_h_r[13]), .PLUS(sp12_h_l[10]));
rm6  R0_12_ ( .MINUS(sp12_h_r[12]), .PLUS(sp12_h_l[11]));
rm6  R0_11_ ( .MINUS(sp12_h_r[11]), .PLUS(sp12_h_l[8]));
rm6  R0_10_ ( .MINUS(sp12_h_r[10]), .PLUS(sp12_h_l[9]));
rm6  R0_9_ ( .MINUS(sp12_h_r[9]), .PLUS(sp12_h_l[6]));
rm6  R0_8_ ( .MINUS(sp12_h_r[8]), .PLUS(sp12_h_l[7]));
rm6  R0_7_ ( .MINUS(sp12_h_r[7]), .PLUS(sp12_h_l[4]));
rm6  R0_6_ ( .MINUS(sp12_h_r[6]), .PLUS(sp12_h_l[5]));
rm6  R0_5_ ( .MINUS(sp12_h_r[5]), .PLUS(sp12_h_l[2]));
rm6  R0_4_ ( .MINUS(sp12_h_r[4]), .PLUS(sp12_h_l[3]));
rm6  R0_3_ ( .MINUS(sp12_h_r[3]), .PLUS(sp12_h_l[0]));
rm6  R0_2_ ( .MINUS(sp12_h_r[2]), .PLUS(sp12_h_l[1]));
rm6  R0_1_ ( .MINUS(sp12_h_r_mid[1]), .PLUS(sp12_h_l[22]));
rm6  R0_0_ ( .MINUS(sp12_h_r_mid[0]), .PLUS(sp12_h_l[23]));
rm7  R2_23_ ( .MINUS(sp12_v_b[23]), .PLUS(sp12_v_t[20]));
rm7  R2_22_ ( .MINUS(sp12_v_b[22]), .PLUS(sp12_v_t[21]));
rm7  R2_21_ ( .MINUS(sp12_v_b[21]), .PLUS(sp12_v_t[18]));
rm7  R2_20_ ( .MINUS(sp12_v_b[20]), .PLUS(sp12_v_t[19]));
rm7  R2_19_ ( .MINUS(sp12_v_b[19]), .PLUS(sp12_v_t[16]));
rm7  R2_18_ ( .MINUS(sp12_v_b[18]), .PLUS(sp12_v_t[17]));
rm7  R2_17_ ( .MINUS(sp12_v_b[17]), .PLUS(sp12_v_t[14]));
rm7  R2_16_ ( .MINUS(sp12_v_b[16]), .PLUS(sp12_v_t[15]));
rm7  R2_15_ ( .MINUS(sp12_v_b[15]), .PLUS(sp12_v_t[12]));
rm7  R2_14_ ( .MINUS(sp12_v_b[14]), .PLUS(sp12_v_t[13]));
rm7  R2_13_ ( .MINUS(sp12_v_b[13]), .PLUS(sp12_v_t[10]));
rm7  R2_12_ ( .MINUS(sp12_v_b[12]), .PLUS(sp12_v_t[11]));
rm7  R2_11_ ( .MINUS(sp12_v_b[11]), .PLUS(sp12_v_t[8]));
rm7  R2_10_ ( .MINUS(sp12_v_b[10]), .PLUS(sp12_v_t[9]));
rm7  R2_9_ ( .MINUS(sp12_v_b[9]), .PLUS(sp12_v_t[6]));
rm7  R2_8_ ( .MINUS(sp12_v_b[8]), .PLUS(sp12_v_t[7]));
rm7  R2_7_ ( .MINUS(sp12_v_b[7]), .PLUS(sp12_v_t[4]));
rm7  R2_6_ ( .MINUS(sp12_v_b[6]), .PLUS(sp12_v_t[5]));
rm7  R2_5_ ( .MINUS(sp12_v_b[5]), .PLUS(sp12_v_t[2]));
rm7  R2_4_ ( .MINUS(sp12_v_b[4]), .PLUS(sp12_v_t[3]));
rm7  R2_3_ ( .MINUS(sp12_v_b[3]), .PLUS(sp12_v_t[0]));
rm7  R2_2_ ( .MINUS(sp12_v_b[2]), .PLUS(sp12_v_t[1]));
rm7  R2_1_ ( .MINUS(sp12_v_b_mid[1]), .PLUS(sp12_v_t[22]));
rm7  R2_0_ ( .MINUS(sp12_v_b_mid[0]), .PLUS(sp12_v_t[23]));
inv_hvt I89 ( .A(progb), .Y(progd));
inv_hvt I90 ( .A(prog), .Y(progb));
gmux_sp12to4 Igmux_sp12to4 ( .vdd_cntl(vdd_cntl[15:0]), .wl(wl[15:0]),
     .top_op(top_op[7:0]), .tnr_op(tnr_op[7:0]), .tnl_op(tnl_op[7:0]),
     .slf_op(slf_op[7:0]), .rgt_op(rgt_op[7:0]), .prog(progd),
     .lft_op(lft_op[7:0]), .bnr_op(bnr_op[7:0]), .bnl_op(bnl_op[7:0]),
     .lc_trk_g0(lc_trk_g0[7:0]), .lc_trk_g3(lc_trk_g3[7:0]),
     .lc_trk_g2(lc_trk_g2[7:0]), .lc_trk_g1(lc_trk_g1[7:0]),
     .bot_op(bot_op[7:0]), .glb2local(net_glb2local[3:0]),
     .reset_b(reset_b[15:0]), .pgate(pgate[15:0]),
     .sp12_v_b(sp12_v_b[23:0]), .bl(bl[25:14]),
     .sp4_r_v_b(sp4_r_v_b[47:0]), .sp12_h_r(sp12_h_r[23:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_r(sp4_h_r[47:0]));
span4 Isp4_sw ( .vdd_cntl(vdd_cntl[15:0]), .sp4_h_r(sp4_h_r[47:0]),
     .sp4_v_b(sp4_v_b[47:0]), .sp4_h_l(sp4_h_l[47:0]),
     .sp4_v_t(sp4_v_t[47:0]), .reset_b(reset_b[15:0]),
     .pgate(pgate[15:0]), .prog(progd), .wl(wl[15:0]), .bl(bl[13:4]));
misc_module4rev Ickmux_sp12to4_sp12sw ( .vdd_cntl(vdd_cntl[15:0]),
     .prog(progd), .carry_in(carry_in), .lc_trk_g0(lc_trk_g0[5:0]),
     .glb_netwk(glb_netwk[7:0]), .lc_trk_g2(lc_trk_g2[5:0]),
     .lc_trk_g3(lc_trk_g3[5:0]), .lc_trk_g1(lc_trk_g1[5:0]),
     .cin2lcl(net174), .wl(wl[15:0]), .S_R(s_r), .clkb(clkb),
     .bl(bl[3:0]), .clk(clk), .sp4(sp4_h_r[23:16]),
     .sp12({sp12_h_r[22], sp12_h_r[20], sp12_h_r[18], sp12_h_r[16],
     sp12_h_r[14], sp12_h_r[12], sp12_h_r[10], sp12_h_r[8]}),
     .reset_b(reset_b[15:0]), .b(sp12_v_b[1:0]), .r(sp12_h_r[1:0]),
     .m(sp12_v_b_mid[1:0]), .l(sp12_h_r_mid[1:0]), .pgate(pgate[15:0]),
     .glb2local(net_glb2local[3:0]), .min2(glb_netwk[7:0]),
     .min1(glb_netwk[7:0]), .min0(glb_netwk[7:0]),
     .min3(glb_netwk[7:0]));

endmodule
// Library - leafcell, Cell - bram_bufferx6, View - schematic
// LAST TIME SAVED: Jun 25 13:45:32 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_bufferx6 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I3 ( .A(in), .Y(net4));
inv_hvt I4 ( .A(net4), .Y(out));

endmodule
// Library - leafcell, Cell - bram_bufferx1, View - schematic
// LAST TIME SAVED: Jun 14 08:59:24 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_bufferx1 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I0 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - leafcell, Cell - bram_4k_buffer, View - schematic
// LAST TIME SAVED: Oct  6 13:53:19 2008
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_buffer ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;

input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



tielo I22 ( .tielo(net055));
bram_bufferx1 I15 ( .in(net055), .out(net49));
bram_bufferx1 I16 ( .in(net49), .out(net52));
bram_bufferx1 I17 ( .in(net52), .out(net53));
bram_bufferx1 I18 ( .in(net53), .out(net55));
bram_bufferx6 I14 ( .in(bm_sdo_i), .out(bm_sdo_o));
bram_bufferx6 I6 ( .in(bm_sdi_i), .out(bm_sdi_o));
bram_bufferx6 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx6 I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx6 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx6 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx6 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx6 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx6 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx6 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx6 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx6 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx6 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx6 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx6 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx6 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx6 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Jun  5 11:34:46 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module leafcell_ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tiehigh, View - schematic
// LAST TIME SAVED: May  8 16:23:56 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module vdd_tiehigh ( vdd_tieh );
inout  vdd_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(vdd_tieh), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - leafcell, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:59 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module ml_mux2_hvt_schematic ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - leafcell, Cell - bram_dff_mux, View - schematic
// LAST TIME SAVED: Jul 25 16:06:22 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_dff_mux ( q, bm_q, bm_sdi, ce, clk, rcapmux_en, rst );
output  q;

input  bm_q, bm_sdi, ce, clk, rcapmux_en, rst;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



leafcell_ml_dff_schematic I2 ( .R(rst), .D(net020), .CLK(clk),
     .QN(net10), .Q(q));
ml_mux2_hvt_schematic I5 ( .in1(net14), .in0(q), .out(net020),
     .sel(ce));
ml_mux2_hvt_schematic I1 ( .in1(bm_q), .in0(bm_sdi), .out(net14),
     .sel(rcapmux_en));

endmodule
// Library - leafcell, Cell - bram_4k_sr_bankout, View - schematic
// LAST TIME SAVED: Jul 25 22:59:22 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_sr_bankout ( bm_dm, bm_sdo, bm_sweb, clk, rcapmux_en,
     rst, bm_q, bm_sdi, wdummymux_en );
output  bm_sdo;

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[0]), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));
leafcell_ml_dff_schematic I29 ( .R(rst), .D(net0151), .CLK(clk),
     .QN(net0160), .Q(bm_sdo));
leafcell_ml_dff_schematic I22 ( .R(rst), .D(bm_dm[14]), .CLK(clk),
     .QN(net165), .Q(rdummy_reg));
ml_mux2_hvt_schematic I21 ( .in1(rdummy_reg), .in0(bm_dm[15]),
     .out(net0151), .sel(rdummymux_en));
nor2_hvt I24 ( .A(bm_swe), .B(rcapmux_en), .Y(net148));
inv_hvt I19 ( .A(bm_sweb), .Y(bm_swe));
inv_hvt I23 ( .A(net148), .Y(rdummymux_en));

endmodule
// Library - leafcell, Cell - bram_4k_bankout, View - schematic
// LAST TIME SAVED: Aug 15 18:09:39 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_bankout ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_ab;
input [7:0]  bm_sa;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [15:0]  bm_dm;



tielo I15 ( .tielo(net092));
tielo I18 ( .tielo(net093));
bram_4k_sr_bankout I12 ( .bm_dm(bm_dm[15:0]), .rst(net093),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]), .bm_sdo(bm_sdo));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM(bm_dm[15:0]), .WEBM(bm_sweb), .WEB(web), .REBM(bm_sreb),
     .REB(reb), .D(bm_d[15:0]), .CLKW(net074), .CLKR(net072),
     .BWEBM({net092, net092, net092, net092, net092, net092, net092,
     net092, net092, net092, net092, net092, net092, net092, net092,
     net092}), .BWEB(bm_bweb[15:0]), .BIST(bm_init), .AMB(bm_sa[7:0]),
     .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]), .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net89), .out(net072));
bram_bufferx6 I8 ( .in(net85), .out(net074));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net85), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net89), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - leafcell, Cell - bram_4kbankout_pbuffer_bot, View -
//schematic
// LAST TIME SAVED: Aug 24 17:34:26 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4kbankout_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;

input [7:0]  bm_aa;
input [15:0]  bm_bweb;
input [7:0]  bm_sa_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sclkrw_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [1:0]  bm_sweb_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankout I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4k_inmux3_0, View - schematic
// LAST TIME SAVED: Aug 23 11:45:13 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_inmux3_0 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_h_r;

input  op, prog;

output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;
output [2:0]  sp4_h_r;
output [1:0]  sp12_v_b;

input [15:0]  min3;
input [15:0]  min0;
input [1:0]  reset_b;
input [1:0]  vdd_cntl;
input [1:0]  wl;
input [15:0]  min1;
input [15:0]  bl;
input [15:0]  min2;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [31:0]  cbitb;

wire  [31:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12_30 Iodrv74 ( .sp12_h_r(sp12_h_r), .sp12_v_b(sp12_v_b[1:0]),
     .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
in_mux in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux7_4, View - schematic
// LAST TIME SAVED: Aug 23 11:44:11 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_inmux7_4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, min0, min1, min2, min3, op,
     pgate, prog, reset_b, vdd_cntl, wl );
output  in0, in1, in2, in3, sp12_v_b;

input  op, prog;

output [1:0]  sp12_h_r;
output [2:0]  sp4_h_r;
output [2:0]  sp4_r_v_b;
output [2:0]  sp4_v_b;

input [15:0]  min3;
input [15:0]  min0;
input [15:0]  bl;
input [1:0]  vdd_cntl;
input [15:0]  min1;
input [1:0]  wl;
input [1:0]  pgate;
input [15:0]  min2;
input [1:0]  reset_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [31:0]  cbit;

wire  [31:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 I0_7_ ( .bl(bl[15:14]), .q_b(cbitb[31:28]), .q(cbit[31:28]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_6_ ( .bl(bl[13:12]), .q_b(cbitb[27:24]), .q(cbit[27:24]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_5_ ( .bl(bl[11:10]), .q_b(cbitb[23:20]), .q(cbit[23:20]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_4_ ( .bl(bl[9:8]), .q_b(cbitb[19:16]), .q(cbit[19:16]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_3_ ( .bl(bl[7:6]), .q_b(cbitb[15:12]), .q(cbit[15:12]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .q(cbit[11:8]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .q(cbit[7:4]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
cram2x2 I0_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .q(cbit[3:0]),
     .wl(wl[1:0]), .pgate(pgate[1:0]), .r_vdd(r_vdd[1:0]),
     .reset(reset_b[1:0]));
odrv12_74 Iodrv74 ( .slfop(op), .prog(prog), .cbitb(cbitb[31:20]),
     .sp4_r_v_b(sp4_r_v_b[2:0]), .sp4_v_b(sp4_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .sp12_v_b(sp12_v_b),
     .sp12_h_r(sp12_h_r[1:0]));
in_mux in3mux ( .prog(prog), .inmuxo(in3), .cbit({cbit[14], cbit[15],
     cbit[18], cbit[11], cbit[9]}), .cbitb({cbitb[14], cbitb[15],
     cbitb[18], cbitb[11], cbitb[9]}), .min(min3[15:0]));
in_mux in2mux ( .prog(prog), .inmuxo(in2), .cbit({cbit[12], cbit[13],
     cbit[16], cbit[19], cbit[17]}), .cbitb({cbitb[12], cbitb[13],
     cbitb[16], cbitb[19], cbitb[17]}), .min(min2[15:0]));
in_mux in0mux ( .prog(prog), .inmuxo(in0), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));
in_mux in1mux ( .prog(prog), .inmuxo(in1), .cbit({cbit[7], cbit[6],
     cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));

endmodule
// Library - leafcell, Cell - bram_4k_inmux_8x4, View - schematic
// LAST TIME SAVED: Aug 29 16:20:56 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_inmux_8x4 ( in0, in1, in2, in3, sp4_h_r, sp4_r_v_b,
     sp4_v_b, sp12_h_r, sp12_v_b, bl, lc_trk_g0, lc_trk_g1, lc_trk_g2,
     lc_trk_g3, op, pgate, prog, reset_b, vdd_cntl, wl );

input  prog;

output [23:0]  sp4_r_v_b;
output [23:0]  sp4_h_r;
output [7:0]  in3;
output [7:0]  in2;
output [7:0]  in1;
output [11:0]  sp12_v_b;
output [11:0]  sp12_h_r;
output [23:0]  sp4_v_b;
output [7:0]  in0;

input [15:0]  bl;
input [7:0]  op;
input [7:0]  lc_trk_g0;
input [7:0]  lc_trk_g2;
input [15:0]  reset_b;
input [7:0]  lc_trk_g1;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [7:0]  lc_trk_g3;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_inmux3_0 I3 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[3]), .sp12_v_b(sp12_v_b[7:6]), .wl(wl[7:6]),
     .reset_b(reset_b[7:6]), .prog(progd), .pgate(pgate[7:6]),
     .op(op[3]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[11:9]), .sp4_r_v_b(sp4_r_v_b[11:9]),
     .sp4_h_r(sp4_h_r[11:9]), .in3(in3[3]), .in2(in2[3]), .in1(in1[3]),
     .in0(in0[3]));
bram_4k_inmux3_0 I2 ( .vdd_cntl(vdd_cntl[5:4]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[2]), .sp12_v_b(sp12_v_b[5:4]), .wl(wl[5:4]),
     .reset_b(reset_b[5:4]), .prog(progd), .pgate(pgate[5:4]),
     .op(op[2]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[8:6]), .sp4_r_v_b(sp4_r_v_b[8:6]),
     .sp4_h_r(sp4_h_r[8:6]), .in3(in3[2]), .in2(in2[2]), .in1(in1[2]),
     .in0(in0[2]));
bram_4k_inmux3_0 I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[1]), .sp12_v_b(sp12_v_b[3:2]), .wl(wl[3:2]),
     .reset_b(reset_b[3:2]), .prog(progd), .pgate(pgate[3:2]),
     .op(op[1]), .min3({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3],
     lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2],
     lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3],
     lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], tiehi}),
     .min2({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min1({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min0({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp4_v_b(sp4_v_b[5:3]), .sp4_r_v_b(sp4_r_v_b[5:3]),
     .sp4_h_r(sp4_h_r[5:3]), .in3(in3[1]), .in2(in2[1]), .in1(in1[1]),
     .in0(in0[1]));
bram_4k_inmux3_0 I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[15:0]),
     .sp12_h_r(sp12_h_r[0]), .sp12_v_b(sp12_v_b[1:0]), .wl(wl[1:0]),
     .reset_b(reset_b[1:0]), .prog(progd), .pgate(pgate[1:0]),
     .op(op[0]), .min3({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2],
     lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3],
     lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2],
     lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], tiehi}),
     .min2({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .min1({lc_trk_g3[6], lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0],
     lc_trk_g2[7], lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1],
     lc_trk_g1[6], lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0],
     lc_trk_g0[7], lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .min0({lc_trk_g3[7], lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1],
     lc_trk_g2[6], lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0],
     lc_trk_g1[7], lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1],
     lc_trk_g0[6], lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp4_v_b(sp4_v_b[2:0]), .sp4_r_v_b(sp4_r_v_b[2:0]),
     .sp4_h_r(sp4_h_r[2:0]), .in3(in3[0]), .in2(in2[0]), .in1(in1[0]),
     .in0(in0[0]));
tiehi I10 ( .tiehi(tiehi));
bram_4k_inmux7_4 I6 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[15:0]),
     .wl(wl[13:12]), .reset_b(reset_b[13:12]), .prog(progd),
     .pgate(pgate[13:12]), .op(op[6]), .min3({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}),
     .sp12_v_b(sp12_v_b[10]), .sp12_h_r(sp12_h_r[9:8]),
     .sp4_v_b(sp4_v_b[20:18]), .sp4_r_v_b(sp4_r_v_b[20:18]),
     .sp4_h_r(sp4_h_r[20:18]), .in3(in3[6]), .in2(in2[6]),
     .in1(in1[6]), .in0(in0[6]));
bram_4k_inmux7_4 I5 ( .vdd_cntl(vdd_cntl[11:10]), .bl(bl[15:0]),
     .wl(wl[11:10]), .reset_b(reset_b[11:10]), .prog(progd),
     .pgate(pgate[11:10]), .op(op[5]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[9]), .sp12_h_r(sp12_h_r[7:6]),
     .sp4_v_b(sp4_v_b[17:15]), .sp4_r_v_b(sp4_r_v_b[17:15]),
     .sp4_h_r(sp4_h_r[17:15]), .in3(in3[5]), .in2(in2[5]),
     .in1(in1[5]), .in0(in0[5]));
bram_4k_inmux7_4 I4 ( .vdd_cntl(vdd_cntl[9:8]), .bl(bl[15:0]),
     .wl(wl[9:8]), .reset_b(reset_b[9:8]), .prog(progd),
     .pgate(pgate[9:8]), .op(op[4]), .min3({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], tiehi}), .min2({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min1({lc_trk_g3[6], lc_trk_g3[4],
     lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7], lc_trk_g2[5],
     lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min0({lc_trk_g3[7], lc_trk_g3[5],
     lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6], lc_trk_g2[4],
     lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .sp12_v_b(sp12_v_b[8]),
     .sp12_h_r(sp12_h_r[5:4]), .sp4_v_b(sp4_v_b[14:12]),
     .sp4_r_v_b(sp4_r_v_b[14:12]), .sp4_h_r(sp4_h_r[14:12]),
     .in3(in3[4]), .in2(in2[4]), .in1(in1[4]), .in0(in0[4]));
bram_4k_inmux7_4 I7 ( .vdd_cntl(vdd_cntl[15:14]), .bl(bl[15:0]),
     .wl(wl[15:14]), .reset_b(reset_b[15:14]), .prog(progd),
     .pgate(pgate[15:14]), .op(op[7]), .min3({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], tiehi}), .min2({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g3[7],
     lc_trk_g3[5], lc_trk_g3[3], lc_trk_g3[1], lc_trk_g2[6],
     lc_trk_g2[4], lc_trk_g2[2], lc_trk_g2[0], lc_trk_g1[7],
     lc_trk_g1[5], lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6],
     lc_trk_g0[4], lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g3[6],
     lc_trk_g3[4], lc_trk_g3[2], lc_trk_g3[0], lc_trk_g2[7],
     lc_trk_g2[5], lc_trk_g2[3], lc_trk_g2[1], lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .sp12_v_b(sp12_v_b[11]), .sp12_h_r(sp12_h_r[11:10]),
     .sp4_v_b(sp4_v_b[23:21]), .sp4_r_v_b(sp4_r_v_b[23:21]),
     .sp4_h_r(sp4_h_r[23:21]), .in3(in3[7]), .in2(in2[7]),
     .in1(in1[7]), .in0(in0[7]));
inv_hvt I81 ( .A(prog), .Y(progb));
inv_hvt I82 ( .A(progb), .Y(progd));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbankout, View -
//schematic
// LAST TIME SAVED: Mar  6 11:33:30 2008
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4kprouting_bbankout ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_top;

inout [47:0]  sp4_h_l_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_h_l_top;
inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_r_bot;

input [7:0]  rgt_op_bot;
input [7:0]  tnl_op_top;
input [1:0]  bm_sdo_i;
input [7:0]  tnr_op_bot;
input [7:0]  bnr_op_top;
input [1:0]  bm_sdi_i;
input [7:0]  lft_op_top;
input [7:0]  top_op_top;
input [7:0]  bot_op_bot;
input [1:0]  bm_sweb_i;
input [7:0]  bnl_op_bot;
input [7:0]  tnl_op_bot;
input [7:0]  bm_sa_i;
input [7:0]  bnr_op_bot;
input [7:0]  lft_op_bot;
input [7:0]  tnr_op_top;
input [7:0]  bnl_op_top;
input [15:0]  wl_top;
input [15:0]  wl_bot;
input [7:0]  glb_netwk;
input [15:0]  reset_b_top;
input [15:0]  pgate_top;
input [1:0]  bm_sclkrw_i;
input [15:0]  vdd_cntl_bot;
input [15:0]  vdd_cntl_top;
input [15:0]  reset_b_bot;
input [15:0]  pgate_bot;
input [7:0]  rgt_op_top;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net284;

wire  [0:7]  net251;

wire  [0:7]  net285;

wire  [0:7]  net254;

wire  [0:7]  net283;

wire  [0:7]  net252;

wire  [0:7]  net286;

wire  [0:7]  net253;

wire  [0:7]  net341;

wire  [0:7]  net320;



bram_routing_tracks4rev I_bot ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}), .s_r(net234),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(tnr_op_bot[7:0]),
     .tnl_op(tnl_op_bot[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net299),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net251[0:7]),
     .lc_trk_g2(net252[0:7]), .lc_trk_g1(net253[0:7]),
     .lc_trk_g0(net254[0:7]), .clk(net255),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev I_top ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}), .s_r(net266),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net298),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net283[0:7]),
     .lc_trk_g2(net284[0:7]), .lc_trk_g1(net285[0:7]),
     .lc_trk_g0(net286[0:7]), .clk(net287),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbankout_pbuffer_bot I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net266), .bm_wen(net234),
     .bm_d(bm_d[15:0]), .bm_clkr(net287), .bm_clkw(net255),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_ab(net341[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net320[0:7]),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
tielo I14 ( .tielo(net298));
tielo I15 ( .tielo(net299));
bram_4k_inmux_8x4 I6 ( .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15],
     vdd_cntl_bot[12], vdd_cntl_bot[13], vdd_cntl_bot[10],
     vdd_cntl_bot[11], vdd_cntl_bot[8], vdd_cntl_bot[9],
     vdd_cntl_bot[6], vdd_cntl_bot[7], vdd_cntl_bot[4],
     vdd_cntl_bot[5], vdd_cntl_bot[2], vdd_cntl_bot[3],
     vdd_cntl_bot[0], vdd_cntl_bot[1]}), .bl(bl[41:26]),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net320[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15],
     vdd_cntl_top[12], vdd_cntl_top[13], vdd_cntl_top[10],
     vdd_cntl_top[11], vdd_cntl_top[8], vdd_cntl_top[9],
     vdd_cntl_top[6], vdd_cntl_top[7], vdd_cntl_top[4],
     vdd_cntl_top[5], vdd_cntl_top[2], vdd_cntl_top[3],
     vdd_cntl_top[0], vdd_cntl_top[1]}), .bl(bl[41:26]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}), .op(slf_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net341[0:7]));

endmodule
// Library - leafcell, Cell - bram_4k_sr, View - schematic
// LAST TIME SAVED: Aug 15 17:41:16 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_sr ( bm_dm, bm_sweb, clk, rcapmux_en, rst, bm_q, bm_sdi,
     wdummymux_en );

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[0]), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));

endmodule
// Library - misc, Cell - eh_io_pup_2_new, View - schematic
// LAST TIME SAVED: Oct  6 15:01:46 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module eh_io_pup_2_new ( por_b, core_por_b, vdd_io );
output  por_b;

input  core_por_b, vdd_io;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_hvt  MP8 ( .D(net104), .B(vdd_), .G(core_por_b), .S(vdd_));
pch_hvt  M4 ( .D(por_b), .B(vdd_), .G(net92), .S(vdd_));
pch_hvt  M1 ( .D(net92), .B(vdd_), .G(net84), .S(vdd_));
pch_hvt  M0 ( .D(net84), .B(vdd_), .G(net104), .S(vdd_));
nch_hvt  M5 ( .D(por_b), .B(gnd_), .G(net92), .S(gnd_));
nch_hvt  M3 ( .D(net92), .B(gnd_), .G(net84), .S(gnd_));
nch_hvt  MN1 ( .D(net80), .B(gnd_), .G(core_por_b), .S(gnd_));
nch_hvt  M2 ( .D(net84), .B(gnd_), .G(net104), .S(gnd_));
pch_25  M6 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  MP11 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
pch_25  MP13 ( .D(net124), .B(vdd_io), .G(net145), .S(net122));
pch_25  MP12 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  M7 ( .D(net122), .B(vdd_io), .G(net122), .S(vdd_io));
pch_25  MP7 ( .D(net104), .B(vdd_), .G(net124), .S(vdd_));
pch_25  MP9 ( .D(vdd_io), .B(vdd_io), .G(vdd_io), .S(vdd_io));
nch_25  MN6 ( .D(net124), .B(gnd_), .G(net145), .S(gnd_));
nch_25  MN38 ( .D(net104), .B(gnd_), .G(net124), .S(net104));
nch_25  M10 ( .D(net124), .B(gnd_), .G(net147), .S(net158));
nch_25  MN39 ( .D(net104), .B(gnd_), .G(net124), .S(net80));
nch_25  M11 ( .D(net140), .B(gnd_), .G(core_por_b), .S(gnd_));
rppolywo_m  R66 ( .MINUS(gnd_), .PLUS(net145), .BULK(gnd_));
vdd_tiehigh I96 ( .vdd_tieh(net147));
nch_na25  M15 ( .D(net154), .B(gnd_), .G(net154), .S(net150));
nch_na25  M16 ( .D(net158), .B(gnd_), .G(net158), .S(net154));
nch_na25  M17 ( .D(net162), .B(gnd_), .G(net162), .S(net166));
nch_na25  M14 ( .D(net150), .B(gnd_), .G(net150), .S(net162));
nch_na25  M18 ( .D(net166), .B(gnd_), .G(net166), .S(net140));

endmodule
// Library - leafcell, Cell - bram_4k, View - schematic
// LAST TIME SAVED: Aug 15 17:44:47 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr, bm_clkw,
     bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk, bm_sclkrw,
     bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_sa;
input [7:0]  bm_ab;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [14:0]  bm_dm;



tielo I15 ( .tielo(net101));
tielo I18 ( .tielo(net102));
bram_4k_sr I12 ( .bm_dm({bm_sdo, bm_dm[14:0]}), .rst(net102),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM({bm_sdo, bm_dm[14:0]}), .WEBM(bm_sweb), .WEB(web),
     .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]), .CLKW(net81),
     .CLKR(net79), .BWEBM({net101, net101, net101, net101, net101,
     net101, net101, net101, net101, net101, net101, net101, net101,
     net101, net101, net101}), .BWEB(bm_bweb[15:0]), .BIST(bm_init),
     .AMB(bm_sa[7:0]), .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]),
     .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net97), .out(net79));
bram_bufferx6 I8 ( .in(net93), .out(net81));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net93), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net97), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - leafcell, Cell - bram_4kbank_pbuffer_bot, View - schematic
// LAST TIME SAVED: Aug 24 17:32:39 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdi_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sdo_o;
output [7:0]  bm_sa_o;

input [15:0]  bm_d;
input [15:0]  bm_bweb;
input [1:0]  bm_sweb_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [1:0]  bm_sclkrw_i;
input [7:0]  bm_sa_i;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbank, View - schematic
// LAST TIME SAVED: Mar  6 12:03:12 2008
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4kprouting_bbank ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_bot;
output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_top;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;

inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [41:0]  bl;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_h_r_top;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_r_bot;
inout [23:0]  sp12_h_r_top;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_v_b_top;

input [7:0]  rgt_op_top;
input [1:0]  bm_sclkrw_i;
input [7:0]  bnl_op_top;
input [1:0]  bm_sweb_i;
input [7:0]  bot_op_bot;
input [7:0]  bnr_op_bot;
input [7:0]  rgt_op_bot;
input [1:0]  bm_sdo_i;
input [7:0]  glb_netwk;
input [7:0]  tnr_op_top;
input [15:0]  reset_b_top;
input [1:0]  bm_sdi_i;
input [15:0]  vdd_cntl_top;
input [7:0]  tnl_op_bot;
input [7:0]  bnl_op_bot;
input [15:0]  vdd_cntl_bot;
input [15:0]  wl_bot;
input [15:0]  pgate_bot;
input [7:0]  tnl_op_top;
input [15:0]  reset_b_bot;
input [7:0]  bm_sa_i;
input [7:0]  top_op_top;
input [15:0]  pgate_top;
input [15:0]  wl_top;
input [7:0]  bnr_op_top;
input [7:0]  lft_op_bot;
input [7:0]  tnr_op_bot;
input [7:0]  lft_op_top;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net260;

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net258;

wire  [0:7]  net261;

wire  [0:7]  net259;

wire  [0:7]  net228;

wire  [0:7]  net227;

wire  [0:7]  net322;

wire  [0:7]  net226;

wire  [0:7]  net343;

wire  [0:7]  net229;



bram_routing_tracks4rev I_bot ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}), .s_r(net210),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(tnr_op_bot[7:0]),
     .tnl_op(tnl_op_bot[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net303),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net226[0:7]),
     .lc_trk_g2(net227[0:7]), .lc_trk_g1(net228[0:7]),
     .lc_trk_g0(net229[0:7]), .clk(net230),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev I_top ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}), .s_r(net242),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net302),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net258[0:7]),
     .lc_trk_g2(net259[0:7]), .lc_trk_g1(net260[0:7]),
     .lc_trk_g0(net261[0:7]), .clk(net262),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbank_pbuffer_bot I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net242), .bm_wen(net210),
     .bm_d(bm_d[15:0]), .bm_clkr(net262), .bm_clkw(net230),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_ab(net343[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net322[0:7]),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
tielo I14 ( .tielo(net302));
tielo I15 ( .tielo(net303));
bram_4k_inmux_8x4 I6 ( .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15],
     vdd_cntl_bot[12], vdd_cntl_bot[13], vdd_cntl_bot[10],
     vdd_cntl_bot[11], vdd_cntl_bot[8], vdd_cntl_bot[9],
     vdd_cntl_bot[6], vdd_cntl_bot[7], vdd_cntl_bot[4],
     vdd_cntl_bot[5], vdd_cntl_bot[2], vdd_cntl_bot[3],
     vdd_cntl_bot[0], vdd_cntl_bot[1]}), .bl(bl[41:26]),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net226[0:7]), .lc_trk_g2(net227[0:7]),
     .lc_trk_g1(net228[0:7]), .lc_trk_g0(net229[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net322[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15],
     vdd_cntl_top[12], vdd_cntl_top[13], vdd_cntl_top[10],
     vdd_cntl_top[11], vdd_cntl_top[8], vdd_cntl_top[9],
     vdd_cntl_top[6], vdd_cntl_top[7], vdd_cntl_top[4],
     vdd_cntl_top[5], vdd_cntl_top[2], vdd_cntl_top[3],
     vdd_cntl_top[0], vdd_cntl_top[1]}), .bl(bl[41:26]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}), .op(slf_op_top[7:0]),
     .lc_trk_g3(net258[0:7]), .lc_trk_g2(net259[0:7]),
     .lc_trk_g1(net260[0:7]), .lc_trk_g0(net261[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net343[0:7]));

endmodule
// Library - leafcell, Cell - bram_4k_sr_bankin, View - schematic
// LAST TIME SAVED: Aug 15 18:05:22 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_sr_bankin ( bm_dm, bm_sweb, clk, rcapmux_en, rst, bm_q,
     bm_sdi, wdummymux_en );

inout  bm_sweb, clk, rcapmux_en, rst;

input  bm_sdi, wdummymux_en;

output [15:0]  bm_dm;

input [15:0]  bm_q;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_dff_mux I0 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[14]), .bm_q(bm_q[15]), .q(bm_dm[15]));
bram_dff_mux I16 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[13]), .bm_q(bm_q[14]), .q(bm_dm[14]));
bram_dff_mux I15 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[12]), .bm_q(bm_q[13]), .q(bm_dm[13]));
bram_dff_mux I14 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[11]), .bm_q(bm_q[12]), .q(bm_dm[12]));
bram_dff_mux I13 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[10]), .bm_q(bm_q[11]), .q(bm_dm[11]));
bram_dff_mux I12 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[9]), .bm_q(bm_q[10]), .q(bm_dm[10]));
bram_dff_mux I11 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[8]), .bm_q(bm_q[9]), .q(bm_dm[9]));
bram_dff_mux I10 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[7]), .bm_q(bm_q[8]), .q(bm_dm[8]));
bram_dff_mux I9 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[6]), .bm_q(bm_q[7]), .q(bm_dm[7]));
bram_dff_mux I8 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[5]), .bm_q(bm_q[6]), .q(bm_dm[6]));
bram_dff_mux I7 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[4]), .bm_q(bm_q[5]), .q(bm_dm[5]));
bram_dff_mux I6 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[3]), .bm_q(bm_q[4]), .q(bm_dm[4]));
bram_dff_mux I5 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[2]), .bm_q(bm_q[3]), .q(bm_dm[3]));
bram_dff_mux I4 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_dm[1]), .bm_q(bm_q[2]), .q(bm_dm[2]));
bram_dff_mux I3 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(net150), .bm_q(bm_q[1]), .q(bm_dm[1]));
bram_dff_mux I2 ( .rst(rst), .ce(bm_sweb), .rcapmux_en(rcapmux_en),
     .clk(clk), .bm_sdi(bm_sdi), .bm_q(bm_q[0]), .q(bm_dm[0]));
ml_mux2_hvt_schematic I20 ( .in1(wdummy_reg), .in0(bm_dm[0]),
     .out(net150), .sel(wdummymux_en));
leafcell_ml_dff_schematic I19 ( .R(rst), .D(bm_sdi), .CLK(clk),
     .QN(net157), .Q(wdummy_reg));

endmodule
// Library - leafcell, Cell - bram_4k_bankin, View - schematic
// LAST TIME SAVED: Aug 15 18:08:05 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4k_bankin ( bm_q, bm_sdo, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init, bm_rcapmux_en, bm_ren, bm_sa, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen );
output  bm_sdo;

input  bm_clkr, bm_clkw, bm_init, bm_rcapmux_en, bm_ren, bm_sclk,
     bm_sclkrw, bm_sdi, bm_sreb, bm_sweb, bm_wdummymux_en, bm_wen;

output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_ab;
input [7:0]  bm_sa;
input [7:0]  bm_aa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [15:0]  q;

wire  [14:0]  bm_dm;



tielo I15 ( .tielo(net102));
tielo I18 ( .tielo(net103));
bram_4k_sr_bankin I12 ( .bm_dm({bm_sdo, bm_dm[14:0]}), .rst(net103),
     .bm_sweb(bm_sweb), .rcapmux_en(bm_rcapmux_en),
     .wdummymux_en(bm_wdummymux_en), .clk(bm_sclk), .bm_sdi(bm_sdi),
     .bm_q(bm_q[15:0]));
bram_bufferx16 I17_15_ ( .in(q[15]), .out(bm_q[15]));
bram_bufferx16 I17_14_ ( .in(q[14]), .out(bm_q[14]));
bram_bufferx16 I17_13_ ( .in(q[13]), .out(bm_q[13]));
bram_bufferx16 I17_12_ ( .in(q[12]), .out(bm_q[12]));
bram_bufferx16 I17_11_ ( .in(q[11]), .out(bm_q[11]));
bram_bufferx16 I17_10_ ( .in(q[10]), .out(bm_q[10]));
bram_bufferx16 I17_9_ ( .in(q[9]), .out(bm_q[9]));
bram_bufferx16 I17_8_ ( .in(q[8]), .out(bm_q[8]));
bram_bufferx16 I17_7_ ( .in(q[7]), .out(bm_q[7]));
bram_bufferx16 I17_6_ ( .in(q[6]), .out(bm_q[6]));
bram_bufferx16 I17_5_ ( .in(q[5]), .out(bm_q[5]));
bram_bufferx16 I17_4_ ( .in(q[4]), .out(bm_q[4]));
bram_bufferx16 I17_3_ ( .in(q[3]), .out(bm_q[3]));
bram_bufferx16 I17_2_ ( .in(q[2]), .out(bm_q[2]));
bram_bufferx16 I17_1_ ( .in(q[1]), .out(bm_q[1]));
bram_bufferx16 I17_0_ ( .in(q[0]), .out(bm_q[0]));
rf_4k I0 ( .DM({bm_sdo, bm_dm[14:0]}), .WEBM(bm_sweb), .WEB(web),
     .REBM(bm_sreb), .REB(reb), .D(bm_d[15:0]), .CLKW(net82),
     .CLKR(net80), .BWEBM({net102, net102, net102, net102, net102,
     net102, net102, net102, net102, net102, net102, net102, net102,
     net102, net102, net102}), .BWEB(bm_bweb[15:0]), .BIST(bm_init),
     .AMB(bm_sa[7:0]), .AMA(bm_sa[7:0]), .AB(bm_ab[7:0]),
     .AA(bm_aa[7:0]), .Q(q[15:0]));
bram_bufferx6 I9 ( .in(net98), .out(net80));
bram_bufferx6 I8 ( .in(net94), .out(net82));
ml_mux2_hvt_schematic I11 ( .in1(bm_sclkrw), .in0(bm_clkw),
     .out(net94), .sel(bm_init));
ml_mux2_hvt_schematic I10 ( .in1(bm_sclkrw), .in0(bm_clkr),
     .out(net98), .sel(bm_init));
inv_hvt I6 ( .A(bm_ren), .Y(reb));
inv_hvt I5 ( .A(bm_wen), .Y(web));

endmodule
// Library - leafcell, Cell - bram_4kbankin_pbuffer_bot, View -
//schematic
// LAST TIME SAVED: Aug 24 17:33:35 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4kbankin_pbuffer_bot ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sreb_i, bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sclkrw_o;

input [7:0]  bm_aa;
input [15:0]  bm_bweb;
input [7:0]  bm_sa_i;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sclkrw_i;
input [1:0]  bm_sdo_i;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [1:0]  bm_sweb_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx6 I18 ( .in(bm_sclkrw_i[1]), .out(bm_sclkrw_o[1]));
bram_bufferx6 I20 ( .in(bm_sweb_i[1]), .out(bm_sweb_o[1]));
bram_bufferx6 I17 ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx6 I16 ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o[0]), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i[0]), .bm_sclkrw_o(bm_sclkrw_o[0]),
     .bm_sdi_o(bm_sdi_o[0]), .bm_sdi_i(bm_sdi_i[0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i[0]),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o[0]), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankin I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o[0]), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i[0]),
     .bm_sclkrw(bm_sclkrw_o[0]), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4kprouting_bbankin, View - schematic
// LAST TIME SAVED: Mar  6 11:28:14 2008
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module bram_4kprouting_bbankin ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [1:0]  bm_sdi_o;
output [7:0]  bm_sa_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_top;
output [7:0]  slf_op_bot;
output [1:0]  bm_sclkrw_o;

inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_h_l_top;
inout [23:0]  sp12_h_r_bot;
inout [41:0]  bl;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_v_b_top;
inout [23:0]  sp12_h_r_top;

input [7:0]  glb_netwk;
input [7:0]  tnr_op_top;
input [7:0]  bnl_op_top;
input [1:0]  bm_sdi_i;
input [7:0]  bnr_op_bot;
input [7:0]  tnl_op_bot;
input [1:0]  bm_sclkrw_i;
input [7:0]  top_op_top;
input [7:0]  tnr_op_bot;
input [7:0]  bnr_op_top;
input [7:0]  lft_op_bot;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_top;
input [15:0]  reset_b_top;
input [15:0]  pgate_top;
input [7:0]  bot_op_bot;
input [7:0]  lft_op_top;
input [1:0]  bm_sweb_i;
input [7:0]  bnl_op_bot;
input [15:0]  vdd_cntl_top;
input [15:0]  wl_top;
input [1:0]  bm_sdo_i;
input [15:0]  pgate_bot;
input [15:0]  vdd_cntl_bot;
input [7:0]  rgt_op_bot;
input [15:0]  wl_bot;
input [15:0]  reset_b_bot;
input [7:0]  rgt_op_top;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net254;

wire  [0:7]  net285;

wire  [0:7]  net284;

wire  [0:7]  net253;

wire  [7:0]  in2_top;

wire  [0:7]  net283;

wire  [0:7]  net252;

wire  [0:7]  net341;

wire  [0:7]  net286;

wire  [0:7]  net320;

wire  [15:0]  bm_bweb;

wire  [0:7]  net251;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;

wire  [23:0]  sp12_v_b_top;



bram_routing_tracks4rev I_bot ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}), .s_r(net234),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(tnr_op_bot[7:0]),
     .tnl_op(tnl_op_bot[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net299),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net251[0:7]),
     .lc_trk_g2(net252[0:7]), .lc_trk_g1(net253[0:7]),
     .lc_trk_g0(net254[0:7]), .clk(net255),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev I_top ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}), .s_r(net266),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net298),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net283[0:7]),
     .lc_trk_g2(net284[0:7]), .lc_trk_g1(net285[0:7]),
     .lc_trk_g0(net286[0:7]), .clk(net287),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbankin_pbuffer_bot I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdi_o(bm_sdi_o[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sclkrw_o(bm_sclkrw_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net266), .bm_wen(net234),
     .bm_d(bm_d[15:0]), .bm_clkr(net287), .bm_clkw(net255),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_ab(net341[0:7]), .bm_sa_i(bm_sa_i[7:0]),
     .bm_sclk_i(bm_sclk_i), .bm_sreb_i(bm_sreb_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net320[0:7]),
     .bm_init_o(bm_init_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_sclk_o(bm_sclk_o), .bm_sreb_o(bm_sreb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15],
     vdd_cntl_bot[12], vdd_cntl_bot[13], vdd_cntl_bot[10],
     vdd_cntl_bot[11], vdd_cntl_bot[8], vdd_cntl_bot[9],
     vdd_cntl_bot[6], vdd_cntl_bot[7], vdd_cntl_bot[4],
     vdd_cntl_bot[5], vdd_cntl_bot[2], vdd_cntl_bot[3],
     vdd_cntl_bot[0], vdd_cntl_bot[1]}), .bl(bl[41:26]),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net251[0:7]), .lc_trk_g2(net252[0:7]),
     .lc_trk_g1(net253[0:7]), .lc_trk_g0(net254[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net320[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15],
     vdd_cntl_top[12], vdd_cntl_top[13], vdd_cntl_top[10],
     vdd_cntl_top[11], vdd_cntl_top[8], vdd_cntl_top[9],
     vdd_cntl_top[6], vdd_cntl_top[7], vdd_cntl_top[4],
     vdd_cntl_top[5], vdd_cntl_top[2], vdd_cntl_top[3],
     vdd_cntl_top[0], vdd_cntl_top[1]}), .bl(bl[41:26]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}), .op(slf_op_top[7:0]),
     .lc_trk_g3(net283[0:7]), .lc_trk_g2(net284[0:7]),
     .lc_trk_g1(net285[0:7]), .lc_trk_g0(net286[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net341[0:7]));
tielo I14 ( .tielo(net298));
tielo I15 ( .tielo(net299));

endmodule
// Library - leafcell, Cell - array_BRAM_1x8bot, View - schematic
// LAST TIME SAVED: Jan 23 13:25:16 2008
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module array_BRAM_1x8bot ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, glb_netwk, slf_op_01, slf_op_02, slf_op_03,
     slf_op_04, slf_op_05, slf_op_06, slf_op_07, slf_op_08, slf_op_09,
     slf_op_10, slf_op_11, slf_op_12, slf_op_13, slf_op_14, slf_op_15,
     slf_op_16, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02, sp4_h_l_03,
     sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07, sp4_h_l_08,
     sp4_h_l_09, sp4_h_l_10, sp4_h_l_11, sp4_h_l_12, sp4_h_l_13,
     sp4_h_l_14, sp4_h_l_15, sp4_h_l_16, sp4_h_r_01, sp4_h_r_02,
     sp4_h_r_03, sp4_h_r_04, sp4_h_r_05, sp4_h_r_06, sp4_h_r_07,
     sp4_h_r_08, sp4_h_r_09, sp4_h_r_10, sp4_h_r_11, sp4_h_r_12,
     sp4_h_r_13, sp4_h_r_14, sp4_h_r_15, sp4_h_r_16, sp4_r_v_b_01,
     sp4_r_v_b_02, sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05,
     sp4_r_v_b_06, sp4_r_v_b_07, sp4_r_v_b_08, sp4_r_v_b_09,
     sp4_r_v_b_10, sp4_r_v_b_11, sp4_r_v_b_12, sp4_r_v_b_13,
     sp4_r_v_b_14, sp4_r_v_b_15, sp4_r_v_b_16, sp4_v_b_01, sp4_v_b_02,
     sp4_v_b_03, sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07,
     sp4_v_b_08, sp4_v_b_09, sp4_v_b_10, sp4_v_b_11, sp4_v_b_12,
     sp4_v_b_13, sp4_v_b_14, sp4_v_b_15, sp4_v_b_16, sp4_v_t_16,
     sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04, sp12_h_l_05,
     sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_l_09, sp12_h_l_10,
     sp12_h_l_11, sp12_h_l_12, sp12_h_l_13, sp12_h_l_14, sp12_h_l_15,
     sp12_h_l_16, sp12_h_r_01, sp12_h_r_02, sp12_h_r_03, sp12_h_r_04,
     sp12_h_r_05, sp12_h_r_06, sp12_h_r_07, sp12_h_r_08, sp12_h_r_09,
     sp12_h_r_10, sp12_h_r_11, sp12_h_r_12, sp12_h_r_13, sp12_h_r_14,
     sp12_h_r_15, sp12_h_r_16, sp12_v_b_01, sp12_v_t_16, vdd_cntl, wl,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i,
     bnl_op_01, bnr_op_01, bot_op_01, glb_netwk_col, lft_op_01,
     lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06, lft_op_07,
     lft_op_08, lft_op_09, lft_op_10, lft_op_11, lft_op_12, lft_op_13,
     lft_op_14, lft_op_15, lft_op_16, prog, rgt_op_01, rgt_op_02,
     rgt_op_03, rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08,
     rgt_op_09, rgt_op_10, rgt_op_11, rgt_op_12, rgt_op_13, rgt_op_14,
     rgt_op_15, rgt_op_16, tnl_op_16, tnr_op_16, top_op_16 );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, prog;

output [7:0]  slf_op_03;
output [7:0]  slf_op_16;
output [7:0]  slf_op_12;
output [7:0]  slf_op_15;
output [7:0]  slf_op_02;
output [7:0]  slf_op_08;
output [1:0]  bm_sclkrw_o;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_01;
output [7:0]  slf_op_04;
output [7:0]  slf_op_14;
output [7:0]  slf_op_11;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_10;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_09;
output [7:0]  slf_op_05;
output [1:0]  bm_sweb_o;
output [7:0]  slf_op_07;
output [7:0]  glb_netwk;
output [7:0]  slf_op_13;
output [7:0]  slf_op_06;

inout [47:0]  sp4_h_r_13;
inout [23:0]  sp12_h_r_12;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_h_r_15;
inout [47:0]  sp4_h_l_14;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_h_r_04;
inout [23:0]  sp12_h_l_11;
inout [47:0]  sp4_h_l_15;
inout [47:0]  sp4_r_v_b_08;
inout [23:0]  sp12_h_l_03;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_h_r_08;
inout [47:0]  sp4_h_r_11;
inout [47:0]  sp4_v_b_06;
inout [47:0]  sp4_h_l_12;
inout [47:0]  sp4_r_v_b_15;
inout [23:0]  sp12_v_b_01;
inout [47:0]  sp4_r_v_b_16;
inout [47:0]  sp4_v_b_11;
inout [47:0]  sp4_h_r_16;
inout [23:0]  sp12_h_l_16;
inout [23:0]  sp12_h_r_08;
inout [23:0]  sp12_h_r_10;
inout [47:0]  sp4_h_l_13;
inout [47:0]  sp4_r_v_b_11;
inout [23:0]  sp12_h_r_09;
inout [23:0]  sp12_h_l_12;
inout [47:0]  sp4_r_v_b_12;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_02;
inout [23:0]  sp12_h_l_01;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_v_t_16;
inout [23:0]  sp12_h_l_10;
inout [23:0]  sp12_h_r_14;
inout [47:0]  sp4_v_b_14;
inout [47:0]  sp4_r_v_b_14;
inout [23:0]  sp12_h_l_05;
inout [47:0]  sp4_v_b_10;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_h_l_16;
inout [47:0]  sp4_r_v_b_03;
inout [47:0]  sp4_v_b_13;
inout [47:0]  sp4_h_l_11;
inout [23:0]  sp12_h_r_15;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_r_v_b_13;
inout [23:0]  sp12_h_r_11;
inout [47:0]  sp4_v_b_04;
inout [23:0]  sp12_h_l_15;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_r_10;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_v_b_15;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_h_l_09;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_v_b_03;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_h_l_04;
inout [47:0]  sp4_h_r_14;
inout [23:0]  sp12_h_r_01;
inout [23:0]  sp12_v_t_16;
inout [47:0]  sp4_h_l_10;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_h_r_12;
inout [47:0]  sp4_v_b_16;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_h_l_03;
inout [47:0]  sp4_v_b_09;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_h_r_16;
inout [23:0]  sp12_h_r_13;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_r_v_b_09;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_v_b_12;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_h_l_02;
inout [47:0]  sp4_r_v_b_05;
inout [23:0]  sp12_h_l_13;
inout [47:0]  sp4_h_l_01;
inout [23:0]  sp12_h_l_09;
inout [47:0]  sp4_h_r_09;
inout [41:0]  bl;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_h_l_08;
inout [47:0]  sp4_v_b_05;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_r_v_b_10;
inout [271:16]  pgate;
inout [271:16]  reset_b;
inout [271:16]  wl;
inout [271:16]  vdd_cntl;
inout [47:0]  sp4_h_l_06;
inout [23:0]  sp12_h_l_14;
inout [47:0]  sp4_r_v_b_04;

input [7:0]  lft_op_15;
input [7:0]  lft_op_08;
input [7:0]  rgt_op_15;
input [7:0]  glb_netwk_col;
input [1:0]  bm_sdi_i;
input [1:0]  bm_sweb_i;
input [7:0]  lft_op_11;
input [7:0]  rgt_op_04;
input [1:0]  bm_sdo_i;
input [7:0]  rgt_op_12;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_09;
input [7:0]  lft_op_04;
input [7:0]  tnl_op_16;
input [7:0]  rgt_op_13;
input [7:0]  lft_op_16;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_02;
input [7:0]  lft_op_09;
input [7:0]  lft_op_02;
input [7:0]  rgt_op_05;
input [7:0]  lft_op_06;
input [7:0]  top_op_16;
input [1:0]  bm_sclkrw_i;
input [7:0]  lft_op_07;
input [7:0]  bnl_op_01;
input [7:0]  lft_op_01;
input [7:0]  rgt_op_10;
input [7:0]  lft_op_10;
input [7:0]  rgt_op_08;
input [7:0]  rgt_op_16;
input [7:0]  tnr_op_16;
input [7:0]  lft_op_14;
input [7:0]  rgt_op_14;
input [7:0]  rgt_op_03;
input [7:0]  lft_op_05;
input [7:0]  lft_op_13;
input [7:0]  rgt_op_11;
input [7:0]  lft_op_03;
input [7:0]  rgt_op_06;
input [7:0]  bot_op_01;
input [7:0]  lft_op_12;
input [7:0]  bnr_op_01;
input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net955;

wire  [0:7]  net944;

wire  [0:1]  net769;

wire  [0:1]  net647;

wire  [0:1]  net1014;

wire  [0:1]  net895;

wire  [0:23]  net924;

wire  [0:1]  net889;

wire  [0:1]  net707;

wire  [0:1]  net890;

wire  [0:1]  net951;

wire  [0:1]  net1013;

wire  [0:7]  net694;

wire  [0:23]  net1043;

wire  [0:1]  net709;

wire  [0:23]  net862;

wire  [0:1]  net957;

wire  [0:23]  net795;

wire  [0:1]  net827;

wire  [0:1]  net641;

wire  [0:23]  net671;

wire  [0:1]  net771;

wire  [0:1]  net1017;

wire  [0:7]  net1006;

wire  [0:1]  net952;

wire  [0:7]  net882;

wire  [0:1]  net1019;

wire  [0:23]  net986;

wire  [0:1]  net828;

wire  [0:1]  net765;

wire  [0:1]  net704;

wire  [0:7]  net821;

wire  [0:1]  net703;

wire  [0:1]  net766;

wire  [0:23]  net733;

wire  [0:1]  net645;

wire  [0:1]  net642;

wire  [0:7]  net759;

wire  [0:1]  net893;

wire  [0:1]  net831;

wire  [0:7]  net1069;

wire  [0:1]  net833;



clk_colbuf8kx8 I107 ( .clko(glb_netwk[7:0]),
     .clki(glb_netwk_col[7:0]));
bram_4kprouting_bbankout I_bram_out_0825_02 ( .bm_sdi_o(net1013[0:1]),
     .bm_sclkrw_o(net1014[0:1]), .bm_sclkrw_i(bm_sclkrw_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sweb_o(net1017[0:1]),
     .bm_sdi_i(bm_sdi_i[1:0]), .bm_sdo_i(net1019[0:1]),
     .bm_sdo_o(bm_sdo_o[1:0]), .slf_op_top(slf_op_02[7:0]),
     .slf_op_bot(slf_op_01[7:0]), .wl_top(wl[47:32]),
     .wl_bot(wl[31:16]), .top_op_top(slf_op_03[7:0]),
     .tnl_op_top(lft_op_03[7:0]), .tnl_op_bot(lft_op_02[7:0]),
     .reset_b_top(reset_b[47:32]), .reset_b_bot(reset_b[31:16]),
     .prog(prog), .pgate_top(pgate[47:32]), .pgate_bot(pgate[31:16]),
     .lft_op_top(lft_op_02[7:0]), .lft_op_bot(lft_op_01[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_01[7:0]), .sp4_h_r_top(sp4_h_r_02[47:0]),
     .bnl_op_top(lft_op_01[7:0]), .bnl_op_bot(bnl_op_01[7:0]),
     .bnr_op_bot(bnr_op_01[7:0]), .sp4_h_r_bot(sp4_h_r_01[47:0]),
     .sp12_v_t_top(net1043[0:23]), .sp12_v_b_bot(sp12_v_b_01[23:0]),
     .bm_init_i(bm_init_i), .sp12_h_l_top(sp12_h_l_02[23:0]),
     .sp12_h_r_bot(sp12_h_r_01[23:0]),
     .sp12_h_l_bot(sp12_h_l_01[23:0]),
     .sp12_h_r_top(sp12_h_r_02[23:0]), .sp4_v_t_top(sp4_v_b_03[47:0]),
     .sp4_v_b_top(sp4_v_b_02[47:0]), .sp4_v_b_bot(sp4_v_b_01[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_01[47:0]),
     .sp4_h_l_top(sp4_h_l_02[47:0]), .tnr_op_top(rgt_op_03[7:0]),
     .sp4_h_l_bot(sp4_h_l_01[47:0]), .tnr_op_bot(rgt_op_02[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .sp4_r_v_b_top(sp4_r_v_b_02[47:0]), .rgt_op_bot(rgt_op_01[7:0]),
     .rgt_op_top(rgt_op_02[7:0]), .bnr_op_top(rgt_op_01[7:0]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(net1067),
     .bm_init_o(net1068), .bm_sa_o(net1069[0:7]), .bm_sclk_o(net1070),
     .bm_sreb_o(net1071), .bm_wdummymux_en_o(net1072),
     .vdd_cntl_top(vdd_cntl[47:32]), .vdd_cntl_bot(vdd_cntl[31:16]));
bram_4kprouting_bbank I_bram_0825_08 ( .bm_sdi_o(net641[0:1]),
     .bm_sclkrw_o(net642[0:1]), .bm_sclkrw_i(net704[0:1]),
     .bm_sweb_i(net707[0:1]), .bm_sweb_o(net645[0:1]),
     .bm_sdi_i(net703[0:1]), .bm_sdo_i(net647[0:1]),
     .bm_sdo_o(net709[0:1]), .slf_op_top(slf_op_08[7:0]),
     .slf_op_bot(slf_op_07[7:0]), .wl_bot(wl[127:112]),
     .top_op_top(slf_op_09[7:0]), .sp12_h_l_bot(sp12_h_l_07[23:0]),
     .sp4_h_l_bot(sp4_h_l_07[47:0]), .tnl_op_top(lft_op_09[7:0]),
     .tnl_op_bot(lft_op_08[7:0]), .reset_b_top(reset_b[143:128]),
     .reset_b_bot(reset_b[127:112]), .vdd_cntl_top(vdd_cntl[143:128]),
     .prog(prog), .pgate_top(pgate[143:128]),
     .pgate_bot(pgate[127:112]), .lft_op_bot(lft_op_07[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(net762),
     .bot_op_bot(slf_op_06[7:0]), .rgt_op_bot(rgt_op_07[7:0]),
     .bnl_op_top(lft_op_07[7:0]), .bnl_op_bot(lft_op_06[7:0]),
     .sp4_h_r_top(sp4_h_r_08[47:0]), .sp12_v_t_top(net671[0:23]),
     .sp12_v_b_bot(net733[0:23]), .bm_init_i(net758),
     .sp4_h_r_bot(sp4_h_r_07[47:0]), .sp12_h_r_bot(sp12_h_r_07[23:0]),
     .sp4_v_t_top(sp4_v_b_09[47:0]), .sp4_v_b_bot(sp4_v_b_07[47:0]),
     .sp12_h_r_top(sp12_h_r_08[23:0]), .tnr_op_bot(rgt_op_08[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net757),
     .sp4_h_l_top(sp4_h_l_08[47:0]), .lft_op_top(lft_op_08[7:0]),
     .wl_top(wl[143:128]), .sp12_h_l_top(sp12_h_l_08[23:0]),
     .sp4_v_b_top(sp4_v_b_08[47:0]), .tnr_op_top(rgt_op_09[7:0]),
     .rgt_op_top(rgt_op_08[7:0]), .bm_sa_i(net759[0:7]),
     .bm_sclk_i(net760), .bm_sreb_i(net761), .bm_rcapmux_en_o(net692),
     .bm_init_o(net693), .bm_sa_o(net694[0:7]), .bm_sclk_o(net695),
     .bm_sreb_o(net696), .bm_wdummymux_en_o(net697),
     .vdd_cntl_bot(vdd_cntl[127:112]), .bnr_op_bot(rgt_op_06[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_07[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_08[47:0]), .bnr_op_top(rgt_op_07[7:0]));
bram_4kprouting_bbank I_bram_0825_06 ( .bm_sdi_o(net703[0:1]),
     .bm_sclkrw_o(net704[0:1]), .bm_sclkrw_i(net766[0:1]),
     .bm_sweb_i(net769[0:1]), .bm_sweb_o(net707[0:1]),
     .bm_sdi_i(net765[0:1]), .bm_sdo_i(net709[0:1]),
     .bm_sdo_o(net771[0:1]), .slf_op_top(slf_op_06[7:0]),
     .slf_op_bot(slf_op_05[7:0]), .wl_top(wl[111:96]),
     .wl_bot(wl[95:80]), .top_op_top(slf_op_07[7:0]),
     .tnl_op_top(lft_op_07[7:0]), .tnl_op_bot(lft_op_06[7:0]),
     .reset_b_top(reset_b[111:96]), .reset_b_bot(reset_b[95:80]),
     .prog(prog), .pgate_top(pgate[111:96]), .pgate_bot(pgate[95:80]),
     .lft_op_top(lft_op_06[7:0]), .lft_op_bot(lft_op_05[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(net824),
     .bot_op_bot(slf_op_04[7:0]), .sp4_h_r_top(sp4_h_r_06[47:0]),
     .bnl_op_top(lft_op_05[7:0]), .bnl_op_bot(lft_op_04[7:0]),
     .bnr_op_bot(rgt_op_04[7:0]), .sp4_h_r_bot(sp4_h_r_05[47:0]),
     .sp12_v_t_top(net733[0:23]), .sp12_v_b_bot(net795[0:23]),
     .bm_init_i(net820), .sp12_h_l_top(sp12_h_l_06[23:0]),
     .sp12_h_r_bot(sp12_h_r_05[23:0]),
     .sp12_h_l_bot(sp12_h_l_05[23:0]),
     .sp12_h_r_top(sp12_h_r_06[23:0]), .sp4_v_t_top(sp4_v_b_07[47:0]),
     .sp4_v_b_top(sp4_v_b_06[47:0]), .sp4_v_b_bot(sp4_v_b_05[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_05[47:0]),
     .sp4_h_l_top(sp4_h_l_06[47:0]), .tnr_op_top(rgt_op_07[7:0]),
     .sp4_h_l_bot(sp4_h_l_05[47:0]), .tnr_op_bot(rgt_op_06[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net819),
     .sp4_r_v_b_top(sp4_r_v_b_06[47:0]), .rgt_op_bot(rgt_op_05[7:0]),
     .rgt_op_top(rgt_op_06[7:0]), .bnr_op_top(rgt_op_05[7:0]),
     .bm_sa_i(net821[0:7]), .bm_sclk_i(net822), .bm_sreb_i(net823),
     .bm_rcapmux_en_o(net757), .bm_init_o(net758),
     .bm_sa_o(net759[0:7]), .bm_sclk_o(net760), .bm_sreb_o(net761),
     .bm_wdummymux_en_o(net762), .vdd_cntl_top(vdd_cntl[111:96]),
     .vdd_cntl_bot(vdd_cntl[95:80]));
bram_4kprouting_bbank I_bram_0825_04 ( .bm_sdi_o(net765[0:1]),
     .bm_sclkrw_o(net766[0:1]), .bm_sclkrw_i(net1014[0:1]),
     .bm_sweb_i(net1017[0:1]), .bm_sweb_o(net769[0:1]),
     .bm_sdi_i(net1013[0:1]), .bm_sdo_i(net771[0:1]),
     .bm_sdo_o(net1019[0:1]), .slf_op_top(slf_op_04[7:0]),
     .slf_op_bot(slf_op_03[7:0]), .wl_top(wl[79:64]),
     .wl_bot(wl[63:48]), .top_op_top(slf_op_05[7:0]),
     .tnl_op_top(lft_op_05[7:0]), .tnl_op_bot(lft_op_04[7:0]),
     .reset_b_top(reset_b[79:64]), .reset_b_bot(reset_b[63:48]),
     .prog(prog), .pgate_top(pgate[79:64]), .pgate_bot(pgate[63:48]),
     .lft_op_top(lft_op_04[7:0]), .lft_op_bot(lft_op_03[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(net1072),
     .bot_op_bot(slf_op_02[7:0]), .sp4_h_r_top(sp4_h_r_04[47:0]),
     .bnl_op_top(lft_op_03[7:0]), .bnl_op_bot(lft_op_02[7:0]),
     .bnr_op_bot(rgt_op_02[7:0]), .sp4_h_r_bot(sp4_h_r_03[47:0]),
     .sp12_v_t_top(net795[0:23]), .sp12_v_b_bot(net1043[0:23]),
     .bm_init_i(net1068), .sp12_h_l_top(sp12_h_l_04[23:0]),
     .sp12_h_r_bot(sp12_h_r_03[23:0]),
     .sp12_h_l_bot(sp12_h_l_03[23:0]),
     .sp12_h_r_top(sp12_h_r_04[23:0]), .sp4_v_t_top(sp4_v_b_05[47:0]),
     .sp4_v_b_top(sp4_v_b_04[47:0]), .sp4_v_b_bot(sp4_v_b_03[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_03[47:0]),
     .sp4_h_l_top(sp4_h_l_04[47:0]), .tnr_op_top(rgt_op_05[7:0]),
     .sp4_h_l_bot(sp4_h_l_03[47:0]), .tnr_op_bot(rgt_op_04[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net1067),
     .sp4_r_v_b_top(sp4_r_v_b_04[47:0]), .rgt_op_bot(rgt_op_03[7:0]),
     .rgt_op_top(rgt_op_04[7:0]), .bnr_op_top(rgt_op_03[7:0]),
     .bm_sa_i(net1069[0:7]), .bm_sclk_i(net1070), .bm_sreb_i(net1071),
     .bm_rcapmux_en_o(net819), .bm_init_o(net820),
     .bm_sa_o(net821[0:7]), .bm_sclk_o(net822), .bm_sreb_o(net823),
     .bm_wdummymux_en_o(net824), .vdd_cntl_top(vdd_cntl[79:64]),
     .vdd_cntl_bot(vdd_cntl[63:48]));
bram_4kprouting_bbank I_bram_0825_12 ( .bm_sdi_o(net827[0:1]),
     .bm_sclkrw_o(net828[0:1]), .bm_sclkrw_i(net890[0:1]),
     .bm_sweb_i(net893[0:1]), .bm_sweb_o(net831[0:1]),
     .bm_sdi_i(net889[0:1]), .bm_sdo_i(net833[0:1]),
     .bm_sdo_o(net895[0:1]), .slf_op_top(slf_op_12[7:0]),
     .sp4_h_l_bot(sp4_h_l_11[47:0]), .slf_op_bot(slf_op_11[7:0]),
     .sp4_r_v_b_top(sp4_r_v_b_12[47:0]),
     .reset_b_top(reset_b[207:192]), .tnl_op_top(lft_op_13[7:0]),
     .top_op_top(slf_op_13[7:0]), .rgt_op_bot(rgt_op_11[7:0]),
     .tnl_op_bot(lft_op_12[7:0]), .prog(prog),
     .lft_op_top(lft_op_12[7:0]), .lft_op_bot(lft_op_11[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bnl_op_top(lft_op_11[7:0]),
     .rgt_op_top(rgt_op_12[7:0]), .bnl_op_bot(lft_op_10[7:0]),
     .sp12_h_l_top(sp12_h_l_12[23:0]), .sp4_v_b_top(sp4_v_b_12[47:0]),
     .bl(bl[41:0]), .bm_wdummymux_en_i(net947),
     .bot_op_bot(slf_op_10[7:0]), .tnr_op_bot(rgt_op_12[7:0]),
     .bnr_op_bot(rgt_op_10[7:0]), .sp4_h_l_top(sp4_h_l_12[47:0]),
     .wl_bot(wl[191:176]), .sp4_r_v_b_bot(sp4_r_v_b_11[47:0]),
     .tnr_op_top(rgt_op_13[7:0]), .sp12_v_t_top(net862[0:23]),
     .sp12_v_b_bot(net924[0:23]), .bm_init_i(net943),
     .sp4_h_r_bot(sp4_h_r_11[47:0]), .pgate_top(pgate[207:192]),
     .sp12_h_r_bot(sp12_h_r_11[23:0]), .sp4_v_t_top(sp4_v_b_13[47:0]),
     .sp12_h_r_top(sp12_h_r_12[23:0]), .sp4_v_b_bot(sp4_v_b_11[47:0]),
     .bnr_op_top(rgt_op_11[7:0]), .reset_b_bot(reset_b[191:176]),
     .wl_top(wl[207:192]), .sp4_h_r_top(sp4_h_r_12[47:0]),
     .bm_rcapmux_en_i(net942), .pgate_bot(pgate[191:176]),
     .bm_sa_i(net944[0:7]), .bm_sclk_i(net945), .bm_sreb_i(net946),
     .bm_rcapmux_en_o(net880), .bm_init_o(net881),
     .bm_sa_o(net882[0:7]), .bm_sclk_o(net883), .bm_sreb_o(net884),
     .bm_wdummymux_en_o(net885), .vdd_cntl_bot(vdd_cntl[191:176]),
     .vdd_cntl_top(vdd_cntl[207:192]),
     .sp12_h_l_bot(sp12_h_l_11[23:0]));
bram_4kprouting_bbank I_bram_0825_10 ( .bm_sdi_o(net889[0:1]),
     .bm_sclkrw_o(net890[0:1]), .bm_sclkrw_i(net642[0:1]),
     .bm_sweb_i(net645[0:1]), .bm_sweb_o(net893[0:1]),
     .bm_sdi_i(net641[0:1]), .bm_sdo_i(net895[0:1]),
     .bm_sdo_o(net647[0:1]), .slf_op_top(slf_op_10[7:0]),
     .sp4_h_l_bot(sp4_h_l_09[47:0]), .slf_op_bot(slf_op_09[7:0]),
     .sp4_r_v_b_top(sp4_r_v_b_10[47:0]),
     .reset_b_top(reset_b[175:160]), .tnl_op_top(lft_op_11[7:0]),
     .top_op_top(slf_op_11[7:0]), .rgt_op_bot(rgt_op_09[7:0]),
     .tnl_op_bot(lft_op_10[7:0]), .prog(prog),
     .lft_op_top(lft_op_10[7:0]), .lft_op_bot(lft_op_09[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bnl_op_top(lft_op_09[7:0]),
     .rgt_op_top(rgt_op_10[7:0]), .bnl_op_bot(lft_op_08[7:0]),
     .sp12_h_l_top(sp12_h_l_10[23:0]), .sp4_v_b_top(sp4_v_b_10[47:0]),
     .bl(bl[41:0]), .bm_wdummymux_en_i(net697),
     .bot_op_bot(slf_op_08[7:0]), .tnr_op_bot(rgt_op_10[7:0]),
     .bnr_op_bot(rgt_op_08[7:0]), .sp4_h_l_top(sp4_h_l_10[47:0]),
     .wl_bot(wl[159:144]), .sp4_r_v_b_bot(sp4_r_v_b_09[47:0]),
     .tnr_op_top(rgt_op_11[7:0]), .sp12_v_t_top(net924[0:23]),
     .sp12_v_b_bot(net671[0:23]), .bm_init_i(net693),
     .sp4_h_r_bot(sp4_h_r_09[47:0]), .pgate_top(pgate[175:160]),
     .sp12_h_r_bot(sp12_h_r_09[23:0]), .sp4_v_t_top(sp4_v_b_11[47:0]),
     .sp12_h_r_top(sp12_h_r_10[23:0]), .sp4_v_b_bot(sp4_v_b_09[47:0]),
     .bnr_op_top(rgt_op_09[7:0]), .reset_b_bot(reset_b[159:144]),
     .wl_top(wl[175:160]), .sp4_h_r_top(sp4_h_r_10[47:0]),
     .bm_rcapmux_en_i(net692), .pgate_bot(pgate[159:144]),
     .bm_sa_i(net694[0:7]), .bm_sclk_i(net695), .bm_sreb_i(net696),
     .bm_rcapmux_en_o(net942), .bm_init_o(net943),
     .bm_sa_o(net944[0:7]), .bm_sclk_o(net945), .bm_sreb_o(net946),
     .bm_wdummymux_en_o(net947), .vdd_cntl_bot(vdd_cntl[159:144]),
     .vdd_cntl_top(vdd_cntl[175:160]),
     .sp12_h_l_bot(sp12_h_l_09[23:0]));
bram_4kprouting_bbank I_bram_0825_14 ( .bm_sdi_o(net951[0:1]),
     .bm_sclkrw_o(net952[0:1]), .bm_sclkrw_i(net828[0:1]),
     .bm_sweb_i(net831[0:1]), .bm_sweb_o(net955[0:1]),
     .bm_sdi_i(net827[0:1]), .bm_sdo_i(net957[0:1]),
     .bm_sdo_o(net833[0:1]), .slf_op_top(slf_op_14[7:0]),
     .sp4_h_l_bot(sp4_h_l_13[47:0]), .slf_op_bot(slf_op_13[7:0]),
     .sp4_r_v_b_top(sp4_r_v_b_14[47:0]),
     .reset_b_top(reset_b[239:224]), .tnl_op_top(lft_op_15[7:0]),
     .top_op_top(slf_op_15[7:0]), .rgt_op_bot(rgt_op_13[7:0]),
     .tnl_op_bot(lft_op_14[7:0]), .prog(prog),
     .lft_op_top(lft_op_14[7:0]), .lft_op_bot(lft_op_13[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bnl_op_top(lft_op_13[7:0]),
     .rgt_op_top(rgt_op_14[7:0]), .bnl_op_bot(lft_op_12[7:0]),
     .sp12_h_l_top(sp12_h_l_14[23:0]), .sp4_v_b_top(sp4_v_b_14[47:0]),
     .bl(bl[41:0]), .bm_wdummymux_en_i(net885),
     .bot_op_bot(slf_op_12[7:0]), .tnr_op_bot(rgt_op_14[7:0]),
     .bnr_op_bot(rgt_op_12[7:0]), .sp4_h_l_top(sp4_h_l_14[47:0]),
     .wl_bot(wl[223:208]), .sp4_r_v_b_bot(sp4_r_v_b_13[47:0]),
     .tnr_op_top(rgt_op_15[7:0]), .sp12_v_t_top(net986[0:23]),
     .sp12_v_b_bot(net862[0:23]), .bm_init_i(net881),
     .sp4_h_r_bot(sp4_h_r_13[47:0]), .pgate_top(pgate[239:224]),
     .sp12_h_r_bot(sp12_h_r_13[23:0]), .sp4_v_t_top(sp4_v_b_15[47:0]),
     .sp12_h_r_top(sp12_h_r_14[23:0]), .sp4_v_b_bot(sp4_v_b_13[47:0]),
     .bnr_op_top(rgt_op_13[7:0]), .reset_b_bot(reset_b[223:208]),
     .wl_top(wl[239:224]), .sp4_h_r_top(sp4_h_r_14[47:0]),
     .bm_rcapmux_en_i(net880), .pgate_bot(pgate[223:208]),
     .bm_sa_i(net882[0:7]), .bm_sclk_i(net883), .bm_sreb_i(net884),
     .bm_rcapmux_en_o(net1004), .bm_init_o(net1005),
     .bm_sa_o(net1006[0:7]), .bm_sclk_o(net1007), .bm_sreb_o(net1008),
     .bm_wdummymux_en_o(net1009), .vdd_cntl_bot(vdd_cntl[223:208]),
     .vdd_cntl_top(vdd_cntl[239:224]),
     .sp12_h_l_bot(sp12_h_l_13[23:0]));
bram_4kprouting_bbankin I_bram_in_0825_16 ( .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sclkrw_i(net952[0:1]),
     .bm_sweb_i(net955[0:1]), .bm_sweb_o(bm_sweb_o[1:0]),
     .bm_sdi_i(net951[0:1]), .bm_sdo_i(bm_sdo_i[1:0]),
     .bm_sdo_o(net957[0:1]), .slf_op_top(slf_op_16[7:0]),
     .slf_op_bot(slf_op_15[7:0]), .wl_bot(wl[255:240]),
     .top_op_top(top_op_16[7:0]), .sp12_h_l_bot(sp12_h_l_15[23:0]),
     .sp4_h_l_bot(sp4_h_l_15[47:0]), .tnl_op_top(tnl_op_16[7:0]),
     .tnl_op_bot(lft_op_16[7:0]), .reset_b_top(reset_b[271:256]),
     .reset_b_bot(reset_b[255:240]), .vdd_cntl_top(vdd_cntl[271:256]),
     .prog(prog), .pgate_top(pgate[271:256]),
     .pgate_bot(pgate[255:240]), .lft_op_bot(lft_op_15[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(net1009),
     .bot_op_bot(slf_op_14[7:0]), .rgt_op_bot(rgt_op_15[7:0]),
     .bnl_op_top(lft_op_15[7:0]), .bnl_op_bot(lft_op_14[7:0]),
     .sp4_h_r_top(sp4_h_r_16[47:0]), .sp12_v_t_top(sp12_v_t_16[23:0]),
     .sp12_v_b_bot(net986[0:23]), .bm_init_i(net1005),
     .sp4_h_r_bot(sp4_h_r_15[47:0]), .sp12_h_r_bot(sp12_h_r_15[23:0]),
     .sp4_v_t_top(sp4_v_t_16[47:0]), .sp4_v_b_bot(sp4_v_b_15[47:0]),
     .sp12_h_r_top(sp12_h_r_16[23:0]), .tnr_op_bot(rgt_op_16[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net1004),
     .sp4_h_l_top(sp4_h_l_16[47:0]), .lft_op_top(lft_op_16[7:0]),
     .wl_top(wl[271:256]), .sp12_h_l_top(sp12_h_l_16[23:0]),
     .sp4_v_b_top(sp4_v_b_16[47:0]), .tnr_op_top(tnr_op_16[7:0]),
     .rgt_op_top(rgt_op_16[7:0]), .bm_sa_i(net1006[0:7]),
     .bm_sclk_i(net1007), .bm_sreb_i(net1008),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .vdd_cntl_bot(vdd_cntl[255:240]), .bnr_op_bot(rgt_op_14[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_15[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_16[47:0]), .bnr_op_top(rgt_op_15[7:0]));

endmodule
// Library - io, Cell - io_odrv4x5, View - schematic
// LAST TIME SAVED: Aug 21 17:59:07 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module io_odrv4x5 ( cbit, sp4_out, bl, pgate, prog,
     reset, slfop, vdd_cntl, wl );


input  prog, slfop;

output [4:0]  sp4_out;
output [7:5]  cbit;

inout [3:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
supply1 vdd_;
supply0 gnd_;

// Buses in the design

wire  [7:0]  cbitb;

wire  [1:0]  r_vdd;

wire [7:0] cbit_int;
assign cbit[7:5] = cbit_int[7:5];

pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv4 I_odrv_4_ ( .cbitb(cbitb[4]), .sp4(sp4_out[4]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_3_ ( .cbitb(cbitb[3]), .sp4(sp4_out[3]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_2_ ( .cbitb(cbitb[2]), .sp4(sp4_out[2]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_1_ ( .cbitb(cbitb[1]), .sp4(sp4_out[1]), .slfop(slfop),
     .prog(prog));
odrv4 I_odrv_0_ ( .cbitb(cbitb[0]), .sp4(sp4_out[0]), .slfop(slfop),
     .prog(prog));
cram2x2 Icram2x2_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]),
     .reset(reset[1:0]), .q(cbit_int[7:4]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));
cram2x2 Icram2x2_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]),
     .reset(reset[1:0]), .q(cbit_int[3:0]), .wl(wl[1:0]),
     .r_vdd(r_vdd[1:0]), .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - io_col_odrv4_x40bare, View - schematic
// LAST TIME SAVED: Jul 31 17:45:40 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module io_col_odrv4_x40bare ( cf, bl, sp4_h_l,
     sp4_v_b, dout0, dout1,
     pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [23:0]  cf;

inout [3:0]  bl;
inout [15:0]  sp4_v_b;
inout [47:0]  sp4_h_l;

input [0:1]  dout0;
input [0:1]  dout1;
input [15:0]  pgate;
input [15:0]  wl;
input [15:0]  reset;
input [15:0]  vdd_cntl;
supply0 gnd_;
supply1 vdd_;



io_odrv4x5 I218 ( cf[20:18], {sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6]}, bl[3:0], pgate[13:12], prog,
     reset[13:12], dout1[1], vdd_cntl[13:12], wl[13:12]);
io_odrv4x5 I217 ( cf[14:12], {sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4]}, bl[3:0], pgate[9:8], prog, reset[9:8],
     dout0[1], vdd_cntl[9:8], wl[9:8]);
io_odrv4x5 I_odrv_4x5_7 ( cf[23:21], {sp4_v_b[15], sp4_v_b[11],
     sp4_v_b[7], sp4_v_b[3], sp4_h_l[46]}, bl[3:0], pgate[15:14], prog,
     reset[15:14], dout1[1], vdd_cntl[15:14], wl[15:14]);
io_odrv4x5 I220 ( cf[11:9], {sp4_v_b[13], sp4_v_b[9], sp4_v_b[5],
     sp4_v_b[1], sp4_h_l[42]}, bl[3:0], pgate[7:6], prog, reset[7:6],
     dout1[0], vdd_cntl[7:6], wl[7:6]);
io_odrv4x5 I221 ( cf[8:6], {sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2]}, bl[3:0], pgate[5:4], prog, reset[5:4],
     dout1[0], vdd_cntl[5:4], wl[5:4]);
io_odrv4x5 I_odrv_4x5_0 ( cf[2:0], {sp4_h_l[32], sp4_h_l[24],
     sp4_h_l[16], sp4_h_l[8], sp4_h_l[0]}, bl[3:0], pgate[1:0], prog,
     reset[1:0], dout0[0], vdd_cntl[1:0], wl[1:0]);
io_odrv4x5 I223 ( cf[5:3], {sp4_v_b[12], sp4_v_b[8], sp4_v_b[4],
     sp4_v_b[0], sp4_h_l[40]}, bl[3:0], pgate[3:2], prog, reset[3:2],
     dout0[0], vdd_cntl[3:2], wl[3:2]);
io_odrv4x5 I215 ( cf[17:15], {sp4_v_b[14], sp4_v_b[10], sp4_v_b[6],
     sp4_v_b[2], sp4_h_l[44]}, bl[3:0], pgate[11:10], prog,
     reset[11:10], dout0[1], vdd_cntl[11:10], wl[11:10]);

endmodule
// Library - misc, Cell - eh_core_pup_2, View - schematic
// LAST TIME SAVED: Jul 11 11:51:16 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module eh_core_pup_2 ( por_b );
output  por_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



rppolywo  R10 ( .MINUS(net130), .PLUS(net109));
rppolywo  R12 ( .MINUS(net154), .PLUS(net157));
rppolywo  R6 ( .MINUS(out_1), .PLUS(net124));
rppolywo  R9 ( .MINUS(net118), .PLUS(net130));
rppolywo  R15 ( .MINUS(net166), .PLUS(div_1));
rppolywo  R13 ( .MINUS(net157), .PLUS(net145));
rppolywo  R1 ( .MINUS(net068), .PLUS(net048));
rppolywo  R2 ( .MINUS(net067), .PLUS(net068));
rppolywo  R4 ( .MINUS(net142), .PLUS(net148));
rppolywo  R5 ( .MINUS(div_1), .PLUS(net142));
rppolywo  R41 ( .MINUS(net039), .PLUS(net042));
rppolywo  R40 ( .MINUS(net042), .PLUS(vdd_));
rppolywo  R11 ( .MINUS(net109), .PLUS(net154));
rppolywo  R0 ( .MINUS(net048), .PLUS(net039));
rppolywo  R8 ( .MINUS(net127), .PLUS(net118));
rppolywo  R14 ( .MINUS(net145), .PLUS(net166));
rppolywo  R3 ( .MINUS(net148), .PLUS(net067));
rppolywo  R7 ( .MINUS(net124), .PLUS(net127));
nch_hvt  M0 ( .D(out_1), .B(gnd_), .G(div_1), .S(gnd_));
nch_hvt  M2 ( .D(out_1), .B(gnd_), .G(out_2), .S(gnd_));
nch_hvt  M6 ( .D(gnd_), .B(gnd_), .G(out_2), .S(gnd_));
inv_hvt I11 ( .A(out_4), .Y(net193));
inv_hvt I2 ( .A(out_3), .Y(out_4));
inv_hvt I7 ( .A(out_1), .Y(out_2));
inv_hvt I9 ( .A(out_2), .Y(out_3));
inv_hvt I6 ( .A(net193), .Y(por_b));

endmodule
// Library - io, Cell - io_gmux_x2, View - schematic
// LAST TIME SAVED: Aug 21 18:00:57 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module io_gmux_x2 ( gout, bl, min0, min1, pgate, prog, reset, vdd_cntl,
     wl );


input  prog;

output [1:0]  gout;

inout [5:0]  bl;

input [15:0]  min1;
input [15:0]  min0;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbit;

wire  [11:0]  cbitb;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
g_mux Ig_upper ( .prog(prog), .inmuxo(gout[1]), .cbit({cbit[7],
     cbit[6], cbit[3], cbit[10], cbit[8]}), .cbitb({cbitb[7], cbitb[6],
     cbitb[3], cbitb[10], cbitb[8]}), .min(min1[15:0]));
g_mux Ig_low ( .prog(prog), .inmuxo(gout[0]), .cbit({cbit[5], cbit[4],
     cbit[1], cbit[2], cbit[0]}), .cbitb({cbitb[5], cbitb[4], cbitb[1],
     cbitb[2], cbitb[0]}), .min(min0[15:0]));

endmodule
// Library - io, Cell - io_gmux_x16bare, View - schematic
// LAST TIME SAVED: Jul 31 17:47:21 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module io_gmux_x16bare ( lc_trk_g0, lc_trk_g1, bl, min0, min1, min2,
     min3, min4, min5, min6, min7, min8, min9, min10, min11, min12,
     min13, min14, min15, pgate, prog, reset, vdd_cntl, wl );


input  prog;

output [7:0]  lc_trk_g1;
output [7:0]  lc_trk_g0;

inout [5:0]  bl;

input [15:0]  min3;
input [15:0]  min9;
input [15:0]  min7;
input [15:0]  min1;
input [15:0]  min13;
input [15:0]  min12;
input [15:0]  min14;
input [15:0]  min6;
input [15:0]  min5;
input [15:0]  min2;
input [15:0]  min10;
input [15:0]  min15;
input [15:0]  vdd_cntl;
input [15:0]  reset;
input [15:0]  wl;
input [15:0]  min11;
input [15:0]  min0;
input [15:0]  min8;
input [15:0]  min4;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



io_gmux_x2 Iio_gmux4 ( .vdd_cntl(vdd_cntl[9:8]), .bl(bl[5:0]),
     .min0(min8[15:0]), .gout(lc_trk_g1[1:0]), .wl(wl[9:8]),
     .reset(reset[9:8]), .pgate(pgate[9:8]), .min1(min9[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux5 ( .vdd_cntl(vdd_cntl[11:10]), .bl(bl[5:0]),
     .min0(min10[15:0]), .gout(lc_trk_g1[3:2]), .wl(wl[11:10]),
     .reset(reset[11:10]), .pgate(pgate[11:10]), .min1(min11[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux6 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]),
     .min0(min12[15:0]), .gout(lc_trk_g1[5:4]), .wl(wl[13:12]),
     .reset(reset[13:12]), .pgate(pgate[13:12]), .min1(min13[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]),
     .min0(min2[15:0]), .gout(lc_trk_g0[3:2]), .wl(wl[3:2]),
     .reset(reset[3:2]), .pgate(pgate[3:2]), .min1(min3[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]),
     .min0(min0[15:0]), .gout(lc_trk_g0[1:0]), .wl(wl[1:0]),
     .reset(reset[1:0]), .pgate(pgate[1:0]), .min1(min1[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux2 ( .vdd_cntl(vdd_cntl[5:4]), .bl(bl[5:0]),
     .min0(min4[15:0]), .gout(lc_trk_g0[5:4]), .wl(wl[5:4]),
     .reset(reset[5:4]), .pgate(pgate[5:4]), .min1(min5[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux3 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]),
     .min0(min6[15:0]), .gout(lc_trk_g0[7:6]), .wl(wl[7:6]),
     .reset(reset[7:6]), .pgate(pgate[7:6]), .min1(min7[15:0]),
     .prog(prog));
io_gmux_x2 Iio_gmux7 ( .vdd_cntl(vdd_cntl[15:14]), .bl(bl[5:0]),
     .min0(min14[15:0]), .gout(lc_trk_g1[7:6]), .wl(wl[15:14]),
     .reset(reset[15:14]), .pgate(pgate[15:14]), .min1(min15[15:0]),
     .prog(prog));

endmodule
// Library - io, Cell - ioin_mux, View - schematic
// LAST TIME SAVED: May 18 11:01:33 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module ioin_mux ( inmuxo, cbit[3], cbit[2], cbit[1], cbit[0], cbitb[3],
     cbitb[2], cbitb[1], cbitb[0], min[7:0], prog );
output  inmuxo;

input  prog;

input [0:3]  cbitb;
input [7:0]  min;
input [0:3]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I278 ( .A(net146), .Y(inmuxo));
nor2_hvt I46 ( .A(prog), .B(cbitb[3]), .Y(en));
nand2_hvt Inand2_muxo ( .A(st2), .Y(net146), .B(en));
txgate_hvt I247 ( .in(min[2]), .out(st01), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I257 ( .in(min[6]), .out(st03), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I254 ( .in(min[3]), .out(st01), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I244 ( .in(min[0]), .out(st00), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I253 ( .in(st02), .out(st11), .pp(cbit[1]), .nn(cbitb[1]));
txgate_hvt I249 ( .in(st01), .out(st10), .pp(cbitb[1]), .nn(cbit[1]));
txgate_hvt I274 ( .in(st03), .out(st11), .pp(cbitb[1]), .nn(cbit[1]));
txgate_hvt I252 ( .in(st11), .out(st2), .pp(cbitb[2]), .nn(cbit[2]));
txgate_hvt I248 ( .in(st00), .out(st10), .pp(cbit[1]), .nn(cbitb[1]));
txgate_hvt I255 ( .in(min[4]), .out(st02), .pp(cbit[0]),
     .nn(cbitb[0]));
txgate_hvt I250 ( .in(st10), .out(st2), .pp(cbit[2]), .nn(cbitb[2]));
txgate_hvt I258 ( .in(min[7]), .out(st03), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I256 ( .in(min[5]), .out(st02), .pp(cbitb[0]),
     .nn(cbit[0]));
txgate_hvt I246 ( .in(min[1]), .out(st00), .pp(cbitb[0]),
     .nn(cbit[0]));

endmodule
// Library - io, Cell - ioinmx2nor2invx2bdlc, View - schematic
// LAST TIME SAVED: Aug 21 18:04:33 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module ioinmx2nor2invx2bdlc ( bankcntl, spi, ti, bl, cdone_in, min0,
     min1, min2, padin, pgate, prog, reset, vdd_cntl, wl );
output  bankcntl;


input  cdone_in, prog;

output [1:0]  ti;
output [1:0]  spi;

inout [5:0]  bl;

input [7:0]  min2;
input [1:0]  vdd_cntl;
input [7:0]  min1;
input [1:0]  reset;
input [1:0]  padin;
input [7:0]  min0;
input [1:0]  pgate;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  spib;

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
nor2_hvt I192_1_ ( .A(padin[1]), .B(cdone_in), .Y(spib[1]));
nor2_hvt I192_0_ ( .A(padin[0]), .B(cdone_in), .Y(spib[0]));
inv_hvt I187_1_ ( .A(spib[1]), .Y(spi[1]));
inv_hvt I187_0_ ( .A(spib[0]), .Y(spi[0]));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
ioin_mux I193 ( bankcntl, {cbit[11], cbit[8], cbit[9], cbit[10]},
     {cbitb[11], cbitb[8], cbitb[9], cbitb[10]}, min2[7:0], prog);
ioin_mux I185 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux I186 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]}, {cbitb[5],
     cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);

endmodule
// Library - io, Cell - ioinmx1mux2, View - schematic
// LAST TIME SAVED: Aug 21 18:09:41 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module ioinmx1mux2 ( clk, mo, ti, bl, cdone_in, ce, ceb, in, min,
     pgate, prog, reset, spi, vdd_cntl, wl );
output  clk, ti;


input  cdone_in, ceb, prog;

output [1:0]  mo;

inout [5:0]  bl;

input [7:0]  min;
input [1:0]  spi;
input [1:0]  wl;
input [1:0]  in;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
input [1:0]  reset;
input [11:0]  ce;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
clk_mux12to1 I298 ( .prog(prog), .min(ce[11:0]), .clk(clk),
     .clkb(net63), .cbitb({cbitb[5], cbitb[9], cbitb[7], cbitb[10],
     cbitb[6], cbitb[4]}), .cbit({cbit[5], cbit[9], cbit[7], cbit[10],
     cbit[6], cbit[4]}), .cenb(ceb));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
mux2x1_hvt Iemux_1_ ( .in1(in[1]), .in0(spi[1]), .out(mo[1]),
     .sel(cdone_in));
mux2x1_hvt Iemux_0_ ( .in1(in[0]), .in0(spi[0]), .out(mo[0]),
     .sel(cdone_in));
ioin_mux I185 ( ti, {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min[7:0], prog);

endmodule
// Library - io, Cell - ioinmx2nand2inv, View - schematic
// LAST TIME SAVED: Sep 26 11:29:24 2007
// NETLIST TIME: Nov 14 16:17:15 2008
`timescale 1ns / 1ns 

module ioinmx2nand2inv ( ceb, ti, updt, bl, bs_en, ce, min0, min1,
     pgate, prog, reset, update, vdd_cntl, wl );
output  ceb, updt;


input  bs_en, prog, update;

output [1:0]  ti;

inout [5:0]  bl;

input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [7:0]  ce;
input [7:0]  min0;
input [1:0]  reset;
input [7:0]  min1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [11:0]  cbit;

wire  [11:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
ce_clkm8to1 I_cemux ( .cbitb({cbitb[11], cbitb[8], cbitb[9],
     cbitb[10]}), .min(ce[7:0]), .cbit({cbit[11], cbit[8], cbit[9],
     cbit[10]}), .moutb(ceb), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
inv_hvt I181 ( .A(update), .Y(bs_enb));
nand2_hvt I180 ( .A(bs_enb), .Y(updt), .B(bs_en));
ioin_mux I185 ( ti[0], {cbit[1], cbit[3], cbit[2], cbit[0]}, {cbitb[1],
     cbitb[3], cbitb[2], cbitb[0]}, min0[7:0], prog);
ioin_mux I186 ( ti[1], {cbit[5], cbit[6], cbit[7], cbit[4]}, {cbitb[5],
     cbitb[6], cbitb[7], cbitb[4]}, min1[7:0], prog);

endmodule
// Library - io, Cell - sbox1mem, View - schematic
// LAST TIME SAVED: Aug 21 18:03:06 2007
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module sbox1mem ( b, bl, l, r, t, pgate, prog, reset, vdd_cntl, wl );
inout  b, l, r, t;

input  prog;

inout [5:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  reset;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [11:0]  cbitb;

wire  [11:0]  cbit;

wire  [1:0]  r_vdd;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
sbox1m3to1 I232 ( .in2(r), .cb({cbitb[3], cbitb[6]}), .op(t), .in0(l),
     .in1(b), .c({cbit[3], cbit[6]}), .prog(prog));
sbox1m3to1 I230 ( .in2(r), .cb({cbitb[1], cbitb[4]}), .op(l), .in0(b),
     .in1(t), .c({cbit[1], cbit[4]}), .prog(prog));
sbox1m3to1 I226 ( .in2(r), .cb({cbitb[8], cbitb[5]}), .op(b), .in0(l),
     .in1(t), .c({cbit[8], cbit[5]}), .prog(prog));
sbox1m3to1 I231 ( .in2(b), .cb({cbitb[10], cbitb[7]}), .op(r), .in0(l),
     .in1(t), .c({cbit[10], cbit[7]}), .prog(prog));
cram2x2 Ixpm_2_ ( .bl(bl[5:4]), .q_b(cbitb[11:8]), .reset(reset[1:0]),
     .q(cbit[11:8]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_1_ ( .bl(bl[3:2]), .q_b(cbitb[7:4]), .reset(reset[1:0]),
     .q(cbit[7:4]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
cram2x2 Ixpm_0_ ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - sbox1_colbdlc, View - schematic
// LAST TIME SAVED: Aug 21 18:09:59 2007
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module sbox1_colbdlc ( fabric_out, inclk, outclk, padeb, pado,
     spi_ss_in_b, ti, updt, bl, l, r, sp4_v_b, t_mid, bs_en, cdone_in,
     ceb_in, clk_in, inclk_in, min0, min1, min2, min3, min4, min5,
     min6, oeb, out, padin, pgate, prog, reset, spioeb, spiout, update,
     vdd_cntl, wl );
output  fabric_out, inclk, outclk, updt;


input  bs_en, cdone_in, prog, update;

output [1:0]  pado;
output [1:0]  padeb;
output [5:0]  ti;
output [1:0]  spi_ss_in_b;

inout [5:0]  bl;
inout [3:0]  r;
inout [3:0]  sp4_v_b;
inout [3:0]  t_mid;
inout [3:0]  l;

input [7:0]  min1;
input [1:0]  spioeb;
input [11:0]  clk_in;
input [7:0]  ceb_in;
input [1:0]  oeb;
input [7:0]  min2;
input [7:0]  min4;
input [7:0]  min0;
input [1:0]  padin;
input [7:0]  min5;
input [7:0]  min3;
input [1:0]  spiout;
input [1:0]  out;
input [7:0]  min6;
input [15:0]  reset;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [11:0]  inclk_in;
input [15:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ioinmx2nor2invx2bdlc I5 ( .vdd_cntl(vdd_cntl[5:4]), .min2(min6[7:0]),
     .bankcntl(fabric_out), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[5:4]), .ti(ti[1:0]), .min0(min0[7:0]),
     .min1(min1[7:0]), .spi(spi_ss_in_b[1:0]), .cdone_in(cdone_in),
     .padin(padin[1:0]), .wl(wl[5:4]), .reset(reset[5:4]));
ioinmx1mux2 I7 ( .vdd_cntl(vdd_cntl[9:8]), .ceb(net169),
     .ce(inclk_in[11:0]), .bl(bl[5:0]), .clk(inclk), .prog(prog),
     .in(out[1:0]), .ti(ti[2]), .min(min2[7:0]), .spi(spiout[1:0]),
     .wl(wl[9:8]), .reset(reset[9:8]), .pgate(pgate[9:8]),
     .cdone_in(cdone_in), .mo(pado[1:0]));
ioinmx1mux2 I6 ( .vdd_cntl(vdd_cntl[15:14]), .ceb(net169),
     .ce(clk_in[11:0]), .bl(bl[5:0]), .clk(outclk), .prog(prog),
     .in(oeb[1:0]), .ti(ti[5]), .min(min5[7:0]), .spi(spioeb[1:0]),
     .wl(wl[15:14]), .reset(reset[15:14]), .pgate(pgate[15:14]),
     .cdone_in(cdone_in), .mo(padeb[1:0]));
ioinmx2nand2inv I4 ( .vdd_cntl(vdd_cntl[11:10]), .ce(ceb_in[7:0]),
     .ceb(net169), .bl(bl[5:0]), .prog(prog), .pgate(pgate[11:10]),
     .ti(ti[4:3]), .min0(min3[7:0]), .min1(min4[7:0]), .update(update),
     .wl(wl[11:10]), .bs_en(bs_en), .reset(reset[11:10]), .updt(updt));
sbox1mem I3 ( .vdd_cntl(vdd_cntl[13:12]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[13:12]), .b(sp4_v_b[3]), .r(r[3]), .t(t_mid[3]),
     .wl(wl[13:12]), .reset(reset[13:12]), .l(l[3]));
sbox1mem I2 ( .vdd_cntl(vdd_cntl[7:6]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[7:6]), .b(sp4_v_b[2]), .r(r[2]), .t(t_mid[2]),
     .wl(wl[7:6]), .reset(reset[7:6]), .l(l[2]));
sbox1mem I1 ( .vdd_cntl(vdd_cntl[3:2]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[3:2]), .b(sp4_v_b[1]), .r(r[1]), .t(t_mid[1]),
     .wl(wl[3:2]), .reset(reset[3:2]), .l(l[1]));
sbox1mem I0 ( .vdd_cntl(vdd_cntl[1:0]), .bl(bl[5:0]), .prog(prog),
     .pgate(pgate[1:0]), .b(sp4_v_b[0]), .r(r[0]), .t(t_mid[0]),
     .wl(wl[1:0]), .reset(reset[1:0]), .l(l[0]));

endmodule
// Library - io, Cell - odrv12x3, View - schematic
// LAST TIME SAVED: Aug 23 11:52:00 2007
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module odrv12x3 ( sp12, bl, pgate, prog, reset, slfop, vdd_cntl, wl );


input  prog;

output [2:0]  sp12;

inout [1:0]  bl;

input [1:0]  pgate;
input [1:0]  wl;
input [1:0]  reset;
input [1:0]  vdd_cntl;
input [2:0]  slfop;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12_2_ ( .slfop(slfop[2]), .cbitb(cbitb[2]),
     .sp12(sp12[2]), .prog(prog));
odrv12 I_odrv12_1_ ( .slfop(slfop[1]), .cbitb(cbitb[1]),
     .sp12(sp12[1]), .prog(prog));
odrv12 I_odrv12_0_ ( .slfop(slfop[0]), .cbitb(cbitb[0]),
     .sp12(sp12[0]), .prog(prog));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - cebdffrqn, View - schematic
// LAST TIME SAVED: Jan 31 09:00:47 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module cebdffrqn ( q, qn, ceb, clk, d, r );
output  q, qn;

input  ceb, clk, d, r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



anor21_hvt I54 ( .A(net62), .B(clk), .Y(clatb), .C(ceb));
nand2_hvt I290 ( .A(clk), .Y(clkb), .B(clatb));
nand2_hvt I42 ( .A(si), .B(rstb), .Y(so));
nor2_hvt INAND2_m ( .A(r), .Y(q), .B(mi));
inv_hvt I39 ( .A(q), .Y(qn));
inv_hvt Iinv_ckfb ( .A(clatb), .Y(net62));
inv_hvt I50 ( .A(clkb), .Y(clkd));
inv_hvt I43 ( .A(so), .Y(low_s));
inv_hvt I40 ( .A(r), .Y(rstb));
txgate_hvt I44 ( .in(d), .out(si), .pp(clkd), .nn(clkb));
txgate_hvt I52 ( .in(so), .out(mi), .pp(clkb), .nn(clkd));
txgate_hvt I51 ( .in(si), .out(low_s), .pp(clkb), .nn(clkd));
txgate_hvt I53 ( .in(mi), .out(qn), .pp(clkd), .nn(clkb));

endmodule
// Library - misc, Cell - SMC_CORE_POR_right, View - schematic
// LAST TIME SAVED: Oct  6 15:00:20 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module SMC_CORE_POR_right ( core_por_b, smc_por_b,
     smc_core_por_bottom1, smc_core_por_bottom2, vddio_rightbank );
output  core_por_b, smc_por_b;

input  smc_core_por_bottom1, smc_core_por_bottom2, vddio_rightbank;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



eh_io_pup_2_new I0 ( .vdd_io(vddio_rightbank), .core_por_b(core_por_b),
     .por_b(net3));
eh_core_pup_2 I1 ( .por_b(core_por_b));
nand4_hvt I2 ( .D(core_por_b), .C(smc_core_por_bottom2), .A(net3),
     .Y(net04), .B(smc_core_por_bottom1));
inv_hvt I3 ( .A(net04), .Y(smc_por_b));

endmodule
// Library - io, Cell - outsel1_hvt, View - schematic
// LAST TIME SAVED: Jul  3 13:08:26 2007
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module outsel1_hvt ( out, clk, in0, in1, in2, sb, sel );
output  out;

input  clk, in0, in1, in2;

input [1:0]  sel;
input [1:0]  sb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I41 ( .A(in1), .Y(net036));
inv_hvt I40 ( .A(clk), .Y(clkb));
txgate_hvt I33 ( .in(whatever), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_hvt I_txgate1 ( .in(net036), .out(whatever), .pp(sb[0]),
     .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(whatever), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(ddr), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_hvt I38 ( .in(in2), .out(ddr), .pp(clkb), .nn(clk));
txgate_hvt I39 ( .in(in1), .out(ddr), .pp(clk), .nn(clkb));

endmodule
// Library - io, Cell - dffrckb, View - schematic
// LAST TIME SAVED: May 11 14:58:52 2007
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module dffrckb ( q, qn, clk, d, e, r );
output  q, qn;

input  clk, d, e, r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



oai21x2_hvt I57 ( .A1(clk), .Y(clat), .A0(clatb), .B0(e));
nor2_hvt I48 ( .B(clat), .A(clk), .Y(clkb));
nand2_hvt I54 ( .A(rstb), .Y(qn), .B(q));
nand2_hvt I42 ( .A(si), .B(rstb), .Y(so));
inv_hvt I55 ( .A(mi), .Y(q));
inv_hvt I50 ( .A(clkb), .Y(clkd));
inv_hvt I56 ( .A(clat), .Y(clatb));
inv_hvt I43 ( .A(so), .Y(low_s));
inv_hvt I40 ( .A(r), .Y(rstb));
txgate_hvt I59 ( .in(d), .out(si), .pp(clkb), .nn(clkd));
txgate_hvt I64 ( .in(low_s), .out(si), .pp(clkd), .nn(clkb));
txgate_hvt I62 ( .in(qn), .out(mi), .pp(clkb), .nn(clkd));
txgate_hvt I60 ( .in(so), .out(mi), .pp(clkd), .nn(clkb));

endmodule
// Library - io, Cell - out_logic_v1, View - schematic
// LAST TIME SAVED: Jan 30 16:41:40 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module out_logic_v1 ( dout, sdo, bs_en, cbit, cbitb, ceb, clk, ddr0,
     ddr1, mode, rstio, sdi, shift, tclk, ud );
output  dout, sdo;

input  bs_en, ceb, clk, ddr0, ddr1, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cebdffrqn Ireg0 ( .ceb(ceb), .clk(mux4clk), .qn(net094), .r(rstio),
     .q(sdo), .d(dd));
outsel1_hvt I169 ( .clk(ddrclk), .in2(udb), .sb(cbitb[1:0]),
     .sel(cbit[1:0]), .in1(net094), .in0(dinb), .out(muxob));
nor2_hvt I179 ( .A(mux4clk), .B(cbit[0]), .Y(ddrclk));
dffrckb Ireg1 ( .e(ud), .clk(mux4clk), .qn(udb), .r(rstio), .q(net44),
     .d(mux4d));
inv_hvt I171 ( .A(doutb), .Y(dout));
inv_hvt I172 ( .A(ddr0), .Y(dinb));
mux2x1_hvt I170 ( .sel(mode), .in1(udb), .in0(muxob), .out(doutb));
mux2x1_hvt I177 ( .in1(tclk), .in0(clk), .out(mux4clk), .sel(bs_en));
mux2x1_hvt I173 ( .in1(sdi), .in0(ddr0), .out(dd), .sel(shift));
mux2x1_hvt I176 ( .in1(sdo), .in0(ddr1), .out(mux4d), .sel(bs_en));

endmodule
// Library - io, Cell - out_logic_v3, View - schematic
// LAST TIME SAVED: Jan 30 16:43:16 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module out_logic_v3 ( dout, sdo, sp12, bl, bs_en, ceb, clk, ddr0, ddr1,
     mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk, ud,
     vdd_cntl, wl );
output  dout, sdo, sp12;


input  bs_en, ceb, clk, ddr0, ddr1, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  vdd_cntl;
input [1:0]  reset;
input [1:0]  pgate;
input [1:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;

wire  [3:0]  cbit;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I181 ( .slfop(slfop), .cbitb(cbitb[1]), .sp12(sp12),
     .prog(prog));
cram2x2 I183 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));
out_logic_v1 I_outlogic_v1 ( .ceb(ceb), .rstio(rstio), .ddr0(ddr0),
     .ddr1(ddr1), .shift(shift), .ud(ud), .clk(clk), .sdo(sdo),
     .sdi(sdi), .cbit({cbit[2], cbit[3]}), .cbitb({cbitb[2],
     cbitb[3]}), .dout(dout), .tclk(tclk), .bs_en(bs_en), .mode(mode));

endmodule
// Library - io, Cell - insel1_hvt, View - schematic
// LAST TIME SAVED: Jul  2 18:38:19 2007
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module insel1_hvt ( out, in0, in1, in2, in3, sb, sel );
output  out;

input  in0, in1, in2, in3;

input [1:0]  sb;
input [1:0]  sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I39 ( .in(in3), .out(net025), .pp(sb[0]), .nn(sel[0]));
txgate_hvt I40 ( .in(in2), .out(net025), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I33 ( .in(net038), .out(out), .pp(sel[1]), .nn(sb[1]));
txgate_hvt I_txgate1 ( .in(in1), .out(net038), .pp(sb[0]),
     .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(net038), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(net025), .out(out), .pp(sb[1]), .nn(sel[1]));

endmodule
// Library - io, Cell - in_logic_v1, View - schematic
// LAST TIME SAVED: Jan 30 16:34:50 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module in_logic_v1 ( dout0, dout1, sdo, bs_en, cbit, cbitb, ceb, clk,
     cntl, din, mode, rstio, sdi, shift, tclk, ud );
output  dout0, dout1, sdo;

input  bs_en, ceb, clk, cntl, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbitb;
input [1:0]  cbit;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cebdffrqn I167 ( .ceb(ceb), .clk(ck2r0), .qn(regb), .r(rstio), .q(sdo),
     .d(dd));
nand2_hvt I184 ( .A(cntl), .Y(cbit1b), .B(cbit[1]));
insel1_hvt I181 ( .in1(dinb), .in0(regb), .out(reg_), .sb({cbit1b,
     cbitb[0]}), .sel({cbit1, cbit[0]}), .in2(net037), .in3(net037));
dffrckb I168 ( .e(ud), .clk(ck2r0), .qn(udd), .r(rstio), .q(net060),
     .d(net056));
inv_hvt I171 ( .A(doutb), .Y(dout0));
inv_hvt I182 ( .A(udd), .Y(dout1));
inv_hvt I185 ( .A(cbit1b), .Y(cbit1));
inv_hvt I186 ( .A(dout0), .Y(net037));
inv_hvt I172 ( .A(din), .Y(dinb));
mux2x1_hvt I170 ( .sel(mode), .in1(udd), .in0(reg_), .out(doutb));
mux2x1_hvt I178 ( .in1(tclk), .in0(clk), .out(ck2r0), .sel(bs_en));
mux2x1_hvt I173 ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
mux2x1_hvt I179 ( .in1(sdo), .in0(din), .out(net056), .sel(bs_en));

endmodule
// Library - io, Cell - in_logic_v3, View - schematic
// LAST TIME SAVED: Jan 30 16:36:21 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module in_logic_v3 ( dout0, dout1, sdo, sp12, bl, bs_en, ceb, clk,
     cntl, din, mode, pgate, prog, reset, rstio, sdi, shift, slfop,
     tclk, ud, vdd_cntl, wl );
output  dout0, dout1, sdo, sp12;


input  bs_en, ceb, clk, cntl, din, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  reset;
input [1:0]  wl;
input [1:0]  vdd_cntl;
input [1:0]  pgate;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  cbit;

wire  [1:0]  r_vdd;

wire  [3:0]  cbitb;



pch_hvt  M0_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]), .S(vdd_));
pch_hvt  M0_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]), .S(vdd_));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[3]), .sp12(sp12),
     .prog(prog));
in_logic_v1 I_in_logic ( .ceb(ceb), .rstio(rstio), .din(din),
     .cntl(cntl), .dout1(dout1), .dout0(dout0), .shift(shift), .ud(ud),
     .clk(clk), .sdo(sdo), .sdi(sdi), .cbit({cbit[0], cbit[1]}),
     .cbitb({cbitb[0], cbitb[1]}), .tclk(tclk), .bs_en(bs_en),
     .mode(mode));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - io, Cell - ioesel_hvt, View - schematic
// LAST TIME SAVED: Aug 21 18:20:13 2007
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module ioesel_hvt ( out, in0, in1, sb, sel );
output  out;

input  in0, in1;

input [1:0]  sel;
input [1:0]  sb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I38 ( .A(sel[0]), .Y(net017));
txgate_hvt I33 ( .in(mid), .out(out), .pp(sb[1]), .nn(sel[1]));
txgate_hvt I_txgate1 ( .in(in1), .out(mid), .pp(sb[0]), .nn(sel[0]));
txgate_hvt I31 ( .in(in0), .out(mid), .pp(sel[0]), .nn(sb[0]));
txgate_hvt I34 ( .in(net017), .out(out), .pp(sel[1]), .nn(sb[1]));

endmodule
// Library - io, Cell - ioe_logic_v1, View - schematic
// LAST TIME SAVED: Jan 30 16:28:17 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module ioe_logic_v1 ( outb, sdo, bs_en, cbit, cbitb, ceb, clk, din,
     mode, rstio, sdi, shift, tclk, ud );
output  outb, sdo;

input  bs_en, ceb, clk, din, mode, rstio, sdi, shift, tclk, ud;

input [1:0]  cbit;
input [1:0]  cbitb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



cebdffrqn I167 ( .ceb(ceb), .clk(net039), .qn(regb), .r(rstio),
     .q(sdo), .d(dd));
dffrckb I168 ( .e(ud), .clk(net039), .qn(udd), .r(rstio), .q(net44),
     .d(sdo));
inv_hvt I172 ( .A(din), .Y(dinb));
mux2x1_hvt I175 ( .in1(tclk), .in0(clk), .out(net039), .sel(bs_en));
mux2x1_hvt I170 ( .sel(mode), .in1(udd), .in0(regmuxb), .out(outb));
mux2x1_hvt I173 ( .in1(sdi), .in0(din), .out(dd), .sel(shift));
ioesel_hvt I_ioe_mux2 ( .sb(cbitb[1:0]), .sel(cbit[1:0]), .in1(regb),
     .in0(dinb), .out(regmuxb));

endmodule
// Library - io, Cell - ioe_logic_v3, View - schematic
// LAST TIME SAVED: Jan 30 16:31:06 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module ioe_logic_v3 ( padeb, sdo, sp12, bl, bs_en, ceb, clk, din,
     hiz_b, mode, pgate, prog, reset, rstio, sdi, shift, slfop, tclk,
     ud, vdd_cntl, wl );
output  padeb, sdo, sp12;


input  bs_en, ceb, clk, din, hiz_b, mode, prog, rstio, sdi, shift,
     slfop, tclk, ud;

inout [1:0]  bl;

input [1:0]  reset;
input [1:0]  wl;
input [1:0]  pgate;
input [1:0]  vdd_cntl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  r_vdd;

wire  [3:0]  cbit;

wire  [3:0]  cbitb;



pch_hvt  vdd_cntrl_1_ ( .D(r_vdd[1]), .B(vdd_), .G(vdd_cntl[1]),
     .S(vdd_));
pch_hvt  vdd_cntrl_0_ ( .D(r_vdd[0]), .B(vdd_), .G(vdd_cntl[0]),
     .S(vdd_));
odrv12 I_odrv12x2 ( .slfop(slfop), .cbitb(cbitb[1]), .sp12(sp12),
     .prog(prog));
nand2_hvt I178 ( .A(oed), .Y(padeb), .B(hiz_b));
inv_hvt I179 ( .A(oeb), .Y(oed));
ioe_logic_v1 I_ioe_logic ( .ceb(ceb), .rstio(rstio), .cbit(cbit[3:2]),
     .cbitb(cbitb[3:2]), .outb(oeb), .bs_en(bs_en), .shift(shift),
     .ud(ud), .clk(clk), .sdo(sdo), .sdi(sdi), .din(din), .tclk(tclk),
     .mode(mode));
cram2x2 Icram2x2 ( .bl(bl[1:0]), .q_b(cbitb[3:0]), .reset(reset[1:0]),
     .q(cbit[3:0]), .wl(wl[1:0]), .r_vdd(r_vdd[1:0]),
     .pgate(pgate[1:0]));

endmodule
// Library - misc, Cell - ml_mux3_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:41 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_mux3_hvt ( out, in0, in1, in2, sel );
output  out;

input  in0, in1, in2;

input [3:0]  sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I25 ( .A(sel[2]), .Y(net26));
inv_hvt I24 ( .A(sel[1]), .Y(net28));
inv_hvt I21 ( .A(sel[0]), .Y(net30));
txgate_hvt I23 ( .in(in1), .out(out), .pp(net28), .nn(sel[1]));
txgate_hvt I20 ( .in(in0), .out(out), .pp(net30), .nn(sel[0]));
txgate_hvt I26 ( .in(in2), .out(out), .pp(net26), .nn(sel[2]));
nch_hvt  MN19 ( .D(out), .B(gnd_), .G(sel[3]), .S(gnd_));

endmodule
// Library - io, Cell - PDIDGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:24:26 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module PDIDGZ ( C, PAD );
output  C;

input  PAD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - io, Cell - ioe_col2, View - schematic
// LAST TIME SAVED: Jan 30 16:46:15 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module ioe_col2 ( dout, padeb, pado, sdo, sp12_h_l, bl, bs_en, ceb,
     hiz_b, hold, inclk, mode, outclk, padin, pgate, prog, reset,
     rstio, sdi, shift, tclk, ti, update, vdd_cntl, wl );
output  sdo;


input  bs_en, ceb, hiz_b, hold, inclk, mode, outclk, prog, rstio, sdi,
     shift, tclk, update;

output [1:0]  padeb;
output [1:0]  pado;
output [23:0]  sp12_h_l;
output [3:0]  dout;

inout [1:0]  bl;

input [1:0]  padin;
input [15:0]  vdd_cntl;
input [5:0]  ti;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  wl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



odrv12x3 I218 ( .vdd_cntl(vdd_cntl[7:6]), .slfop({dout[1], dout[1],
     dout[1]}), .sp12({sp12_h_l[18], sp12_h_l[10], sp12_h_l[2]}),
     .bl(bl[1:0]), .wl(wl[7:6]), .reset(reset[7:6]),
     .pgate(pgate[7:6]), .prog(prog));
odrv12x3 I217 ( .vdd_cntl(vdd_cntl[9:8]), .slfop({dout[2], dout[2],
     dout[2]}), .sp12({sp12_h_l[20], sp12_h_l[12], sp12_h_l[4]}),
     .bl(bl[1:0]), .wl(wl[9:8]), .reset(reset[9:8]),
     .pgate(pgate[9:8]), .prog(prog));
out_logic_v3 I_out0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[1:0]),
     .ddr0(ti[1]), .ddr1(ti[2]), .rstio(rstio), .slfop(dout[0]),
     .sp12(sp12_h_l[0]), .dout(pado[0]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[1:0]),
     .reset(reset[1:0]), .sdo(s0), .sdi(sdi), .pgate(pgate[1:0]),
     .tclk(tclk), .bs_en(bs_en), .mode(mode));
out_logic_v3 I_out1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[11:10]),
     .ddr0(ti[4]), .ddr1(ti[5]), .rstio(rstio), .slfop(dout[3]),
     .sp12(sp12_h_l[6]), .dout(pado[1]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[11:10]),
     .reset(reset[11:10]), .sdo(s3), .sdi(s2), .pgate(pgate[11:10]),
     .tclk(tclk), .bs_en(bs_en), .mode(mode));
in_logic_v3 I_in0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[3:2]), .rstio(rstio),
     .slfop(dout[0]), .sp12(sp12_h_l[8]), .shift(shift),
     .dout1(dout[1]), .ud(update), .bl(bl[1:0]), .prog(prog),
     .clk(inclk), .dout0(dout[0]), .wl(wl[3:2]), .reset(reset[3:2]),
     .sdo(s1), .sdi(s0), .pgate(pgate[3:2]), .din(padin[0]),
     .tclk(tclk), .bs_en(bs_en), .cntl(hold), .mode(mode));
in_logic_v3 I_in1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[13:12]),
     .rstio(rstio), .slfop(dout[3]), .sp12(sp12_h_l[14]),
     .shift(shift), .dout1(dout[3]), .ud(update), .bl(bl[1:0]),
     .prog(prog), .clk(inclk), .dout0(dout[2]), .wl(wl[13:12]),
     .reset(reset[13:12]), .sdo(s4), .sdi(s3), .pgate(pgate[13:12]),
     .din(padin[1]), .tclk(tclk), .bs_en(bs_en), .cntl(hold),
     .mode(mode));
ioe_logic_v3 I_ioe0 ( .ceb(ceb), .vdd_cntl(vdd_cntl[5:4]),
     .rstio(rstio), .slfop(dout[0]), .sp12(sp12_h_l[16]),
     .hiz_b(hiz_b), .padeb(padeb[0]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[5:4]),
     .reset(reset[5:4]), .sdo(s2), .sdi(s1), .pgate(pgate[5:4]),
     .din(ti[0]), .tclk(tclk), .bs_en(bs_en), .mode(mode));
ioe_logic_v3 I_ioe1 ( .ceb(ceb), .vdd_cntl(vdd_cntl[15:14]),
     .rstio(rstio), .slfop(dout[3]), .sp12(sp12_h_l[22]),
     .hiz_b(hiz_b), .padeb(padeb[1]), .shift(shift), .ud(update),
     .bl(bl[1:0]), .prog(prog), .clk(outclk), .wl(wl[15:14]),
     .reset(reset[15:14]), .sdo(sdo), .sdi(s4), .pgate(pgate[15:14]),
     .din(ti[3]), .tclk(tclk), .bs_en(bs_en), .mode(mode));

endmodule
// Library - io, Cell - io_col4_BRAM_BOT, View - schematic
// LAST TIME SAVED: Feb  5 08:38:27 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module io_col4_BRAM_BOT ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [1:0]  spi_ss_in_b;
output [1:0]  padeb;
output [3:0]  slf_op;
output [23:0]  cf;

inout [15:0]  sp4_v_t;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_b;
inout [17:0]  bl;

input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  wl;
input [1:0]  padin;
input [7:0]  glb_netwk;
input [1:0]  spioeb;
input [7:0]  lft_op;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [15:0]  vdd_cntl;
input [1:0]  spiout;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net128));
rm6  R14_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R14_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R14_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R14_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R14_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R14_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R14_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R14_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R14_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R14_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R14_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R14_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R14_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R14_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R14_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R14_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net128, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(net128),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net128));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net128), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));

endmodule
// Library - io, Cell - io_col4_BOT, View - schematic
// LAST TIME SAVED: Feb  5 08:37:42 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module io_col4_BOT ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [1:0]  spi_ss_in_b;
output [1:0]  padeb;
output [23:0]  cf;
output [3:0]  slf_op;

inout [15:0]  sp4_v_t;
inout [17:0]  bl;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;

input [1:0]  spioeb;
input [1:0]  padin;
input [1:0]  spiout;
input [15:0]  pgate;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [7:0]  glb_netwk;
input [15:0]  reset;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [3:0]  t_mid;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net0214));
rm6  R14_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R14_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R14_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R14_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R14_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R14_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R14_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R14_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R14_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R14_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R14_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R14_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R14_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R14_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R14_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R14_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net0214, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(net0214),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net0214));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net0214), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));

endmodule
// Library - leafcell, Cell - preio_bot_l, View - schematic
// LAST TIME SAVED: Oct 16 14:34:39 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module preio_bot_l ( bs_en_o, ceb_o, cf_b, fabric_out_16_00, hiz_b_o,
     mode_o, padeb_b, padin_80, pado_b, r_o, sdo, shift_o,
     slf_op_01_00, slf_op_02_00, slf_op_03_00, slf_op_04_00,
     slf_op_05_00, slf_op_06_00, slf_op_07_00, slf_op_08_00,
     slf_op_09_00, slf_op_10_00, slf_op_11_00, slf_op_12_00,
     slf_op_13_00, slf_op_14_00, slf_op_15_00, slf_op_16_00, tclk_o,
     update_o, bl_01, bl_02, bl_03, bl_04, bl_05, bl_06, bl_07, bl_08,
     bl_09, bl_10, bl_11, bl_12, bl_13, bl_14, bl_15, bl_16,
     sp4_h_l_01_00, sp4_h_l_02_00, sp4_h_l_03_00, sp4_h_l_04_00,
     sp4_h_l_05_00, sp4_h_l_06_00, sp4_h_l_07_00, sp4_h_l_08_00,
     sp4_h_l_09_00, sp4_h_l_10_00, sp4_h_l_11_00, sp4_h_l_12_00,
     sp4_h_l_13_00, sp4_h_l_14_00, sp4_h_l_15_00, sp4_h_l_16_00,
     sp4_h_r_16_00, sp4_v_t_00_01, sp12_h_l_01_00, sp12_h_l_02_00,
     sp12_h_l_03_00, sp12_h_l_04_00, sp12_h_l_05_00, sp12_h_l_06_00,
     sp12_h_l_07_00, sp12_h_l_08_00, sp12_h_l_09_00, sp12_h_l_10_00,
     sp12_h_l_11_00, sp12_h_l_12_00, sp12_h_l_13_00, sp12_h_l_14_00,
     sp12_h_l_15_00, sp12_h_l_16_00, bs_en_i, ceb_i, glb_net_01,
     glb_net_02, glb_net_03, glb_net_04, glb_net_05, glb_net_06,
     glb_net_07, glb_net_08, glb_net_09, glb_net_10, glb_net_11,
     glb_net_12, glb_net_13, glb_net_14, glb_net_15, glb_net_16,
     hiz_b_i, hold_b_l, lft_op_01_00, lft_op_02_00, lft_op_03_00,
     lft_op_04_00, lft_op_05_00, lft_op_06_00, lft_op_07_00,
     lft_op_08_00, lft_op_09_00, lft_op_10_00, lft_op_11_00,
     lft_op_12_00, lft_op_13_00, lft_op_14_00, lft_op_15_00,
     lft_op_16_00, mode_i, padin_b, pgate_l, prog, r_i, reset_l, sdi,
     shift_i, tclk_i, tiegnd, tievdd, tnl_op_01_00, tnr_op_16_00,
     update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_16_00, hiz_b_o, mode_o, padin_80,
     r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, tiegnd, tievdd, update_i;

output [3:0]  slf_op_02_00;
output [3:0]  slf_op_14_00;
output [3:0]  slf_op_11_00;
output [3:0]  slf_op_09_00;
output [3:0]  slf_op_12_00;
output [3:0]  slf_op_04_00;
output [3:0]  slf_op_16_00;
output [3:0]  slf_op_15_00;
output [3:0]  slf_op_08_00;
output [3:0]  slf_op_03_00;
output [3:0]  slf_op_07_00;
output [383:0]  cf_b;
output [3:0]  slf_op_05_00;
output [3:0]  slf_op_10_00;
output [3:0]  slf_op_06_00;
output [3:0]  slf_op_01_00;
output [29:0]  pado_b;
output [3:0]  slf_op_13_00;
output [29:0]  padeb_b;

inout [23:0]  sp12_h_l_14_00;
inout [23:0]  sp12_h_l_09_00;
inout [47:0]  sp4_h_l_09_00;
inout [47:0]  sp4_h_l_11_00;
inout [47:0]  sp4_h_l_03_00;
inout [23:0]  sp12_h_l_08_00;
inout [23:0]  sp12_h_l_07_00;
inout [47:0]  sp4_h_l_06_00;
inout [23:0]  sp12_h_l_12_00;
inout [23:0]  sp12_h_l_11_00;
inout [15:0]  sp4_v_t_00_01;
inout [23:0]  sp12_h_l_01_00;
inout [53:0]  bl_01;
inout [53:0]  bl_02;
inout [53:0]  bl_05;
inout [53:0]  bl_07;
inout [53:0]  bl_11;
inout [47:0]  sp4_h_l_04_00;
inout [47:0]  sp4_h_l_14_00;
inout [47:0]  sp4_h_l_02_00;
inout [53:0]  bl_03;
inout [53:0]  bl_06;
inout [23:0]  sp12_h_l_16_00;
inout [23:0]  sp12_h_l_02_00;
inout [47:0]  sp4_h_l_05_00;
inout [53:0]  bl_16;
inout [53:0]  bl_14;
inout [23:0]  sp12_h_l_13_00;
inout [47:0]  sp4_h_l_10_00;
inout [53:0]  bl_15;
inout [23:0]  sp12_h_l_10_00;
inout [47:0]  sp4_h_l_12_00;
inout [53:0]  bl_10;
inout [41:0]  bl_08;
inout [47:0]  sp4_h_l_01_00;
inout [23:0]  sp12_h_l_15_00;
inout [53:0]  bl_04;
inout [47:0]  sp4_h_l_08_00;
inout [47:0]  sp4_h_l_07_00;
inout [23:0]  sp12_h_l_05_00;
inout [23:0]  sp12_h_l_04_00;
inout [15:0]  sp4_h_r_16_00;
inout [23:0]  sp12_h_l_06_00;
inout [53:0]  bl_12;
inout [47:0]  sp4_h_l_15_00;
inout [53:0]  bl_13;
inout [47:0]  sp4_h_l_16_00;
inout [47:0]  sp4_h_l_13_00;
inout [53:0]  bl_09;
inout [23:0]  sp12_h_l_03_00;

input [7:0]  tnr_op_16_00;
input [7:0]  glb_net_01;
input [7:0]  lft_op_07_00;
input [7:0]  glb_net_03;
input [7:0]  lft_op_05_00;
input [7:0]  glb_net_07;
input [7:0]  glb_net_10;
input [7:0]  glb_net_12;
input [7:0]  glb_net_09;
input [7:0]  lft_op_16_00;
input [7:0]  glb_net_02;
input [15:0]  pgate_l;
input [7:0]  glb_net_13;
input [7:0]  glb_net_05;
input [7:0]  lft_op_09_00;
input [7:0]  lft_op_01_00;
input [7:0]  lft_op_11_00;
input [7:0]  glb_net_04;
input [7:0]  glb_net_11;
input [7:0]  glb_net_14;
input [7:0]  lft_op_06_00;
input [7:0]  lft_op_13_00;
input [7:0]  glb_net_15;
input [7:0]  glb_net_16;
input [7:0]  lft_op_12_00;
input [7:0]  lft_op_02_00;
input [7:0]  lft_op_03_00;
input [29:0]  padin_b;
input [7:0]  lft_op_04_00;
input [7:0]  tnl_op_01_00;
input [7:0]  glb_net_06;
input [15:0]  wl_l;
input [7:0]  lft_op_15_00;
input [7:0]  lft_op_10_00;
input [7:0]  lft_op_08_00;
input [7:0]  lft_op_14_00;
input [7:0]  glb_net_08;
input [15:0]  reset_l;
input [15:0]  vdd_cntl_l;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net1007;

wire  [0:1]  net1133;

wire  [0:15]  net867;

wire  [0:15]  net692;

wire  [0:1]  net1209;

wire  [0:1]  net1223;

wire  [0:15]  net797;

wire  [0:1]  net1198;

wire  [0:15]  net1112;

wire  [0:1]  net1217;

wire  [0:1]  net1200;

wire  [0:15]  net1042;

wire  [0:15]  net972;

wire  [0:1]  net993;

wire  [0:1]  net744;

wire  [0:15]  net727;

wire  [0:1]  net1215;

wire  [0:15]  net1147;

wire  [0:1]  net1210;

wire  [0:1]  net1206;

wire  [0:15]  net937;

wire  [0:1]  net1028;

wire  [0:15]  net1077;

wire  [0:15]  net657;

wire  [0:15]  net902;

wire  [0:15]  net762;

wire  [0:1]  net1203;

wire  [0:1]  net1219;

wire  [0:1]  net1207;

wire  [0:1]  net1213;

wire  [0:1]  net1216;

wire  [0:15]  net832;

wire  [0:1]  net742;



bram_bufferx4x6 I268 ( .in(sdi), .out(net0614));
lowla_modified I267 ( .clk(tclk_i), .min(net0614), .lao(net618));
tckbufx16 I242 ( .in(tclk_i), .out(tclk_o));
fabric_buf8k I264 ( .f_in(padin_b[29]), .f_out(padin_80));
fabric_buf8k I265 ( .f_in(net1180), .f_out(fabric_out_16_00));
io_col4_BRAM_BOT I_IO_08_00bram ( .ceb(ceb_o), .bl({bl_08[5], bl_08[4],
     bl_08[37], bl_08[36], bl_08[35], bl_08[34], bl_08[33], bl_08[32],
     bl_08[14], bl_08[20], bl_08[19], bl_08[18], bl_08[17], bl_08[16],
     bl_08[27], bl_08[26], bl_08[25], bl_08[23]}), .sdo(net625),
     .sdi(net870), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[13:12]), .pado(pado_b[13:12]),
     .padeb(padeb_b[13:12]), .sp4_h_l(sp4_h_l_08_00[47:0]),
     .sp12_h_l(sp12_h_l_08_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1216[0:1]), .tnl_op(lft_op_07_00[7:0]),
     .lft_op(lft_op_08_00[7:0]), .bnl_op(lft_op_09_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[191:168]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_08_00[3:0]), .glb_netwk(glb_net_08[7:0]),
     .hold(hold_b_l), .fabric_out(net1208), .sp4_v_t(net902[0:15]),
     .sp4_v_b(net657[0:15]));
io_col4_BOT I_IO_02_00 ( .ceb(ceb_o), .bl({bl_02[5], bl_02[4],
     bl_02[37], bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32],
     bl_02[14], bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16],
     bl_02[27], bl_02[26], bl_02[25], bl_02[23]}), .sdo(net660),
     .sdi(net730), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[1:0]), .pado(pado_b[1:0]),
     .padeb(padeb_b[1:0]), .sp4_h_l(sp4_h_l_02_00[47:0]),
     .sp12_h_l(sp12_h_l_02_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1207[0:1]), .tnl_op(lft_op_01_00[7:0]),
     .lft_op(lft_op_02_00[7:0]), .bnl_op(lft_op_03_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[47:24]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_00[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_b_l), .fabric_out(net1220), .sp4_v_t(net762[0:15]),
     .sp4_v_b(net692[0:15]));
io_col4_BOT I_IO_11_00 ( .ceb(ceb_o), .bl({bl_11[5], bl_11[4],
     bl_11[37], bl_11[36], bl_11[35], bl_11[34], bl_11[33], bl_11[32],
     bl_11[14], bl_11[20], bl_11[19], bl_11[18], bl_11[17], bl_11[16],
     bl_11[27], bl_11[26], bl_11[25], bl_11[23]}), .sdo(net695),
     .sdi(net765), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[19:18]), .pado(pado_b[19:18]),
     .padeb(padeb_b[19:18]), .sp4_h_l(sp4_h_l_11_00[47:0]),
     .sp12_h_l(sp12_h_l_11_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1217[0:1]), .tnl_op(lft_op_10_00[7:0]),
     .lft_op(lft_op_11_00[7:0]), .bnl_op(lft_op_12_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[263:240]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_11_00[3:0]), .glb_netwk(glb_net_11[7:0]),
     .hold(hold_b_l), .fabric_out(net1221), .sp4_v_t(net797[0:15]),
     .sp4_v_b(net727[0:15]));
io_col4_BOT I_IO_01_00 ( .ceb(ceb_o), .bl({bl_01[5], bl_01[4],
     bl_01[37], bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32],
     bl_01[14], bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16],
     bl_01[27], bl_01[26], bl_01[25], bl_01[23]}), .sdo(net730),
     .sdi(net618), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(net742[0:1]), .pado(net742[0:1]),
     .padeb(net744[0:1]), .sp4_h_l(sp4_h_l_01_00[47:0]),
     .sp12_h_l(sp12_h_l_01_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1210[0:1]), .tnl_op(tnl_op_01_00[7:0]),
     .lft_op(lft_op_01_00[7:0]), .bnl_op(lft_op_02_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[23:0]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_00[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_b_l), .fabric_out(net1222),
     .sp4_v_t(sp4_v_t_00_01[15:0]), .sp4_v_b(net762[0:15]));
io_col4_BOT I_IO_10_00 ( .ceb(ceb_o), .bl({bl_10[5], bl_10[4],
     bl_10[37], bl_10[36], bl_10[35], bl_10[34], bl_10[33], bl_10[32],
     bl_10[14], bl_10[20], bl_10[19], bl_10[18], bl_10[17], bl_10[16],
     bl_10[27], bl_10[26], bl_10[25], bl_10[23]}), .sdo(net765),
     .sdi(net1115), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[17:16]), .pado(pado_b[17:16]),
     .padeb(padeb_b[17:16]), .sp4_h_l(sp4_h_l_10_00[47:0]),
     .sp12_h_l(sp12_h_l_10_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1213[0:1]), .tnl_op(lft_op_09_00[7:0]),
     .lft_op(lft_op_10_00[7:0]), .bnl_op(lft_op_11_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[239:216]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_10_00[3:0]), .glb_netwk(glb_net_10[7:0]),
     .hold(hold_b_l), .fabric_out(net1204), .sp4_v_t(net1147[0:15]),
     .sp4_v_b(net797[0:15]));
io_col4_BOT I_IO_15_00 ( .ceb(ceb_o), .bl({bl_15[5], bl_15[4],
     bl_15[37], bl_15[36], bl_15[35], bl_15[34], bl_15[33], bl_15[32],
     bl_15[14], bl_15[20], bl_15[19], bl_15[18], bl_15[17], bl_15[16],
     bl_15[27], bl_15[26], bl_15[25], bl_15[23]}), .sdo(net800),
     .sdi(net1045), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[27:26]), .pado(pado_b[27:26]),
     .padeb(padeb_b[27:26]), .sp4_h_l(sp4_h_l_15_00[47:0]),
     .sp12_h_l(sp12_h_l_15_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1223[0:1]), .tnl_op(lft_op_14_00[7:0]),
     .lft_op(lft_op_15_00[7:0]), .bnl_op(lft_op_16_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[359:336]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_15_00[3:0]), .glb_netwk(glb_net_15[7:0]),
     .hold(hold_b_l), .fabric_out(net1224), .sp4_v_t(net1077[0:15]),
     .sp4_v_b(net832[0:15]));
io_col4_BOT I_IO_05_00 ( .ceb(ceb_o), .bl({bl_05[5], bl_05[4],
     bl_05[37], bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32],
     bl_05[14], bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16],
     bl_05[27], bl_05[26], bl_05[25], bl_05[23]}), .sdo(net835),
     .sdi(net1080), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[7:6]), .pado(pado_b[7:6]),
     .padeb(padeb_b[7:6]), .sp4_h_l(sp4_h_l_05_00[47:0]),
     .sp12_h_l(sp12_h_l_05_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1219[0:1]), .tnl_op(lft_op_04_00[7:0]),
     .lft_op(lft_op_05_00[7:0]), .bnl_op(lft_op_06_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[119:96]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_00[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_b_l), .fabric_out(net1212), .sp4_v_t(net1112[0:15]),
     .sp4_v_b(net867[0:15]));
io_col4_BOT I_IO_07_00 ( .ceb(ceb_o), .bl({bl_07[5], bl_07[4],
     bl_07[37], bl_07[36], bl_07[35], bl_07[34], bl_07[33], bl_07[32],
     bl_07[14], bl_07[20], bl_07[19], bl_07[18], bl_07[17], bl_07[16],
     bl_07[27], bl_07[26], bl_07[25], bl_07[23]}), .sdo(net870),
     .sdi(net905), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[11:10]), .pado(pado_b[11:10]),
     .padeb(padeb_b[11:10]), .sp4_h_l(sp4_h_l_07_00[47:0]),
     .sp12_h_l(sp12_h_l_07_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1203[0:1]), .tnl_op(lft_op_06_00[7:0]),
     .lft_op(lft_op_07_00[7:0]), .bnl_op(lft_op_08_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[167:144]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_07_00[3:0]), .glb_netwk(glb_net_07[7:0]),
     .hold(hold_b_l), .fabric_out(net1202), .sp4_v_t(net937[0:15]),
     .sp4_v_b(net902[0:15]));
io_col4_BOT I_IO_06_00 ( .ceb(ceb_o), .bl({bl_06[5], bl_06[4],
     bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33], bl_06[32],
     bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17], bl_06[16],
     bl_06[27], bl_06[26], bl_06[25], bl_06[23]}), .sdo(net905),
     .sdi(net835), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[9:8]), .pado(pado_b[9:8]),
     .padeb(padeb_b[9:8]), .sp4_h_l(sp4_h_l_06_00[47:0]),
     .sp12_h_l(sp12_h_l_06_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1209[0:1]), .tnl_op(lft_op_05_00[7:0]),
     .lft_op(lft_op_06_00[7:0]), .bnl_op(lft_op_07_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[143:120]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_00[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_b_l), .fabric_out(net1205), .sp4_v_t(net867[0:15]),
     .sp4_v_b(net937[0:15]));
io_col4_BOT I_IO_03_00 ( .ceb(ceb_o), .bl({bl_03[5], bl_03[4],
     bl_03[37], bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32],
     bl_03[14], bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16],
     bl_03[27], bl_03[26], bl_03[25], bl_03[23]}), .sdo(net940),
     .sdi(net660), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[3:2]), .pado(pado_b[3:2]),
     .padeb(padeb_b[3:2]), .sp4_h_l(sp4_h_l_03_00[47:0]),
     .sp12_h_l(sp12_h_l_03_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1215[0:1]), .tnl_op(lft_op_02_00[7:0]),
     .lft_op(lft_op_03_00[7:0]), .bnl_op(lft_op_04_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[71:48]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_00[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_b_l), .fabric_out(net1211), .sp4_v_t(net692[0:15]),
     .sp4_v_b(net972[0:15]));
io_col4_BOT I_IO_13_00 ( .ceb(ceb_o), .bl({bl_13[5], bl_13[4],
     bl_13[37], bl_13[36], bl_13[35], bl_13[34], bl_13[33], bl_13[32],
     bl_13[14], bl_13[20], bl_13[19], bl_13[18], bl_13[17], bl_13[16],
     bl_13[27], bl_13[26], bl_13[25], bl_13[23]}), .sdo(net975),
     .sdi(net1010), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[23:22]), .pado(pado_b[23:22]),
     .padeb(padeb_b[23:22]), .sp4_h_l(sp4_h_l_13_00[47:0]),
     .sp12_h_l(sp12_h_l_13_00[23:0]), .prog(prog),
     .spi_ss_in_b(net993[0:1]), .tnl_op(lft_op_12_00[7:0]),
     .lft_op(lft_op_13_00[7:0]), .bnl_op(lft_op_14_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[311:288]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_13_00[3:0]), .glb_netwk(glb_net_13[7:0]),
     .hold(hold_b_l), .fabric_out(net1005), .sp4_v_t(net1042[0:15]),
     .sp4_v_b(net1007[0:15]));
io_col4_BOT I_IO_12_00 ( .ceb(ceb_o), .bl({bl_12[5], bl_12[4],
     bl_12[37], bl_12[36], bl_12[35], bl_12[34], bl_12[33], bl_12[32],
     bl_12[14], bl_12[20], bl_12[19], bl_12[18], bl_12[17], bl_12[16],
     bl_12[27], bl_12[26], bl_12[25], bl_12[23]}), .sdo(net1010),
     .sdi(net695), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[21:20]), .pado(pado_b[21:20]),
     .padeb(padeb_b[21:20]), .sp4_h_l(sp4_h_l_12_00[47:0]),
     .sp12_h_l(sp12_h_l_12_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1028[0:1]), .tnl_op(lft_op_11_00[7:0]),
     .lft_op(lft_op_12_00[7:0]), .bnl_op(lft_op_13_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[287:264]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_12_00[3:0]), .glb_netwk(glb_net_12[7:0]),
     .hold(hold_b_l), .fabric_out(net1228), .sp4_v_t(net727[0:15]),
     .sp4_v_b(net1042[0:15]));
io_col4_BOT I_IO_14_00 ( .ceb(ceb_o), .bl({bl_14[5], bl_14[4],
     bl_14[37], bl_14[36], bl_14[35], bl_14[34], bl_14[33], bl_14[32],
     bl_14[14], bl_14[20], bl_14[19], bl_14[18], bl_14[17], bl_14[16],
     bl_14[27], bl_14[26], bl_14[25], bl_14[23]}), .sdo(net1045),
     .sdi(net975), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[25:24]), .pado(pado_b[25:24]),
     .padeb(padeb_b[25:24]), .sp4_h_l(sp4_h_l_14_00[47:0]),
     .sp12_h_l(sp12_h_l_14_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1198[0:1]), .tnl_op(lft_op_13_00[7:0]),
     .lft_op(lft_op_14_00[7:0]), .bnl_op(lft_op_15_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[335:312]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_14_00[3:0]), .glb_netwk(glb_net_14[7:0]),
     .hold(hold_b_l), .fabric_out(net1227), .sp4_v_t(net1007[0:15]),
     .sp4_v_b(net1077[0:15]));
io_col4_BOT I_IO_04_00 ( .ceb(ceb_o), .bl({bl_04[5], bl_04[4],
     bl_04[37], bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32],
     bl_04[14], bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16],
     bl_04[27], bl_04[26], bl_04[25], bl_04[23]}), .sdo(net1080),
     .sdi(net940), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[5:4]), .pado(pado_b[5:4]),
     .padeb(padeb_b[5:4]), .sp4_h_l(sp4_h_l_04_00[47:0]),
     .sp12_h_l(sp12_h_l_04_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1206[0:1]), .tnl_op(lft_op_03_00[7:0]),
     .lft_op(lft_op_04_00[7:0]), .bnl_op(lft_op_05_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[95:72]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_00[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_b_l), .fabric_out(net1110), .sp4_v_t(net972[0:15]),
     .sp4_v_b(net1112[0:15]));
io_col4_BOT I_IO_09_00 ( .ceb(ceb_o), .bl({bl_09[5], bl_09[4],
     bl_09[37], bl_09[36], bl_09[35], bl_09[34], bl_09[33], bl_09[32],
     bl_09[14], bl_09[20], bl_09[19], bl_09[18], bl_09[17], bl_09[16],
     bl_09[27], bl_09[26], bl_09[25], bl_09[23]}), .sdo(net1115),
     .sdi(net625), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[15:14]), .pado(pado_b[15:14]),
     .padeb(padeb_b[15:14]), .sp4_h_l(sp4_h_l_09_00[47:0]),
     .sp12_h_l(sp12_h_l_09_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1133[0:1]), .tnl_op(lft_op_08_00[7:0]),
     .lft_op(lft_op_09_00[7:0]), .bnl_op(lft_op_10_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[215:192]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_09_00[3:0]), .glb_netwk(glb_net_09[7:0]),
     .hold(hold_b_l), .fabric_out(net1145), .sp4_v_t(net657[0:15]),
     .sp4_v_b(net1147[0:15]));
io_col4_BOT I_IO_16_00 ( .ceb(ceb_o), .bl({bl_16[5], bl_16[4],
     bl_16[37], bl_16[36], bl_16[35], bl_16[34], bl_16[33], bl_16[32],
     bl_16[14], bl_16[20], bl_16[19], bl_16[18], bl_16[17], bl_16[16],
     bl_16[27], bl_16[26], bl_16[25], bl_16[23]}), .sdo(sdo),
     .sdi(net800), .spiout({tiegnd, tiegnd}), .cdone_in(tievdd),
     .spioeb({tievdd, tievdd}), .mode(mode_o), .shift(shift_o),
     .hiz_b(hiz_b_o), .r(r_o), .bs_en(bs_en_o), .tclk(tclk_o),
     .update(update_o), .padin(padin_b[29:28]), .pado(pado_b[29:28]),
     .padeb(padeb_b[29:28]), .sp4_h_l(sp4_h_l_16_00[47:0]),
     .sp12_h_l(sp12_h_l_16_00[23:0]), .prog(prog),
     .spi_ss_in_b(net1200[0:1]), .tnl_op(lft_op_15_00[7:0]),
     .lft_op(lft_op_16_00[7:0]), .bnl_op(tnr_op_16_00[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_b[383:360]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_16_00[3:0]), .glb_netwk(glb_net_16[7:0]),
     .hold(hold_b_l), .fabric_out(net1180), .sp4_v_t(net832[0:15]),
     .sp4_v_b(sp4_h_r_16_00[15:0]));
bram_bufferx4 I266 ( .in(ceb_i), .out(ceb_o));
bram_bufferx4 I244 ( .in(mode_i), .out(mode_o));
bram_bufferx4 I249 ( .in(r_i), .out(r_o));
bram_bufferx4 I246 ( .in(shift_i), .out(shift_o));
bram_bufferx4 I247 ( .in(bs_en_i), .out(bs_en_o));
bram_bufferx4 I245 ( .in(update_i), .out(update_o));
bram_bufferx4 I250 ( .in(hiz_b_i), .out(hiz_b_o));

endmodule
// Library - io, Cell - io_col4_LFT, View - schematic
// LAST TIME SAVED: Feb  5 08:40:04 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module io_col4_LFT ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  padeb;
output [1:0]  spi_ss_in_b;
output [23:0]  cf;
output [1:0]  pado;
output [3:0]  slf_op;

inout [15:0]  sp4_v_t;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;

input [1:0]  spioeb;
input [1:0]  padin;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [1:0]  spiout;
input [15:0]  pgate;
input [7:0]  tnl_op;
input [7:0]  lft_op;
input [7:0]  bnl_op;
input [7:0]  glb_netwk;
input [15:0]  reset;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net127));
rm7  R14_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7  R14_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7  R14_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7  R14_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7  R14_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7  R14_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7  R14_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7  R14_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7  R14_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7  R14_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7  R14_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7  R14_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7  R14_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7  R14_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7  R14_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7  R14_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net127, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(net127),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net127));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net127), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));

endmodule
// Library - leafcell, Cell - array_LFT_IO_1x16, View - schematic
// LAST TIME SAVED: Feb  4 15:28:36 2008
// NETLIST TIME: Nov 14 16:17:16 2008
`timescale 1ns / 1ns 

module array_LFT_IO_1x16 ( cf_l, fabric_out_01, fabric_out_02,
     fabric_out_03, fabric_out_04, fabric_out_05, fabric_out_06,
     fabric_out_07, fabric_out_08, fabric_out_09, fabric_out_10,
     fabric_out_11, fabric_out_12, fabric_out_13, fabric_out_14,
     fabric_out_15, fabric_out_16, padeb, pado, sdo, slf_op_01,
     slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07,
     slf_op_08, slf_op_09, slf_op_10, slf_op_11, slf_op_12, slf_op_13,
     slf_op_14, slf_op_15, slf_op_16, spi_ss_in_b, SP4_h_l_01,
     SP4_h_l_02, SP4_h_l_03, SP4_h_l_04, SP4_h_l_05, SP4_h_l_06,
     SP4_h_l_07, SP4_h_l_08, SP4_h_l_09, SP4_h_l_10, SP4_h_l_11,
     SP4_h_l_12, SP4_h_l_13, SP4_h_l_14, SP4_h_l_15, SP4_h_l_16,
     SP12_h_l_01, SP12_h_l_02, SP12_h_l_03, SP12_h_l_04, SP12_h_l_05,
     SP12_h_l_06, SP12_h_l_07, SP12_h_l_08, SP12_h_l_09, SP12_h_l_10,
     SP12_h_l_11, SP12_h_l_12, SP12_h_l_13, SP12_h_l_14, SP12_h_l_15,
     SP12_h_l_16, bl, pgate, reset_b, sp4_v_b_01, sp4_v_t_16, vdd_cntl,
     wl, bnl_op_01, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     mode, padin, prog, r, rgt_op_01, rgt_op_02, rgt_op_03, rgt_op_04,
     rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, rgt_op_09, rgt_op_10,
     rgt_op_11, rgt_op_12, rgt_op_13, rgt_op_14, rgt_op_15, rgt_op_16,
     sdi, shift, spioeb, spiout, tclk, tnl_op_16, update );
output  fabric_out_01, fabric_out_02, fabric_out_03, fabric_out_04,
     fabric_out_05, fabric_out_06, fabric_out_07, fabric_out_08,
     fabric_out_09, fabric_out_10, fabric_out_11, fabric_out_12,
     fabric_out_13, fabric_out_14, fabric_out_15, fabric_out_16, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_16;
output [3:0]  slf_op_15;
output [3:0]  slf_op_10;
output [3:0]  slf_op_03;
output [3:0]  slf_op_09;
output [3:0]  slf_op_12;
output [3:0]  slf_op_13;
output [3:0]  slf_op_02;
output [3:0]  slf_op_06;
output [3:0]  slf_op_14;
output [3:0]  slf_op_07;
output [3:0]  slf_op_05;
output [31:0]  spi_ss_in_b;
output [3:0]  slf_op_08;
output [3:0]  slf_op_11;
output [23:0]  pado;
output [3:0]  slf_op_04;
output [23:0]  padeb;
output [3:0]  slf_op_01;
output [383:0]  cf_l;

inout [23:0]  SP12_h_l_04;
inout [23:0]  SP12_h_l_09;
inout [47:0]  SP4_h_l_12;
inout [23:0]  SP12_h_l_01;
inout [47:0]  SP4_h_l_15;
inout [23:0]  SP12_h_l_07;
inout [23:0]  SP12_h_l_08;
inout [47:0]  SP4_h_l_04;
inout [23:0]  SP12_h_l_13;
inout [23:0]  SP12_h_l_10;
inout [23:0]  SP12_h_l_05;
inout [23:0]  SP12_h_l_02;
inout [47:0]  SP4_h_l_11;
inout [47:0]  SP4_h_l_01;
inout [23:0]  SP12_h_l_16;
inout [47:0]  SP4_h_l_07;
inout [15:0]  sp4_v_t_16;
inout [47:0]  SP4_h_l_06;
inout [23:0]  SP12_h_l_03;
inout [23:0]  SP12_h_l_12;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_08;
inout [47:0]  SP4_h_l_10;
inout [23:0]  SP12_h_l_14;
inout [47:0]  SP4_h_l_16;
inout [23:0]  SP12_h_l_06;
inout [47:0]  SP4_h_l_09;
inout [23:0]  SP12_h_l_15;
inout [47:0]  SP4_h_l_05;
inout [47:0]  SP4_h_l_03;
inout [47:0]  SP4_h_l_14;
inout [15:0]  sp4_v_b_01;
inout [47:0]  SP4_h_l_02;
inout [255:0]  pgate;
inout [255:0]  vdd_cntl;
inout [47:0]  SP4_h_l_13;
inout [23:0]  SP12_h_l_11;
inout [255:0]  reset_b;
inout [255:0]  wl;

input [7:0]  bnl_op_01;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_15;
input [7:0]  rgt_op_13;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_09;
input [7:0]  rgt_op_01;
input [7:0]  rgt_op_04;
input [7:0]  rgt_op_14;
input [7:0]  rgt_op_06;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_02;
input [7:0]  tnl_op_16;
input [7:0]  rgt_op_08;
input [7:0]  rgt_op_10;
input [7:0]  rgt_op_16;
input [7:0]  rgt_op_11;
input [31:0]  spiout;
input [23:0]  padin;
input [7:0]  rgt_op_03;
input [31:0]  spioeb;
input [15:0]  cdone_in;
input [7:0]  rgt_op_12;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net966;

wire  [0:15]  net830;

wire  [0:15]  net1000;

wire  [7:0]  glb_netwk;

wire  [0:15]  net1068;

wire  [0:15]  net796;

wire  [0:15]  net864;

wire  [0:1]  net930;

wire  [0:15]  net932;

wire  [0:1]  net1032;

wire  [0:1]  net931;

wire  [0:15]  net728;

wire  [0:15]  net1170;

wire  [0:1]  net0757;

wire  [0:15]  net694;

wire  [0:15]  net1102;

wire  [0:15]  net1034;

wire  [0:1]  net641;

wire  [0:1]  net1033;

wire  [0:15]  net1136;

wire  [0:1]  net0758;

wire  [0:15]  net762;

wire  [0:15]  net660;

wire  [0:1]  net998;



clk_colbuf8kx8 I109 ( .clko(glb_netwk[7:0]),
     .clki(glb_netwk_col[7:0]));
io_col4_LFT I_io_00_09 ( .ceb(ceb), .sdo(net680), .sdi(net646),
     .spiout(spiout[17:16]), .cdone_in(cdone_in[8]),
     .spioeb(spioeb[17:16]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[11:10]), .pado(pado[11:10]), .padeb(padeb[11:10]),
     .sp4_v_t(net660[0:15]), .spi_ss_in_b(spi_ss_in_b[17:16]),
     .reset(reset_b[143:128]), .sp4_v_b(net694[0:15]),
     .cf(cf_l[215:192]), .bl(bl[17:0]), .slf_op(slf_op_09[3:0]),
     .hold(hold), .fabric_out(fabric_out_09), .prog(prog),
     .lft_op(rgt_op_09[7:0]), .sp12_h_l(SP12_h_l_09[23:0]),
     .sp4_h_l(SP4_h_l_09[47:0]), .wl(wl[143:128]),
     .vdd_cntl(vdd_cntl[143:128]), .glb_netwk(glb_netwk[7:0]),
     .pgate(pgate[143:128]), .bnl_op(rgt_op_08[7:0]),
     .tnl_op(rgt_op_10[7:0]));
io_col4_LFT I_io_00_08 ( .ceb(ceb), .sdo(net714), .sdi(net680),
     .spiout(spiout[15:14]), .cdone_in(cdone_in[7]),
     .spioeb(spioeb[15:14]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[9:8]), .pado(pado[9:8]), .padeb(padeb[9:8]),
     .sp4_v_t(net694[0:15]), .sp4_h_l(SP4_h_l_08[47:0]),
     .sp12_h_l(SP12_h_l_08[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[15:14]), .tnl_op(rgt_op_09[7:0]),
     .lft_op(rgt_op_08[7:0]), .bnl_op(rgt_op_07[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net728[0:15]), .wl(wl[127:112]), .cf(cf_l[191:168]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_08[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_08));
io_col4_LFT I_io_00_07 ( .ceb(ceb), .sdo(net952), .sdi(net714),
     .spiout(spiout[13:12]), .cdone_in(cdone_in[6]),
     .spioeb(spioeb[13:12]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[7:6]), .pado(pado[7:6]), .padeb(padeb[7:6]),
     .sp4_v_t(net728[0:15]), .sp4_h_l(SP4_h_l_07[47:0]),
     .sp12_h_l(SP12_h_l_07[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[13:12]), .tnl_op(rgt_op_08[7:0]),
     .lft_op(rgt_op_07[7:0]), .bnl_op(rgt_op_06[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net966[0:15]), .wl(wl[111:96]), .cf(cf_l[167:144]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_07[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_07));
io_col4_LFT I_io_00_15 ( .ceb(ceb), .sdo(net782), .sdi(net748),
     .spiout(spiout[29:28]), .cdone_in(cdone_in[14]),
     .spioeb(spioeb[29:28]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net0757[0:1]), .pado(net0757[0:1]), .padeb(net0758[0:1]),
     .sp4_v_t(net762[0:15]), .sp4_h_l(SP4_h_l_15[47:0]),
     .sp12_h_l(SP12_h_l_15[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[29:28]), .tnl_op(rgt_op_16[7:0]),
     .lft_op(rgt_op_15[7:0]), .bnl_op(rgt_op_14[7:0]),
     .pgate(pgate[239:224]), .reset(reset_b[239:224]),
     .sp4_v_b(net796[0:15]), .wl(wl[239:224]), .cf(cf_l[359:336]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[239:224]),
     .slf_op(slf_op_15[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_15));
io_col4_LFT I_io_00_14 ( .ceb(ceb), .sdo(net816), .sdi(net782),
     .spiout(spiout[27:26]), .cdone_in(cdone_in[13]),
     .spioeb(spioeb[27:26]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[21:20]), .pado(pado[21:20]), .padeb(padeb[21:20]),
     .sp4_v_t(net796[0:15]), .sp4_h_l(SP4_h_l_14[47:0]),
     .sp12_h_l(SP12_h_l_14[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[27:26]), .tnl_op(rgt_op_15[7:0]),
     .lft_op(rgt_op_14[7:0]), .bnl_op(rgt_op_13[7:0]),
     .pgate(pgate[223:208]), .reset(reset_b[223:208]),
     .sp4_v_b(net830[0:15]), .wl(wl[223:208]), .cf(cf_l[335:312]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[223:208]),
     .slf_op(slf_op_14[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_14));
io_col4_LFT I_io_00_13 ( .ceb(ceb), .sdo(net850), .sdi(net816),
     .spiout(spiout[25:24]), .cdone_in(cdone_in[12]),
     .spioeb(spioeb[25:24]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[19:18]), .pado(pado[19:18]), .padeb(padeb[19:18]),
     .sp4_v_t(net830[0:15]), .sp4_h_l(SP4_h_l_13[47:0]),
     .sp12_h_l(SP12_h_l_13[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[25:24]), .tnl_op(rgt_op_14[7:0]),
     .lft_op(rgt_op_13[7:0]), .bnl_op(rgt_op_12[7:0]),
     .pgate(pgate[207:192]), .reset(reset_b[207:192]),
     .sp4_v_b(net864[0:15]), .wl(wl[207:192]), .cf(cf_l[311:288]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[207:192]),
     .slf_op(slf_op_13[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_13));
io_col4_LFT I_io_00_12 ( .ceb(ceb), .sdo(net1156), .sdi(net850),
     .spiout(spiout[23:22]), .cdone_in(cdone_in[11]),
     .spioeb(spioeb[23:22]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[17:16]), .pado(pado[17:16]), .padeb(padeb[17:16]),
     .sp4_v_t(net864[0:15]), .sp4_h_l(SP4_h_l_12[47:0]),
     .sp12_h_l(SP12_h_l_12[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[23:22]), .tnl_op(rgt_op_13[7:0]),
     .lft_op(rgt_op_12[7:0]), .bnl_op(rgt_op_11[7:0]),
     .pgate(pgate[191:176]), .reset(reset_b[191:176]),
     .sp4_v_b(net1170[0:15]), .wl(wl[191:176]), .cf(cf_l[287:264]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[191:176]),
     .slf_op(slf_op_12[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_12));
io_col4_LFT I_io_00_16 ( .ceb(ceb), .sdo(net748), .sdi(sdi),
     .spiout(spiout[31:30]), .cdone_in(cdone_in[15]),
     .spioeb(spioeb[31:30]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[23:22]), .pado(pado[23:22]), .padeb(padeb[23:22]),
     .sp4_v_t(sp4_v_t_16[15:0]), .sp4_h_l(SP4_h_l_16[47:0]),
     .sp12_h_l(SP12_h_l_16[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[31:30]), .tnl_op(tnl_op_16[7:0]),
     .lft_op(rgt_op_16[7:0]), .bnl_op(rgt_op_15[7:0]),
     .pgate(pgate[255:240]), .reset(reset_b[255:240]),
     .sp4_v_b(net762[0:15]), .wl(wl[255:240]), .cf(cf_l[383:360]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[255:240]),
     .slf_op(slf_op_16[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_16));
io_col4_LFT I_io_00_05 ( .ceb(ceb), .sdo(net1088), .sdi(net918),
     .spiout(spiout[9:8]), .cdone_in(cdone_in[4]),
     .spioeb(spioeb[9:8]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net930[0:1]), .pado(net930[0:1]), .padeb(net931[0:1]),
     .sp4_v_t(net932[0:15]), .sp4_h_l(SP4_h_l_05[47:0]),
     .sp12_h_l(SP12_h_l_05[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[9:8]), .tnl_op(rgt_op_06[7:0]),
     .lft_op(rgt_op_05[7:0]), .bnl_op(rgt_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net1102[0:15]), .wl(wl[79:64]), .cf(cf_l[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_05));
io_col4_LFT I_io_00_06 ( .ceb(ceb), .sdo(net918), .sdi(net952),
     .spiout(spiout[11:10]), .cdone_in(cdone_in[5]),
     .spioeb(spioeb[11:10]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[5:4]), .pado(pado[5:4]), .padeb(padeb[5:4]),
     .sp4_v_t(net966[0:15]), .sp4_h_l(SP4_h_l_06[47:0]),
     .sp12_h_l(SP12_h_l_06[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[11:10]), .tnl_op(rgt_op_07[7:0]),
     .lft_op(rgt_op_06[7:0]), .bnl_op(rgt_op_05[7:0]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net932[0:15]), .wl(wl[95:80]), .cf(cf_l[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_06));
io_col4_LFT I_io_00_02 ( .ceb(ceb), .sdo(net1020), .sdi(net986),
     .spiout(spiout[3:2]), .cdone_in(cdone_in[1]),
     .spioeb(spioeb[3:2]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net998[0:1]), .pado(net998[0:1]), .padeb(net641[0:1]),
     .sp4_v_t(net1000[0:15]), .sp4_h_l(SP4_h_l_02[47:0]),
     .sp12_h_l(SP12_h_l_02[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[3:2]), .tnl_op(rgt_op_03[7:0]),
     .lft_op(rgt_op_02[7:0]), .bnl_op(rgt_op_01[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(net1034[0:15]), .wl(wl[31:16]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_02));
io_col4_LFT I_io_00_01 ( .ceb(ceb), .sdo(sdo), .sdi(net1020),
     .spiout(spiout[1:0]), .cdone_in(cdone_in[0]),
     .spioeb(spioeb[1:0]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net1032[0:1]), .pado(net1032[0:1]), .padeb(net1033[0:1]),
     .sp4_v_t(net1034[0:15]), .sp4_h_l(SP4_h_l_01[47:0]),
     .sp12_h_l(SP12_h_l_01[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .tnl_op(rgt_op_02[7:0]),
     .lft_op(rgt_op_01[7:0]), .bnl_op(bnl_op_01[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_v_b_01[15:0]), .wl(wl[15:0]), .cf(cf_l[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_01));
io_col4_LFT I_io_00_03 ( .ceb(ceb), .sdo(net986), .sdi(net1054),
     .spiout(spiout[5:4]), .cdone_in(cdone_in[2]),
     .spioeb(spioeb[5:4]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[1:0]), .pado(pado[1:0]), .padeb(padeb[1:0]),
     .sp4_v_t(net1068[0:15]), .sp4_h_l(SP4_h_l_03[47:0]),
     .sp12_h_l(SP12_h_l_03[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[5:4]), .tnl_op(rgt_op_04[7:0]),
     .lft_op(rgt_op_03[7:0]), .bnl_op(rgt_op_02[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net1000[0:15]), .wl(wl[47:32]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_03));
io_col4_LFT I_io_00_04 ( .ceb(ceb), .sdo(net1054), .sdi(net1088),
     .spiout(spiout[7:6]), .cdone_in(cdone_in[3]),
     .spioeb(spioeb[7:6]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[3:2]), .pado(pado[3:2]), .padeb(padeb[3:2]),
     .sp4_v_t(net1102[0:15]), .sp4_h_l(SP4_h_l_04[47:0]),
     .sp12_h_l(SP12_h_l_04[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[7:6]), .tnl_op(rgt_op_05[7:0]),
     .lft_op(rgt_op_04[7:0]), .bnl_op(rgt_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net1068[0:15]), .wl(wl[63:48]), .cf(cf_l[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_04));
io_col4_LFT I_io_00_10 ( .ceb(ceb), .sdo(net646), .sdi(net1122),
     .spiout(spiout[19:18]), .cdone_in(cdone_in[9]),
     .spioeb(spioeb[19:18]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[13:12]), .pado(pado[13:12]), .padeb(padeb[13:12]),
     .sp4_v_t(net1136[0:15]), .sp4_h_l(SP4_h_l_10[47:0]),
     .sp12_h_l(SP12_h_l_10[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[19:18]), .tnl_op(rgt_op_11[7:0]),
     .lft_op(rgt_op_10[7:0]), .bnl_op(rgt_op_09[7:0]),
     .pgate(pgate[159:144]), .reset(reset_b[159:144]),
     .sp4_v_b(net660[0:15]), .wl(wl[159:144]), .cf(cf_l[239:216]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[159:144]),
     .slf_op(slf_op_10[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_10));
io_col4_LFT I_io_00_11 ( .ceb(ceb), .sdo(net1122), .sdi(net1156),
     .spiout(spiout[21:20]), .cdone_in(cdone_in[10]),
     .spioeb(spioeb[21:20]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[15:14]), .pado(pado[15:14]), .padeb(padeb[15:14]),
     .sp4_v_t(net1170[0:15]), .sp4_h_l(SP4_h_l_11[47:0]),
     .sp12_h_l(SP12_h_l_11[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[21:20]), .tnl_op(rgt_op_12[7:0]),
     .lft_op(rgt_op_11[7:0]), .bnl_op(rgt_op_10[7:0]),
     .pgate(pgate[175:160]), .reset(reset_b[175:160]),
     .sp4_v_b(net1136[0:15]), .wl(wl[175:160]), .cf(cf_l[263:240]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[175:160]),
     .slf_op(slf_op_11[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_11));

endmodule
// Library - leafcell, Cell - quad_bl_ice8, View - schematic
// LAST TIME SAVED: Oct 16 14:36:40 2008
// NETLIST TIME: Nov 14 16:17:17 2008
`timescale 1ns / 1ns 

module quad_bl_ice8 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_16, carry_out_02_16,
     carry_out_03_16, carry_out_04_16, carry_out_05_16,
     carry_out_06_16, carry_out_07_16, carry_out_09_16,
     carry_out_10_16, carry_out_11_16, carry_out_12_16,
     carry_out_13_16, carry_out_14_16, carry_out_15_16,
     carry_out_16_16, ceb_o, cf_b, cf_l, fabric_out_00_15,
     fabric_out_00_16, fabric_out_16_00, hiz_b_o, mode_o, padeb_b,
     padeb_l, padin_27, padin_80, pado_b, pado_l, r_o, sdo, shift_o,
     slf_op_00_16, slf_op_01_16, slf_op_02_16, slf_op_03_16,
     slf_op_04_16, slf_op_05_16, slf_op_06_16, slf_op_07_16,
     slf_op_08_16, slf_op_09_16, slf_op_10_16, slf_op_11_16,
     slf_op_12_16, slf_op_13_16, slf_op_14_16, slf_op_15_16,
     slf_op_16_00, slf_op_16_01, slf_op_16_02, slf_op_16_03,
     slf_op_16_04, slf_op_16_05, slf_op_16_06, slf_op_16_07,
     slf_op_16_08, slf_op_16_09, slf_op_16_10, slf_op_16_11,
     slf_op_16_12, slf_op_16_13, slf_op_16_14, slf_op_16_15,
     slf_op_16_16, spi_ss_in_l, tclk_o, update_o, bl, pgate_l, reset_l,
     sp4_h_r_16_00, sp4_h_r_16_01, sp4_h_r_16_02, sp4_h_r_16_03,
     sp4_h_r_16_04, sp4_h_r_16_05, sp4_h_r_16_06, sp4_h_r_16_07,
     sp4_h_r_16_08, sp4_h_r_16_09, sp4_h_r_16_10, sp4_h_r_16_11,
     sp4_h_r_16_12, sp4_h_r_16_13, sp4_h_r_16_14, sp4_h_r_16_15,
     sp4_h_r_16_16, sp4_r_v_b_16_01, sp4_r_v_b_16_02, sp4_r_v_b_16_03,
     sp4_r_v_b_16_04, sp4_r_v_b_16_05, sp4_r_v_b_16_06,
     sp4_r_v_b_16_07, sp4_r_v_b_16_08, sp4_r_v_b_16_09,
     sp4_r_v_b_16_10, sp4_r_v_b_16_11, sp4_r_v_b_16_12,
     sp4_r_v_b_16_13, sp4_r_v_b_16_14, sp4_r_v_b_16_15,
     sp4_r_v_b_16_16, sp4_v_t_00_16, sp4_v_t_01_16, sp4_v_t_02_16,
     sp4_v_t_03_16, sp4_v_t_04_16, sp4_v_t_05_16, sp4_v_t_06_16,
     sp4_v_t_07_16, sp4_v_t_08_16, sp4_v_t_09_16, sp4_v_t_10_16,
     sp4_v_t_11_16, sp4_v_t_12_16, sp4_v_t_13_16, sp4_v_t_14_16,
     sp4_v_t_15_16, sp4_v_t_16_16, sp12_h_r_16_01, sp12_h_r_16_02,
     sp12_h_r_16_03, sp12_h_r_16_04, sp12_h_r_16_05, sp12_h_r_16_06,
     sp12_h_r_16_07, sp12_h_r_16_08, sp12_h_r_16_09, sp12_h_r_16_10,
     sp12_h_r_16_11, sp12_h_r_16_12, sp12_h_r_16_13, sp12_h_r_16_14,
     sp12_h_r_16_15, sp12_h_r_16_16, sp12_v_t_01_16, sp12_v_t_02_16,
     sp12_v_t_03_16, sp12_v_t_04_16, sp12_v_t_05_16, sp12_v_t_06_16,
     sp12_v_t_07_16, sp12_v_t_08_16, sp12_v_t_09_16, sp12_v_t_10_16,
     sp12_v_t_11_16, sp12_v_t_12_16, sp12_v_t_13_16, sp12_v_t_14_16,
     sp12_v_t_15_16, sp12_v_t_16_16, vdd_cntl_l, wl_l, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnr_op_16_01,
     bs_en_i, ceb_i, end_of_startup_lft_b, glb_in, hiz_b_i, hold_b_l,
     hold_l_b, mode_i, padin_b, padin_l, prog, purst, r_i,
     rgt_op_16_01, rgt_op_16_02, rgt_op_16_03, rgt_op_16_04,
     rgt_op_16_05, rgt_op_16_06, rgt_op_16_07, rgt_op_16_08,
     rgt_op_16_09, rgt_op_16_10, rgt_op_16_11, rgt_op_16_12,
     rgt_op_16_13, rgt_op_16_14, rgt_op_16_15, rgt_op_16_16, sdi,
     shift_i, spioeb_l, spiout_l, tclk_i, tiegnd, tievdd, tnl_op_01_16,
     tnl_op_02_16, tnl_op_03_16, tnl_op_04_16, tnl_op_05_16,
     tnl_op_06_16, tnl_op_07_16, tnl_op_08_16, tnl_op_09_16,
     tnl_op_10_16, tnl_op_11_16, tnl_op_12_16, tnl_op_13_16,
     tnl_op_14_16, tnl_op_15_16, tnl_op_16_16, tnr_op_00_16,
     tnr_op_01_16, tnr_op_02_16, tnr_op_03_16, tnr_op_04_16,
     tnr_op_05_16, tnr_op_06_16, tnr_op_07_16, tnr_op_08_16,
     tnr_op_09_16, tnr_op_10_16, tnr_op_11_16, tnr_op_12_16,
     tnr_op_13_16, tnr_op_14_16, tnr_op_15_16, tnr_op_16_16,
     top_op_01_16, top_op_02_16, top_op_03_16, top_op_04_16,
     top_op_05_16, top_op_06_16, top_op_07_16, top_op_08_16,
     top_op_09_16, top_op_10_16, top_op_11_16, top_op_12_16,
     top_op_13_16, top_op_14_16, top_op_15_16, top_op_16_16, update_i
     );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_01_16, carry_out_02_16,
     carry_out_03_16, carry_out_04_16, carry_out_05_16,
     carry_out_06_16, carry_out_07_16, carry_out_09_16,
     carry_out_10_16, carry_out_11_16, carry_out_12_16,
     carry_out_13_16, carry_out_14_16, carry_out_15_16,
     carry_out_16_16, ceb_o, fabric_out_00_15, fabric_out_00_16,
     fabric_out_16_00, hiz_b_o, mode_o, padin_27, padin_80, r_o, sdo,
     shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, ceb_i, hiz_b_i, hold_b_l, hold_l_b,
     mode_i, prog, purst, r_i, sdi, shift_i, tclk_i, tiegnd, tievdd,
     update_i;

output [1:0]  bm_sweb_o;
output [7:0]  slf_op_13_16;
output [7:0]  slf_op_10_16;
output [7:0]  slf_op_07_16;
output [7:0]  slf_op_16_11;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_16_04;
output [7:0]  slf_op_02_16;
output [7:0]  slf_op_09_16;
output [7:0]  slf_op_16_15;
output [23:0]  padeb_l;
output [7:0]  slf_op_01_16;
output [7:0]  slf_op_08_16;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_05_16;
output [1:0]  bm_sdi_o;
output [7:0]  slf_op_11_16;
output [7:0]  slf_op_16_05;
output [7:0]  slf_op_16_06;
output [7:0]  slf_op_16_01;
output [7:0]  slf_op_03_16;
output [29:0]  pado_b;
output [7:0]  slf_op_16_08;
output [29:0]  padeb_b;
output [7:0]  slf_op_16_03;
output [7:0]  slf_op_16_14;
output [1:0]  bm_sclkrw_o;
output [31:0]  spi_ss_in_l;
output [383:0]  cf_b;
output [7:0]  slf_op_16_07;
output [383:0]  cf_l;
output [3:0]  slf_op_16_00;
output [3:0]  slf_op_00_16;
output [7:0]  slf_op_14_16;
output [7:0]  slf_op_06_16;
output [7:0]  slf_op_12_16;
output [7:0]  slf_op_16_02;
output [7:0]  slf_op_04_16;
output [7:0]  slf_op_16_12;
output [7:0]  slf_op_15_16;
output [23:0]  pado_l;
output [7:0]  slf_op_16_09;
output [7:0]  slf_op_16_10;
output [7:0]  slf_op_16_16;
output [7:0]  slf_op_16_13;

inout [47:0]  sp4_h_r_16_09;
inout [23:0]  sp12_h_r_16_14;
inout [47:0]  sp4_h_r_16_14;
inout [47:0]  sp4_r_v_b_16_09;
inout [23:0]  sp12_h_r_16_09;
inout [47:0]  sp4_h_r_16_01;
inout [47:0]  sp4_r_v_b_16_02;
inout [47:0]  sp4_v_t_06_16;
inout [23:0]  sp12_v_t_06_16;
inout [23:0]  sp12_h_r_16_16;
inout [23:0]  sp12_h_r_16_06;
inout [47:0]  sp4_r_v_b_16_16;
inout [23:0]  sp12_v_t_09_16;
inout [47:0]  sp4_v_t_04_16;
inout [47:0]  sp4_r_v_b_16_13;
inout [47:0]  sp4_r_v_b_16_08;
inout [23:0]  sp12_v_t_03_16;
inout [15:0]  sp4_v_t_00_16;
inout [47:0]  sp4_r_v_b_16_11;
inout [47:0]  sp4_v_t_15_16;
inout [47:0]  sp4_h_r_16_08;
inout [47:0]  sp4_v_t_03_16;
inout [47:0]  sp4_r_v_b_16_15;
inout [23:0]  sp12_v_t_01_16;
inout [47:0]  sp4_r_v_b_16_03;
inout [47:0]  sp4_v_t_14_16;
inout [47:0]  sp4_h_r_16_12;
inout [47:0]  sp4_v_t_11_16;
inout [47:0]  sp4_v_t_01_16;
inout [23:0]  sp12_v_t_07_16;
inout [47:0]  sp4_h_r_16_15;
inout [47:0]  sp4_r_v_b_16_01;
inout [23:0]  sp12_h_r_16_08;
inout [23:0]  sp12_h_r_16_05;
inout [23:0]  sp12_v_t_15_16;
inout [47:0]  sp4_v_t_12_16;
inout [23:0]  sp12_v_t_05_16;
inout [23:0]  sp12_h_r_16_03;
inout [23:0]  sp12_h_r_16_04;
inout [23:0]  sp12_h_r_16_13;
inout [47:0]  sp4_r_v_b_16_04;
inout [23:0]  sp12_h_r_16_12;
inout [47:0]  sp4_h_r_16_13;
inout [271:0]  pgate_l;
inout [23:0]  sp12_v_t_12_16;
inout [47:0]  sp4_h_r_16_16;
inout [47:0]  sp4_h_r_16_02;
inout [47:0]  sp4_r_v_b_16_06;
inout [47:0]  sp4_h_r_16_10;
inout [23:0]  sp12_h_r_16_15;
inout [47:0]  sp4_h_r_16_06;
inout [23:0]  sp12_v_t_14_16;
inout [23:0]  sp12_h_r_16_10;
inout [47:0]  sp4_v_t_13_16;
inout [47:0]  sp4_r_v_b_16_12;
inout [23:0]  sp12_v_t_16_16;
inout [23:0]  sp12_v_t_10_16;
inout [47:0]  sp4_h_r_16_03;
inout [47:0]  sp4_v_t_02_16;
inout [271:0]  wl_l;
inout [271:0]  reset_l;
inout [47:0]  sp4_h_r_16_07;
inout [23:0]  sp12_v_t_11_16;
inout [271:0]  vdd_cntl_l;
inout [47:0]  sp4_h_r_16_04;
inout [23:0]  sp12_h_r_16_02;
inout [23:0]  sp12_h_r_16_11;
inout [869:0]  bl;
inout [47:0]  sp4_h_r_16_05;
inout [23:0]  sp12_v_t_08_16;
inout [47:0]  sp4_v_t_16_16;
inout [47:0]  sp4_v_t_10_16;
inout [47:0]  sp4_r_v_b_16_14;
inout [47:0]  sp4_v_t_05_16;
inout [47:0]  sp4_v_t_07_16;
inout [23:0]  sp12_v_t_13_16;
inout [47:0]  sp4_r_v_b_16_07;
inout [47:0]  sp4_v_t_08_16;
inout [47:0]  sp4_r_v_b_16_10;
inout [15:0]  sp4_h_r_16_00;
inout [23:0]  sp12_v_t_04_16;
inout [47:0]  sp4_v_t_09_16;
inout [23:0]  sp12_h_r_16_01;
inout [23:0]  sp12_h_r_16_07;
inout [47:0]  sp4_r_v_b_16_05;
inout [23:0]  sp12_v_t_02_16;
inout [47:0]  sp4_h_r_16_11;

input [31:0]  spiout_l;
input [7:0]  rgt_op_16_15;
input [7:0]  top_op_09_16;
input [7:0]  glb_in;
input [7:0]  tnl_op_07_16;
input [7:0]  tnl_op_05_16;
input [1:0]  bm_sdo_i;
input [7:0]  tnl_op_01_16;
input [7:0]  tnr_op_15_16;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_06_16;
input [7:0]  tnr_op_02_16;
input [1:0]  bm_sdi_i;
input [31:0]  spioeb_l;
input [7:0]  top_op_03_16;
input [7:0]  rgt_op_16_05;
input [7:0]  tnr_op_04_16;
input [7:0]  tnl_op_08_16;
input [7:0]  tnr_op_14_16;
input [7:0]  rgt_op_16_11;
input [7:0]  top_op_10_16;
input [7:0]  top_op_01_16;
input [7:0]  top_op_04_16;
input [7:0]  tnr_op_06_16;
input [7:0]  tnl_op_03_16;
input [7:0]  tnr_op_00_16;
input [7:0]  rgt_op_16_09;
input [7:0]  tnl_op_09_16;
input [7:0]  top_op_12_16;
input [1:0]  bm_sclkrw_i;
input [7:0]  top_op_02_16;
input [7:0]  tnl_op_10_16;
input [7:0]  top_op_16_16;
input [7:0]  rgt_op_16_06;
input [7:0]  tnl_op_14_16;
input [1:0]  bm_sweb_i;
input [7:0]  rgt_op_16_10;
input [7:0]  tnr_op_01_16;
input [7:0]  tnr_op_12_16;
input [16:1]  end_of_startup_lft_b;
input [7:0]  tnl_op_02_16;
input [7:0]  rgt_op_16_13;
input [7:0]  rgt_op_16_08;
input [7:0]  top_op_14_16;
input [7:0]  tnr_op_05_16;
input [7:0]  tnr_op_08_16;
input [7:0]  top_op_08_16;
input [7:0]  top_op_13_16;
input [7:0]  tnl_op_16_16;
input [23:0]  padin_l;
input [7:0]  tnr_op_13_16;
input [7:0]  rgt_op_16_01;
input [7:0]  top_op_11_16;
input [7:0]  tnl_op_15_16;
input [7:0]  tnl_op_12_16;
input [3:0]  bnr_op_16_01;
input [7:0]  rgt_op_16_07;
input [7:0]  tnl_op_11_16;
input [7:0]  rgt_op_16_02;
input [7:0]  rgt_op_16_14;
input [7:0]  tnl_op_13_16;
input [7:0]  tnr_op_03_16;
input [7:0]  tnr_op_11_16;
input [7:0]  top_op_15_16;
input [7:0]  rgt_op_16_03;
input [7:0]  tnr_op_07_16;
input [7:0]  tnr_op_10_16;
input [7:0]  rgt_op_16_16;
input [7:0]  tnr_op_09_16;
input [7:0]  rgt_op_16_12;
input [29:0]  padin_b;
input [7:0]  top_op_07_16;
input [7:0]  top_op_06_16;
input [7:0]  tnl_op_04_16;
input [7:0]  rgt_op_16_04;
input [7:0]  top_op_05_16;
input [7:0]  tnr_op_16_16;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:47]  net4199;

wire  [0:47]  net4005;

wire  [0:47]  net3463;

wire  [0:7]  net4912;

wire  [0:23]  net2406;

wire  [0:7]  net4920;

wire  [0:47]  net3186;

wire  [0:7]  net4669;

wire  [0:7]  net3206;

wire  [0:7]  net2260;

wire  [0:47]  net4850;

wire  [0:47]  net4037;

wire  [0:7]  net2815;

wire  [0:47]  net2694;

wire  [0:23]  net4893;

wire  [0:7]  net4674;

wire  [0:23]  net4632;

wire  [0:23]  net2278;

wire  [0:47]  net2313;

wire  [0:47]  net4898;

wire  [0:7]  net4807;

wire  [0:23]  net3225;

wire  [0:23]  net3983;

wire  [0:7]  net3962;

wire  [0:47]  net4442;

wire  [0:7]  net3533;

wire  [0:7]  net2222;

wire  [0:47]  net3433;

wire  [0:23]  net2736;

wire  [0:47]  net3183;

wire  [0:47]  net3185;

wire  [0:23]  net2408;

wire  [0:23]  net4082;

wire  [0:23]  net2933;

wire  [0:7]  net3242;

wire  [0:47]  net4090;

wire  [0:7]  net2326;

wire  [0:47]  net2121;

wire  [0:47]  net4195;

wire  [0:23]  net2670;

wire  [0:47]  net3925;

wire  [0:47]  net3660;

wire  [0:47]  net4584;

wire  [0:7]  net4766;

wire  [0:47]  net4497;

wire  [0:47]  net4900;

wire  [0:47]  net4948;

wire  [0:23]  net3817;

wire  [0:23]  net4931;

wire  [0:47]  net3346;

wire  [0:47]  net4860;

wire  [0:47]  net3005;

wire  [0:47]  net3624;

wire  [0:23]  net2343;

wire  [0:7]  net4062;

wire  [0:23]  net2344;

wire  [0:47]  net4938;

wire  [0:7]  net4760;

wire  [0:47]  net2124;

wire  [0:47]  net3434;

wire  [0:47]  net3824;

wire  [0:7]  net4126;

wire  [0:7]  net4799;

wire  [0:47]  net4498;

wire  [0:7]  net3367;

wire  [0:23]  net4081;

wire  [0:23]  net2769;

wire  [0:7]  net3145;

wire  [0:23]  net2835;

wire  [0:7]  net3634;

wire  [0:47]  net2558;

wire  [0:47]  net2838;

wire  [0:47]  net2942;

wire  [0:47]  net3764;

wire  [0:47]  net2395;

wire  [0:47]  net3541;

wire  [0:47]  net3169;

wire  [0:7]  net4764;

wire  [0:47]  net3298;

wire  [0:47]  net4585;

wire  [0:7]  net4672;

wire  [0:23]  net3164;

wire  [0:47]  net4695;

wire  [0:47]  net3546;

wire  [0:47]  net2350;

wire  [0:47]  net3049;

wire  [0:47]  net2805;

wire  [0:23]  net2178;

wire  [0:47]  net3512;

wire  [0:7]  net4763;

wire  [0:23]  net4211;

wire  [0:47]  net2366;

wire  [0:47]  net4526;

wire  [0:7]  net4515;

wire  [0:23]  net3227;

wire  [0:47]  net2890;

wire  [0:47]  net2346;

wire  [0:7]  net4517;

wire  [0:47]  net3842;

wire  [0:7]  net3310;

wire  [0:23]  net4045;

wire  [0:47]  net2640;

wire  [0:47]  net3330;

wire  [0:47]  net4481;

wire  [0:47]  net2511;

wire  [0:47]  net4154;

wire  [0:7]  net2096;

wire  [0:23]  net3391;

wire  [0:23]  net3592;

wire  [0:7]  net3042;

wire  [0:7]  net3470;

wire  [0:47]  net2182;

wire  [0:47]  net4853;

wire  [0:7]  net2162;

wire  [0:47]  net4903;

wire  [0:7]  net4909;

wire  [0:23]  net4641;

wire  [0:23]  net4924;

wire  [0:23]  net3061;

wire  [0:23]  net2902;

wire  [0:47]  net2777;

wire  [0:47]  net3601;

wire  [0:47]  net3002;

wire  [0:47]  net4088;

wire  [0:23]  net4830;

wire  [0:23]  net3883;

wire  [0:47]  net2530;

wire  [0:7]  net3898;

wire  [0:47]  net3673;

wire  [0:47]  net4689;

wire  [0:47]  net2560;

wire  [0:47]  net3767;

wire  [0:47]  net3295;

wire  [0:47]  net2723;

wire  [0:47]  net2971;

wire  [0:47]  net4116;

wire  [0:7]  net4761;

wire  [0:47]  net2474;

wire  [0:23]  net4474;

wire  [0:23]  net3229;

wire  [0:47]  net4848;

wire  [0:47]  net3627;

wire  [0:47]  net2347;

wire  [0:7]  net3530;

wire  [0:23]  net2999;

wire  [0:47]  net2515;

wire  [0:7]  net2432;

wire  [0:7]  net3966;

wire  [0:47]  net4683;

wire  [0:23]  net2996;

wire  [0:7]  net4072;

wire  [0:7]  net4129;

wire  [0:47]  net3513;

wire  [0:47]  net2781;

wire  [0:7]  net4456;

wire  [0:47]  net2858;

wire  [0:23]  net2833;

wire  [0:23]  net4048;

wire  [0:23]  net2991;

wire  [0:47]  net4004;

wire  [0:23]  net3918;

wire  [0:47]  net2454;

wire  [0:7]  net4455;

wire  [0:47]  net3707;

wire  [0:47]  net2562;

wire  [0:7]  net2327;

wire  [0:47]  net4577;

wire  [0:47]  net3761;

wire  [0:7]  net4810;

wire  [0:23]  net2898;

wire  [0:47]  net2200;

wire  [0:23]  net2836;

wire  [0:47]  net3350;

wire  [0:47]  net3931;

wire  [0:23]  net3492;

wire  [0:47]  net3381;

wire  [0:7]  net2981;

wire  [0:47]  net3436;

wire  [0:47]  net2361;

wire  [0:7]  net4801;

wire  [0:47]  net4851;

wire  [0:23]  net3390;

wire  [0:7]  net3146;

wire  [0:23]  net2442;

wire  [0:47]  net4201;

wire  [0:47]  net4494;

wire  [0:47]  net2940;

wire  [0:7]  net4187;

wire  [0:23]  net3886;

wire  [0:23]  net3881;

wire  [0:23]  net4932;

wire  [0:47]  net3382;

wire  [0:47]  net2693;

wire  [0:47]  net4157;

wire  [0:47]  net4901;

wire  [0:47]  net2125;

wire  [0:7]  net3205;

wire  [0:7]  net4805;

wire  [0:23]  net3656;

wire  [0:23]  net3328;

wire  [0:47]  net4681;

wire  [0:47]  net3213;

wire  [0:47]  net4856;

wire  [0:47]  net3603;

wire  [0:23]  net4476;

wire  [0:23]  net4829;

wire  [0:23]  net4139;

wire  [0:7]  net2982;

wire  [0:47]  net2186;

wire  [0:47]  net2452;

wire  [0:7]  net2760;

wire  [0:23]  net3326;

wire  [0:47]  net2291;

wire  [0:47]  net3788;

wire  [0:47]  net3597;

wire  [0:7]  net3472;

wire  [0:7]  net4752;

wire  [0:47]  net3345;

wire  [0:47]  net4160;

wire  [0:47]  net4118;

wire  [0:47]  net4423;

wire  [0:47]  net2724;

wire  [0:47]  net3706;

wire  [0:47]  net3331;

wire  [0:47]  net3825;

wire  [0:47]  net4899;

wire  [0:7]  net4754;

wire  [0:47]  net4688;

wire  [0:7]  net4064;

wire  [0:47]  net3104;

wire  [0:7]  net2878;

wire  [0:47]  net3823;

wire  [0:7]  net3744;

wire  [0:47]  net4422;

wire  [0:23]  net3652;

wire  [0:23]  net4084;

wire  [0:47]  net4447;

wire  [0:47]  net2476;

wire  [0:47]  net4573;

wire  [0:23]  net4209;

wire  [0:23]  net3753;

wire  [0:47]  net2726;

wire  [0:47]  net2514;

wire  [0:7]  net3204;

wire  [0:47]  net3787;

wire  [0:47]  net3870;

wire  [0:23]  net3394;

wire  [0:47]  net2616;

wire  [0:23]  net4212;

wire  [0:47]  net4587;

wire  [0:47]  net4165;

wire  [0:23]  net4928;

wire  [0:23]  net4923;

wire  [0:23]  net3489;

wire  [0:47]  net3273;

wire  [0:7]  net3408;

wire  [0:47]  net4001;

wire  [0:7]  net2486;

wire  [0:23]  net3553;

wire  [0:47]  net3674;

wire  [3:0]  slf_op_00_01;

wire  [3:0]  slf_op_00_07;

wire  [0:47]  net2148;

wire  [3:0]  slf_op_00_03;

wire  [0:47]  net3462;

wire  [0:47]  net3432;

wire  [0:47]  net4151;

wire  [0:7]  net3531;

wire  [0:7]  net4914;

wire  [0:7]  net4024;

wire  [0:23]  net4542;

wire  [0:7]  net2914;

wire  [0:23]  net3820;

wire  [0:7]  net3088;

wire  [0:23]  net3556;

wire  [0:23]  net4841;

wire  [0:7]  net4916;

wire  [0:47]  net3216;

wire  [0:47]  net4846;

wire  [0:7]  net4755;

wire  [0:7]  net3862;

wire  [0:47]  net3018;

wire  [0:47]  net3827;

wire  [0:47]  net3052;

wire  [0:23]  net4842;

wire  [0:47]  net3622;

wire  [0:7]  net2814;

wire  [0:47]  net3661;

wire  [0:7]  net3078;

wire  [0:7]  net4759;

wire  [0:7]  net3473;

wire  [0:47]  net3333;

wire  [0:47]  net3678;

wire  [0:23]  net2241;

wire  [0:47]  net2126;

wire  [0:47]  net4170;

wire  [0:47]  net2398;

wire  [0:47]  net4684;

wire  [0:47]  net3871;

wire  [0:23]  net4838;

wire  [0:23]  net4146;

wire  [0:47]  net2802;

wire  [0:7]  net3963;

wire  [0:7]  net4883;

wire  [0:47]  net3987;

wire  [0:47]  net4527;

wire  [0:47]  net2677;

wire  [0:7]  net4130;

wire  [0:23]  net3063;

wire  [0:47]  net2310;

wire  [0:7]  net3369;

wire  [0:7]  net3534;

wire  [0:47]  net3596;

wire  [0:47]  net3498;

wire  [0:23]  net4473;

wire  [0:47]  net3053;

wire  [0:47]  net2455;

wire  [0:47]  net2453;

wire  [0:47]  net4105;

wire  [0:7]  net2817;

wire  [0:7]  net2490;

wire  [0:47]  net2691;

wire  [0:23]  net2936;

wire  [0:7]  net4806;

wire  [0:47]  net2314;

wire  [0:47]  net4158;

wire  [0:47]  net2968;

wire  [0:47]  net3348;

wire  [0:47]  net3110;

wire  [0:23]  net2998;

wire  [0:23]  net2444;

wire  [0:47]  net3297;

wire  [0:47]  net4167;

wire  [0:47]  net2941;

wire  [0:47]  net3499;

wire  [0:47]  net3928;

wire  [0:47]  net3299;

wire  [0:47]  net4033;

wire  [0:47]  net4006;

wire  [0:23]  net4935;

wire  [0:47]  net2396;

wire  [0:7]  net4765;

wire  [0:7]  net3964;

wire  [0:23]  net4412;

wire  [0:47]  net3132;

wire  [0:47]  net4198;

wire  [0:7]  net4186;

wire  [0:47]  net2290;

wire  [0:23]  net2504;

wire  [0:47]  net4445;

wire  [0:23]  net4831;

wire  [0:7]  net4666;

wire  [0:7]  net2220;

wire  [0:47]  net3708;

wire  [0:47]  net3184;

wire  [0:23]  net4933;

wire  [0:47]  net4528;

wire  [0:23]  net3160;

wire  [0:7]  net3475;

wire  [0:47]  net3438;

wire  [0:7]  net4905;

wire  [0:7]  net4128;

wire  [0:7]  net4026;

wire  [0:47]  net4576;

wire  [0:23]  net3818;

wire  [0:23]  net2506;

wire  [0:47]  net2967;

wire  [0:23]  net3097;

wire  [0:23]  net3819;

wire  [0:47]  net3869;

wire  [0:47]  net4117;

wire  [0:7]  net3858;

wire  [0:7]  net2488;

wire  [0:47]  net2183;

wire  [0:7]  net4458;

wire  [0:47]  net3494;

wire  [0:23]  net4472;

wire  [0:23]  net3098;

wire  [0:47]  net2722;

wire  [0:47]  net4952;

wire  [0:23]  net4621;

wire  [0:47]  net2230;

wire  [0:23]  net2834;

wire  [0:23]  net2573;

wire  [0:47]  net3272;

wire  [0:23]  net4633;

wire  [0:23]  net4636;

wire  [0:23]  net4832;

wire  [0:47]  net4035;

wire  [0:47]  net2725;

wire  [0:47]  net2855;

wire  [0:23]  net4638;

wire  [0:47]  net4444;

wire  [0:7]  net4459;

wire  [0:47]  net4155;

wire  [0:47]  net2393;

wire  [0:47]  net4849;

wire  [0:47]  net4583;

wire  [0:7]  net3694;

wire  [0:23]  net2409;

wire  [0:47]  net3837;

wire  [0:47]  net4034;

wire  [0:47]  net2526;

wire  [0:47]  net2149;

wire  [0:23]  net3882;

wire  [0:23]  net4835;

wire  [0:47]  net3181;

wire  [0:47]  net2311;

wire  [0:47]  net2397;

wire  [0:23]  net3647;

wire  [0:47]  net3050;

wire  [0:47]  net3790;

wire  [0:7]  net2487;

wire  [0:47]  net3294;

wire  [0:23]  net2180;

wire  [0:23]  net4538;

wire  [0:47]  net2561;

wire  [0:23]  net2570;

wire  [0:7]  net3471;

wire  [0:7]  net4758;

wire  [0:7]  net4022;

wire  [0:47]  net2803;

wire  [0:23]  net3655;

wire  [0:7]  net3800;

wire  [0:7]  net3734;

wire  [0:7]  net4664;

wire  [0:7]  net3041;

wire  [0:47]  net4496;

wire  [0:47]  net2853;

wire  [0:47]  net2559;

wire  [0:47]  net2202;

wire  [0:47]  net4152;

wire  [0:23]  net3590;

wire  [0:23]  net2572;

wire  [0:23]  net2897;

wire  [0:23]  net3066;

wire  [0:7]  net3965;

wire  [0:47]  net4692;

wire  [0:47]  net3990;

wire  [0:23]  net2771;

wire  [0:7]  net3801;

wire  [0:23]  net3488;

wire  [0:47]  net2151;

wire  [0:7]  net2158;

wire  [0:23]  net2832;

wire  [0:23]  net4537;

wire  [0:7]  net3803;

wire  [0:7]  net2268;

wire  [0:7]  net2325;

wire  [0:23]  net2441;

wire  [0:23]  net2901;

wire  [0:23]  net2663;

wire  [0:7]  net3203;

wire  [0:47]  net3988;

wire  [0:23]  net2243;

wire  [0:47]  net4095;

wire  [0:47]  net3296;

wire  [0:47]  net2839;

wire  [0:23]  net4922;

wire  [0:7]  net3900;

wire  [0:47]  net4682;

wire  [0:23]  net2772;

wire  [0:23]  net3263;

wire  [0:47]  net2201;

wire  [0:47]  net2889;

wire  [0:47]  net3926;

wire  [0:47]  net2885;

wire  [0:23]  net4145;

wire  [0:23]  net2507;

wire  [0:23]  net2279;

wire  [0:47]  net3275;

wire  [0:47]  net2315;

wire  [0:7]  net2546;

wire  [0:47]  net4589;

wire  [0:47]  net3269;

wire  [0:47]  net4950;

wire  [0:47]  net4094;

wire  [0:47]  net3497;

wire  [0:23]  net4050;

wire  [0:7]  net4676;

wire  [0:47]  net4529;

wire  [0:47]  net4416;

wire  [0:47]  net2232;

wire  [0:23]  net2900;

wire  [0:23]  net2607;

wire  [0:47]  net4579;

wire  [0:47]  net3544;

wire  [7:0]  clk_tree_drv;

wire  [0:47]  net4119;

wire  [0:47]  net2364;

wire  [0:7]  net4390;

wire  [0:47]  net2857;

wire  [0:47]  net3130;

wire  [0:23]  net3491;

wire  [0:7]  net4911;

wire  [0:47]  net2612;

wire  [0:7]  net3142;

wire  [0:7]  net3416;

wire  [0:47]  net3459;

wire  [0:23]  net4467;

wire  [0:47]  net2231;

wire  [0:7]  net3406;

wire  [0:7]  net3908;

wire  [0:7]  net4753;

wire  [0:23]  net3721;

wire  [0:47]  net4161;

wire  [3:0]  slf_op_01_00;

wire  [3:0]  slf_op_13_00;

wire  [0:7]  net3144;

wire  [0:47]  net3929;

wire  [0:47]  net3105;

wire  [3:0]  slf_op_15_00;

wire  [3:0]  slf_op_10_00;

wire  [3:0]  slf_op_03_00;

wire  [3:0]  slf_op_07_00;

wire  [3:0]  slf_op_09_00;

wire  [3:0]  slf_op_00_11;

wire  [3:0]  slf_op_00_14;

wire  [3:0]  slf_op_00_13;

wire  [3:0]  slf_op_00_09;

wire  [3:0]  slf_op_00_12;

wire  [3:0]  slf_op_00_04;

wire  [3:0]  slf_op_00_15;

wire  [3:0]  slf_op_00_05;

wire  [3:0]  slf_op_00_06;

wire  [0:23]  net3754;

wire  [0:7]  net2159;

wire  [0:47]  net3950;

wire  [3:0]  slf_op_00_02;

wire  [0:47]  net2234;

wire  [0:23]  net4148;

wire  [0:7]  net3696;

wire  [0:23]  net3327;

wire  [0:7]  net3202;

wire  [3:0]  slf_op_05_00;

wire  [3:0]  slf_op_02_00;

wire  [3:0]  slf_op_00_08;

wire  [3:0]  slf_op_00_10;

wire  [0:7]  net4919;

wire  [0:23]  net4927;

wire  [0:47]  net2944;

wire  [0:47]  net3051;

wire  [0:47]  net3658;

wire  [0:47]  net3134;

wire  [0:47]  net3510;

wire  [3:0]  slf_op_04_00;

wire  [3:0]  slf_op_08_00;

wire  [3:0]  slf_op_12_00;

wire  [3:0]  slf_op_14_00;

wire  [3:0]  slf_op_11_00;

wire  [3:0]  slf_op_06_00;

wire  [0:47]  net4418;

wire  [0:47]  net3677;

wire  [0:7]  net4751;

wire  [0:7]  net4800;

wire  [0:7]  net2816;

wire  [0:47]  net2678;

wire  [0:23]  net2735;

wire  [0:47]  net3765;

wire  [0:47]  net2479;

wire  [0:23]  net2899;

wire  [0:23]  net3920;

wire  [0:47]  net3705;

wire  [0:7]  net3307;

wire  [0:47]  net3675;

wire  [0:47]  net2528;

wire  [0:47]  net2614;

wire  [0:23]  net3000;

wire  [0:47]  net4169;

wire  [0:47]  net4694;

wire  [0:23]  net4837;

wire  [0:23]  net3654;

wire  [0:23]  net3228;

wire  [0:47]  net4089;

wire  [0:47]  net3600;

wire  [0:47]  net3131;

wire  [0:47]  net2692;

wire  [0:47]  net3171;

wire  [0:47]  net3270;

wire  [0:7]  net2980;

wire  [0:47]  net2842;

wire  [0:7]  net4803;

wire  [0:47]  net3268;

wire  [0:47]  net2120;

wire  [0:23]  net2280;

wire  [0:47]  net3274;

wire  [0:47]  net2966;

wire  [0:23]  net2113;

wire  [0:47]  net3214;

wire  [0:23]  net2669;

wire  [0:23]  net2571;

wire  [0:7]  net2877;

wire  [0:7]  net3861;

wire  [0:47]  net3020;

wire  [0:47]  net3439;

wire  [0:47]  net4847;

wire  [0:47]  net4443;

wire  [0:23]  net3483;

wire  [0:23]  net2179;

wire  [0:47]  net2284;

wire  [0:47]  net2639;

wire  [0:47]  net2197;

wire  [0:7]  net4804;

wire  [0:23]  net3884;

wire  [0:23]  net2340;

wire  [0:23]  net4637;

wire  [0:47]  net3840;

wire  [0:23]  net3557;

wire  [0:47]  net2478;

wire  [0:7]  net4514;

wire  [0:47]  net2365;

wire  [0:47]  net2289;

wire  [0:23]  net2114;

wire  [0:7]  net2322;

wire  [0:47]  net3106;

wire  [0:23]  net2171;

wire  [0:7]  net4665;

wire  [0:47]  net4104;

wire  [0:7]  net2916;

wire  [0:47]  net4685;

wire  [0:23]  net4834;

wire  [0:47]  net3991;

wire  [0:23]  net2246;

wire  [0:47]  net3762;

wire  [0:47]  net2362;

wire  [0:7]  net3370;

wire  [0:47]  net4530;

wire  [0:47]  net2840;

wire  [0:7]  net3638;

wire  [0:23]  net2245;

wire  [0:7]  net4811;

wire  [0:7]  net4797;

wire  [0:47]  net3108;

wire  [0:23]  net2606;

wire  [0:47]  net2689;

wire  [0:47]  net4192;

wire  [0:47]  net2184;

wire  [0:47]  net2690;

wire  [0:23]  net2508;

wire  [0:23]  net3554;

wire  [0:23]  net3980;

wire  [0:47]  net2886;

wire  [0:47]  net3839;

wire  [0:47]  net4446;

wire  [0:23]  net4833;

wire  [0:47]  net3542;

wire  [0:7]  net2978;

wire  [0:23]  net3811;

wire  [0:23]  net2505;

wire  [0:23]  net4475;

wire  [0:7]  net4809;

wire  [0:7]  net2752;

wire  [0:7]  net2382;

wire  [0:47]  net3509;

wire  [0:23]  net3325;

wire  [0:23]  net3155;

wire  [0:47]  net2122;

wire  [0:47]  net2619;

wire  [0:47]  net3019;

wire  [0:23]  net3389;

wire  [0:23]  net4635;

wire  [0:47]  net3511;

wire  [0:47]  net2642;

wire  [0:23]  net3162;

wire  [0:23]  net4926;

wire  [0:23]  net4214;

wire  [0:47]  net2843;

wire  [0:23]  net3065;

wire  [0:7]  net4802;

wire  [0:47]  net2199;

wire  [0:23]  net2407;

wire  [0:23]  net3490;

wire  [0:47]  net3109;

wire  [0:7]  net2874;

wire  [0:23]  net3099;

wire  [0:23]  net3717;

wire  [0:23]  net3722;

wire  [0:7]  net3636;

wire  [0:23]  net3062;

wire  [0:47]  net4417;

wire  [0:47]  net2782;

wire  [0:47]  net3460;

wire  [0:47]  net2198;

wire  [0:47]  net4482;

wire  [0:47]  net3662;

wire  [0:47]  net3182;

wire  [0:7]  net3639;

wire  [0:23]  net3425;

wire  [0:47]  net3461;

wire  [0:7]  net3244;

wire  [0:47]  net2512;

wire  [0:23]  net4622;

wire  [0:7]  net4756;

wire  [0:47]  net2946;

wire  [0:47]  net3826;

wire  [0:7]  net2323;

wire  [0:47]  net3989;

wire  [0:7]  net4025;

wire  [0:7]  net3859;

wire  [0:23]  net2733;

wire  [0:7]  net4808;

wire  [0:47]  net3514;

wire  [0:23]  net2410;

wire  [0:23]  net3982;

wire  [0:47]  net3017;

wire  [0:47]  net2288;

wire  [0:47]  net3347;

wire  [0:47]  net4197;

wire  [0:47]  net3133;

wire  [0:47]  net3766;

wire  [0:7]  net3080;

wire  [0:23]  net3226;

wire  [0:47]  net2721;

wire  [0:47]  net2617;

wire  [0:47]  net3874;

wire  [0:23]  net3981;

wire  [0:7]  net2491;

wire  [0:47]  net2285;

wire  [0:47]  net3602;

wire  [0:23]  net2734;

wire  [0:23]  net4843;

wire  [0:47]  net2841;

wire  [0:23]  net2335;

wire  [0:23]  net3064;

wire  [0:47]  net3930;

wire  [0:23]  net3720;

wire  [0:23]  net3392;

wire  [0:47]  net2856;

wire  [0:47]  net2854;

wire  [0:7]  net4454;

wire  [0:47]  net2348;

wire  [0:47]  net2187;

wire  [0:47]  net3335;

wire  [0:23]  net4844;

wire  [0:23]  net3426;

wire  [0:47]  net4582;

wire  [0:23]  net3816;

wire  [0:47]  net3952;

wire  [0:47]  net4845;

wire  [0:47]  net4194;

wire  [0:23]  net3589;

wire  [0:47]  net2525;

wire  [0:47]  net3760;

wire  [0:47]  net4687;

wire  [0:7]  net4913;

wire  [0:23]  net4925;

wire  [0:47]  net2448;

wire  [0:23]  net3324;

wire  [0:23]  net3427;

wire  [0:47]  net3986;

wire  [0:23]  net3261;

wire  [0:23]  net4046;

wire  [0:47]  net3951;

wire  [0:23]  net3163;

wire  [0:47]  net3167;

wire  [0:47]  net3625;

wire  [0:23]  net3428;

wire  [0:7]  net3039;

wire  [0:7]  net3736;

wire  [0:47]  net3111;

wire  [0:7]  net4671;

wire  [0:47]  net2613;

wire  [0:23]  net4540;

wire  [0:23]  net4049;

wire  [0:23]  net2672;

wire  [0:47]  net4478;

wire  [0:23]  net4541;

wire  [0:47]  net2638;

wire  [0:7]  net3580;

wire  [0:7]  net2219;

wire  [0:47]  net3135;

wire  [0:23]  net2997;

wire  [0:47]  net4480;

wire  [0:7]  net2422;

wire  [0:23]  net2341;

wire  [0:23]  net2668;

wire  [0:47]  net3873;

wire  [0:47]  net3659;

wire  [0:47]  net3663;

wire  [0:7]  net2550;

wire  [0:47]  net2780;

wire  [0:23]  net3718;

wire  [0:23]  net3555;

wire  [0:47]  net4191;

wire  [0:47]  net4580;

wire  [0:23]  net4411;

wire  [0:47]  net2146;

wire  [0:7]  net3038;

wire  [0:7]  net2094;

wire  [0:47]  net3378;

wire  [0:7]  net2549;

wire  [0:47]  net2449;

wire  [0:47]  net2185;

wire  [0:47]  net2970;

wire  [0:7]  net3798;

wire  [0:23]  net2935;

wire  [0:47]  net4581;

wire  [0:23]  net4210;

wire  [0:47]  net3786;

wire  [0:23]  net2934;

wire  [0:47]  net3841;

wire  [0:23]  net4639;

wire  [0:47]  net3349;

wire  [0:47]  net2618;

wire  [0:23]  net3653;

wire  [0:47]  net4483;

wire  [0:7]  net4908;

wire  [0:47]  net4586;

wire  [0:47]  net3377;

wire  [0:7]  net3697;

wire  [0:47]  net4493;

wire  [0:47]  net2229;

wire  [0:7]  net3366;

wire  [0:23]  net4625;

wire  [0:47]  net3166;

wire  [0:47]  net3022;

wire  [0:47]  net3822;

wire  [0:23]  net2737;

wire  [0:47]  net3379;

wire  [0:47]  net2557;

wire  [0:23]  net3756;

wire  [0:47]  net4588;

wire  [0:7]  net4904;

wire  [0:7]  net3572;

wire  [0:47]  net4852;

wire  [0:7]  net2218;

wire  [0:23]  net2176;

wire  [0:23]  net3984;

wire  [0:47]  net4946;

wire  [0:47]  net3003;

wire  [0:7]  net3967;

wire  [0:23]  net4561;

wire  [0:47]  net4858;

wire  [0:7]  net3570;

wire  [0:47]  net2312;

wire  [0:7]  net2383;

wire  [0:7]  net3860;

wire  [0:47]  net3217;

wire  [0:47]  net4003;

wire  [0:47]  net2778;

wire  [0:7]  net3474;

wire  [0:7]  net4663;

wire  [0:47]  net4944;

wire  [0:7]  net3635;

wire  [0:23]  net4539;

wire  [0:47]  net2349;

wire  [0:47]  net4525;

wire  [0:23]  net4929;

wire  [0:23]  net4147;

wire  [0:47]  net4196;

wire  [0:47]  net3953;

wire  [0:7]  net3040;

wire  [0:23]  net3919;

wire  [0:7]  net2384;

wire  [0:47]  net4479;

wire  [0:47]  net2475;

wire  [0:47]  net4156;

wire  [0:7]  net4400;

wire  [0:47]  net3218;

wire  [0:23]  net4839;

wire  [0:7]  net2548;

wire  [0:47]  net3543;

wire  [0:23]  net3591;

wire  [0:23]  net2605;

wire  [0:7]  net4668;

wire  [0:47]  net3006;

wire  [0:7]  net2424;

wire  [0:47]  net2641;

wire  [0:47]  net4106;

wire  [0:47]  net3954;

wire  [0:23]  net4840;

wire  [0:47]  net2643;

wire  [0:47]  net4859;

wire  [0:47]  net3437;

wire  [0:47]  net4854;

wire  [0:23]  net4410;

wire  [0:7]  net4516;

wire  [0:47]  net4115;

wire  [0:47]  net2450;

wire  [0:47]  net3004;

wire  [0:7]  net4667;

wire  [0:23]  net4626;

wire  [0:7]  net3308;

wire  [0:7]  net2221;

wire  [0:23]  net3264;

wire  [0:47]  net3623;

wire  [0:47]  net4202;

wire  [0:47]  net4168;

wire  [0:23]  net4634;

wire  [0:23]  net4047;

wire  [0:7]  net3252;

wire  [0:23]  net2770;

wire  [0:7]  net3799;

wire  [0:47]  net3054;

wire  [0:23]  net2671;

wire  [0:15]  net4910;

wire  [0:47]  net4150;

wire  [0:7]  net3695;

wire  [0:23]  net2608;

wire  [0:7]  net3306;

wire  [0:47]  net4038;

wire  [0:7]  net4189;

wire  [0:47]  net3545;

wire  [0:47]  net2351;

wire  [0:47]  net3626;

wire  [0:7]  net4127;

wire  [0:23]  net4836;

wire  [0:47]  net3676;

wire  [0:47]  net3495;

wire  [0:23]  net2277;

wire  [0:47]  net2477;

wire  [0:23]  net4144;

wire  [0:47]  net4686;

wire  [0:47]  net2675;

wire  [0:47]  net4855;

wire  [0:23]  net4934;

wire  [0:47]  net3872;

wire  [0:23]  net3885;

wire  [0:47]  net2887;

wire  [0:47]  net2676;

wire  [0:7]  net2160;

wire  [0:7]  net3698;

wire  [0:23]  net3975;

wire  [0:47]  net4495;

wire  [0:47]  net4200;

wire  [0:23]  net4083;

wire  [0:23]  net2574;

wire  [0:47]  net3955;

wire  [0:7]  net2818;

wire  [0:23]  net2405;

wire  [0:7]  net2979;

wire  [0:7]  net2876;

wire  [0:47]  net2529;

wire  [0:47]  net3789;

wire  [0:7]  net3637;

wire  [0:47]  net3710;

wire  [0:47]  net4002;

wire  [0:47]  net4949;

wire  [0:47]  net4857;

wire  [0:47]  net2147;

wire  [0:47]  net4153;

wire  [0:7]  net4188;

wire  [0:23]  net3917;

wire  [0:47]  net2783;

wire  [0:7]  net2258;

wire  [0:47]  net2527;

wire  [0:7]  net2386;

wire  [0:47]  net2150;

wire  [0:47]  net4951;

wire  [0:7]  net2489;

wire  [0:7]  net2161;

wire  [0:7]  net2547;

wire  [0:23]  net2177;

wire  [0:7]  net2819;

wire  [0:7]  net3368;

wire  [0:47]  net4902;

wire  [0:47]  net3215;

wire  [0:47]  net4578;

wire  [0:7]  net3532;

wire  [0:47]  net4590;

wire  [0:7]  net3143;

wire  [0:23]  net2738;

wire  [0:47]  net2674;

wire  [0:47]  net2947;

wire  [0:47]  net2233;

wire  [0:47]  net3021;

wire  [0:7]  net4907;

wire  [0:7]  net4673;

wire  [0:7]  net4762;

wire  [0:7]  net3802;

wire  [0:47]  net2806;

wire  [0:23]  net3262;

wire  [0:47]  net4166;

wire  [0:23]  net3558;

wire  [0:47]  net4036;

wire  [0:7]  net3309;

wire  [0:47]  net4690;

wire  [0:47]  net4092;

wire  [0:47]  net4945;

wire  [0:23]  net2242;

wire  [0:47]  net3007;

wire  [0:23]  net2827;

wire  [0:47]  net2945;

wire  [0:23]  net3100;

wire  [0:47]  net4691;

wire  [0:7]  net2163;

wire  [0:7]  net4518;

wire  [0:47]  net3709;

wire  [0:47]  net3598;

wire  [0:7]  net2104;

wire  [0:23]  net4936;

wire  [0:23]  net2569;

wire  [0:47]  net2969;

wire  [0:23]  net2115;

wire  [0:47]  net3458;

wire  [0:23]  net4409;

wire  [0:47]  net2394;

wire  [0:7]  net2750;

wire  [0:23]  net2342;

wire  [0:7]  net2385;

wire  [0:47]  net3170;

wire  [0:47]  net4947;

wire  [0:47]  net4159;

wire  [0:23]  net3319;

wire  [0:7]  net4675;

wire  [0:23]  net4631;

wire  [0:47]  net3924;

wire  [0:7]  net4798;

wire  [0:7]  net4131;

wire  [0:47]  net2888;

wire  [0:23]  net3755;

wire  [0:47]  net4093;

wire  [0:23]  net3393;

wire  [0:47]  net2679;

wire  [0:47]  net3791;

wire  [0:47]  net4420;

wire  [0:47]  net2776;

wire  [0:7]  net4757;

wire  [0:23]  net2443;

wire  [0:7]  net2324;

wire  [0:7]  net4670;

wire  [0:23]  net3161;

wire  [0:47]  net2807;

wire  [0:7]  net2924;

wire  [0:47]  net2127;

wire  [0:47]  net3168;

wire  [0:7]  net4392;

wire  [0:23]  net4930;

wire  [0:7]  net2875;

wire  [0:7]  net3147;

wire  [0:47]  net4193;

wire  [0:47]  net3334;

wire  [0:47]  net2363;

wire  [0:47]  net2513;

wire  [0:47]  net2804;

wire  [0:23]  net3719;

wire  [0:47]  net4693;

wire  [0:23]  net3230;

wire  [0:23]  net2116;

wire  [0:47]  net2286;

wire  [0:47]  net3838;

wire  [0:7]  net2983;

wire  [0:7]  net4023;

wire  [0:7]  net4190;

wire  [0:47]  net3332;

wire  [0:23]  net2244;

wire  [0:47]  net4421;

wire  [0:23]  net2499;

wire  [0:23]  net4213;

wire  [0:47]  net3496;

wire  [0:47]  net2510;

wire  [0:7]  net4457;

wire  [0:23]  net4640;

wire  [0:47]  net4114;

wire  [0:7]  net4915;

wire  [0:7]  net3311;

wire  [0:47]  net3380;



lowla_modified I294 ( .clk(tclk_i), .min(net02076), .lao(net2079));
bram_bufferx4x6 I295 ( .in(sdi), .out(net02076));
tckbufx16 I242 ( .in(tclk_i), .out(net2076));
clk_colbuf8kx8 I346 ( .clko(clk_tree_drv[7:0]), .clki(glb_in[7:0]));
fabric_buf8k I290 ( .f_in(padin_l[23]), .f_out(padin_27));
fabric_buf8k I291 ( .f_in(net2084), .f_out(fabric_out_00_16));
fabric_buf8k I292 ( .f_in(net2086), .f_out(fabric_out_00_15));
array_LT1x16 I_it_05_bot ( .sp12_v_b_01(net4840[0:23]),
     .glb_netwk(net4755[0:7]), .bot_op_01({slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0],
     slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0]}), .sp12_v_t_16(sp12_v_t_05_16[23:0]),
     .rgt_op_16(slf_op_06_16[7:0]), .top_op_16(top_op_05_16[7:0]),
     .rgt_op_03(net2094[0:7]), .slf_op_02(net4392[0:7]),
     .rgt_op_02(net2096[0:7]), .rgt_op_01(net4806[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2924[0:7]), .lft_op_03(net2914[0:7]),
     .lft_op_02(net2916[0:7]), .lft_op_01(net4808[0:7]),
     .rgt_op_04(net2104[0:7]), .carry_in(net4996),
     .bnl_op_01({slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0], slf_op_04_00[3], slf_op_04_00[2],
     slf_op_04_00[1], slf_op_04_00[0]}), .slf_op_04(net4400[0:7]),
     .slf_op_03(net4390[0:7]), .slf_op_01(net4807[0:7]),
     .sp4_h_l_04(net4420[0:47]), .carry_out(carry_out_05_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net2113[0:23]),
     .sp12_h_r_03(net2114[0:23]), .sp12_h_r_02(net2115[0:23]),
     .sp12_h_r_01(net2116[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_05_16[7:0]), .sp4_v_b_01(net4856[0:47]),
     .sp4_r_v_b_04(net2120[0:47]), .sp4_r_v_b_03(net2121[0:47]),
     .sp4_r_v_b_02(net2122[0:47]), .sp4_r_v_b_01(net4855[0:47]),
     .sp4_h_r_04(net2124[0:47]), .sp4_h_r_03(net2125[0:47]),
     .sp4_h_r_02(net2126[0:47]), .sp4_h_r_01(net2127[0:47]),
     .sp4_h_l_03(net4421[0:47]), .sp4_h_l_02(net4422[0:47]),
     .sp4_h_l_01(net4423[0:47]), .bl(bl[287:234]),
     .sp12_h_l_01(net4412[0:23]), .sp12_h_l_02(net4411[0:23]),
     .sp12_h_l_03(net4410[0:23]), .sp12_h_l_04(net4409[0:23]),
     .sp4_v_b_04(net4416[0:47]), .sp4_v_b_03(net4417[0:47]),
     .sp4_v_b_02(net4418[0:47]), .bnr_op_01({slf_op_06_00[3],
     slf_op_06_00[2], slf_op_06_00[1], slf_op_06_00[0],
     slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0]}), .sp4_h_l_05(net4447[0:47]),
     .sp4_h_l_06(net4446[0:47]), .sp4_h_l_07(net4445[0:47]),
     .sp4_h_l_08(net4444[0:47]), .sp4_h_l_09(net4443[0:47]),
     .sp4_h_l_10(net4442[0:47]), .sp4_h_r_10(net2146[0:47]),
     .sp4_h_r_09(net2147[0:47]), .sp4_h_r_08(net2148[0:47]),
     .sp4_h_r_07(net2149[0:47]), .sp4_h_r_06(net2150[0:47]),
     .sp4_h_r_05(net2151[0:47]), .slf_op_05(net4459[0:7]),
     .slf_op_06(net4458[0:7]), .slf_op_07(net4457[0:7]),
     .slf_op_08(net4456[0:7]), .slf_op_09(net4455[0:7]),
     .slf_op_10(net4454[0:7]), .rgt_op_10(net2158[0:7]),
     .rgt_op_09(net2159[0:7]), .rgt_op_08(net2160[0:7]),
     .rgt_op_07(net2161[0:7]), .rgt_op_06(net2162[0:7]),
     .rgt_op_05(net2163[0:7]), .lft_op_10(net2978[0:7]),
     .lft_op_09(net2979[0:7]), .lft_op_08(net2980[0:7]),
     .lft_op_07(net2981[0:7]), .lft_op_06(net2982[0:7]),
     .lft_op_05(net2983[0:7]), .sp12_h_l_10(net4467[0:23]),
     .sp12_h_r_10(net2171[0:23]), .sp12_h_l_09(net4476[0:23]),
     .sp12_h_l_08(net4475[0:23]), .sp12_h_l_07(net4474[0:23]),
     .sp12_h_l_06(net4473[0:23]), .sp12_h_r_05(net2176[0:23]),
     .sp12_h_r_06(net2177[0:23]), .sp12_h_r_07(net2178[0:23]),
     .sp12_h_r_08(net2179[0:23]), .sp12_h_r_09(net2180[0:23]),
     .sp12_h_l_05(net4472[0:23]), .sp4_r_v_b_05(net2182[0:47]),
     .sp4_r_v_b_06(net2183[0:47]), .sp4_r_v_b_07(net2184[0:47]),
     .sp4_r_v_b_08(net2185[0:47]), .sp4_r_v_b_09(net2186[0:47]),
     .sp4_r_v_b_10(net2187[0:47]), .sp4_v_b_10(net4483[0:47]),
     .sp4_v_b_09(net4482[0:47]), .sp4_v_b_08(net4481[0:47]),
     .sp4_v_b_07(net4480[0:47]), .sp4_v_b_06(net4479[0:47]),
     .sp4_v_b_05(net4478[0:47]), .sp4_v_t_16(sp4_v_t_05_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net2197[0:47]), .sp4_h_r_12(net2198[0:47]),
     .sp4_h_r_13(net2199[0:47]), .sp4_h_r_14(net2200[0:47]),
     .sp4_h_r_15(net2201[0:47]), .sp4_h_r_16(net2202[0:47]),
     .sp4_h_l_16(net4498[0:47]), .sp4_h_l_15(net4497[0:47]),
     .sp4_h_l_14(net4496[0:47]), .sp4_h_l_13(net4495[0:47]),
     .sp4_h_l_12(net4494[0:47]), .sp4_h_l_11(net4493[0:47]),
     .tnr_op_16(tnr_op_05_16[7:0]), .tnl_op_16(tnl_op_05_16[7:0]),
     .lft_op_16(slf_op_04_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net4515[0:7]), .slf_op_14(net4514[0:7]),
     .slf_op_13(net4517[0:7]), .slf_op_12(net4516[0:7]),
     .slf_op_11(net4518[0:7]), .rgt_op_14(net2218[0:7]),
     .rgt_op_15(net2219[0:7]), .rgt_op_12(net2220[0:7]),
     .rgt_op_13(net2221[0:7]), .rgt_op_11(net2222[0:7]),
     .sp4_v_b_16(net4525[0:47]), .sp4_v_b_14(net4528[0:47]),
     .sp4_v_b_15(net4526[0:47]), .sp4_v_b_13(net4527[0:47]),
     .sp4_v_b_11(net4530[0:47]), .sp4_v_b_12(net4529[0:47]),
     .sp4_r_v_b_16(net2229[0:47]), .sp4_r_v_b_15(net2230[0:47]),
     .sp4_r_v_b_13(net2231[0:47]), .sp4_r_v_b_14(net2232[0:47]),
     .sp4_r_v_b_12(net2233[0:47]), .sp4_r_v_b_11(net2234[0:47]),
     .sp12_h_l_16(net4537[0:23]), .sp12_h_l_15(net4539[0:23]),
     .sp12_h_l_14(net4538[0:23]), .sp12_h_l_13(net4541[0:23]),
     .sp12_h_l_12(net4540[0:23]), .sp12_h_l_11(net4542[0:23]),
     .sp12_h_r_16(net2241[0:23]), .sp12_h_r_14(net2242[0:23]),
     .sp12_h_r_15(net2243[0:23]), .sp12_h_r_12(net2244[0:23]),
     .sp12_h_r_13(net2245[0:23]), .sp12_h_r_11(net2246[0:23]),
     .lft_op_14(net3038[0:7]), .lft_op_15(net3039[0:7]),
     .lft_op_12(net3040[0:7]), .lft_op_11(net3042[0:7]),
     .lft_op_13(net3041[0:7]));
array_LT1x16 I_it_11_bot ( .sp12_v_b_01(net4834[0:23]),
     .glb_netwk(net4761[0:7]), .bot_op_01({slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0],
     slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0]}), .sp12_v_t_16(sp12_v_t_11_16[23:0]),
     .rgt_op_16(slf_op_12_16[7:0]), .top_op_16(top_op_11_16[7:0]),
     .rgt_op_03(net2258[0:7]), .slf_op_02(net2424[0:7]),
     .rgt_op_02(net2260[0:7]), .rgt_op_01(net4800[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3744[0:7]), .lft_op_03(net3734[0:7]),
     .lft_op_02(net3736[0:7]), .lft_op_01(net4802[0:7]),
     .rgt_op_04(net2268[0:7]), .carry_in(net4989),
     .bnl_op_01({slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0], slf_op_10_00[3], slf_op_10_00[2],
     slf_op_10_00[1], slf_op_10_00[0]}), .slf_op_04(net2432[0:7]),
     .slf_op_03(net2422[0:7]), .slf_op_01(net4801[0:7]),
     .sp4_h_l_04(net2452[0:47]), .carry_out(carry_out_11_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net2277[0:23]),
     .sp12_h_r_03(net2278[0:23]), .sp12_h_r_02(net2279[0:23]),
     .sp12_h_r_01(net2280[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_11_16[7:0]), .sp4_v_b_01(net4850[0:47]),
     .sp4_r_v_b_04(net2284[0:47]), .sp4_r_v_b_03(net2285[0:47]),
     .sp4_r_v_b_02(net2286[0:47]), .sp4_r_v_b_01(net4849[0:47]),
     .sp4_h_r_04(net2288[0:47]), .sp4_h_r_03(net2289[0:47]),
     .sp4_h_r_02(net2290[0:47]), .sp4_h_r_01(net2291[0:47]),
     .sp4_h_l_03(net2453[0:47]), .sp4_h_l_02(net2454[0:47]),
     .sp4_h_l_01(net2455[0:47]), .bl(bl[599:546]),
     .sp12_h_l_01(net2444[0:23]), .sp12_h_l_02(net2443[0:23]),
     .sp12_h_l_03(net2442[0:23]), .sp12_h_l_04(net2441[0:23]),
     .sp4_v_b_04(net2448[0:47]), .sp4_v_b_03(net2449[0:47]),
     .sp4_v_b_02(net2450[0:47]), .bnr_op_01({slf_op_12_00[3],
     slf_op_12_00[2], slf_op_12_00[1], slf_op_12_00[0],
     slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0]}), .sp4_h_l_05(net2479[0:47]),
     .sp4_h_l_06(net2478[0:47]), .sp4_h_l_07(net2477[0:47]),
     .sp4_h_l_08(net2476[0:47]), .sp4_h_l_09(net2475[0:47]),
     .sp4_h_l_10(net2474[0:47]), .sp4_h_r_10(net2310[0:47]),
     .sp4_h_r_09(net2311[0:47]), .sp4_h_r_08(net2312[0:47]),
     .sp4_h_r_07(net2313[0:47]), .sp4_h_r_06(net2314[0:47]),
     .sp4_h_r_05(net2315[0:47]), .slf_op_05(net2491[0:7]),
     .slf_op_06(net2490[0:7]), .slf_op_07(net2489[0:7]),
     .slf_op_08(net2488[0:7]), .slf_op_09(net2487[0:7]),
     .slf_op_10(net2486[0:7]), .rgt_op_10(net2322[0:7]),
     .rgt_op_09(net2323[0:7]), .rgt_op_08(net2324[0:7]),
     .rgt_op_07(net2325[0:7]), .rgt_op_06(net2326[0:7]),
     .rgt_op_05(net2327[0:7]), .lft_op_10(net3798[0:7]),
     .lft_op_09(net3799[0:7]), .lft_op_08(net3800[0:7]),
     .lft_op_07(net3801[0:7]), .lft_op_06(net3802[0:7]),
     .lft_op_05(net3803[0:7]), .sp12_h_l_10(net2499[0:23]),
     .sp12_h_r_10(net2335[0:23]), .sp12_h_l_09(net2508[0:23]),
     .sp12_h_l_08(net2507[0:23]), .sp12_h_l_07(net2506[0:23]),
     .sp12_h_l_06(net2505[0:23]), .sp12_h_r_05(net2340[0:23]),
     .sp12_h_r_06(net2341[0:23]), .sp12_h_r_07(net2342[0:23]),
     .sp12_h_r_08(net2343[0:23]), .sp12_h_r_09(net2344[0:23]),
     .sp12_h_l_05(net2504[0:23]), .sp4_r_v_b_05(net2346[0:47]),
     .sp4_r_v_b_06(net2347[0:47]), .sp4_r_v_b_07(net2348[0:47]),
     .sp4_r_v_b_08(net2349[0:47]), .sp4_r_v_b_09(net2350[0:47]),
     .sp4_r_v_b_10(net2351[0:47]), .sp4_v_b_10(net2515[0:47]),
     .sp4_v_b_09(net2514[0:47]), .sp4_v_b_08(net2513[0:47]),
     .sp4_v_b_07(net2512[0:47]), .sp4_v_b_06(net2511[0:47]),
     .sp4_v_b_05(net2510[0:47]), .sp4_v_t_16(sp4_v_t_11_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net2361[0:47]), .sp4_h_r_12(net2362[0:47]),
     .sp4_h_r_13(net2363[0:47]), .sp4_h_r_14(net2364[0:47]),
     .sp4_h_r_15(net2365[0:47]), .sp4_h_r_16(net2366[0:47]),
     .sp4_h_l_16(net2530[0:47]), .sp4_h_l_15(net2529[0:47]),
     .sp4_h_l_14(net2528[0:47]), .sp4_h_l_13(net2527[0:47]),
     .sp4_h_l_12(net2526[0:47]), .sp4_h_l_11(net2525[0:47]),
     .tnr_op_16(tnr_op_11_16[7:0]), .tnl_op_16(tnl_op_11_16[7:0]),
     .lft_op_16(slf_op_10_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net2547[0:7]), .slf_op_14(net2546[0:7]),
     .slf_op_13(net2549[0:7]), .slf_op_12(net2548[0:7]),
     .slf_op_11(net2550[0:7]), .rgt_op_14(net2382[0:7]),
     .rgt_op_15(net2383[0:7]), .rgt_op_12(net2384[0:7]),
     .rgt_op_13(net2385[0:7]), .rgt_op_11(net2386[0:7]),
     .sp4_v_b_16(net2557[0:47]), .sp4_v_b_14(net2560[0:47]),
     .sp4_v_b_15(net2558[0:47]), .sp4_v_b_13(net2559[0:47]),
     .sp4_v_b_11(net2562[0:47]), .sp4_v_b_12(net2561[0:47]),
     .sp4_r_v_b_16(net2393[0:47]), .sp4_r_v_b_15(net2394[0:47]),
     .sp4_r_v_b_13(net2395[0:47]), .sp4_r_v_b_14(net2396[0:47]),
     .sp4_r_v_b_12(net2397[0:47]), .sp4_r_v_b_11(net2398[0:47]),
     .sp12_h_l_16(net2569[0:23]), .sp12_h_l_15(net2571[0:23]),
     .sp12_h_l_14(net2570[0:23]), .sp12_h_l_13(net2573[0:23]),
     .sp12_h_l_12(net2572[0:23]), .sp12_h_l_11(net2574[0:23]),
     .sp12_h_r_16(net2405[0:23]), .sp12_h_r_14(net2406[0:23]),
     .sp12_h_r_15(net2407[0:23]), .sp12_h_r_12(net2408[0:23]),
     .sp12_h_r_13(net2409[0:23]), .sp12_h_r_11(net2410[0:23]),
     .lft_op_14(net3858[0:7]), .lft_op_15(net3859[0:7]),
     .lft_op_12(net3860[0:7]), .lft_op_11(net3862[0:7]),
     .lft_op_13(net3861[0:7]));
array_LT1x16 I_it_10_bot ( .sp12_v_b_01(net4835[0:23]),
     .glb_netwk(net4760[0:7]), .bot_op_01({slf_op_10_00[3],
     slf_op_10_00[2], slf_op_10_00[1], slf_op_10_00[0],
     slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0]}), .sp12_v_t_16(sp12_v_t_10_16[23:0]),
     .rgt_op_16(slf_op_11_16[7:0]), .top_op_16(top_op_10_16[7:0]),
     .rgt_op_03(net2422[0:7]), .slf_op_02(net3736[0:7]),
     .rgt_op_02(net2424[0:7]), .rgt_op_01(net4801[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4665[0:7]), .lft_op_03(net4664[0:7]),
     .lft_op_02(net4663[0:7]), .lft_op_01(net4803[0:7]),
     .rgt_op_04(net2432[0:7]), .carry_in(net5023),
     .bnl_op_01({slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0], slf_op_09_00[3], slf_op_09_00[2],
     slf_op_09_00[1], slf_op_09_00[0]}), .slf_op_04(net3744[0:7]),
     .slf_op_03(net3734[0:7]), .slf_op_01(net4802[0:7]),
     .sp4_h_l_04(net3764[0:47]), .carry_out(carry_out_10_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net2441[0:23]),
     .sp12_h_r_03(net2442[0:23]), .sp12_h_r_02(net2443[0:23]),
     .sp12_h_r_01(net2444[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_10_16[7:0]), .sp4_v_b_01(net4851[0:47]),
     .sp4_r_v_b_04(net2448[0:47]), .sp4_r_v_b_03(net2449[0:47]),
     .sp4_r_v_b_02(net2450[0:47]), .sp4_r_v_b_01(net4850[0:47]),
     .sp4_h_r_04(net2452[0:47]), .sp4_h_r_03(net2453[0:47]),
     .sp4_h_r_02(net2454[0:47]), .sp4_h_r_01(net2455[0:47]),
     .sp4_h_l_03(net3765[0:47]), .sp4_h_l_02(net3766[0:47]),
     .sp4_h_l_01(net3767[0:47]), .bl(bl[545:492]),
     .sp12_h_l_01(net3756[0:23]), .sp12_h_l_02(net3755[0:23]),
     .sp12_h_l_03(net3754[0:23]), .sp12_h_l_04(net3753[0:23]),
     .sp4_v_b_04(net3760[0:47]), .sp4_v_b_03(net3761[0:47]),
     .sp4_v_b_02(net3762[0:47]), .bnr_op_01({slf_op_11_00[3],
     slf_op_11_00[2], slf_op_11_00[1], slf_op_11_00[0],
     slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0]}), .sp4_h_l_05(net3791[0:47]),
     .sp4_h_l_06(net3790[0:47]), .sp4_h_l_07(net3789[0:47]),
     .sp4_h_l_08(net3788[0:47]), .sp4_h_l_09(net3787[0:47]),
     .sp4_h_l_10(net3786[0:47]), .sp4_h_r_10(net2474[0:47]),
     .sp4_h_r_09(net2475[0:47]), .sp4_h_r_08(net2476[0:47]),
     .sp4_h_r_07(net2477[0:47]), .sp4_h_r_06(net2478[0:47]),
     .sp4_h_r_05(net2479[0:47]), .slf_op_05(net3803[0:7]),
     .slf_op_06(net3802[0:7]), .slf_op_07(net3801[0:7]),
     .slf_op_08(net3800[0:7]), .slf_op_09(net3799[0:7]),
     .slf_op_10(net3798[0:7]), .rgt_op_10(net2486[0:7]),
     .rgt_op_09(net2487[0:7]), .rgt_op_08(net2488[0:7]),
     .rgt_op_07(net2489[0:7]), .rgt_op_06(net2490[0:7]),
     .rgt_op_05(net2491[0:7]), .lft_op_10(net4671[0:7]),
     .lft_op_09(net4670[0:7]), .lft_op_08(net4669[0:7]),
     .lft_op_07(net4668[0:7]), .lft_op_06(net4667[0:7]),
     .lft_op_05(net4666[0:7]), .sp12_h_l_10(net3811[0:23]),
     .sp12_h_r_10(net2499[0:23]), .sp12_h_l_09(net3820[0:23]),
     .sp12_h_l_08(net3819[0:23]), .sp12_h_l_07(net3818[0:23]),
     .sp12_h_l_06(net3817[0:23]), .sp12_h_r_05(net2504[0:23]),
     .sp12_h_r_06(net2505[0:23]), .sp12_h_r_07(net2506[0:23]),
     .sp12_h_r_08(net2507[0:23]), .sp12_h_r_09(net2508[0:23]),
     .sp12_h_l_05(net3816[0:23]), .sp4_r_v_b_05(net2510[0:47]),
     .sp4_r_v_b_06(net2511[0:47]), .sp4_r_v_b_07(net2512[0:47]),
     .sp4_r_v_b_08(net2513[0:47]), .sp4_r_v_b_09(net2514[0:47]),
     .sp4_r_v_b_10(net2515[0:47]), .sp4_v_b_10(net3827[0:47]),
     .sp4_v_b_09(net3826[0:47]), .sp4_v_b_08(net3825[0:47]),
     .sp4_v_b_07(net3824[0:47]), .sp4_v_b_06(net3823[0:47]),
     .sp4_v_b_05(net3822[0:47]), .sp4_v_t_16(sp4_v_t_10_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net2525[0:47]), .sp4_h_r_12(net2526[0:47]),
     .sp4_h_r_13(net2527[0:47]), .sp4_h_r_14(net2528[0:47]),
     .sp4_h_r_15(net2529[0:47]), .sp4_h_r_16(net2530[0:47]),
     .sp4_h_l_16(net3842[0:47]), .sp4_h_l_15(net3841[0:47]),
     .sp4_h_l_14(net3840[0:47]), .sp4_h_l_13(net3839[0:47]),
     .sp4_h_l_12(net3838[0:47]), .sp4_h_l_11(net3837[0:47]),
     .tnr_op_16(tnr_op_10_16[7:0]), .tnl_op_16(tnl_op_10_16[7:0]),
     .lft_op_16(slf_op_09_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net3859[0:7]), .slf_op_14(net3858[0:7]),
     .slf_op_13(net3861[0:7]), .slf_op_12(net3860[0:7]),
     .slf_op_11(net3862[0:7]), .rgt_op_14(net2546[0:7]),
     .rgt_op_15(net2547[0:7]), .rgt_op_12(net2548[0:7]),
     .rgt_op_13(net2549[0:7]), .rgt_op_11(net2550[0:7]),
     .sp4_v_b_16(net3869[0:47]), .sp4_v_b_14(net3872[0:47]),
     .sp4_v_b_15(net3870[0:47]), .sp4_v_b_13(net3871[0:47]),
     .sp4_v_b_11(net3874[0:47]), .sp4_v_b_12(net3873[0:47]),
     .sp4_r_v_b_16(net2557[0:47]), .sp4_r_v_b_15(net2558[0:47]),
     .sp4_r_v_b_13(net2559[0:47]), .sp4_r_v_b_14(net2560[0:47]),
     .sp4_r_v_b_12(net2561[0:47]), .sp4_r_v_b_11(net2562[0:47]),
     .sp12_h_l_16(net3881[0:23]), .sp12_h_l_15(net3883[0:23]),
     .sp12_h_l_14(net3882[0:23]), .sp12_h_l_13(net3885[0:23]),
     .sp12_h_l_12(net3884[0:23]), .sp12_h_l_11(net3886[0:23]),
     .sp12_h_r_16(net2569[0:23]), .sp12_h_r_14(net2570[0:23]),
     .sp12_h_r_15(net2571[0:23]), .sp12_h_r_12(net2572[0:23]),
     .sp12_h_r_13(net2573[0:23]), .sp12_h_r_11(net2574[0:23]),
     .lft_op_14(net4675[0:7]), .lft_op_15(net4676[0:7]),
     .lft_op_12(net4673[0:7]), .lft_op_11(net4672[0:7]),
     .lft_op_13(net4674[0:7]));
array_LT1x16 I_it_15_bot ( .sp12_v_b_01(net4830[0:23]),
     .glb_netwk(net4765[0:7]), .bot_op_01({slf_op_15_00[3],
     slf_op_15_00[2], slf_op_15_00[1], slf_op_15_00[0],
     slf_op_15_00[3], slf_op_15_00[2], slf_op_15_00[1],
     slf_op_15_00[0]}), .sp12_v_t_16(sp12_v_t_15_16[23:0]),
     .rgt_op_16(slf_op_16_16[7:0]), .top_op_16(top_op_15_16[7:0]),
     .rgt_op_03(slf_op_16_03[7:0]), .slf_op_02(net3080[0:7]),
     .rgt_op_02(slf_op_16_02[7:0]), .rgt_op_01(slf_op_16_01[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net3580[0:7]),
     .lft_op_03(net3570[0:7]), .lft_op_02(net3572[0:7]),
     .lft_op_01(net4798[0:7]), .rgt_op_04(slf_op_16_04[7:0]),
     .carry_in(net2597), .bnl_op_01({slf_op_14_00[3], slf_op_14_00[2],
     slf_op_14_00[1], slf_op_14_00[0], slf_op_14_00[3],
     slf_op_14_00[2], slf_op_14_00[1], slf_op_14_00[0]}),
     .slf_op_04(net3088[0:7]), .slf_op_03(net3078[0:7]),
     .slf_op_01(net4797[0:7]), .sp4_h_l_04(net3108[0:47]),
     .carry_out(carry_out_15_16), .vdd_cntl(vdd_cntl_l[271:16]),
     .sp12_h_r_04(net2605[0:23]), .sp12_h_r_03(net2606[0:23]),
     .sp12_h_r_02(net2607[0:23]), .sp12_h_r_01(net2608[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(slf_op_15_16[7:0]),
     .sp4_v_b_01(net4846[0:47]), .sp4_r_v_b_04(net2612[0:47]),
     .sp4_r_v_b_03(net2613[0:47]), .sp4_r_v_b_02(net2614[0:47]),
     .sp4_r_v_b_01(net4845[0:47]), .sp4_h_r_04(net2616[0:47]),
     .sp4_h_r_03(net2617[0:47]), .sp4_h_r_02(net2618[0:47]),
     .sp4_h_r_01(net2619[0:47]), .sp4_h_l_03(net3109[0:47]),
     .sp4_h_l_02(net3110[0:47]), .sp4_h_l_01(net3111[0:47]),
     .bl(bl[815:762]), .sp12_h_l_01(net3100[0:23]),
     .sp12_h_l_02(net3099[0:23]), .sp12_h_l_03(net3098[0:23]),
     .sp12_h_l_04(net3097[0:23]), .sp4_v_b_04(net3104[0:47]),
     .sp4_v_b_03(net3105[0:47]), .sp4_v_b_02(net3106[0:47]),
     .bnr_op_01({slf_op_16_00[3], slf_op_16_00[2], slf_op_16_00[1],
     slf_op_16_00[0], slf_op_16_00[3], slf_op_16_00[2],
     slf_op_16_00[1], slf_op_16_00[0]}), .sp4_h_l_05(net3135[0:47]),
     .sp4_h_l_06(net3134[0:47]), .sp4_h_l_07(net3133[0:47]),
     .sp4_h_l_08(net3132[0:47]), .sp4_h_l_09(net3131[0:47]),
     .sp4_h_l_10(net3130[0:47]), .sp4_h_r_10(net2638[0:47]),
     .sp4_h_r_09(net2639[0:47]), .sp4_h_r_08(net2640[0:47]),
     .sp4_h_r_07(net2641[0:47]), .sp4_h_r_06(net2642[0:47]),
     .sp4_h_r_05(net2643[0:47]), .slf_op_05(net3147[0:7]),
     .slf_op_06(net3146[0:7]), .slf_op_07(net3145[0:7]),
     .slf_op_08(net3144[0:7]), .slf_op_09(net3143[0:7]),
     .slf_op_10(net3142[0:7]), .rgt_op_10(slf_op_16_10[7:0]),
     .rgt_op_09(slf_op_16_09[7:0]), .rgt_op_08(slf_op_16_08[7:0]),
     .rgt_op_07(slf_op_16_07[7:0]), .rgt_op_06(slf_op_16_06[7:0]),
     .rgt_op_05(slf_op_16_05[7:0]), .lft_op_10(net3634[0:7]),
     .lft_op_09(net3635[0:7]), .lft_op_08(net3636[0:7]),
     .lft_op_07(net3637[0:7]), .lft_op_06(net3638[0:7]),
     .lft_op_05(net3639[0:7]), .sp12_h_l_10(net3155[0:23]),
     .sp12_h_r_10(net2663[0:23]), .sp12_h_l_09(net3164[0:23]),
     .sp12_h_l_08(net3163[0:23]), .sp12_h_l_07(net3162[0:23]),
     .sp12_h_l_06(net3161[0:23]), .sp12_h_r_05(net2668[0:23]),
     .sp12_h_r_06(net2669[0:23]), .sp12_h_r_07(net2670[0:23]),
     .sp12_h_r_08(net2671[0:23]), .sp12_h_r_09(net2672[0:23]),
     .sp12_h_l_05(net3160[0:23]), .sp4_r_v_b_05(net2674[0:47]),
     .sp4_r_v_b_06(net2675[0:47]), .sp4_r_v_b_07(net2676[0:47]),
     .sp4_r_v_b_08(net2677[0:47]), .sp4_r_v_b_09(net2678[0:47]),
     .sp4_r_v_b_10(net2679[0:47]), .sp4_v_b_10(net3171[0:47]),
     .sp4_v_b_09(net3170[0:47]), .sp4_v_b_08(net3169[0:47]),
     .sp4_v_b_07(net3168[0:47]), .sp4_v_b_06(net3167[0:47]),
     .sp4_v_b_05(net3166[0:47]), .sp4_v_t_16(sp4_v_t_15_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net2689[0:47]), .sp4_h_r_12(net2690[0:47]),
     .sp4_h_r_13(net2691[0:47]), .sp4_h_r_14(net2692[0:47]),
     .sp4_h_r_15(net2693[0:47]), .sp4_h_r_16(net2694[0:47]),
     .sp4_h_l_16(net3186[0:47]), .sp4_h_l_15(net3185[0:47]),
     .sp4_h_l_14(net3184[0:47]), .sp4_h_l_13(net3183[0:47]),
     .sp4_h_l_12(net3182[0:47]), .sp4_h_l_11(net3181[0:47]),
     .tnr_op_16(tnr_op_15_16[7:0]), .tnl_op_16(tnl_op_15_16[7:0]),
     .lft_op_16(slf_op_14_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net3203[0:7]), .slf_op_14(net3202[0:7]),
     .slf_op_13(net3205[0:7]), .slf_op_12(net3204[0:7]),
     .slf_op_11(net3206[0:7]), .rgt_op_14(slf_op_16_14[7:0]),
     .rgt_op_15(slf_op_16_15[7:0]), .rgt_op_12(slf_op_16_12[7:0]),
     .rgt_op_13(slf_op_16_13[7:0]), .rgt_op_11(slf_op_16_11[7:0]),
     .sp4_v_b_16(net3213[0:47]), .sp4_v_b_14(net3216[0:47]),
     .sp4_v_b_15(net3214[0:47]), .sp4_v_b_13(net3215[0:47]),
     .sp4_v_b_11(net3218[0:47]), .sp4_v_b_12(net3217[0:47]),
     .sp4_r_v_b_16(net2721[0:47]), .sp4_r_v_b_15(net2722[0:47]),
     .sp4_r_v_b_13(net2723[0:47]), .sp4_r_v_b_14(net2724[0:47]),
     .sp4_r_v_b_12(net2725[0:47]), .sp4_r_v_b_11(net2726[0:47]),
     .sp12_h_l_16(net3225[0:23]), .sp12_h_l_15(net3227[0:23]),
     .sp12_h_l_14(net3226[0:23]), .sp12_h_l_13(net3229[0:23]),
     .sp12_h_l_12(net3228[0:23]), .sp12_h_l_11(net3230[0:23]),
     .sp12_h_r_16(net2733[0:23]), .sp12_h_r_14(net2734[0:23]),
     .sp12_h_r_15(net2735[0:23]), .sp12_h_r_12(net2736[0:23]),
     .sp12_h_r_13(net2737[0:23]), .sp12_h_r_11(net2738[0:23]),
     .lft_op_14(net3694[0:7]), .lft_op_15(net3695[0:7]),
     .lft_op_12(net3696[0:7]), .lft_op_11(net3698[0:7]),
     .lft_op_13(net3697[0:7]));
array_LT1x16 I_it_06_bot ( .sp12_v_b_01(net4839[0:23]),
     .glb_netwk(net4756[0:7]), .bot_op_01({slf_op_06_00[3],
     slf_op_06_00[2], slf_op_06_00[1], slf_op_06_00[0],
     slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0]}), .sp12_v_t_16(sp12_v_t_06_16[23:0]),
     .rgt_op_16(slf_op_07_16[7:0]), .top_op_16(top_op_06_16[7:0]),
     .rgt_op_03(net2750[0:7]), .slf_op_02(net2096[0:7]),
     .rgt_op_02(net2752[0:7]), .rgt_op_01(net4805[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4400[0:7]), .lft_op_03(net4390[0:7]),
     .lft_op_02(net4392[0:7]), .lft_op_01(net4807[0:7]),
     .rgt_op_04(net2760[0:7]), .carry_in(net4986),
     .bnl_op_01({slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0], slf_op_05_00[3], slf_op_05_00[2],
     slf_op_05_00[1], slf_op_05_00[0]}), .slf_op_04(net2104[0:7]),
     .slf_op_03(net2094[0:7]), .slf_op_01(net4806[0:7]),
     .sp4_h_l_04(net2124[0:47]), .carry_out(carry_out_06_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net2769[0:23]),
     .sp12_h_r_03(net2770[0:23]), .sp12_h_r_02(net2771[0:23]),
     .sp12_h_r_01(net2772[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_06_16[7:0]), .sp4_v_b_01(net4855[0:47]),
     .sp4_r_v_b_04(net2776[0:47]), .sp4_r_v_b_03(net2777[0:47]),
     .sp4_r_v_b_02(net2778[0:47]), .sp4_r_v_b_01(net4854[0:47]),
     .sp4_h_r_04(net2780[0:47]), .sp4_h_r_03(net2781[0:47]),
     .sp4_h_r_02(net2782[0:47]), .sp4_h_r_01(net2783[0:47]),
     .sp4_h_l_03(net2125[0:47]), .sp4_h_l_02(net2126[0:47]),
     .sp4_h_l_01(net2127[0:47]), .bl(bl[341:288]),
     .sp12_h_l_01(net2116[0:23]), .sp12_h_l_02(net2115[0:23]),
     .sp12_h_l_03(net2114[0:23]), .sp12_h_l_04(net2113[0:23]),
     .sp4_v_b_04(net2120[0:47]), .sp4_v_b_03(net2121[0:47]),
     .sp4_v_b_02(net2122[0:47]), .bnr_op_01({slf_op_07_00[3],
     slf_op_07_00[2], slf_op_07_00[1], slf_op_07_00[0],
     slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0]}), .sp4_h_l_05(net2151[0:47]),
     .sp4_h_l_06(net2150[0:47]), .sp4_h_l_07(net2149[0:47]),
     .sp4_h_l_08(net2148[0:47]), .sp4_h_l_09(net2147[0:47]),
     .sp4_h_l_10(net2146[0:47]), .sp4_h_r_10(net2802[0:47]),
     .sp4_h_r_09(net2803[0:47]), .sp4_h_r_08(net2804[0:47]),
     .sp4_h_r_07(net2805[0:47]), .sp4_h_r_06(net2806[0:47]),
     .sp4_h_r_05(net2807[0:47]), .slf_op_05(net2163[0:7]),
     .slf_op_06(net2162[0:7]), .slf_op_07(net2161[0:7]),
     .slf_op_08(net2160[0:7]), .slf_op_09(net2159[0:7]),
     .slf_op_10(net2158[0:7]), .rgt_op_10(net2814[0:7]),
     .rgt_op_09(net2815[0:7]), .rgt_op_08(net2816[0:7]),
     .rgt_op_07(net2817[0:7]), .rgt_op_06(net2818[0:7]),
     .rgt_op_05(net2819[0:7]), .lft_op_10(net4454[0:7]),
     .lft_op_09(net4455[0:7]), .lft_op_08(net4456[0:7]),
     .lft_op_07(net4457[0:7]), .lft_op_06(net4458[0:7]),
     .lft_op_05(net4459[0:7]), .sp12_h_l_10(net2171[0:23]),
     .sp12_h_r_10(net2827[0:23]), .sp12_h_l_09(net2180[0:23]),
     .sp12_h_l_08(net2179[0:23]), .sp12_h_l_07(net2178[0:23]),
     .sp12_h_l_06(net2177[0:23]), .sp12_h_r_05(net2832[0:23]),
     .sp12_h_r_06(net2833[0:23]), .sp12_h_r_07(net2834[0:23]),
     .sp12_h_r_08(net2835[0:23]), .sp12_h_r_09(net2836[0:23]),
     .sp12_h_l_05(net2176[0:23]), .sp4_r_v_b_05(net2838[0:47]),
     .sp4_r_v_b_06(net2839[0:47]), .sp4_r_v_b_07(net2840[0:47]),
     .sp4_r_v_b_08(net2841[0:47]), .sp4_r_v_b_09(net2842[0:47]),
     .sp4_r_v_b_10(net2843[0:47]), .sp4_v_b_10(net2187[0:47]),
     .sp4_v_b_09(net2186[0:47]), .sp4_v_b_08(net2185[0:47]),
     .sp4_v_b_07(net2184[0:47]), .sp4_v_b_06(net2183[0:47]),
     .sp4_v_b_05(net2182[0:47]), .sp4_v_t_16(sp4_v_t_06_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net2853[0:47]), .sp4_h_r_12(net2854[0:47]),
     .sp4_h_r_13(net2855[0:47]), .sp4_h_r_14(net2856[0:47]),
     .sp4_h_r_15(net2857[0:47]), .sp4_h_r_16(net2858[0:47]),
     .sp4_h_l_16(net2202[0:47]), .sp4_h_l_15(net2201[0:47]),
     .sp4_h_l_14(net2200[0:47]), .sp4_h_l_13(net2199[0:47]),
     .sp4_h_l_12(net2198[0:47]), .sp4_h_l_11(net2197[0:47]),
     .tnr_op_16(tnr_op_06_16[7:0]), .tnl_op_16(tnl_op_06_16[7:0]),
     .lft_op_16(slf_op_05_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net2219[0:7]), .slf_op_14(net2218[0:7]),
     .slf_op_13(net2221[0:7]), .slf_op_12(net2220[0:7]),
     .slf_op_11(net2222[0:7]), .rgt_op_14(net2874[0:7]),
     .rgt_op_15(net2875[0:7]), .rgt_op_12(net2876[0:7]),
     .rgt_op_13(net2877[0:7]), .rgt_op_11(net2878[0:7]),
     .sp4_v_b_16(net2229[0:47]), .sp4_v_b_14(net2232[0:47]),
     .sp4_v_b_15(net2230[0:47]), .sp4_v_b_13(net2231[0:47]),
     .sp4_v_b_11(net2234[0:47]), .sp4_v_b_12(net2233[0:47]),
     .sp4_r_v_b_16(net2885[0:47]), .sp4_r_v_b_15(net2886[0:47]),
     .sp4_r_v_b_13(net2887[0:47]), .sp4_r_v_b_14(net2888[0:47]),
     .sp4_r_v_b_12(net2889[0:47]), .sp4_r_v_b_11(net2890[0:47]),
     .sp12_h_l_16(net2241[0:23]), .sp12_h_l_15(net2243[0:23]),
     .sp12_h_l_14(net2242[0:23]), .sp12_h_l_13(net2245[0:23]),
     .sp12_h_l_12(net2244[0:23]), .sp12_h_l_11(net2246[0:23]),
     .sp12_h_r_16(net2897[0:23]), .sp12_h_r_14(net2898[0:23]),
     .sp12_h_r_15(net2899[0:23]), .sp12_h_r_12(net2900[0:23]),
     .sp12_h_r_13(net2901[0:23]), .sp12_h_r_11(net2902[0:23]),
     .lft_op_14(net4514[0:7]), .lft_op_15(net4515[0:7]),
     .lft_op_12(net4516[0:7]), .lft_op_11(net4518[0:7]),
     .lft_op_13(net4517[0:7]));
array_LT1x16 I_it_03_bot ( .sp12_v_b_01(net4842[0:23]),
     .glb_netwk(net4753[0:7]), .bot_op_01({slf_op_03_00[3],
     slf_op_03_00[2], slf_op_03_00[1], slf_op_03_00[0],
     slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0]}), .sp12_v_t_16(sp12_v_t_03_16[23:0]),
     .rgt_op_16(slf_op_04_16[7:0]), .top_op_16(top_op_03_16[7:0]),
     .rgt_op_03(net2914[0:7]), .slf_op_02(net3900[0:7]),
     .rgt_op_02(net2916[0:7]), .rgt_op_01(net4808[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4072[0:7]), .lft_op_03(net4062[0:7]),
     .lft_op_02(net4064[0:7]), .lft_op_01(net4810[0:7]),
     .rgt_op_04(net2924[0:7]), .carry_in(net5052),
     .bnl_op_01({slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0], slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0]}), .slf_op_04(net3908[0:7]),
     .slf_op_03(net3898[0:7]), .slf_op_01(net4809[0:7]),
     .sp4_h_l_04(net3928[0:47]), .carry_out(carry_out_03_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net2933[0:23]),
     .sp12_h_r_03(net2934[0:23]), .sp12_h_r_02(net2935[0:23]),
     .sp12_h_r_01(net2936[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_03_16[7:0]), .sp4_v_b_01(net4858[0:47]),
     .sp4_r_v_b_04(net2940[0:47]), .sp4_r_v_b_03(net2941[0:47]),
     .sp4_r_v_b_02(net2942[0:47]), .sp4_r_v_b_01(net4857[0:47]),
     .sp4_h_r_04(net2944[0:47]), .sp4_h_r_03(net2945[0:47]),
     .sp4_h_r_02(net2946[0:47]), .sp4_h_r_01(net2947[0:47]),
     .sp4_h_l_03(net3929[0:47]), .sp4_h_l_02(net3930[0:47]),
     .sp4_h_l_01(net3931[0:47]), .bl(bl[179:126]),
     .sp12_h_l_01(net3920[0:23]), .sp12_h_l_02(net3919[0:23]),
     .sp12_h_l_03(net3918[0:23]), .sp12_h_l_04(net3917[0:23]),
     .sp4_v_b_04(net3924[0:47]), .sp4_v_b_03(net3925[0:47]),
     .sp4_v_b_02(net3926[0:47]), .bnr_op_01({slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0],
     slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0]}), .sp4_h_l_05(net3955[0:47]),
     .sp4_h_l_06(net3954[0:47]), .sp4_h_l_07(net3953[0:47]),
     .sp4_h_l_08(net3952[0:47]), .sp4_h_l_09(net3951[0:47]),
     .sp4_h_l_10(net3950[0:47]), .sp4_h_r_10(net2966[0:47]),
     .sp4_h_r_09(net2967[0:47]), .sp4_h_r_08(net2968[0:47]),
     .sp4_h_r_07(net2969[0:47]), .sp4_h_r_06(net2970[0:47]),
     .sp4_h_r_05(net2971[0:47]), .slf_op_05(net3967[0:7]),
     .slf_op_06(net3966[0:7]), .slf_op_07(net3965[0:7]),
     .slf_op_08(net3964[0:7]), .slf_op_09(net3963[0:7]),
     .slf_op_10(net3962[0:7]), .rgt_op_10(net2978[0:7]),
     .rgt_op_09(net2979[0:7]), .rgt_op_08(net2980[0:7]),
     .rgt_op_07(net2981[0:7]), .rgt_op_06(net2982[0:7]),
     .rgt_op_05(net2983[0:7]), .lft_op_10(net4126[0:7]),
     .lft_op_09(net4127[0:7]), .lft_op_08(net4128[0:7]),
     .lft_op_07(net4129[0:7]), .lft_op_06(net4130[0:7]),
     .lft_op_05(net4131[0:7]), .sp12_h_l_10(net3975[0:23]),
     .sp12_h_r_10(net2991[0:23]), .sp12_h_l_09(net3984[0:23]),
     .sp12_h_l_08(net3983[0:23]), .sp12_h_l_07(net3982[0:23]),
     .sp12_h_l_06(net3981[0:23]), .sp12_h_r_05(net2996[0:23]),
     .sp12_h_r_06(net2997[0:23]), .sp12_h_r_07(net2998[0:23]),
     .sp12_h_r_08(net2999[0:23]), .sp12_h_r_09(net3000[0:23]),
     .sp12_h_l_05(net3980[0:23]), .sp4_r_v_b_05(net3002[0:47]),
     .sp4_r_v_b_06(net3003[0:47]), .sp4_r_v_b_07(net3004[0:47]),
     .sp4_r_v_b_08(net3005[0:47]), .sp4_r_v_b_09(net3006[0:47]),
     .sp4_r_v_b_10(net3007[0:47]), .sp4_v_b_10(net3991[0:47]),
     .sp4_v_b_09(net3990[0:47]), .sp4_v_b_08(net3989[0:47]),
     .sp4_v_b_07(net3988[0:47]), .sp4_v_b_06(net3987[0:47]),
     .sp4_v_b_05(net3986[0:47]), .sp4_v_t_16(sp4_v_t_03_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net3017[0:47]), .sp4_h_r_12(net3018[0:47]),
     .sp4_h_r_13(net3019[0:47]), .sp4_h_r_14(net3020[0:47]),
     .sp4_h_r_15(net3021[0:47]), .sp4_h_r_16(net3022[0:47]),
     .sp4_h_l_16(net4006[0:47]), .sp4_h_l_15(net4005[0:47]),
     .sp4_h_l_14(net4004[0:47]), .sp4_h_l_13(net4003[0:47]),
     .sp4_h_l_12(net4002[0:47]), .sp4_h_l_11(net4001[0:47]),
     .tnr_op_16(tnr_op_03_16[7:0]), .tnl_op_16(tnl_op_03_16[7:0]),
     .lft_op_16(slf_op_02_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net4023[0:7]), .slf_op_14(net4022[0:7]),
     .slf_op_13(net4025[0:7]), .slf_op_12(net4024[0:7]),
     .slf_op_11(net4026[0:7]), .rgt_op_14(net3038[0:7]),
     .rgt_op_15(net3039[0:7]), .rgt_op_12(net3040[0:7]),
     .rgt_op_13(net3041[0:7]), .rgt_op_11(net3042[0:7]),
     .sp4_v_b_16(net4033[0:47]), .sp4_v_b_14(net4036[0:47]),
     .sp4_v_b_15(net4034[0:47]), .sp4_v_b_13(net4035[0:47]),
     .sp4_v_b_11(net4038[0:47]), .sp4_v_b_12(net4037[0:47]),
     .sp4_r_v_b_16(net3049[0:47]), .sp4_r_v_b_15(net3050[0:47]),
     .sp4_r_v_b_13(net3051[0:47]), .sp4_r_v_b_14(net3052[0:47]),
     .sp4_r_v_b_12(net3053[0:47]), .sp4_r_v_b_11(net3054[0:47]),
     .sp12_h_l_16(net4045[0:23]), .sp12_h_l_15(net4047[0:23]),
     .sp12_h_l_14(net4046[0:23]), .sp12_h_l_13(net4049[0:23]),
     .sp12_h_l_12(net4048[0:23]), .sp12_h_l_11(net4050[0:23]),
     .sp12_h_r_16(net3061[0:23]), .sp12_h_r_14(net3062[0:23]),
     .sp12_h_r_15(net3063[0:23]), .sp12_h_r_12(net3064[0:23]),
     .sp12_h_r_13(net3065[0:23]), .sp12_h_r_11(net3066[0:23]),
     .lft_op_14(net4186[0:7]), .lft_op_15(net4187[0:7]),
     .lft_op_12(net4188[0:7]), .lft_op_11(net4190[0:7]),
     .lft_op_13(net4189[0:7]));
array_LT1x16 I_it_14_bot ( .sp12_v_b_01(net4831[0:23]),
     .glb_netwk(net4764[0:7]), .bot_op_01({slf_op_14_00[3],
     slf_op_14_00[2], slf_op_14_00[1], slf_op_14_00[0],
     slf_op_14_00[3], slf_op_14_00[2], slf_op_14_00[1],
     slf_op_14_00[0]}), .sp12_v_t_16(sp12_v_t_14_16[23:0]),
     .rgt_op_16(slf_op_15_16[7:0]), .top_op_16(top_op_14_16[7:0]),
     .rgt_op_03(net3078[0:7]), .slf_op_02(net3572[0:7]),
     .rgt_op_02(net3080[0:7]), .rgt_op_01(net4797[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3252[0:7]), .lft_op_03(net3242[0:7]),
     .lft_op_02(net3244[0:7]), .lft_op_01(net4799[0:7]),
     .rgt_op_04(net3088[0:7]), .carry_in(net4987),
     .bnl_op_01({slf_op_13_00[3], slf_op_13_00[2], slf_op_13_00[1],
     slf_op_13_00[0], slf_op_13_00[3], slf_op_13_00[2],
     slf_op_13_00[1], slf_op_13_00[0]}), .slf_op_04(net3580[0:7]),
     .slf_op_03(net3570[0:7]), .slf_op_01(net4798[0:7]),
     .sp4_h_l_04(net3600[0:47]), .carry_out(carry_out_14_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net3097[0:23]),
     .sp12_h_r_03(net3098[0:23]), .sp12_h_r_02(net3099[0:23]),
     .sp12_h_r_01(net3100[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_14_16[7:0]), .sp4_v_b_01(net4847[0:47]),
     .sp4_r_v_b_04(net3104[0:47]), .sp4_r_v_b_03(net3105[0:47]),
     .sp4_r_v_b_02(net3106[0:47]), .sp4_r_v_b_01(net4846[0:47]),
     .sp4_h_r_04(net3108[0:47]), .sp4_h_r_03(net3109[0:47]),
     .sp4_h_r_02(net3110[0:47]), .sp4_h_r_01(net3111[0:47]),
     .sp4_h_l_03(net3601[0:47]), .sp4_h_l_02(net3602[0:47]),
     .sp4_h_l_01(net3603[0:47]), .bl(bl[761:708]),
     .sp12_h_l_01(net3592[0:23]), .sp12_h_l_02(net3591[0:23]),
     .sp12_h_l_03(net3590[0:23]), .sp12_h_l_04(net3589[0:23]),
     .sp4_v_b_04(net3596[0:47]), .sp4_v_b_03(net3597[0:47]),
     .sp4_v_b_02(net3598[0:47]), .bnr_op_01({slf_op_15_00[3],
     slf_op_15_00[2], slf_op_15_00[1], slf_op_15_00[0],
     slf_op_15_00[3], slf_op_15_00[2], slf_op_15_00[1],
     slf_op_15_00[0]}), .sp4_h_l_05(net3627[0:47]),
     .sp4_h_l_06(net3626[0:47]), .sp4_h_l_07(net3625[0:47]),
     .sp4_h_l_08(net3624[0:47]), .sp4_h_l_09(net3623[0:47]),
     .sp4_h_l_10(net3622[0:47]), .sp4_h_r_10(net3130[0:47]),
     .sp4_h_r_09(net3131[0:47]), .sp4_h_r_08(net3132[0:47]),
     .sp4_h_r_07(net3133[0:47]), .sp4_h_r_06(net3134[0:47]),
     .sp4_h_r_05(net3135[0:47]), .slf_op_05(net3639[0:7]),
     .slf_op_06(net3638[0:7]), .slf_op_07(net3637[0:7]),
     .slf_op_08(net3636[0:7]), .slf_op_09(net3635[0:7]),
     .slf_op_10(net3634[0:7]), .rgt_op_10(net3142[0:7]),
     .rgt_op_09(net3143[0:7]), .rgt_op_08(net3144[0:7]),
     .rgt_op_07(net3145[0:7]), .rgt_op_06(net3146[0:7]),
     .rgt_op_05(net3147[0:7]), .lft_op_10(net3306[0:7]),
     .lft_op_09(net3307[0:7]), .lft_op_08(net3308[0:7]),
     .lft_op_07(net3309[0:7]), .lft_op_06(net3310[0:7]),
     .lft_op_05(net3311[0:7]), .sp12_h_l_10(net3647[0:23]),
     .sp12_h_r_10(net3155[0:23]), .sp12_h_l_09(net3656[0:23]),
     .sp12_h_l_08(net3655[0:23]), .sp12_h_l_07(net3654[0:23]),
     .sp12_h_l_06(net3653[0:23]), .sp12_h_r_05(net3160[0:23]),
     .sp12_h_r_06(net3161[0:23]), .sp12_h_r_07(net3162[0:23]),
     .sp12_h_r_08(net3163[0:23]), .sp12_h_r_09(net3164[0:23]),
     .sp12_h_l_05(net3652[0:23]), .sp4_r_v_b_05(net3166[0:47]),
     .sp4_r_v_b_06(net3167[0:47]), .sp4_r_v_b_07(net3168[0:47]),
     .sp4_r_v_b_08(net3169[0:47]), .sp4_r_v_b_09(net3170[0:47]),
     .sp4_r_v_b_10(net3171[0:47]), .sp4_v_b_10(net3663[0:47]),
     .sp4_v_b_09(net3662[0:47]), .sp4_v_b_08(net3661[0:47]),
     .sp4_v_b_07(net3660[0:47]), .sp4_v_b_06(net3659[0:47]),
     .sp4_v_b_05(net3658[0:47]), .sp4_v_t_16(sp4_v_t_14_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net3181[0:47]), .sp4_h_r_12(net3182[0:47]),
     .sp4_h_r_13(net3183[0:47]), .sp4_h_r_14(net3184[0:47]),
     .sp4_h_r_15(net3185[0:47]), .sp4_h_r_16(net3186[0:47]),
     .sp4_h_l_16(net3678[0:47]), .sp4_h_l_15(net3677[0:47]),
     .sp4_h_l_14(net3676[0:47]), .sp4_h_l_13(net3675[0:47]),
     .sp4_h_l_12(net3674[0:47]), .sp4_h_l_11(net3673[0:47]),
     .tnr_op_16(tnr_op_14_16[7:0]), .tnl_op_16(tnl_op_14_16[7:0]),
     .lft_op_16(slf_op_13_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net3695[0:7]), .slf_op_14(net3694[0:7]),
     .slf_op_13(net3697[0:7]), .slf_op_12(net3696[0:7]),
     .slf_op_11(net3698[0:7]), .rgt_op_14(net3202[0:7]),
     .rgt_op_15(net3203[0:7]), .rgt_op_12(net3204[0:7]),
     .rgt_op_13(net3205[0:7]), .rgt_op_11(net3206[0:7]),
     .sp4_v_b_16(net3705[0:47]), .sp4_v_b_14(net3708[0:47]),
     .sp4_v_b_15(net3706[0:47]), .sp4_v_b_13(net3707[0:47]),
     .sp4_v_b_11(net3710[0:47]), .sp4_v_b_12(net3709[0:47]),
     .sp4_r_v_b_16(net3213[0:47]), .sp4_r_v_b_15(net3214[0:47]),
     .sp4_r_v_b_13(net3215[0:47]), .sp4_r_v_b_14(net3216[0:47]),
     .sp4_r_v_b_12(net3217[0:47]), .sp4_r_v_b_11(net3218[0:47]),
     .sp12_h_l_16(net3717[0:23]), .sp12_h_l_15(net3719[0:23]),
     .sp12_h_l_14(net3718[0:23]), .sp12_h_l_13(net3721[0:23]),
     .sp12_h_l_12(net3720[0:23]), .sp12_h_l_11(net3722[0:23]),
     .sp12_h_r_16(net3225[0:23]), .sp12_h_r_14(net3226[0:23]),
     .sp12_h_r_15(net3227[0:23]), .sp12_h_r_12(net3228[0:23]),
     .sp12_h_r_13(net3229[0:23]), .sp12_h_r_11(net3230[0:23]),
     .lft_op_14(net3366[0:7]), .lft_op_15(net3367[0:7]),
     .lft_op_12(net3368[0:7]), .lft_op_11(net3370[0:7]),
     .lft_op_13(net3369[0:7]));
array_LT1x16 I_it_12_bot ( .sp12_v_b_01(net4833[0:23]),
     .glb_netwk(net4762[0:7]), .bot_op_01({slf_op_12_00[3],
     slf_op_12_00[2], slf_op_12_00[1], slf_op_12_00[0],
     slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0]}), .sp12_v_t_16(sp12_v_t_12_16[23:0]),
     .rgt_op_16(slf_op_13_16[7:0]), .top_op_16(top_op_12_16[7:0]),
     .rgt_op_03(net3242[0:7]), .slf_op_02(net2260[0:7]),
     .rgt_op_02(net3244[0:7]), .rgt_op_01(net4799[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2432[0:7]), .lft_op_03(net2422[0:7]),
     .lft_op_02(net2424[0:7]), .lft_op_01(net4801[0:7]),
     .rgt_op_04(net3252[0:7]), .carry_in(net5055),
     .bnl_op_01({slf_op_11_00[3], slf_op_11_00[2], slf_op_11_00[1],
     slf_op_11_00[0], slf_op_11_00[3], slf_op_11_00[2],
     slf_op_11_00[1], slf_op_11_00[0]}), .slf_op_04(net2268[0:7]),
     .slf_op_03(net2258[0:7]), .slf_op_01(net4800[0:7]),
     .sp4_h_l_04(net2288[0:47]), .carry_out(carry_out_12_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net3261[0:23]),
     .sp12_h_r_03(net3262[0:23]), .sp12_h_r_02(net3263[0:23]),
     .sp12_h_r_01(net3264[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_12_16[7:0]), .sp4_v_b_01(net4849[0:47]),
     .sp4_r_v_b_04(net3268[0:47]), .sp4_r_v_b_03(net3269[0:47]),
     .sp4_r_v_b_02(net3270[0:47]), .sp4_r_v_b_01(net4848[0:47]),
     .sp4_h_r_04(net3272[0:47]), .sp4_h_r_03(net3273[0:47]),
     .sp4_h_r_02(net3274[0:47]), .sp4_h_r_01(net3275[0:47]),
     .sp4_h_l_03(net2289[0:47]), .sp4_h_l_02(net2290[0:47]),
     .sp4_h_l_01(net2291[0:47]), .bl(bl[653:600]),
     .sp12_h_l_01(net2280[0:23]), .sp12_h_l_02(net2279[0:23]),
     .sp12_h_l_03(net2278[0:23]), .sp12_h_l_04(net2277[0:23]),
     .sp4_v_b_04(net2284[0:47]), .sp4_v_b_03(net2285[0:47]),
     .sp4_v_b_02(net2286[0:47]), .bnr_op_01({slf_op_13_00[3],
     slf_op_13_00[2], slf_op_13_00[1], slf_op_13_00[0],
     slf_op_13_00[3], slf_op_13_00[2], slf_op_13_00[1],
     slf_op_13_00[0]}), .sp4_h_l_05(net2315[0:47]),
     .sp4_h_l_06(net2314[0:47]), .sp4_h_l_07(net2313[0:47]),
     .sp4_h_l_08(net2312[0:47]), .sp4_h_l_09(net2311[0:47]),
     .sp4_h_l_10(net2310[0:47]), .sp4_h_r_10(net3294[0:47]),
     .sp4_h_r_09(net3295[0:47]), .sp4_h_r_08(net3296[0:47]),
     .sp4_h_r_07(net3297[0:47]), .sp4_h_r_06(net3298[0:47]),
     .sp4_h_r_05(net3299[0:47]), .slf_op_05(net2327[0:7]),
     .slf_op_06(net2326[0:7]), .slf_op_07(net2325[0:7]),
     .slf_op_08(net2324[0:7]), .slf_op_09(net2323[0:7]),
     .slf_op_10(net2322[0:7]), .rgt_op_10(net3306[0:7]),
     .rgt_op_09(net3307[0:7]), .rgt_op_08(net3308[0:7]),
     .rgt_op_07(net3309[0:7]), .rgt_op_06(net3310[0:7]),
     .rgt_op_05(net3311[0:7]), .lft_op_10(net2486[0:7]),
     .lft_op_09(net2487[0:7]), .lft_op_08(net2488[0:7]),
     .lft_op_07(net2489[0:7]), .lft_op_06(net2490[0:7]),
     .lft_op_05(net2491[0:7]), .sp12_h_l_10(net2335[0:23]),
     .sp12_h_r_10(net3319[0:23]), .sp12_h_l_09(net2344[0:23]),
     .sp12_h_l_08(net2343[0:23]), .sp12_h_l_07(net2342[0:23]),
     .sp12_h_l_06(net2341[0:23]), .sp12_h_r_05(net3324[0:23]),
     .sp12_h_r_06(net3325[0:23]), .sp12_h_r_07(net3326[0:23]),
     .sp12_h_r_08(net3327[0:23]), .sp12_h_r_09(net3328[0:23]),
     .sp12_h_l_05(net2340[0:23]), .sp4_r_v_b_05(net3330[0:47]),
     .sp4_r_v_b_06(net3331[0:47]), .sp4_r_v_b_07(net3332[0:47]),
     .sp4_r_v_b_08(net3333[0:47]), .sp4_r_v_b_09(net3334[0:47]),
     .sp4_r_v_b_10(net3335[0:47]), .sp4_v_b_10(net2351[0:47]),
     .sp4_v_b_09(net2350[0:47]), .sp4_v_b_08(net2349[0:47]),
     .sp4_v_b_07(net2348[0:47]), .sp4_v_b_06(net2347[0:47]),
     .sp4_v_b_05(net2346[0:47]), .sp4_v_t_16(sp4_v_t_12_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net3345[0:47]), .sp4_h_r_12(net3346[0:47]),
     .sp4_h_r_13(net3347[0:47]), .sp4_h_r_14(net3348[0:47]),
     .sp4_h_r_15(net3349[0:47]), .sp4_h_r_16(net3350[0:47]),
     .sp4_h_l_16(net2366[0:47]), .sp4_h_l_15(net2365[0:47]),
     .sp4_h_l_14(net2364[0:47]), .sp4_h_l_13(net2363[0:47]),
     .sp4_h_l_12(net2362[0:47]), .sp4_h_l_11(net2361[0:47]),
     .tnr_op_16(tnr_op_12_16[7:0]), .tnl_op_16(tnl_op_12_16[7:0]),
     .lft_op_16(slf_op_11_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net2383[0:7]), .slf_op_14(net2382[0:7]),
     .slf_op_13(net2385[0:7]), .slf_op_12(net2384[0:7]),
     .slf_op_11(net2386[0:7]), .rgt_op_14(net3366[0:7]),
     .rgt_op_15(net3367[0:7]), .rgt_op_12(net3368[0:7]),
     .rgt_op_13(net3369[0:7]), .rgt_op_11(net3370[0:7]),
     .sp4_v_b_16(net2393[0:47]), .sp4_v_b_14(net2396[0:47]),
     .sp4_v_b_15(net2394[0:47]), .sp4_v_b_13(net2395[0:47]),
     .sp4_v_b_11(net2398[0:47]), .sp4_v_b_12(net2397[0:47]),
     .sp4_r_v_b_16(net3377[0:47]), .sp4_r_v_b_15(net3378[0:47]),
     .sp4_r_v_b_13(net3379[0:47]), .sp4_r_v_b_14(net3380[0:47]),
     .sp4_r_v_b_12(net3381[0:47]), .sp4_r_v_b_11(net3382[0:47]),
     .sp12_h_l_16(net2405[0:23]), .sp12_h_l_15(net2407[0:23]),
     .sp12_h_l_14(net2406[0:23]), .sp12_h_l_13(net2409[0:23]),
     .sp12_h_l_12(net2408[0:23]), .sp12_h_l_11(net2410[0:23]),
     .sp12_h_r_16(net3389[0:23]), .sp12_h_r_14(net3390[0:23]),
     .sp12_h_r_15(net3391[0:23]), .sp12_h_r_12(net3392[0:23]),
     .sp12_h_r_13(net3393[0:23]), .sp12_h_r_11(net3394[0:23]),
     .lft_op_14(net2546[0:7]), .lft_op_15(net2547[0:7]),
     .lft_op_12(net2548[0:7]), .lft_op_11(net2550[0:7]),
     .lft_op_13(net2549[0:7]));
array_LT1x16 I_it_07_bot ( .sp12_v_b_01(net4838[0:23]),
     .glb_netwk(net4757[0:7]), .bot_op_01({slf_op_07_00[3],
     slf_op_07_00[2], slf_op_07_00[1], slf_op_07_00[0],
     slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0]}), .sp12_v_t_16(sp12_v_t_07_16[23:0]),
     .rgt_op_16(slf_op_08_16[7:0]), .top_op_16(top_op_07_16[7:0]),
     .rgt_op_03(net3406[0:7]), .slf_op_02(net2752[0:7]),
     .rgt_op_02(net3408[0:7]), .rgt_op_01(net4804[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2104[0:7]), .lft_op_03(net2094[0:7]),
     .lft_op_02(net2096[0:7]), .lft_op_01(net4806[0:7]),
     .rgt_op_04(net3416[0:7]), .carry_in(net5051),
     .bnl_op_01({slf_op_06_00[3], slf_op_06_00[2], slf_op_06_00[1],
     slf_op_06_00[0], slf_op_06_00[3], slf_op_06_00[2],
     slf_op_06_00[1], slf_op_06_00[0]}), .slf_op_04(net2760[0:7]),
     .slf_op_03(net2750[0:7]), .slf_op_01(net4805[0:7]),
     .sp4_h_l_04(net2780[0:47]), .carry_out(carry_out_07_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net3425[0:23]),
     .sp12_h_r_03(net3426[0:23]), .sp12_h_r_02(net3427[0:23]),
     .sp12_h_r_01(net3428[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_07_16[7:0]), .sp4_v_b_01(net4854[0:47]),
     .sp4_r_v_b_04(net3432[0:47]), .sp4_r_v_b_03(net3433[0:47]),
     .sp4_r_v_b_02(net3434[0:47]), .sp4_r_v_b_01(net4853[0:47]),
     .sp4_h_r_04(net3436[0:47]), .sp4_h_r_03(net3437[0:47]),
     .sp4_h_r_02(net3438[0:47]), .sp4_h_r_01(net3439[0:47]),
     .sp4_h_l_03(net2781[0:47]), .sp4_h_l_02(net2782[0:47]),
     .sp4_h_l_01(net2783[0:47]), .bl(bl[395:342]),
     .sp12_h_l_01(net2772[0:23]), .sp12_h_l_02(net2771[0:23]),
     .sp12_h_l_03(net2770[0:23]), .sp12_h_l_04(net2769[0:23]),
     .sp4_v_b_04(net2776[0:47]), .sp4_v_b_03(net2777[0:47]),
     .sp4_v_b_02(net2778[0:47]), .bnr_op_01({slf_op_08_00[3],
     slf_op_08_00[2], slf_op_08_00[1], slf_op_08_00[0],
     slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0]}), .sp4_h_l_05(net2807[0:47]),
     .sp4_h_l_06(net2806[0:47]), .sp4_h_l_07(net2805[0:47]),
     .sp4_h_l_08(net2804[0:47]), .sp4_h_l_09(net2803[0:47]),
     .sp4_h_l_10(net2802[0:47]), .sp4_h_r_10(net3458[0:47]),
     .sp4_h_r_09(net3459[0:47]), .sp4_h_r_08(net3460[0:47]),
     .sp4_h_r_07(net3461[0:47]), .sp4_h_r_06(net3462[0:47]),
     .sp4_h_r_05(net3463[0:47]), .slf_op_05(net2819[0:7]),
     .slf_op_06(net2818[0:7]), .slf_op_07(net2817[0:7]),
     .slf_op_08(net2816[0:7]), .slf_op_09(net2815[0:7]),
     .slf_op_10(net2814[0:7]), .rgt_op_10(net3470[0:7]),
     .rgt_op_09(net3471[0:7]), .rgt_op_08(net3472[0:7]),
     .rgt_op_07(net3473[0:7]), .rgt_op_06(net3474[0:7]),
     .rgt_op_05(net3475[0:7]), .lft_op_10(net2158[0:7]),
     .lft_op_09(net2159[0:7]), .lft_op_08(net2160[0:7]),
     .lft_op_07(net2161[0:7]), .lft_op_06(net2162[0:7]),
     .lft_op_05(net2163[0:7]), .sp12_h_l_10(net2827[0:23]),
     .sp12_h_r_10(net3483[0:23]), .sp12_h_l_09(net2836[0:23]),
     .sp12_h_l_08(net2835[0:23]), .sp12_h_l_07(net2834[0:23]),
     .sp12_h_l_06(net2833[0:23]), .sp12_h_r_05(net3488[0:23]),
     .sp12_h_r_06(net3489[0:23]), .sp12_h_r_07(net3490[0:23]),
     .sp12_h_r_08(net3491[0:23]), .sp12_h_r_09(net3492[0:23]),
     .sp12_h_l_05(net2832[0:23]), .sp4_r_v_b_05(net3494[0:47]),
     .sp4_r_v_b_06(net3495[0:47]), .sp4_r_v_b_07(net3496[0:47]),
     .sp4_r_v_b_08(net3497[0:47]), .sp4_r_v_b_09(net3498[0:47]),
     .sp4_r_v_b_10(net3499[0:47]), .sp4_v_b_10(net2843[0:47]),
     .sp4_v_b_09(net2842[0:47]), .sp4_v_b_08(net2841[0:47]),
     .sp4_v_b_07(net2840[0:47]), .sp4_v_b_06(net2839[0:47]),
     .sp4_v_b_05(net2838[0:47]), .sp4_v_t_16(sp4_v_t_07_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net3509[0:47]), .sp4_h_r_12(net3510[0:47]),
     .sp4_h_r_13(net3511[0:47]), .sp4_h_r_14(net3512[0:47]),
     .sp4_h_r_15(net3513[0:47]), .sp4_h_r_16(net3514[0:47]),
     .sp4_h_l_16(net2858[0:47]), .sp4_h_l_15(net2857[0:47]),
     .sp4_h_l_14(net2856[0:47]), .sp4_h_l_13(net2855[0:47]),
     .sp4_h_l_12(net2854[0:47]), .sp4_h_l_11(net2853[0:47]),
     .tnr_op_16(tnr_op_07_16[7:0]), .tnl_op_16(tnl_op_07_16[7:0]),
     .lft_op_16(slf_op_06_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net2875[0:7]), .slf_op_14(net2874[0:7]),
     .slf_op_13(net2877[0:7]), .slf_op_12(net2876[0:7]),
     .slf_op_11(net2878[0:7]), .rgt_op_14(net3530[0:7]),
     .rgt_op_15(net3531[0:7]), .rgt_op_12(net3532[0:7]),
     .rgt_op_13(net3533[0:7]), .rgt_op_11(net3534[0:7]),
     .sp4_v_b_16(net2885[0:47]), .sp4_v_b_14(net2888[0:47]),
     .sp4_v_b_15(net2886[0:47]), .sp4_v_b_13(net2887[0:47]),
     .sp4_v_b_11(net2890[0:47]), .sp4_v_b_12(net2889[0:47]),
     .sp4_r_v_b_16(net3541[0:47]), .sp4_r_v_b_15(net3542[0:47]),
     .sp4_r_v_b_13(net3543[0:47]), .sp4_r_v_b_14(net3544[0:47]),
     .sp4_r_v_b_12(net3545[0:47]), .sp4_r_v_b_11(net3546[0:47]),
     .sp12_h_l_16(net2897[0:23]), .sp12_h_l_15(net2899[0:23]),
     .sp12_h_l_14(net2898[0:23]), .sp12_h_l_13(net2901[0:23]),
     .sp12_h_l_12(net2900[0:23]), .sp12_h_l_11(net2902[0:23]),
     .sp12_h_r_16(net3553[0:23]), .sp12_h_r_14(net3554[0:23]),
     .sp12_h_r_15(net3555[0:23]), .sp12_h_r_12(net3556[0:23]),
     .sp12_h_r_13(net3557[0:23]), .sp12_h_r_11(net3558[0:23]),
     .lft_op_14(net2218[0:7]), .lft_op_15(net2219[0:7]),
     .lft_op_12(net2220[0:7]), .lft_op_11(net2222[0:7]),
     .lft_op_13(net2221[0:7]));
array_LT1x16 I_it_13_bot ( .sp12_v_b_01(net4832[0:23]),
     .glb_netwk(net4763[0:7]), .bot_op_01({slf_op_13_00[3],
     slf_op_13_00[2], slf_op_13_00[1], slf_op_13_00[0],
     slf_op_13_00[3], slf_op_13_00[2], slf_op_13_00[1],
     slf_op_13_00[0]}), .sp12_v_t_16(sp12_v_t_13_16[23:0]),
     .rgt_op_16(slf_op_14_16[7:0]), .top_op_16(top_op_13_16[7:0]),
     .rgt_op_03(net3570[0:7]), .slf_op_02(net3244[0:7]),
     .rgt_op_02(net3572[0:7]), .rgt_op_01(net4798[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2268[0:7]), .lft_op_03(net2258[0:7]),
     .lft_op_02(net2260[0:7]), .lft_op_01(net4800[0:7]),
     .rgt_op_04(net3580[0:7]), .carry_in(net4994),
     .bnl_op_01({slf_op_12_00[3], slf_op_12_00[2], slf_op_12_00[1],
     slf_op_12_00[0], slf_op_12_00[3], slf_op_12_00[2],
     slf_op_12_00[1], slf_op_12_00[0]}), .slf_op_04(net3252[0:7]),
     .slf_op_03(net3242[0:7]), .slf_op_01(net4799[0:7]),
     .sp4_h_l_04(net3272[0:47]), .carry_out(carry_out_13_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net3589[0:23]),
     .sp12_h_r_03(net3590[0:23]), .sp12_h_r_02(net3591[0:23]),
     .sp12_h_r_01(net3592[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_13_16[7:0]), .sp4_v_b_01(net4848[0:47]),
     .sp4_r_v_b_04(net3596[0:47]), .sp4_r_v_b_03(net3597[0:47]),
     .sp4_r_v_b_02(net3598[0:47]), .sp4_r_v_b_01(net4847[0:47]),
     .sp4_h_r_04(net3600[0:47]), .sp4_h_r_03(net3601[0:47]),
     .sp4_h_r_02(net3602[0:47]), .sp4_h_r_01(net3603[0:47]),
     .sp4_h_l_03(net3273[0:47]), .sp4_h_l_02(net3274[0:47]),
     .sp4_h_l_01(net3275[0:47]), .bl(bl[707:654]),
     .sp12_h_l_01(net3264[0:23]), .sp12_h_l_02(net3263[0:23]),
     .sp12_h_l_03(net3262[0:23]), .sp12_h_l_04(net3261[0:23]),
     .sp4_v_b_04(net3268[0:47]), .sp4_v_b_03(net3269[0:47]),
     .sp4_v_b_02(net3270[0:47]), .bnr_op_01({slf_op_14_00[3],
     slf_op_14_00[2], slf_op_14_00[1], slf_op_14_00[0],
     slf_op_14_00[3], slf_op_14_00[2], slf_op_14_00[1],
     slf_op_14_00[0]}), .sp4_h_l_05(net3299[0:47]),
     .sp4_h_l_06(net3298[0:47]), .sp4_h_l_07(net3297[0:47]),
     .sp4_h_l_08(net3296[0:47]), .sp4_h_l_09(net3295[0:47]),
     .sp4_h_l_10(net3294[0:47]), .sp4_h_r_10(net3622[0:47]),
     .sp4_h_r_09(net3623[0:47]), .sp4_h_r_08(net3624[0:47]),
     .sp4_h_r_07(net3625[0:47]), .sp4_h_r_06(net3626[0:47]),
     .sp4_h_r_05(net3627[0:47]), .slf_op_05(net3311[0:7]),
     .slf_op_06(net3310[0:7]), .slf_op_07(net3309[0:7]),
     .slf_op_08(net3308[0:7]), .slf_op_09(net3307[0:7]),
     .slf_op_10(net3306[0:7]), .rgt_op_10(net3634[0:7]),
     .rgt_op_09(net3635[0:7]), .rgt_op_08(net3636[0:7]),
     .rgt_op_07(net3637[0:7]), .rgt_op_06(net3638[0:7]),
     .rgt_op_05(net3639[0:7]), .lft_op_10(net2322[0:7]),
     .lft_op_09(net2323[0:7]), .lft_op_08(net2324[0:7]),
     .lft_op_07(net2325[0:7]), .lft_op_06(net2326[0:7]),
     .lft_op_05(net2327[0:7]), .sp12_h_l_10(net3319[0:23]),
     .sp12_h_r_10(net3647[0:23]), .sp12_h_l_09(net3328[0:23]),
     .sp12_h_l_08(net3327[0:23]), .sp12_h_l_07(net3326[0:23]),
     .sp12_h_l_06(net3325[0:23]), .sp12_h_r_05(net3652[0:23]),
     .sp12_h_r_06(net3653[0:23]), .sp12_h_r_07(net3654[0:23]),
     .sp12_h_r_08(net3655[0:23]), .sp12_h_r_09(net3656[0:23]),
     .sp12_h_l_05(net3324[0:23]), .sp4_r_v_b_05(net3658[0:47]),
     .sp4_r_v_b_06(net3659[0:47]), .sp4_r_v_b_07(net3660[0:47]),
     .sp4_r_v_b_08(net3661[0:47]), .sp4_r_v_b_09(net3662[0:47]),
     .sp4_r_v_b_10(net3663[0:47]), .sp4_v_b_10(net3335[0:47]),
     .sp4_v_b_09(net3334[0:47]), .sp4_v_b_08(net3333[0:47]),
     .sp4_v_b_07(net3332[0:47]), .sp4_v_b_06(net3331[0:47]),
     .sp4_v_b_05(net3330[0:47]), .sp4_v_t_16(sp4_v_t_13_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net3673[0:47]), .sp4_h_r_12(net3674[0:47]),
     .sp4_h_r_13(net3675[0:47]), .sp4_h_r_14(net3676[0:47]),
     .sp4_h_r_15(net3677[0:47]), .sp4_h_r_16(net3678[0:47]),
     .sp4_h_l_16(net3350[0:47]), .sp4_h_l_15(net3349[0:47]),
     .sp4_h_l_14(net3348[0:47]), .sp4_h_l_13(net3347[0:47]),
     .sp4_h_l_12(net3346[0:47]), .sp4_h_l_11(net3345[0:47]),
     .tnr_op_16(tnr_op_13_16[7:0]), .tnl_op_16(tnl_op_13_16[7:0]),
     .lft_op_16(slf_op_12_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net3367[0:7]), .slf_op_14(net3366[0:7]),
     .slf_op_13(net3369[0:7]), .slf_op_12(net3368[0:7]),
     .slf_op_11(net3370[0:7]), .rgt_op_14(net3694[0:7]),
     .rgt_op_15(net3695[0:7]), .rgt_op_12(net3696[0:7]),
     .rgt_op_13(net3697[0:7]), .rgt_op_11(net3698[0:7]),
     .sp4_v_b_16(net3377[0:47]), .sp4_v_b_14(net3380[0:47]),
     .sp4_v_b_15(net3378[0:47]), .sp4_v_b_13(net3379[0:47]),
     .sp4_v_b_11(net3382[0:47]), .sp4_v_b_12(net3381[0:47]),
     .sp4_r_v_b_16(net3705[0:47]), .sp4_r_v_b_15(net3706[0:47]),
     .sp4_r_v_b_13(net3707[0:47]), .sp4_r_v_b_14(net3708[0:47]),
     .sp4_r_v_b_12(net3709[0:47]), .sp4_r_v_b_11(net3710[0:47]),
     .sp12_h_l_16(net3389[0:23]), .sp12_h_l_15(net3391[0:23]),
     .sp12_h_l_14(net3390[0:23]), .sp12_h_l_13(net3393[0:23]),
     .sp12_h_l_12(net3392[0:23]), .sp12_h_l_11(net3394[0:23]),
     .sp12_h_r_16(net3717[0:23]), .sp12_h_r_14(net3718[0:23]),
     .sp12_h_r_15(net3719[0:23]), .sp12_h_r_12(net3720[0:23]),
     .sp12_h_r_13(net3721[0:23]), .sp12_h_r_11(net3722[0:23]),
     .lft_op_14(net2382[0:7]), .lft_op_15(net2383[0:7]),
     .lft_op_12(net2384[0:7]), .lft_op_11(net2386[0:7]),
     .lft_op_13(net2385[0:7]));
array_LT1x16 I_it_09_bot ( .sp12_v_b_01(net4836[0:23]),
     .glb_netwk(net4759[0:7]), .bot_op_01({slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0],
     slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0]}), .sp12_v_t_16(sp12_v_t_09_16[23:0]),
     .rgt_op_16(slf_op_10_16[7:0]), .top_op_16(top_op_09_16[7:0]),
     .rgt_op_03(net3734[0:7]), .slf_op_02(net4663[0:7]),
     .rgt_op_02(net3736[0:7]), .rgt_op_01(net4802[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3416[0:7]), .lft_op_03(net3406[0:7]),
     .lft_op_02(net3408[0:7]), .lft_op_01(net4804[0:7]),
     .rgt_op_04(net3744[0:7]), .carry_in(net4999),
     .bnl_op_01({slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0], slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0]}), .slf_op_04(net4665[0:7]),
     .slf_op_03(net4664[0:7]), .slf_op_01(net4803[0:7]),
     .sp4_h_l_04(net4684[0:47]), .carry_out(carry_out_09_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net3753[0:23]),
     .sp12_h_r_03(net3754[0:23]), .sp12_h_r_02(net3755[0:23]),
     .sp12_h_r_01(net3756[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_09_16[7:0]), .sp4_v_b_01(net4852[0:47]),
     .sp4_r_v_b_04(net3760[0:47]), .sp4_r_v_b_03(net3761[0:47]),
     .sp4_r_v_b_02(net3762[0:47]), .sp4_r_v_b_01(net4851[0:47]),
     .sp4_h_r_04(net3764[0:47]), .sp4_h_r_03(net3765[0:47]),
     .sp4_h_r_02(net3766[0:47]), .sp4_h_r_01(net3767[0:47]),
     .sp4_h_l_03(net4683[0:47]), .sp4_h_l_02(net4682[0:47]),
     .sp4_h_l_01(net4681[0:47]), .bl(bl[491:438]),
     .sp12_h_l_01(net4561[0:23]), .sp12_h_l_02(net4641[0:23]),
     .sp12_h_l_03(net4640[0:23]), .sp12_h_l_04(net4639[0:23]),
     .sp4_v_b_04(net4578[0:47]), .sp4_v_b_03(net4577[0:47]),
     .sp4_v_b_02(net4576[0:47]), .bnr_op_01({slf_op_10_00[3],
     slf_op_10_00[2], slf_op_10_00[1], slf_op_10_00[0],
     slf_op_10_00[3], slf_op_10_00[2], slf_op_10_00[1],
     slf_op_10_00[0]}), .sp4_h_l_05(net4685[0:47]),
     .sp4_h_l_06(net4686[0:47]), .sp4_h_l_07(net4687[0:47]),
     .sp4_h_l_08(net4688[0:47]), .sp4_h_l_09(net4573[0:47]),
     .sp4_h_l_10(net4689[0:47]), .sp4_h_r_10(net3786[0:47]),
     .sp4_h_r_09(net3787[0:47]), .sp4_h_r_08(net3788[0:47]),
     .sp4_h_r_07(net3789[0:47]), .sp4_h_r_06(net3790[0:47]),
     .sp4_h_r_05(net3791[0:47]), .slf_op_05(net4666[0:7]),
     .slf_op_06(net4667[0:7]), .slf_op_07(net4668[0:7]),
     .slf_op_08(net4669[0:7]), .slf_op_09(net4670[0:7]),
     .slf_op_10(net4671[0:7]), .rgt_op_10(net3798[0:7]),
     .rgt_op_09(net3799[0:7]), .rgt_op_08(net3800[0:7]),
     .rgt_op_07(net3801[0:7]), .rgt_op_06(net3802[0:7]),
     .rgt_op_05(net3803[0:7]), .lft_op_10(net3470[0:7]),
     .lft_op_09(net3471[0:7]), .lft_op_08(net3472[0:7]),
     .lft_op_07(net3473[0:7]), .lft_op_06(net3474[0:7]),
     .lft_op_05(net3475[0:7]), .sp12_h_l_10(net4621[0:23]),
     .sp12_h_r_10(net3811[0:23]), .sp12_h_l_09(net4634[0:23]),
     .sp12_h_l_08(net4635[0:23]), .sp12_h_l_07(net4636[0:23]),
     .sp12_h_l_06(net4637[0:23]), .sp12_h_r_05(net3816[0:23]),
     .sp12_h_r_06(net3817[0:23]), .sp12_h_r_07(net3818[0:23]),
     .sp12_h_r_08(net3819[0:23]), .sp12_h_r_09(net3820[0:23]),
     .sp12_h_l_05(net4638[0:23]), .sp4_r_v_b_05(net3822[0:47]),
     .sp4_r_v_b_06(net3823[0:47]), .sp4_r_v_b_07(net3824[0:47]),
     .sp4_r_v_b_08(net3825[0:47]), .sp4_r_v_b_09(net3826[0:47]),
     .sp4_r_v_b_10(net3827[0:47]), .sp4_v_b_10(net4584[0:47]),
     .sp4_v_b_09(net4583[0:47]), .sp4_v_b_08(net4582[0:47]),
     .sp4_v_b_07(net4581[0:47]), .sp4_v_b_06(net4580[0:47]),
     .sp4_v_b_05(net4579[0:47]), .sp4_v_t_16(sp4_v_t_09_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net3837[0:47]), .sp4_h_r_12(net3838[0:47]),
     .sp4_h_r_13(net3839[0:47]), .sp4_h_r_14(net3840[0:47]),
     .sp4_h_r_15(net3841[0:47]), .sp4_h_r_16(net3842[0:47]),
     .sp4_h_l_16(net4695[0:47]), .sp4_h_l_15(net4694[0:47]),
     .sp4_h_l_14(net4693[0:47]), .sp4_h_l_13(net4692[0:47]),
     .sp4_h_l_12(net4691[0:47]), .sp4_h_l_11(net4690[0:47]),
     .tnr_op_16(tnr_op_09_16[7:0]), .tnl_op_16(tnl_op_09_16[7:0]),
     .lft_op_16(slf_op_08_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net4676[0:7]), .slf_op_14(net4675[0:7]),
     .slf_op_13(net4674[0:7]), .slf_op_12(net4673[0:7]),
     .slf_op_11(net4672[0:7]), .rgt_op_14(net3858[0:7]),
     .rgt_op_15(net3859[0:7]), .rgt_op_12(net3860[0:7]),
     .rgt_op_13(net3861[0:7]), .rgt_op_11(net3862[0:7]),
     .sp4_v_b_16(net4589[0:47]), .sp4_v_b_14(net4588[0:47]),
     .sp4_v_b_15(net4590[0:47]), .sp4_v_b_13(net4587[0:47]),
     .sp4_v_b_11(net4585[0:47]), .sp4_v_b_12(net4586[0:47]),
     .sp4_r_v_b_16(net3869[0:47]), .sp4_r_v_b_15(net3870[0:47]),
     .sp4_r_v_b_13(net3871[0:47]), .sp4_r_v_b_14(net3872[0:47]),
     .sp4_r_v_b_12(net3873[0:47]), .sp4_r_v_b_11(net3874[0:47]),
     .sp12_h_l_16(net4626[0:23]), .sp12_h_l_15(net4622[0:23]),
     .sp12_h_l_14(net4625[0:23]), .sp12_h_l_13(net4631[0:23]),
     .sp12_h_l_12(net4632[0:23]), .sp12_h_l_11(net4633[0:23]),
     .sp12_h_r_16(net3881[0:23]), .sp12_h_r_14(net3882[0:23]),
     .sp12_h_r_15(net3883[0:23]), .sp12_h_r_12(net3884[0:23]),
     .sp12_h_r_13(net3885[0:23]), .sp12_h_r_11(net3886[0:23]),
     .lft_op_14(net3530[0:7]), .lft_op_15(net3531[0:7]),
     .lft_op_12(net3532[0:7]), .lft_op_11(net3534[0:7]),
     .lft_op_13(net3533[0:7]));
array_LT1x16 I_lt_02bot ( .sp12_v_b_01(net4843[0:23]),
     .glb_netwk(net4752[0:7]), .bot_op_01({slf_op_02_00[3],
     slf_op_02_00[2], slf_op_02_00[1], slf_op_02_00[0],
     slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0]}), .sp12_v_t_16(sp12_v_t_02_16[23:0]),
     .rgt_op_16(slf_op_03_16[7:0]), .top_op_16(top_op_02_16[7:0]),
     .rgt_op_03(net3898[0:7]), .slf_op_02(net4064[0:7]),
     .rgt_op_02(net3900[0:7]), .rgt_op_01(net4809[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4920[0:7]), .lft_op_03(net4919[0:7]),
     .lft_op_02(net4883[0:7]), .lft_op_01(net4811[0:7]),
     .rgt_op_04(net3908[0:7]), .carry_in(net5058),
     .bnl_op_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}), .slf_op_04(net4072[0:7]),
     .slf_op_03(net4062[0:7]), .slf_op_01(net4810[0:7]),
     .sp4_h_l_04(net4092[0:47]), .carry_out(carry_out_02_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net3917[0:23]),
     .sp12_h_r_03(net3918[0:23]), .sp12_h_r_02(net3919[0:23]),
     .sp12_h_r_01(net3920[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_02_16[7:0]), .sp4_v_b_01(net4859[0:47]),
     .sp4_r_v_b_04(net3924[0:47]), .sp4_r_v_b_03(net3925[0:47]),
     .sp4_r_v_b_02(net3926[0:47]), .sp4_r_v_b_01(net4858[0:47]),
     .sp4_h_r_04(net3928[0:47]), .sp4_h_r_03(net3929[0:47]),
     .sp4_h_r_02(net3930[0:47]), .sp4_h_r_01(net3931[0:47]),
     .sp4_h_l_03(net4093[0:47]), .sp4_h_l_02(net4094[0:47]),
     .sp4_h_l_01(net4095[0:47]), .bl(bl[125:72]),
     .sp12_h_l_01(net4084[0:23]), .sp12_h_l_02(net4083[0:23]),
     .sp12_h_l_03(net4082[0:23]), .sp12_h_l_04(net4081[0:23]),
     .sp4_v_b_04(net4088[0:47]), .sp4_v_b_03(net4089[0:47]),
     .sp4_v_b_02(net4090[0:47]), .bnr_op_01({slf_op_03_00[3],
     slf_op_03_00[2], slf_op_03_00[1], slf_op_03_00[0],
     slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0]}), .sp4_h_l_05(net4119[0:47]),
     .sp4_h_l_06(net4118[0:47]), .sp4_h_l_07(net4117[0:47]),
     .sp4_h_l_08(net4116[0:47]), .sp4_h_l_09(net4115[0:47]),
     .sp4_h_l_10(net4114[0:47]), .sp4_h_r_10(net3950[0:47]),
     .sp4_h_r_09(net3951[0:47]), .sp4_h_r_08(net3952[0:47]),
     .sp4_h_r_07(net3953[0:47]), .sp4_h_r_06(net3954[0:47]),
     .sp4_h_r_05(net3955[0:47]), .slf_op_05(net4131[0:7]),
     .slf_op_06(net4130[0:7]), .slf_op_07(net4129[0:7]),
     .slf_op_08(net4128[0:7]), .slf_op_09(net4127[0:7]),
     .slf_op_10(net4126[0:7]), .rgt_op_10(net3962[0:7]),
     .rgt_op_09(net3963[0:7]), .rgt_op_08(net3964[0:7]),
     .rgt_op_07(net3965[0:7]), .rgt_op_06(net3966[0:7]),
     .rgt_op_05(net3967[0:7]), .lft_op_10(net4914[0:7]),
     .lft_op_09(net4913[0:7]), .lft_op_08(net4908[0:7]),
     .lft_op_07(net4916[0:7]), .lft_op_06(net4915[0:7]),
     .lft_op_05(net4909[0:7]), .sp12_h_l_10(net4139[0:23]),
     .sp12_h_r_10(net3975[0:23]), .sp12_h_l_09(net4148[0:23]),
     .sp12_h_l_08(net4147[0:23]), .sp12_h_l_07(net4146[0:23]),
     .sp12_h_l_06(net4145[0:23]), .sp12_h_r_05(net3980[0:23]),
     .sp12_h_r_06(net3981[0:23]), .sp12_h_r_07(net3982[0:23]),
     .sp12_h_r_08(net3983[0:23]), .sp12_h_r_09(net3984[0:23]),
     .sp12_h_l_05(net4144[0:23]), .sp4_r_v_b_05(net3986[0:47]),
     .sp4_r_v_b_06(net3987[0:47]), .sp4_r_v_b_07(net3988[0:47]),
     .sp4_r_v_b_08(net3989[0:47]), .sp4_r_v_b_09(net3990[0:47]),
     .sp4_r_v_b_10(net3991[0:47]), .sp4_v_b_10(net4155[0:47]),
     .sp4_v_b_09(net4154[0:47]), .sp4_v_b_08(net4153[0:47]),
     .sp4_v_b_07(net4152[0:47]), .sp4_v_b_06(net4151[0:47]),
     .sp4_v_b_05(net4150[0:47]), .sp4_v_t_16(sp4_v_t_02_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net4001[0:47]), .sp4_h_r_12(net4002[0:47]),
     .sp4_h_r_13(net4003[0:47]), .sp4_h_r_14(net4004[0:47]),
     .sp4_h_r_15(net4005[0:47]), .sp4_h_r_16(net4006[0:47]),
     .sp4_h_l_16(net4170[0:47]), .sp4_h_l_15(net4169[0:47]),
     .sp4_h_l_14(net4168[0:47]), .sp4_h_l_13(net4167[0:47]),
     .sp4_h_l_12(net4166[0:47]), .sp4_h_l_11(net4165[0:47]),
     .tnr_op_16(tnr_op_02_16[7:0]), .tnl_op_16(tnl_op_02_16[7:0]),
     .lft_op_16(slf_op_01_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net4187[0:7]), .slf_op_14(net4186[0:7]),
     .slf_op_13(net4189[0:7]), .slf_op_12(net4188[0:7]),
     .slf_op_11(net4190[0:7]), .rgt_op_14(net4022[0:7]),
     .rgt_op_15(net4023[0:7]), .rgt_op_12(net4024[0:7]),
     .rgt_op_13(net4025[0:7]), .rgt_op_11(net4026[0:7]),
     .sp4_v_b_16(net4197[0:47]), .sp4_v_b_14(net4200[0:47]),
     .sp4_v_b_15(net4198[0:47]), .sp4_v_b_13(net4199[0:47]),
     .sp4_v_b_11(net4202[0:47]), .sp4_v_b_12(net4201[0:47]),
     .sp4_r_v_b_16(net4033[0:47]), .sp4_r_v_b_15(net4034[0:47]),
     .sp4_r_v_b_13(net4035[0:47]), .sp4_r_v_b_14(net4036[0:47]),
     .sp4_r_v_b_12(net4037[0:47]), .sp4_r_v_b_11(net4038[0:47]),
     .sp12_h_l_16(net4209[0:23]), .sp12_h_l_15(net4211[0:23]),
     .sp12_h_l_14(net4210[0:23]), .sp12_h_l_13(net4213[0:23]),
     .sp12_h_l_12(net4212[0:23]), .sp12_h_l_11(net4214[0:23]),
     .sp12_h_r_16(net4045[0:23]), .sp12_h_r_14(net4046[0:23]),
     .sp12_h_r_15(net4047[0:23]), .sp12_h_r_12(net4048[0:23]),
     .sp12_h_r_13(net4049[0:23]), .sp12_h_r_11(net4050[0:23]),
     .lft_op_14(net4904[0:7]), .lft_op_15(net4905[0:7]),
     .lft_op_12(net4911[0:7]), .lft_op_11(net4907[0:7]),
     .lft_op_13(net4912[0:7]));
array_LT1x16 I_lt_01bot ( .sp12_v_b_01(net4844[0:23]),
     .glb_netwk(net4751[0:7]), .bot_op_01({slf_op_01_00[3],
     slf_op_01_00[2], slf_op_01_00[1], slf_op_01_00[0],
     slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0]}), .sp12_v_t_16(sp12_v_t_01_16[23:0]),
     .rgt_op_16(slf_op_02_16[7:0]), .top_op_16(top_op_01_16[7:0]),
     .rgt_op_03(net4062[0:7]), .slf_op_02(net4883[0:7]),
     .rgt_op_02(net4064[0:7]), .rgt_op_01(net4810[0:7]), .purst(purst),
     .prog(prog), .lft_op_04({slf_op_00_04[3], slf_op_00_04[2],
     slf_op_00_04[1], slf_op_00_04[0], slf_op_00_04[3],
     slf_op_00_04[2], slf_op_00_04[1], slf_op_00_04[0]}),
     .lft_op_03({slf_op_00_03[3], slf_op_00_03[2], slf_op_00_03[1],
     slf_op_00_03[0], slf_op_00_03[3], slf_op_00_03[2],
     slf_op_00_03[1], slf_op_00_03[0]}), .lft_op_02({slf_op_00_02[3],
     slf_op_00_02[2], slf_op_00_02[1], slf_op_00_02[0],
     slf_op_00_02[3], slf_op_00_02[2], slf_op_00_02[1],
     slf_op_00_02[0]}), .lft_op_01({slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0], slf_op_00_01[3],
     slf_op_00_01[2], slf_op_00_01[1], slf_op_00_01[0]}),
     .rgt_op_04(net4072[0:7]), .carry_in(net5037), .bnl_op_01({tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .slf_op_04(net4920[0:7]), .slf_op_03(net4919[0:7]),
     .slf_op_01(net4811[0:7]), .sp4_h_l_04(net4900[0:47]),
     .carry_out(carry_out_01_16), .vdd_cntl(vdd_cntl_l[271:16]),
     .sp12_h_r_04(net4081[0:23]), .sp12_h_r_03(net4082[0:23]),
     .sp12_h_r_02(net4083[0:23]), .sp12_h_r_01(net4084[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(slf_op_01_16[7:0]),
     .sp4_v_b_01(net4860[0:47]), .sp4_r_v_b_04(net4088[0:47]),
     .sp4_r_v_b_03(net4089[0:47]), .sp4_r_v_b_02(net4090[0:47]),
     .sp4_r_v_b_01(net4859[0:47]), .sp4_h_r_04(net4092[0:47]),
     .sp4_h_r_03(net4093[0:47]), .sp4_h_r_02(net4094[0:47]),
     .sp4_h_r_01(net4095[0:47]), .sp4_h_l_03(net4903[0:47]),
     .sp4_h_l_02(net4902[0:47]), .sp4_h_l_01(net4952[0:47]),
     .bl(bl[71:18]), .sp12_h_l_01(net4893[0:23]),
     .sp12_h_l_02(net4936[0:23]), .sp12_h_l_03(net4935[0:23]),
     .sp12_h_l_04(net4934[0:23]), .sp4_v_b_04(net4104[0:47]),
     .sp4_v_b_03(net4105[0:47]), .sp4_v_b_02(net4106[0:47]),
     .bnr_op_01({slf_op_02_00[3], slf_op_02_00[2], slf_op_02_00[1],
     slf_op_02_00[0], slf_op_02_00[3], slf_op_02_00[2],
     slf_op_02_00[1], slf_op_02_00[0]}), .sp4_h_l_05(net4901[0:47]),
     .sp4_h_l_06(net4898[0:47]), .sp4_h_l_07(net4899[0:47]),
     .sp4_h_l_08(net4951[0:47]), .sp4_h_l_09(net4950[0:47]),
     .sp4_h_l_10(net4949[0:47]), .sp4_h_r_10(net4114[0:47]),
     .sp4_h_r_09(net4115[0:47]), .sp4_h_r_08(net4116[0:47]),
     .sp4_h_r_07(net4117[0:47]), .sp4_h_r_06(net4118[0:47]),
     .sp4_h_r_05(net4119[0:47]), .slf_op_05(net4909[0:7]),
     .slf_op_06(net4915[0:7]), .slf_op_07(net4916[0:7]),
     .slf_op_08(net4908[0:7]), .slf_op_09(net4913[0:7]),
     .slf_op_10(net4914[0:7]), .rgt_op_10(net4126[0:7]),
     .rgt_op_09(net4127[0:7]), .rgt_op_08(net4128[0:7]),
     .rgt_op_07(net4129[0:7]), .rgt_op_06(net4130[0:7]),
     .rgt_op_05(net4131[0:7]), .lft_op_10({slf_op_00_10[3],
     slf_op_00_10[2], slf_op_00_10[1], slf_op_00_10[0],
     slf_op_00_10[3], slf_op_00_10[2], slf_op_00_10[1],
     slf_op_00_10[0]}), .lft_op_09({slf_op_00_09[3], slf_op_00_09[2],
     slf_op_00_09[1], slf_op_00_09[0], slf_op_00_09[3],
     slf_op_00_09[2], slf_op_00_09[1], slf_op_00_09[0]}),
     .lft_op_08({slf_op_00_08[3], slf_op_00_08[2], slf_op_00_08[1],
     slf_op_00_08[0], slf_op_00_08[3], slf_op_00_08[2],
     slf_op_00_08[1], slf_op_00_08[0]}), .lft_op_07({slf_op_00_07[3],
     slf_op_00_07[2], slf_op_00_07[1], slf_op_00_07[0],
     slf_op_00_07[3], slf_op_00_07[2], slf_op_00_07[1],
     slf_op_00_07[0]}), .lft_op_06({slf_op_00_06[3], slf_op_00_06[2],
     slf_op_00_06[1], slf_op_00_06[0], slf_op_00_06[3],
     slf_op_00_06[2], slf_op_00_06[1], slf_op_00_06[0]}),
     .lft_op_05({slf_op_00_05[3], slf_op_00_05[2], slf_op_00_05[1],
     slf_op_00_05[0], slf_op_00_05[3], slf_op_00_05[2],
     slf_op_00_05[1], slf_op_00_05[0]}), .sp12_h_l_10(net4928[0:23]),
     .sp12_h_r_10(net4139[0:23]), .sp12_h_l_09(net4929[0:23]),
     .sp12_h_l_08(net4930[0:23]), .sp12_h_l_07(net4931[0:23]),
     .sp12_h_l_06(net4932[0:23]), .sp12_h_r_05(net4144[0:23]),
     .sp12_h_r_06(net4145[0:23]), .sp12_h_r_07(net4146[0:23]),
     .sp12_h_r_08(net4147[0:23]), .sp12_h_r_09(net4148[0:23]),
     .sp12_h_l_05(net4933[0:23]), .sp4_r_v_b_05(net4150[0:47]),
     .sp4_r_v_b_06(net4151[0:47]), .sp4_r_v_b_07(net4152[0:47]),
     .sp4_r_v_b_08(net4153[0:47]), .sp4_r_v_b_09(net4154[0:47]),
     .sp4_r_v_b_10(net4155[0:47]), .sp4_v_b_10(net4156[0:47]),
     .sp4_v_b_09(net4157[0:47]), .sp4_v_b_08(net4158[0:47]),
     .sp4_v_b_07(net4159[0:47]), .sp4_v_b_06(net4160[0:47]),
     .sp4_v_b_05(net4161[0:47]), .sp4_v_t_16(sp4_v_t_01_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net4165[0:47]), .sp4_h_r_12(net4166[0:47]),
     .sp4_h_r_13(net4167[0:47]), .sp4_h_r_14(net4168[0:47]),
     .sp4_h_r_15(net4169[0:47]), .sp4_h_r_16(net4170[0:47]),
     .sp4_h_l_16(net4938[0:47]), .sp4_h_l_15(net4944[0:47]),
     .sp4_h_l_14(net4945[0:47]), .sp4_h_l_13(net4946[0:47]),
     .sp4_h_l_12(net4947[0:47]), .sp4_h_l_11(net4948[0:47]),
     .tnr_op_16(tnr_op_01_16[7:0]), .tnl_op_16(tnl_op_01_16[7:0]),
     .lft_op_16({slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0], slf_op_00_16[3], slf_op_00_16[2],
     slf_op_00_16[1], slf_op_00_16[0]}), .wl(wl_l[271:16]),
     .slf_op_15(net4905[0:7]), .slf_op_14(net4904[0:7]),
     .slf_op_13(net4912[0:7]), .slf_op_12(net4911[0:7]),
     .slf_op_11(net4907[0:7]), .rgt_op_14(net4186[0:7]),
     .rgt_op_15(net4187[0:7]), .rgt_op_12(net4188[0:7]),
     .rgt_op_13(net4189[0:7]), .rgt_op_11(net4190[0:7]),
     .sp4_v_b_16(net4191[0:47]), .sp4_v_b_14(net4192[0:47]),
     .sp4_v_b_15(net4193[0:47]), .sp4_v_b_13(net4194[0:47]),
     .sp4_v_b_11(net4195[0:47]), .sp4_v_b_12(net4196[0:47]),
     .sp4_r_v_b_16(net4197[0:47]), .sp4_r_v_b_15(net4198[0:47]),
     .sp4_r_v_b_13(net4199[0:47]), .sp4_r_v_b_14(net4200[0:47]),
     .sp4_r_v_b_12(net4201[0:47]), .sp4_r_v_b_11(net4202[0:47]),
     .sp12_h_l_16(net4922[0:23]), .sp12_h_l_15(net4923[0:23]),
     .sp12_h_l_14(net4924[0:23]), .sp12_h_l_13(net4925[0:23]),
     .sp12_h_l_12(net4926[0:23]), .sp12_h_l_11(net4927[0:23]),
     .sp12_h_r_16(net4209[0:23]), .sp12_h_r_14(net4210[0:23]),
     .sp12_h_r_15(net4211[0:23]), .sp12_h_r_12(net4212[0:23]),
     .sp12_h_r_13(net4213[0:23]), .sp12_h_r_11(net4214[0:23]),
     .lft_op_14({slf_op_00_14[3], slf_op_00_14[2], slf_op_00_14[1],
     slf_op_00_14[0], slf_op_00_14[3], slf_op_00_14[2],
     slf_op_00_14[1], slf_op_00_14[0]}), .lft_op_15({slf_op_00_15[3],
     slf_op_00_15[2], slf_op_00_15[1], slf_op_00_15[0],
     slf_op_00_15[3], slf_op_00_15[2], slf_op_00_15[1],
     slf_op_00_15[0]}), .lft_op_12({slf_op_00_12[3], slf_op_00_12[2],
     slf_op_00_12[1], slf_op_00_12[0], slf_op_00_12[3],
     slf_op_00_12[2], slf_op_00_12[1], slf_op_00_12[0]}),
     .lft_op_11({slf_op_00_11[3], slf_op_00_11[2], slf_op_00_11[1],
     slf_op_00_11[0], slf_op_00_11[3], slf_op_00_11[2],
     slf_op_00_11[1], slf_op_00_11[0]}), .lft_op_13({slf_op_00_13[3],
     slf_op_00_13[2], slf_op_00_13[1], slf_op_00_13[0],
     slf_op_00_13[3], slf_op_00_13[2], slf_op_00_13[1],
     slf_op_00_13[0]}));
array_LT1x16 I_it_16_bot ( .sp12_v_b_01(net4829[0:23]),
     .glb_netwk(net4766[0:7]), .bot_op_01({slf_op_16_00[3],
     slf_op_16_00[2], slf_op_16_00[1], slf_op_16_00[0],
     slf_op_16_00[3], slf_op_16_00[2], slf_op_16_00[1],
     slf_op_16_00[0]}), .sp12_v_t_16(sp12_v_t_16_16[23:0]),
     .rgt_op_16(rgt_op_16_16[7:0]), .top_op_16(top_op_16_16[7:0]),
     .rgt_op_03(rgt_op_16_03[7:0]), .slf_op_02(slf_op_16_02[7:0]),
     .rgt_op_02(rgt_op_16_02[7:0]), .rgt_op_01(rgt_op_16_01[7:0]),
     .purst(purst), .prog(prog), .lft_op_04(net3088[0:7]),
     .lft_op_03(net3078[0:7]), .lft_op_02(net3080[0:7]),
     .lft_op_01(net4797[0:7]), .rgt_op_04(rgt_op_16_04[7:0]),
     .carry_in(net4985), .bnl_op_01({slf_op_15_00[3], slf_op_15_00[2],
     slf_op_15_00[1], slf_op_15_00[0], slf_op_15_00[3],
     slf_op_15_00[2], slf_op_15_00[1], slf_op_15_00[0]}),
     .slf_op_04(slf_op_16_04[7:0]), .slf_op_03(slf_op_16_03[7:0]),
     .slf_op_01(slf_op_16_01[7:0]), .sp4_h_l_04(net2616[0:47]),
     .carry_out(carry_out_16_16), .vdd_cntl(vdd_cntl_l[271:16]),
     .sp12_h_r_04(sp12_h_r_16_04[23:0]),
     .sp12_h_r_03(sp12_h_r_16_03[23:0]),
     .sp12_h_r_02(sp12_h_r_16_02[23:0]),
     .sp12_h_r_01(sp12_h_r_16_01[23:0]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(slf_op_16_16[7:0]),
     .sp4_v_b_01(net4845[0:47]), .sp4_r_v_b_04(sp4_r_v_b_16_04[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_16_03[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_16_02[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_16_01[47:0]),
     .sp4_h_r_04(sp4_h_r_16_04[47:0]),
     .sp4_h_r_03(sp4_h_r_16_03[47:0]),
     .sp4_h_r_02(sp4_h_r_16_02[47:0]),
     .sp4_h_r_01(sp4_h_r_16_01[47:0]), .sp4_h_l_03(net2617[0:47]),
     .sp4_h_l_02(net2618[0:47]), .sp4_h_l_01(net2619[0:47]),
     .bl(bl[869:816]), .sp12_h_l_01(net2608[0:23]),
     .sp12_h_l_02(net2607[0:23]), .sp12_h_l_03(net2606[0:23]),
     .sp12_h_l_04(net2605[0:23]), .sp4_v_b_04(net2612[0:47]),
     .sp4_v_b_03(net2613[0:47]), .sp4_v_b_02(net2614[0:47]),
     .bnr_op_01({bnr_op_16_01[3], bnr_op_16_01[2], bnr_op_16_01[1],
     bnr_op_16_01[0], bnr_op_16_01[3], bnr_op_16_01[2],
     bnr_op_16_01[1], bnr_op_16_01[0]}), .sp4_h_l_05(net2643[0:47]),
     .sp4_h_l_06(net2642[0:47]), .sp4_h_l_07(net2641[0:47]),
     .sp4_h_l_08(net2640[0:47]), .sp4_h_l_09(net2639[0:47]),
     .sp4_h_l_10(net2638[0:47]), .sp4_h_r_10(sp4_h_r_16_10[47:0]),
     .sp4_h_r_09(sp4_h_r_16_09[47:0]),
     .sp4_h_r_08(sp4_h_r_16_08[47:0]),
     .sp4_h_r_07(sp4_h_r_16_07[47:0]),
     .sp4_h_r_06(sp4_h_r_16_06[47:0]),
     .sp4_h_r_05(sp4_h_r_16_05[47:0]), .slf_op_05(slf_op_16_05[7:0]),
     .slf_op_06(slf_op_16_06[7:0]), .slf_op_07(slf_op_16_07[7:0]),
     .slf_op_08(slf_op_16_08[7:0]), .slf_op_09(slf_op_16_09[7:0]),
     .slf_op_10(slf_op_16_10[7:0]), .rgt_op_10(rgt_op_16_10[7:0]),
     .rgt_op_09(rgt_op_16_09[7:0]), .rgt_op_08(rgt_op_16_08[7:0]),
     .rgt_op_07(rgt_op_16_07[7:0]), .rgt_op_06(rgt_op_16_06[7:0]),
     .rgt_op_05(rgt_op_16_05[7:0]), .lft_op_10(net3142[0:7]),
     .lft_op_09(net3143[0:7]), .lft_op_08(net3144[0:7]),
     .lft_op_07(net3145[0:7]), .lft_op_06(net3146[0:7]),
     .lft_op_05(net3147[0:7]), .sp12_h_l_10(net2663[0:23]),
     .sp12_h_r_10(sp12_h_r_16_10[23:0]), .sp12_h_l_09(net2672[0:23]),
     .sp12_h_l_08(net2671[0:23]), .sp12_h_l_07(net2670[0:23]),
     .sp12_h_l_06(net2669[0:23]), .sp12_h_r_05(sp12_h_r_16_05[23:0]),
     .sp12_h_r_06(sp12_h_r_16_06[23:0]),
     .sp12_h_r_07(sp12_h_r_16_07[23:0]),
     .sp12_h_r_08(sp12_h_r_16_08[23:0]),
     .sp12_h_r_09(sp12_h_r_16_09[23:0]), .sp12_h_l_05(net2668[0:23]),
     .sp4_r_v_b_05(sp4_r_v_b_16_05[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_16_06[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_16_07[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_16_08[47:0]),
     .sp4_r_v_b_09(sp4_r_v_b_16_09[47:0]),
     .sp4_r_v_b_10(sp4_r_v_b_16_10[47:0]), .sp4_v_b_10(net2679[0:47]),
     .sp4_v_b_09(net2678[0:47]), .sp4_v_b_08(net2677[0:47]),
     .sp4_v_b_07(net2676[0:47]), .sp4_v_b_06(net2675[0:47]),
     .sp4_v_b_05(net2674[0:47]), .sp4_v_t_16(sp4_v_t_16_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(sp4_h_r_16_11[47:0]),
     .sp4_h_r_12(sp4_h_r_16_12[47:0]),
     .sp4_h_r_13(sp4_h_r_16_13[47:0]),
     .sp4_h_r_14(sp4_h_r_16_14[47:0]),
     .sp4_h_r_15(sp4_h_r_16_15[47:0]),
     .sp4_h_r_16(sp4_h_r_16_16[47:0]), .sp4_h_l_16(net2694[0:47]),
     .sp4_h_l_15(net2693[0:47]), .sp4_h_l_14(net2692[0:47]),
     .sp4_h_l_13(net2691[0:47]), .sp4_h_l_12(net2690[0:47]),
     .sp4_h_l_11(net2689[0:47]), .tnr_op_16(tnr_op_16_16[7:0]),
     .tnl_op_16(tnl_op_16_16[7:0]), .lft_op_16(slf_op_15_16[7:0]),
     .wl(wl_l[271:16]), .slf_op_15(slf_op_16_15[7:0]),
     .slf_op_14(slf_op_16_14[7:0]), .slf_op_13(slf_op_16_13[7:0]),
     .slf_op_12(slf_op_16_12[7:0]), .slf_op_11(slf_op_16_11[7:0]),
     .rgt_op_14(rgt_op_16_14[7:0]), .rgt_op_15(rgt_op_16_15[7:0]),
     .rgt_op_12(rgt_op_16_12[7:0]), .rgt_op_13(rgt_op_16_13[7:0]),
     .rgt_op_11(rgt_op_16_11[7:0]), .sp4_v_b_16(net2721[0:47]),
     .sp4_v_b_14(net2724[0:47]), .sp4_v_b_15(net2722[0:47]),
     .sp4_v_b_13(net2723[0:47]), .sp4_v_b_11(net2726[0:47]),
     .sp4_v_b_12(net2725[0:47]), .sp4_r_v_b_16(sp4_r_v_b_16_16[47:0]),
     .sp4_r_v_b_15(sp4_r_v_b_16_15[47:0]),
     .sp4_r_v_b_13(sp4_r_v_b_16_13[47:0]),
     .sp4_r_v_b_14(sp4_r_v_b_16_14[47:0]),
     .sp4_r_v_b_12(sp4_r_v_b_16_12[47:0]),
     .sp4_r_v_b_11(sp4_r_v_b_16_11[47:0]), .sp12_h_l_16(net2733[0:23]),
     .sp12_h_l_15(net2735[0:23]), .sp12_h_l_14(net2734[0:23]),
     .sp12_h_l_13(net2737[0:23]), .sp12_h_l_12(net2736[0:23]),
     .sp12_h_l_11(net2738[0:23]), .sp12_h_r_16(sp12_h_r_16_16[23:0]),
     .sp12_h_r_14(sp12_h_r_16_14[23:0]),
     .sp12_h_r_15(sp12_h_r_16_15[23:0]),
     .sp12_h_r_12(sp12_h_r_16_12[23:0]),
     .sp12_h_r_13(sp12_h_r_16_13[23:0]),
     .sp12_h_r_11(sp12_h_r_16_11[23:0]), .lft_op_14(net3202[0:7]),
     .lft_op_15(net3203[0:7]), .lft_op_12(net3204[0:7]),
     .lft_op_11(net3206[0:7]), .lft_op_13(net3205[0:7]));
array_LT1x16 I_it_04_bot ( .sp12_v_b_01(net4841[0:23]),
     .glb_netwk(net4754[0:7]), .bot_op_01({slf_op_04_00[3],
     slf_op_04_00[2], slf_op_04_00[1], slf_op_04_00[0],
     slf_op_04_00[3], slf_op_04_00[2], slf_op_04_00[1],
     slf_op_04_00[0]}), .sp12_v_t_16(sp12_v_t_04_16[23:0]),
     .rgt_op_16(slf_op_05_16[7:0]), .top_op_16(top_op_04_16[7:0]),
     .rgt_op_03(net4390[0:7]), .slf_op_02(net2916[0:7]),
     .rgt_op_02(net4392[0:7]), .rgt_op_01(net4807[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3908[0:7]), .lft_op_03(net3898[0:7]),
     .lft_op_02(net3900[0:7]), .lft_op_01(net4809[0:7]),
     .rgt_op_04(net4400[0:7]), .carry_in(net5057),
     .bnl_op_01({slf_op_03_00[3], slf_op_03_00[2], slf_op_03_00[1],
     slf_op_03_00[0], slf_op_03_00[3], slf_op_03_00[2],
     slf_op_03_00[1], slf_op_03_00[0]}), .slf_op_04(net2924[0:7]),
     .slf_op_03(net2914[0:7]), .slf_op_01(net4808[0:7]),
     .sp4_h_l_04(net2944[0:47]), .carry_out(carry_out_04_16),
     .vdd_cntl(vdd_cntl_l[271:16]), .sp12_h_r_04(net4409[0:23]),
     .sp12_h_r_03(net4410[0:23]), .sp12_h_r_02(net4411[0:23]),
     .sp12_h_r_01(net4412[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_04_16[7:0]), .sp4_v_b_01(net4857[0:47]),
     .sp4_r_v_b_04(net4416[0:47]), .sp4_r_v_b_03(net4417[0:47]),
     .sp4_r_v_b_02(net4418[0:47]), .sp4_r_v_b_01(net4856[0:47]),
     .sp4_h_r_04(net4420[0:47]), .sp4_h_r_03(net4421[0:47]),
     .sp4_h_r_02(net4422[0:47]), .sp4_h_r_01(net4423[0:47]),
     .sp4_h_l_03(net2945[0:47]), .sp4_h_l_02(net2946[0:47]),
     .sp4_h_l_01(net2947[0:47]), .bl(bl[233:180]),
     .sp12_h_l_01(net2936[0:23]), .sp12_h_l_02(net2935[0:23]),
     .sp12_h_l_03(net2934[0:23]), .sp12_h_l_04(net2933[0:23]),
     .sp4_v_b_04(net2940[0:47]), .sp4_v_b_03(net2941[0:47]),
     .sp4_v_b_02(net2942[0:47]), .bnr_op_01({slf_op_05_00[3],
     slf_op_05_00[2], slf_op_05_00[1], slf_op_05_00[0],
     slf_op_05_00[3], slf_op_05_00[2], slf_op_05_00[1],
     slf_op_05_00[0]}), .sp4_h_l_05(net2971[0:47]),
     .sp4_h_l_06(net2970[0:47]), .sp4_h_l_07(net2969[0:47]),
     .sp4_h_l_08(net2968[0:47]), .sp4_h_l_09(net2967[0:47]),
     .sp4_h_l_10(net2966[0:47]), .sp4_h_r_10(net4442[0:47]),
     .sp4_h_r_09(net4443[0:47]), .sp4_h_r_08(net4444[0:47]),
     .sp4_h_r_07(net4445[0:47]), .sp4_h_r_06(net4446[0:47]),
     .sp4_h_r_05(net4447[0:47]), .slf_op_05(net2983[0:7]),
     .slf_op_06(net2982[0:7]), .slf_op_07(net2981[0:7]),
     .slf_op_08(net2980[0:7]), .slf_op_09(net2979[0:7]),
     .slf_op_10(net2978[0:7]), .rgt_op_10(net4454[0:7]),
     .rgt_op_09(net4455[0:7]), .rgt_op_08(net4456[0:7]),
     .rgt_op_07(net4457[0:7]), .rgt_op_06(net4458[0:7]),
     .rgt_op_05(net4459[0:7]), .lft_op_10(net3962[0:7]),
     .lft_op_09(net3963[0:7]), .lft_op_08(net3964[0:7]),
     .lft_op_07(net3965[0:7]), .lft_op_06(net3966[0:7]),
     .lft_op_05(net3967[0:7]), .sp12_h_l_10(net2991[0:23]),
     .sp12_h_r_10(net4467[0:23]), .sp12_h_l_09(net3000[0:23]),
     .sp12_h_l_08(net2999[0:23]), .sp12_h_l_07(net2998[0:23]),
     .sp12_h_l_06(net2997[0:23]), .sp12_h_r_05(net4472[0:23]),
     .sp12_h_r_06(net4473[0:23]), .sp12_h_r_07(net4474[0:23]),
     .sp12_h_r_08(net4475[0:23]), .sp12_h_r_09(net4476[0:23]),
     .sp12_h_l_05(net2996[0:23]), .sp4_r_v_b_05(net4478[0:47]),
     .sp4_r_v_b_06(net4479[0:47]), .sp4_r_v_b_07(net4480[0:47]),
     .sp4_r_v_b_08(net4481[0:47]), .sp4_r_v_b_09(net4482[0:47]),
     .sp4_r_v_b_10(net4483[0:47]), .sp4_v_b_10(net3007[0:47]),
     .sp4_v_b_09(net3006[0:47]), .sp4_v_b_08(net3005[0:47]),
     .sp4_v_b_07(net3004[0:47]), .sp4_v_b_06(net3003[0:47]),
     .sp4_v_b_05(net3002[0:47]), .sp4_v_t_16(sp4_v_t_04_16[47:0]),
     .pgate(pgate_l[271:16]), .reset_b(reset_l[271:16]),
     .sp4_h_r_11(net4493[0:47]), .sp4_h_r_12(net4494[0:47]),
     .sp4_h_r_13(net4495[0:47]), .sp4_h_r_14(net4496[0:47]),
     .sp4_h_r_15(net4497[0:47]), .sp4_h_r_16(net4498[0:47]),
     .sp4_h_l_16(net3022[0:47]), .sp4_h_l_15(net3021[0:47]),
     .sp4_h_l_14(net3020[0:47]), .sp4_h_l_13(net3019[0:47]),
     .sp4_h_l_12(net3018[0:47]), .sp4_h_l_11(net3017[0:47]),
     .tnr_op_16(tnr_op_04_16[7:0]), .tnl_op_16(tnl_op_04_16[7:0]),
     .lft_op_16(slf_op_03_16[7:0]), .wl(wl_l[271:16]),
     .slf_op_15(net3039[0:7]), .slf_op_14(net3038[0:7]),
     .slf_op_13(net3041[0:7]), .slf_op_12(net3040[0:7]),
     .slf_op_11(net3042[0:7]), .rgt_op_14(net4514[0:7]),
     .rgt_op_15(net4515[0:7]), .rgt_op_12(net4516[0:7]),
     .rgt_op_13(net4517[0:7]), .rgt_op_11(net4518[0:7]),
     .sp4_v_b_16(net3049[0:47]), .sp4_v_b_14(net3052[0:47]),
     .sp4_v_b_15(net3050[0:47]), .sp4_v_b_13(net3051[0:47]),
     .sp4_v_b_11(net3054[0:47]), .sp4_v_b_12(net3053[0:47]),
     .sp4_r_v_b_16(net4525[0:47]), .sp4_r_v_b_15(net4526[0:47]),
     .sp4_r_v_b_13(net4527[0:47]), .sp4_r_v_b_14(net4528[0:47]),
     .sp4_r_v_b_12(net4529[0:47]), .sp4_r_v_b_11(net4530[0:47]),
     .sp12_h_l_16(net3061[0:23]), .sp12_h_l_15(net3063[0:23]),
     .sp12_h_l_14(net3062[0:23]), .sp12_h_l_13(net3065[0:23]),
     .sp12_h_l_12(net3064[0:23]), .sp12_h_l_11(net3066[0:23]),
     .sp12_h_r_16(net4537[0:23]), .sp12_h_r_14(net4538[0:23]),
     .sp12_h_r_15(net4539[0:23]), .sp12_h_r_12(net4540[0:23]),
     .sp12_h_r_13(net4541[0:23]), .sp12_h_r_11(net4542[0:23]),
     .lft_op_14(net4022[0:7]), .lft_op_15(net4023[0:7]),
     .lft_op_12(net4024[0:7]), .lft_op_11(net4026[0:7]),
     .lft_op_13(net4025[0:7]));
array_BRAM_1x8bot I_bram_08_bot ( .glb_netwk(net4758[0:7]),
     .wl(wl_l[271:16]), .pgate(pgate_l[271:16]),
     .vdd_cntl(vdd_cntl_l[271:16]), .reset_b(reset_l[271:16]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sdo_i(bm_sdo_i[1:0]),
     .sp12_h_r_01(net4561[0:23]), .lft_op_10(net2814[0:7]),
     .sp4_h_l_04(net3436[0:47]), .sp4_h_l_06(net3462[0:47]),
     .lft_op_09(net2815[0:7]), .lft_op_08(net2816[0:7]),
     .lft_op_06(net2818[0:7]), .lft_op_07(net2817[0:7]),
     .lft_op_05(net2819[0:7]), .lft_op_03(net2750[0:7]),
     .lft_op_04(net2760[0:7]), .lft_op_02(net2752[0:7]),
     .sp4_h_r_09(net4573[0:47]), .bnr_op_01({slf_op_09_00[3],
     slf_op_09_00[2], slf_op_09_00[1], slf_op_09_00[0],
     slf_op_09_00[3], slf_op_09_00[2], slf_op_09_00[1],
     slf_op_09_00[0]}), .sp4_r_v_b_01(net4852[0:47]),
     .sp4_r_v_b_02(net4576[0:47]), .sp4_r_v_b_03(net4577[0:47]),
     .sp4_r_v_b_04(net4578[0:47]), .sp4_r_v_b_05(net4579[0:47]),
     .sp4_r_v_b_06(net4580[0:47]), .sp4_r_v_b_07(net4581[0:47]),
     .sp4_r_v_b_08(net4582[0:47]), .sp4_r_v_b_09(net4583[0:47]),
     .sp4_r_v_b_10(net4584[0:47]), .sp4_r_v_b_11(net4585[0:47]),
     .sp4_r_v_b_12(net4586[0:47]), .sp4_r_v_b_13(net4587[0:47]),
     .sp4_r_v_b_14(net4588[0:47]), .sp4_r_v_b_16(net4589[0:47]),
     .sp4_r_v_b_15(net4590[0:47]), .bnl_op_01({slf_op_07_00[3],
     slf_op_07_00[2], slf_op_07_00[1], slf_op_07_00[0],
     slf_op_07_00[3], slf_op_07_00[2], slf_op_07_00[1],
     slf_op_07_00[0]}), .lft_op_01(net4805[0:7]),
     .bot_op_01({slf_op_08_00[3], slf_op_08_00[2], slf_op_08_00[1],
     slf_op_08_00[0], slf_op_08_00[3], slf_op_08_00[2],
     slf_op_08_00[1], slf_op_08_00[0]}), .sp12_v_b_01(net4837[0:23]),
     .sp4_v_b_16(net3541[0:47]), .sp4_v_b_15(net3542[0:47]),
     .sp4_v_b_14(net3544[0:47]), .sp4_v_b_13(net3543[0:47]),
     .sp4_v_b_12(net3545[0:47]), .sp4_v_b_11(net3546[0:47]),
     .sp4_v_b_10(net3499[0:47]), .sp4_v_b_09(net3498[0:47]),
     .sp4_v_b_08(net3497[0:47]), .sp4_v_b_07(net3496[0:47]),
     .sp4_v_b_06(net3495[0:47]), .sp4_v_b_05(net3494[0:47]),
     .sp4_v_b_04(net3432[0:47]), .sp4_v_b_03(net3433[0:47]),
     .sp4_v_b_02(net3434[0:47]), .sp4_v_b_01(net4853[0:47]),
     .sp12_h_l_10(net3483[0:23]), .sp12_h_l_09(net3492[0:23]),
     .sp12_h_l_08(net3491[0:23]), .sp12_h_l_07(net3490[0:23]),
     .sp12_h_l_06(net3489[0:23]), .sp12_h_l_05(net3488[0:23]),
     .sp12_h_l_04(net3425[0:23]), .sp12_h_l_03(net3426[0:23]),
     .sp12_h_l_02(net3427[0:23]), .sp12_h_l_01(net3428[0:23]),
     .sp12_h_r_10(net4621[0:23]), .sp12_h_r_15(net4622[0:23]),
     .sp12_h_l_15(net3555[0:23]), .sp12_h_l_14(net3554[0:23]),
     .sp12_h_r_14(net4625[0:23]), .sp12_h_r_16(net4626[0:23]),
     .sp12_h_l_16(net3553[0:23]), .sp12_h_l_13(net3557[0:23]),
     .sp12_h_l_12(net3556[0:23]), .sp12_h_l_11(net3558[0:23]),
     .sp12_h_r_13(net4631[0:23]), .sp12_h_r_12(net4632[0:23]),
     .sp12_h_r_11(net4633[0:23]), .sp12_h_r_09(net4634[0:23]),
     .sp12_h_r_08(net4635[0:23]), .sp12_h_r_07(net4636[0:23]),
     .sp12_h_r_06(net4637[0:23]), .sp12_h_r_05(net4638[0:23]),
     .sp12_h_r_04(net4639[0:23]), .sp12_h_r_03(net4640[0:23]),
     .sp12_h_r_02(net4641[0:23]), .lft_op_14(net2874[0:7]),
     .lft_op_13(net2877[0:7]), .lft_op_12(net2876[0:7]),
     .lft_op_11(net2878[0:7]), .lft_op_15(net2875[0:7]),
     .slf_op_15(net3531[0:7]), .slf_op_14(net3530[0:7]),
     .slf_op_13(net3533[0:7]), .slf_op_12(net3532[0:7]),
     .slf_op_11(net3534[0:7]), .slf_op_10(net3470[0:7]),
     .slf_op_09(net3471[0:7]), .slf_op_08(net3472[0:7]),
     .slf_op_07(net3473[0:7]), .slf_op_06(net3474[0:7]),
     .slf_op_05(net3475[0:7]), .slf_op_04(net3416[0:7]),
     .slf_op_03(net3406[0:7]), .slf_op_01(net4804[0:7]),
     .slf_op_02(net3408[0:7]), .rgt_op_01(net4803[0:7]),
     .rgt_op_02(net4663[0:7]), .rgt_op_03(net4664[0:7]),
     .rgt_op_04(net4665[0:7]), .rgt_op_05(net4666[0:7]),
     .rgt_op_06(net4667[0:7]), .rgt_op_07(net4668[0:7]),
     .rgt_op_08(net4669[0:7]), .rgt_op_09(net4670[0:7]),
     .rgt_op_10(net4671[0:7]), .rgt_op_11(net4672[0:7]),
     .rgt_op_12(net4673[0:7]), .rgt_op_13(net4674[0:7]),
     .rgt_op_14(net4675[0:7]), .rgt_op_15(net4676[0:7]),
     .sp4_h_l_05(net3463[0:47]), .sp4_h_l_02(net3438[0:47]),
     .sp4_h_l_03(net3437[0:47]), .sp4_h_l_01(net3439[0:47]),
     .sp4_h_r_01(net4681[0:47]), .sp4_h_r_02(net4682[0:47]),
     .sp4_h_r_03(net4683[0:47]), .sp4_h_r_04(net4684[0:47]),
     .sp4_h_r_05(net4685[0:47]), .sp4_h_r_06(net4686[0:47]),
     .sp4_h_r_07(net4687[0:47]), .sp4_h_r_08(net4688[0:47]),
     .sp4_h_r_10(net4689[0:47]), .sp4_h_r_11(net4690[0:47]),
     .sp4_h_r_12(net4691[0:47]), .sp4_h_r_13(net4692[0:47]),
     .sp4_h_r_14(net4693[0:47]), .sp4_h_r_15(net4694[0:47]),
     .sp4_h_r_16(net4695[0:47]), .lft_op_16(slf_op_07_16[7:0]),
     .tnl_op_16(tnl_op_08_16[7:0]), .sp4_v_t_16(sp4_v_t_08_16[47:0]),
     .top_op_16(top_op_08_16[7:0]), .slf_op_16(slf_op_08_16[7:0]),
     .tnr_op_16(tnr_op_08_16[7:0]), .sp12_v_t_16(sp12_v_t_08_16[23:0]),
     .rgt_op_16(slf_op_09_16[7:0]), .sp4_h_l_16(net3514[0:47]),
     .sp4_h_l_14(net3512[0:47]), .sp4_h_l_15(net3513[0:47]),
     .sp4_h_l_13(net3511[0:47]), .sp4_h_l_12(net3510[0:47]),
     .sp4_h_l_11(net3509[0:47]), .sp4_h_l_10(net3458[0:47]),
     .sp4_h_l_09(net3459[0:47]), .sp4_h_l_08(net3460[0:47]),
     .sp4_h_l_07(net3461[0:47]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_sreb_o(bm_sreb_o), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .bl(bl[437:396]), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]));
preio_bot_l I_preIO_1to16_00 ( .ceb_o(ceb_o), .ceb_i(net4863),
     .tnr_op_16_00(rgt_op_16_01[7:0]),
     .fabric_out_16_00(fabric_out_16_00), .padin_80(padin_80),
     .sp4_h_r_16_00(sp4_h_r_16_00[15:0]), .bs_en_i(net4980),
     .r_i(net4976), .hiz_b_i(net4958), .update_i(net4961),
     .shift_i(net4954), .mode_i(net4956), .tclk_i(net2076),
     .hold_b_l(hold_b_l), .bs_en_o(bs_en_o), .r_o(r_o),
     .hiz_b_o(hiz_b_o), .update_o(update_o), .shift_o(shift_o),
     .mode_o(mode_o), .tclk_o(tclk_o), .bl_04(bl[233:180]),
     .glb_net_01(net4751[0:7]), .glb_net_02(net4752[0:7]),
     .glb_net_03(net4753[0:7]), .glb_net_04(net4754[0:7]),
     .glb_net_05(net4755[0:7]), .glb_net_06(net4756[0:7]),
     .glb_net_07(net4757[0:7]), .glb_net_08(net4758[0:7]),
     .glb_net_09(net4759[0:7]), .glb_net_10(net4760[0:7]),
     .glb_net_11(net4761[0:7]), .glb_net_12(net4762[0:7]),
     .glb_net_13(net4763[0:7]), .glb_net_14(net4764[0:7]),
     .glb_net_15(net4765[0:7]), .glb_net_16(net4766[0:7]),
     .sp4_v_t_00_01(net4910[0:15]), .tievdd(tievdd), .tiegnd(tiegnd),
     .cf_b(cf_b[383:0]), .padeb_b(padeb_b[29:0]),
     .pado_b(pado_b[29:0]), .padin_b(padin_b[29:0]),
     .pgate_l({pgate_l[1], pgate_l[0], pgate_l[2], pgate_l[3],
     pgate_l[5], pgate_l[4], pgate_l[6], pgate_l[7], pgate_l[9],
     pgate_l[8], pgate_l[10], pgate_l[11], pgate_l[13], pgate_l[12],
     pgate_l[14], pgate_l[15]}), .reset_l({reset_l[1], reset_l[0],
     reset_l[2], reset_l[3], reset_l[5], reset_l[4], reset_l[6],
     reset_l[7], reset_l[9], reset_l[8], reset_l[10], reset_l[11],
     reset_l[13], reset_l[12], reset_l[14], reset_l[15]}),
     .vdd_cntl_l({vdd_cntl_l[1], vdd_cntl_l[0], vdd_cntl_l[2],
     vdd_cntl_l[3], vdd_cntl_l[5], vdd_cntl_l[4], vdd_cntl_l[6],
     vdd_cntl_l[7], vdd_cntl_l[9], vdd_cntl_l[8], vdd_cntl_l[10],
     vdd_cntl_l[11], vdd_cntl_l[13], vdd_cntl_l[12], vdd_cntl_l[14],
     vdd_cntl_l[15]}), .wl_l({wl_l[1], wl_l[0], wl_l[2], wl_l[3],
     wl_l[5], wl_l[4], wl_l[6], wl_l[7], wl_l[9], wl_l[8], wl_l[10],
     wl_l[11], wl_l[13], wl_l[12], wl_l[14], wl_l[15]}),
     .bl_16(bl[869:816]), .bl_15(bl[815:762]), .bl_14(bl[761:708]),
     .bl_13(bl[707:654]), .bl_12(bl[653:600]), .bl_11(bl[599:546]),
     .bl_10(bl[545:492]), .bl_09(bl[491:438]), .bl_08(bl[437:396]),
     .bl_07(bl[395:342]), .bl_06(bl[341:288]), .bl_05(bl[287:234]),
     .bl_03(bl[179:126]), .bl_02(bl[125:72]), .bl_01(bl[71:18]),
     .tnl_op_01_00({slf_op_00_01[3], slf_op_00_01[2], slf_op_00_01[1],
     slf_op_00_01[0], slf_op_00_01[3], slf_op_00_01[2],
     slf_op_00_01[1], slf_op_00_01[0]}), .sdi(net4965), .prog(prog),
     .lft_op_16_00(slf_op_16_01[7:0]), .lft_op_15_00(net4797[0:7]),
     .lft_op_14_00(net4798[0:7]), .lft_op_13_00(net4799[0:7]),
     .lft_op_12_00(net4800[0:7]), .lft_op_11_00(net4801[0:7]),
     .lft_op_10_00(net4802[0:7]), .lft_op_09_00(net4803[0:7]),
     .lft_op_08_00(net4804[0:7]), .lft_op_07_00(net4805[0:7]),
     .lft_op_06_00(net4806[0:7]), .lft_op_05_00(net4807[0:7]),
     .lft_op_04_00(net4808[0:7]), .lft_op_03_00(net4809[0:7]),
     .lft_op_02_00(net4810[0:7]), .lft_op_01_00(net4811[0:7]),
     .slf_op_16_00(slf_op_16_00[3:0]),
     .slf_op_15_00(slf_op_15_00[3:0]),
     .slf_op_14_00(slf_op_14_00[3:0]),
     .slf_op_13_00(slf_op_13_00[3:0]),
     .slf_op_12_00(slf_op_12_00[3:0]),
     .slf_op_11_00(slf_op_11_00[3:0]),
     .slf_op_10_00(slf_op_10_00[3:0]),
     .slf_op_09_00(slf_op_09_00[3:0]),
     .slf_op_08_00(slf_op_08_00[3:0]),
     .slf_op_07_00(slf_op_07_00[3:0]),
     .slf_op_06_00(slf_op_06_00[3:0]),
     .slf_op_05_00(slf_op_05_00[3:0]),
     .slf_op_04_00(slf_op_04_00[3:0]),
     .slf_op_03_00(slf_op_03_00[3:0]),
     .slf_op_02_00(slf_op_02_00[3:0]),
     .slf_op_01_00(slf_op_01_00[3:0]), .sdo(sdo),
     .sp12_h_l_16_00(net4829[0:23]), .sp12_h_l_15_00(net4830[0:23]),
     .sp12_h_l_14_00(net4831[0:23]), .sp12_h_l_13_00(net4832[0:23]),
     .sp12_h_l_12_00(net4833[0:23]), .sp12_h_l_11_00(net4834[0:23]),
     .sp12_h_l_10_00(net4835[0:23]), .sp12_h_l_09_00(net4836[0:23]),
     .sp12_h_l_08_00(net4837[0:23]), .sp12_h_l_07_00(net4838[0:23]),
     .sp12_h_l_06_00(net4839[0:23]), .sp12_h_l_05_00(net4840[0:23]),
     .sp12_h_l_04_00(net4841[0:23]), .sp12_h_l_03_00(net4842[0:23]),
     .sp12_h_l_02_00(net4843[0:23]), .sp12_h_l_01_00(net4844[0:23]),
     .sp4_h_l_16_00(net4845[0:47]), .sp4_h_l_15_00(net4846[0:47]),
     .sp4_h_l_14_00(net4847[0:47]), .sp4_h_l_13_00(net4848[0:47]),
     .sp4_h_l_12_00(net4849[0:47]), .sp4_h_l_11_00(net4850[0:47]),
     .sp4_h_l_10_00(net4851[0:47]), .sp4_h_l_09_00(net4852[0:47]),
     .sp4_h_l_08_00(net4853[0:47]), .sp4_h_l_07_00(net4854[0:47]),
     .sp4_h_l_06_00(net4855[0:47]), .sp4_h_l_05_00(net4856[0:47]),
     .sp4_h_l_04_00(net4857[0:47]), .sp4_h_l_03_00(net4858[0:47]),
     .sp4_h_l_02_00(net4859[0:47]), .sp4_h_l_01_00(net4860[0:47]));
array_LFT_IO_1x16 I_io_00bot ( .tnl_op_16(tnr_op_00_16[7:0]),
     .bnl_op_01({slf_op_01_00[3], slf_op_01_00[2], slf_op_01_00[1],
     slf_op_01_00[0], slf_op_01_00[3], slf_op_01_00[2],
     slf_op_01_00[1], slf_op_01_00[0]}), .ceb(net4863),
     .pado(pado_l[23:0]), .padin(padin_l[23:0]), .padeb(padeb_l[23:0]),
     .fabric_out_16(net2084), .fabric_out_15(net2086),
     .fabric_out_14(net4993), .fabric_out_13(net4997),
     .fabric_out_12(net4992), .fabric_out_11(net5038),
     .fabric_out_01(net4988), .fabric_out_02(net5048),
     .fabric_out_03(net4991), .fabric_out_04(net5049),
     .fabric_out_05(net4995), .fabric_out_06(net4998),
     .fabric_out_07(net5024), .fabric_out_08(net4990),
     .fabric_out_09(net5036), .fabric_out_10(net5050),
     .rgt_op_02(net4883[0:7]), .slf_op_16(slf_op_00_16[3:0]),
     .slf_op_12(slf_op_00_12[3:0]), .sp4_v_t_16(sp4_v_t_00_16[15:0]),
     .reset_b(reset_l[271:16]), .slf_op_11(slf_op_00_11[3:0]),
     .slf_op_09(slf_op_00_09[3:0]), .slf_op_08(slf_op_00_08[3:0]),
     .slf_op_06(slf_op_00_06[3:0]), .slf_op_05(slf_op_00_05[3:0]),
     .SP12_h_l_01(net4893[0:23]), .slf_op_10(slf_op_00_10[3:0]),
     .slf_op_07(slf_op_00_07[3:0]), .slf_op_04(slf_op_00_04[3:0]),
     .wl(wl_l[271:16]), .SP4_h_l_06(net4898[0:47]),
     .SP4_h_l_07(net4899[0:47]), .SP4_h_l_04(net4900[0:47]),
     .SP4_h_l_05(net4901[0:47]), .SP4_h_l_02(net4902[0:47]),
     .SP4_h_l_03(net4903[0:47]), .rgt_op_14(net4904[0:7]),
     .rgt_op_15(net4905[0:7]), .rgt_op_16(slf_op_01_16[7:0]),
     .rgt_op_11(net4907[0:7]), .rgt_op_08(net4908[0:7]),
     .rgt_op_05(net4909[0:7]), .sp4_v_b_01(net4910[0:15]),
     .rgt_op_12(net4911[0:7]), .rgt_op_13(net4912[0:7]),
     .rgt_op_09(net4913[0:7]), .rgt_op_10(net4914[0:7]),
     .rgt_op_06(net4915[0:7]), .rgt_op_07(net4916[0:7]),
     .slf_op_02(slf_op_00_02[3:0]), .slf_op_03(slf_op_00_03[3:0]),
     .rgt_op_03(net4919[0:7]), .rgt_op_04(net4920[0:7]),
     .pgate(pgate_l[271:16]), .SP12_h_l_16(net4922[0:23]),
     .SP12_h_l_15(net4923[0:23]), .SP12_h_l_14(net4924[0:23]),
     .SP12_h_l_13(net4925[0:23]), .SP12_h_l_12(net4926[0:23]),
     .SP12_h_l_11(net4927[0:23]), .SP12_h_l_10(net4928[0:23]),
     .SP12_h_l_09(net4929[0:23]), .SP12_h_l_08(net4930[0:23]),
     .SP12_h_l_07(net4931[0:23]), .SP12_h_l_06(net4932[0:23]),
     .SP12_h_l_05(net4933[0:23]), .SP12_h_l_04(net4934[0:23]),
     .SP12_h_l_03(net4935[0:23]), .SP12_h_l_02(net4936[0:23]),
     .slf_op_01(slf_op_00_01[3:0]), .SP4_h_l_16(net4938[0:47]),
     .rgt_op_01(net4811[0:7]), .cdone_in(end_of_startup_lft_b[16:1]),
     .slf_op_13(slf_op_00_13[3:0]), .slf_op_14(slf_op_00_14[3:0]),
     .slf_op_15(slf_op_00_15[3:0]), .SP4_h_l_15(net4944[0:47]),
     .SP4_h_l_14(net4945[0:47]), .SP4_h_l_13(net4946[0:47]),
     .SP4_h_l_12(net4947[0:47]), .SP4_h_l_11(net4948[0:47]),
     .SP4_h_l_10(net4949[0:47]), .SP4_h_l_09(net4950[0:47]),
     .SP4_h_l_08(net4951[0:47]), .SP4_h_l_01(net4952[0:47]),
     .vdd_cntl(vdd_cntl_l[271:16]), .shift(net4954), .bs_en(net4980),
     .mode(net4956), .sdi(net2079), .hiz_b(net4958), .prog(prog),
     .hold(hold_l_b), .update(net4961),
     .glb_netwk_col(clk_tree_drv[7:0]), .r(net4976),
     .spi_ss_in_b(spi_ss_in_l[31:0]), .sdo(net4965), .bl({bl[0], bl[1],
     bl[2], bl[3], bl[4], bl[5], bl[6], bl[7], bl[8], bl[9], bl[10],
     bl[11], bl[12], bl[13], bl[14], bl[15], bl[16], bl[17]}),
     .tclk(net2076), .cf_l(cf_l[383:0]), .spioeb(spioeb_l[31:0]),
     .spiout(spiout_l[31:0]));
bram_bufferx4 I293 ( .in(ceb_i), .out(net4863));
bram_bufferx4 I244 ( .in(mode_i), .out(net4956));
bram_bufferx4 I249 ( .in(r_i), .out(net4976));
bram_bufferx4 I246 ( .in(shift_i), .out(net4954));
bram_bufferx4 I247 ( .in(bs_en_i), .out(net4980));
bram_bufferx4 I245 ( .in(update_i), .out(net4961));
bram_bufferx4 I250 ( .in(hiz_b_i), .out(net4958));

endmodule
// Library - leafcell, Cell - preio_bot_r, View - schematic
// LAST TIME SAVED: Oct 30 14:31:43 2008
// NETLIST TIME: Nov 14 16:17:17 2008
`timescale 1ns / 1ns 

module preio_bot_r ( cf_b, fabric_out_17_00, fabric_out_18_00,
     fabric_out_32_00, padeb_b, padin_81, pado_b, sdo_pad,
     slf_op_17_00, slf_op_18_00, slf_op_19_00, slf_op_20_00,
     slf_op_21_00, slf_op_22_00, slf_op_23_00, slf_op_24_00,
     slf_op_25_00, slf_op_26_00, slf_op_27_00, slf_op_28_00,
     slf_op_29_00, slf_op_30_00, slf_op_31_00, slf_op_32_00,
     spi_ss_in_b, bl_17, bl_18, bl_19, bl_20, bl_21, bl_22, bl_23,
     bl_24, bl_25, bl_26, bl_27, bl_28, bl_29, bl_30, bl_31, bl_32,
     sp4_h_l_17_00, sp4_h_r_32_00, sp4_v_t_17_00, sp4_v_t_18_00,
     sp4_v_t_19_00, sp4_v_t_20_00, sp4_v_t_21_00, sp4_v_t_22_00,
     sp4_v_t_23_00, sp4_v_t_24_00, sp4_v_t_25_00, sp4_v_t_26_00,
     sp4_v_t_27_00, sp4_v_t_28_00, sp4_v_t_29_00, sp4_v_t_30_00,
     sp4_v_t_31_00, sp4_v_t_32_00, sp12_v_t_17_00, sp12_v_t_18_00,
     sp12_v_t_19_00, sp12_v_t_20_00, sp12_v_t_21_00, sp12_v_t_22_00,
     sp12_v_t_23_00, sp12_v_t_24_00, sp12_v_t_25_00, sp12_v_t_26_00,
     sp12_v_t_27_00, sp12_v_t_28_00, sp12_v_t_29_00, sp12_v_t_30_00,
     sp12_v_t_31_00, sp12_v_t_32_00, bs_en_i, ceb_i,
     end_of_startup_bot_r, glb_net_17, glb_net_18, glb_net_19,
     glb_net_20, glb_net_21, glb_net_22, glb_net_23, glb_net_24,
     glb_net_25, glb_net_26, glb_net_27, glb_net_28, glb_net_29,
     glb_net_30, glb_net_31, glb_net_32, hiz_b_i, hold_b_r,
     lft_op_17_00, lft_op_18_00, lft_op_19_00, lft_op_20_00,
     lft_op_21_00, lft_op_22_00, lft_op_23_00, lft_op_24_00,
     lft_op_25_00, lft_op_26_00, lft_op_27_00, lft_op_28_00,
     lft_op_29_00, lft_op_30_00, lft_op_31_00, lft_op_32_00, mode_i,
     padin_b, pgate_r, prog, r_i, reset_r, sdi, shift_i, spioeb_b,
     spiout_b, tclk_i, tnl_op_17_00, tnr_op_32_00, update_i,
     vdd_cntl_r, wl_r );
output  fabric_out_17_00, fabric_out_18_00, fabric_out_32_00, padin_81,
     sdo_pad;


input  bs_en_i, ceb_i, hiz_b_i, hold_b_r, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, update_i;

output [3:0]  slf_op_27_00;
output [3:0]  slf_op_25_00;
output [3:0]  slf_op_21_00;
output [3:0]  slf_op_18_00;
output [3:0]  slf_op_28_00;
output [3:0]  slf_op_19_00;
output [3:0]  slf_op_23_00;
output [3:0]  slf_op_26_00;
output [3:0]  slf_op_31_00;
output [3:0]  slf_op_30_00;
output [3:0]  slf_op_22_00;
output [3:0]  slf_op_17_00;
output [383:0]  cf_b;
output [56:30]  pado_b;
output [63:32]  spi_ss_in_b;
output [3:0]  slf_op_32_00;
output [3:0]  slf_op_29_00;
output [3:0]  slf_op_24_00;
output [56:30]  padeb_b;
output [3:0]  slf_op_20_00;

inout [23:0]  sp12_v_t_30_00;
inout [47:0]  sp4_v_t_28_00;
inout [47:0]  sp4_v_t_27_00;
inout [15:0]  sp4_h_l_17_00;
inout [47:0]  sp4_v_t_26_00;
inout [15:0]  sp4_h_r_32_00;
inout [47:0]  sp4_v_t_22_00;
inout [23:0]  sp12_v_t_21_00;
inout [47:0]  sp4_v_t_30_00;
inout [23:0]  sp12_v_t_20_00;
inout [47:0]  sp4_v_t_20_00;
inout [23:0]  sp12_v_t_22_00;
inout [53:0]  bl_29;
inout [23:0]  sp12_v_t_19_00;
inout [47:0]  sp4_v_t_25_00;
inout [53:0]  bl_28;
inout [47:0]  sp4_v_t_24_00;
inout [47:0]  sp4_v_t_17_00;
inout [23:0]  sp12_v_t_28_00;
inout [47:0]  sp4_v_t_21_00;
inout [47:0]  sp4_v_t_29_00;
inout [23:0]  sp12_v_t_29_00;
inout [47:0]  sp4_v_t_31_00;
inout [47:0]  sp4_v_t_18_00;
inout [23:0]  sp12_v_t_23_00;
inout [23:0]  sp12_v_t_25_00;
inout [23:0]  sp12_v_t_24_00;
inout [23:0]  sp12_v_t_18_00;
inout [23:0]  sp12_v_t_31_00;
inout [47:0]  sp4_v_t_19_00;
inout [23:0]  sp12_v_t_27_00;
inout [53:0]  bl_26;
inout [53:0]  bl_27;
inout [53:0]  bl_18;
inout [53:0]  bl_31;
inout [53:0]  bl_30;
inout [53:0]  bl_17;
inout [53:0]  bl_32;
inout [53:0]  bl_24;
inout [47:0]  sp4_v_t_32_00;
inout [53:0]  bl_23;
inout [41:0]  bl_25;
inout [47:0]  sp4_v_t_23_00;
inout [53:0]  bl_19;
inout [23:0]  sp12_v_t_32_00;
inout [23:0]  sp12_v_t_26_00;
inout [23:0]  sp12_v_t_17_00;
inout [53:0]  bl_20;
inout [53:0]  bl_21;
inout [53:0]  bl_22;

input [7:0]  glb_net_26;
input [7:0]  glb_net_17;
input [7:0]  glb_net_23;
input [7:0]  lft_op_18_00;
input [7:0]  glb_net_24;
input [7:0]  glb_net_28;
input [7:0]  lft_op_25_00;
input [7:0]  glb_net_19;
input [7:0]  glb_net_18;
input [7:0]  glb_net_22;
input [7:0]  glb_net_20;
input [7:0]  glb_net_27;
input [7:0]  glb_net_21;
input [7:0]  glb_net_25;
input [15:0]  reset_r;
input [7:0]  lft_op_26_00;
input [7:0]  glb_net_29;
input [15:0]  wl_r;
input [7:0]  lft_op_30_00;
input [7:0]  lft_op_20_00;
input [7:0]  lft_op_28_00;
input [7:0]  tnr_op_32_00;
input [7:0]  lft_op_29_00;
input [7:0]  lft_op_17_00;
input [7:0]  lft_op_21_00;
input [7:0]  lft_op_31_00;
input [7:0]  lft_op_19_00;
input [7:0]  glb_net_30;
input [56:30]  padin_b;
input [7:0]  lft_op_32_00;
input [15:0]  vdd_cntl_r;
input [7:0]  lft_op_22_00;
input [15:0]  pgate_r;
input [7:0]  lft_op_27_00;
input [63:32]  spioeb_b;
input [7:0]  glb_net_31;
input [7:0]  lft_op_24_00;
input [63:32]  spiout_b;
input [7:0]  lft_op_23_00;
input [7:0]  tnl_op_17_00;
input [7:0]  glb_net_32;
input [31:16]  end_of_startup_bot_r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net1206;

wire  [0:15]  net1036;

wire  [0:1]  net710;

wire  [0:15]  net696;

wire  [0:15]  net1070;

wire  [0:1]  net846;

wire  [0:15]  net934;

wire  [0:15]  net832;

wire  [0:1]  net1241;

wire  [0:1]  net1254;

wire  [0:15]  net764;

wire  [0:15]  net1138;

wire  [0:15]  net968;

wire  [0:15]  net1172;

wire  [0:15]  net1002;

wire  [0:15]  net1104;

wire  [0:15]  net730;

wire  [0:15]  net798;

wire  [0:15]  net893;



tckbufx16 I888 ( .in(tclk_i), .out(endtck));
lowla_modified I292 ( .clk(endtck), .min(net0677), .lao(sdo_pad));
lowla_modified I293 ( .clk(tclk_i), .min(net0681), .lao(net1224));
bram_bufferx4x6 I294 ( .in(net0866), .out(net0677));
bram_bufferx4x6 I295 ( .in(sdi), .out(net0681));
fabric_buf8k I287 ( .f_in(padin_b[30]), .f_out(padin_81));
fabric_buf8k I290 ( .f_in(net1207), .f_out(fabric_out_32_00));
fabric_buf8k I288 ( .f_in(net1209), .f_out(fabric_out_17_00));
fabric_buf8k I289 ( .f_in(net1217), .f_out(fabric_out_18_00));
io_col4_BRAM_BOT I_IO_25_00bram ( .ceb(net01234), .bl({bl_25[5],
     bl_25[4], bl_25[37], bl_25[36], bl_25[35], bl_25[34], bl_25[33],
     bl_25[32], bl_25[14], bl_25[20], bl_25[19], bl_25[18], bl_25[17],
     bl_25[16], bl_25[27], bl_25[26], bl_25[25], bl_25[23]}),
     .sdo(net664), .sdi(net868), .spiout(spiout_b[49:48]),
     .cdone_in(end_of_startup_bot_r[24]), .spioeb(spioeb_b[49:48]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[45:44]), .pado(pado_b[45:44]),
     .padeb(padeb_b[45:44]), .sp4_h_l(sp4_v_t_25_00[47:0]),
     .sp12_h_l(sp12_v_t_25_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[49:48]), .tnl_op(lft_op_24_00[7:0]),
     .lft_op(lft_op_25_00[7:0]), .bnl_op(lft_op_26_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[215:192]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_25_00[3:0]), .glb_netwk(glb_net_25[7:0]),
     .hold(hold_b_r), .fabric_out(net1246), .sp4_v_t(net893[0:15]),
     .sp4_v_b(net696[0:15]));
io_col4_BOT I_IO_18_00 ( .ceb(net01234), .bl({bl_18[5], bl_18[4],
     bl_18[37], bl_18[36], bl_18[35], bl_18[34], bl_18[33], bl_18[32],
     bl_18[14], bl_18[20], bl_18[19], bl_18[18], bl_18[17], bl_18[16],
     bl_18[27], bl_18[26], bl_18[25], bl_18[23]}), .sdo(net698),
     .sdi(net766), .spiout(spiout_b[35:34]),
     .cdone_in(end_of_startup_bot_r[17]), .spioeb(spioeb_b[35:34]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(net710[0:1]), .pado(net710[0:1]), .padeb(net1254[0:1]),
     .sp4_h_l(sp4_v_t_18_00[47:0]), .sp12_h_l(sp12_v_t_18_00[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[35:34]),
     .tnl_op(lft_op_17_00[7:0]), .lft_op(lft_op_18_00[7:0]),
     .bnl_op(lft_op_19_00[7:0]), .pgate(pgate_r[15:0]),
     .reset(reset_r[15:0]), .wl(wl_r[15:0]), .cf(cf_b[47:24]),
     .vdd_cntl(vdd_cntl_r[15:0]), .slf_op(slf_op_18_00[3:0]),
     .glb_netwk(glb_net_18[7:0]), .hold(hold_b_r),
     .fabric_out(net1217), .sp4_v_t(net798[0:15]),
     .sp4_v_b(net730[0:15]));
io_col4_BOT I_IO_28_00 ( .ceb(net01234), .bl({bl_28[5], bl_28[4],
     bl_28[37], bl_28[36], bl_28[35], bl_28[34], bl_28[33], bl_28[32],
     bl_28[14], bl_28[20], bl_28[19], bl_28[18], bl_28[17], bl_28[16],
     bl_28[27], bl_28[26], bl_28[25], bl_28[23]}), .sdo(net732),
     .sdi(net800), .spiout(spiout_b[55:54]),
     .cdone_in(end_of_startup_bot_r[27]), .spioeb(spioeb_b[55:54]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238), .padin({n_short,
     padin_b[50]}), .pado({n_short, pado_b[50]}), .padeb({n_idle,
     padeb_b[50]}), .sp4_h_l(sp4_v_t_28_00[47:0]),
     .sp12_h_l(sp12_v_t_28_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[55:54]), .tnl_op(lft_op_27_00[7:0]),
     .lft_op(lft_op_28_00[7:0]), .bnl_op(lft_op_29_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[287:264]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_28_00[3:0]), .glb_netwk(glb_net_28[7:0]),
     .hold(hold_b_r), .fabric_out(net1250), .sp4_v_t(net832[0:15]),
     .sp4_v_b(net764[0:15]));
io_col4_BOT I_IO_17_00 ( .ceb(net01234), .bl({bl_17[5], bl_17[4],
     bl_17[37], bl_17[36], bl_17[35], bl_17[34], bl_17[33], bl_17[32],
     bl_17[14], bl_17[20], bl_17[19], bl_17[18], bl_17[17], bl_17[16],
     bl_17[27], bl_17[26], bl_17[25], bl_17[23]}), .sdo(net766),
     .sdi(net1224), .spiout(spiout_b[33:32]),
     .cdone_in(end_of_startup_bot_r[16]), .spioeb(spioeb_b[33:32]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[31:30]), .pado(pado_b[31:30]),
     .padeb(padeb_b[31:30]), .sp4_h_l(sp4_v_t_17_00[47:0]),
     .sp12_h_l(sp12_v_t_17_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[33:32]), .tnl_op(tnl_op_17_00[7:0]),
     .lft_op(lft_op_17_00[7:0]), .bnl_op(lft_op_18_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[23:0]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_17_00[3:0]), .glb_netwk(glb_net_17[7:0]),
     .hold(hold_b_r), .fabric_out(net1209),
     .sp4_v_t(sp4_h_l_17_00[15:0]), .sp4_v_b(net798[0:15]));
io_col4_BOT I_IO_27_00 ( .ceb(net01234), .bl({bl_27[5], bl_27[4],
     bl_27[37], bl_27[36], bl_27[35], bl_27[34], bl_27[33], bl_27[32],
     bl_27[14], bl_27[20], bl_27[19], bl_27[18], bl_27[17], bl_27[16],
     bl_27[27], bl_27[26], bl_27[25], bl_27[23]}), .sdo(net800),
     .sdi(net1174), .spiout(spiout_b[53:52]),
     .cdone_in(end_of_startup_bot_r[26]), .spioeb(spioeb_b[53:52]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[49:48]), .pado(pado_b[49:48]),
     .padeb(padeb_b[49:48]), .sp4_h_l(sp4_v_t_27_00[47:0]),
     .sp12_h_l(sp12_v_t_27_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[53:52]), .tnl_op(lft_op_26_00[7:0]),
     .lft_op(lft_op_27_00[7:0]), .bnl_op(lft_op_28_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[263:240]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_27_00[3:0]), .glb_netwk(glb_net_27[7:0]),
     .hold(hold_b_r), .fabric_out(net1243), .sp4_v_t(net1206[0:15]),
     .sp4_v_b(net832[0:15]));
io_col4_BOT I_IO_32_00 ( .ceb(net01234), .bl({bl_32[5], bl_32[4],
     bl_32[37], bl_32[36], bl_32[35], bl_32[34], bl_32[33], bl_32[32],
     bl_32[14], bl_32[20], bl_32[19], bl_32[18], bl_32[17], bl_32[16],
     bl_32[27], bl_32[26], bl_32[25], bl_32[23]}), .sdo(net0866),
     .sdi(net1106), .spiout(spiout_b[63:62]),
     .cdone_in(end_of_startup_bot_r[31]), .spioeb(spioeb_b[63:62]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(net846[0:1]), .pado(net846[0:1]), .padeb(net1241[0:1]),
     .sp4_h_l(sp4_v_t_32_00[47:0]), .sp12_h_l(sp12_v_t_32_00[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[63:62]),
     .tnl_op(lft_op_31_00[7:0]), .lft_op(lft_op_32_00[7:0]),
     .bnl_op(tnr_op_32_00[7:0]), .pgate(pgate_r[15:0]),
     .reset(reset_r[15:0]), .wl(wl_r[15:0]), .cf(cf_b[383:360]),
     .vdd_cntl(vdd_cntl_r[15:0]), .slf_op(slf_op_32_00[3:0]),
     .glb_netwk(glb_net_32[7:0]), .hold(hold_b_r), .fabric_out(net864),
     .sp4_v_t(net1138[0:15]), .sp4_v_b(sp4_h_r_32_00[15:0]));
io_col4_BOT I_IO_24_00 ( .ceb(net01234), .bl({bl_24[5], bl_24[4],
     bl_24[37], bl_24[36], bl_24[35], bl_24[34], bl_24[33], bl_24[32],
     bl_24[14], bl_24[20], bl_24[19], bl_24[18], bl_24[17], bl_24[16],
     bl_24[27], bl_24[26], bl_24[25], bl_24[23]}), .sdo(net868),
     .sdi(net936), .spiout(spiout_b[47:46]),
     .cdone_in(end_of_startup_bot_r[23]), .spioeb(spioeb_b[47:46]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[43:42]), .pado(pado_b[43:42]),
     .padeb(padeb_b[43:42]), .sp4_v_t(net968[0:15]),
     .sp4_h_l(sp4_v_t_24_00[47:0]), .sp12_h_l(sp12_v_t_24_00[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[47:46]),
     .tnl_op(lft_op_23_00[7:0]), .lft_op(lft_op_24_00[7:0]),
     .bnl_op(lft_op_25_00[7:0]), .pgate(pgate_r[15:0]),
     .reset(reset_r[15:0]), .sp4_v_b(net893[0:15]), .wl(wl_r[15:0]),
     .cf(cf_b[191:168]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_24_00[3:0]), .glb_netwk(glb_net_24[7:0]),
     .hold(hold_b_r), .fabric_out(net1252));
io_col4_BOT I_IO_21_00 ( .ceb(net01234), .bl({bl_21[5], bl_21[4],
     bl_21[37], bl_21[36], bl_21[35], bl_21[34], bl_21[33], bl_21[32],
     bl_21[14], bl_21[20], bl_21[19], bl_21[18], bl_21[17], bl_21[16],
     bl_21[27], bl_21[26], bl_21[25], bl_21[23]}), .sdo(net902),
     .sdi(net1140), .spiout(spiout_b[41:40]),
     .cdone_in(end_of_startup_bot_r[20]), .spioeb(spioeb_b[41:40]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[37:36]), .pado(pado_b[37:36]),
     .padeb(padeb_b[37:36]), .sp4_h_l(sp4_v_t_21_00[47:0]),
     .sp12_h_l(sp12_v_t_21_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[41:40]), .tnl_op(lft_op_20_00[7:0]),
     .lft_op(lft_op_21_00[7:0]), .bnl_op(lft_op_22_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[119:96]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_21_00[3:0]), .glb_netwk(glb_net_21[7:0]),
     .hold(hold_b_r), .fabric_out(net932), .sp4_v_t(net1172[0:15]),
     .sp4_v_b(net934[0:15]));
io_col4_BOT I_IO_23_00 ( .ceb(net01234), .bl({bl_23[5], bl_23[4],
     bl_23[37], bl_23[36], bl_23[35], bl_23[34], bl_23[33], bl_23[32],
     bl_23[14], bl_23[20], bl_23[19], bl_23[18], bl_23[17], bl_23[16],
     bl_23[27], bl_23[26], bl_23[25], bl_23[23]}), .sdo(net936),
     .sdi(net970), .spiout(spiout_b[45:44]),
     .cdone_in(end_of_startup_bot_r[22]), .spioeb(spioeb_b[45:44]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[41:40]), .pado(pado_b[41:40]),
     .padeb(padeb_b[41:40]), .sp4_h_l(sp4_v_t_23_00[47:0]),
     .sp12_h_l(sp12_v_t_23_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[45:44]), .tnl_op(lft_op_22_00[7:0]),
     .lft_op(lft_op_23_00[7:0]), .bnl_op(lft_op_24_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[167:144]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_23_00[3:0]), .glb_netwk(glb_net_23[7:0]),
     .hold(hold_b_r), .fabric_out(net966), .sp4_v_t(net1002[0:15]),
     .sp4_v_b(net968[0:15]));
io_col4_BOT I_IO_22_00 ( .ceb(net01234), .bl({bl_22[5], bl_22[4],
     bl_22[37], bl_22[36], bl_22[35], bl_22[34], bl_22[33], bl_22[32],
     bl_22[14], bl_22[20], bl_22[19], bl_22[18], bl_22[17], bl_22[16],
     bl_22[27], bl_22[26], bl_22[25], bl_22[23]}), .sdo(net970),
     .sdi(net902), .spiout(spiout_b[43:42]),
     .cdone_in(end_of_startup_bot_r[21]), .spioeb(spioeb_b[43:42]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[39:38]), .pado(pado_b[39:38]),
     .padeb(padeb_b[39:38]), .sp4_h_l(sp4_v_t_22_00[47:0]),
     .sp12_h_l(sp12_v_t_22_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[43:42]), .tnl_op(lft_op_21_00[7:0]),
     .lft_op(lft_op_22_00[7:0]), .bnl_op(lft_op_23_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[143:120]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_22_00[3:0]), .glb_netwk(glb_net_22[7:0]),
     .hold(hold_b_r), .fabric_out(net1000), .sp4_v_t(net934[0:15]),
     .sp4_v_b(net1002[0:15]));
io_col4_BOT I_IO_19_00 ( .ceb(net01234), .bl({bl_19[5], bl_19[4],
     bl_19[37], bl_19[36], bl_19[35], bl_19[34], bl_19[33], bl_19[32],
     bl_19[14], bl_19[20], bl_19[19], bl_19[18], bl_19[17], bl_19[16],
     bl_19[27], bl_19[26], bl_19[25], bl_19[23]}), .sdo(net1004),
     .sdi(net698), .spiout(spiout_b[37:36]),
     .cdone_in(end_of_startup_bot_r[18]), .spioeb(spioeb_b[37:36]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[33:32]), .pado(pado_b[33:32]),
     .padeb(padeb_b[33:32]), .sp4_h_l(sp4_v_t_19_00[47:0]),
     .sp12_h_l(sp12_v_t_19_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[37:36]), .tnl_op(lft_op_18_00[7:0]),
     .lft_op(lft_op_19_00[7:0]), .bnl_op(lft_op_20_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[71:48]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_19_00[3:0]), .glb_netwk(glb_net_19[7:0]),
     .hold(hold_b_r), .fabric_out(net1034), .sp4_v_t(net730[0:15]),
     .sp4_v_b(net1036[0:15]));
io_col4_BOT I_IO_30_00 ( .ceb(net01234), .bl({bl_30[5], bl_30[4],
     bl_30[37], bl_30[36], bl_30[35], bl_30[34], bl_30[33], bl_30[32],
     bl_30[14], bl_30[20], bl_30[19], bl_30[18], bl_30[17], bl_30[16],
     bl_30[27], bl_30[26], bl_30[25], bl_30[23]}), .sdo(net1038),
     .sdi(net1072), .spiout(spiout_b[59:58]),
     .cdone_in(end_of_startup_bot_r[29]), .spioeb(spioeb_b[59:58]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[54:53]), .pado(pado_b[54:53]),
     .padeb(padeb_b[54:53]), .sp4_h_l(sp4_v_t_30_00[47:0]),
     .sp12_h_l(sp12_v_t_30_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[59:58]), .tnl_op(lft_op_29_00[7:0]),
     .lft_op(lft_op_30_00[7:0]), .bnl_op(lft_op_31_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[335:312]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_30_00[3:0]), .glb_netwk(glb_net_30[7:0]),
     .hold(hold_b_r), .fabric_out(net1251), .sp4_v_t(net1104[0:15]),
     .sp4_v_b(net1070[0:15]));
io_col4_BOT I_IO_29_00 ( .ceb(net01234), .bl({bl_29[5], bl_29[4],
     bl_29[37], bl_29[36], bl_29[35], bl_29[34], bl_29[33], bl_29[32],
     bl_29[14], bl_29[20], bl_29[19], bl_29[18], bl_29[17], bl_29[16],
     bl_29[27], bl_29[26], bl_29[25], bl_29[23]}), .sdo(net1072),
     .sdi(net732), .spiout(spiout_b[57:56]),
     .cdone_in(end_of_startup_bot_r[28]), .spioeb(spioeb_b[57:56]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[52:51]), .pado(pado_b[52:51]),
     .padeb(padeb_b[52:51]), .sp4_h_l(sp4_v_t_29_00[47:0]),
     .sp12_h_l(sp12_v_t_29_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[57:56]), .tnl_op(lft_op_28_00[7:0]),
     .lft_op(lft_op_29_00[7:0]), .bnl_op(lft_op_30_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[311:288]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_29_00[3:0]), .glb_netwk(glb_net_29[7:0]),
     .hold(hold_b_r), .fabric_out(net1253), .sp4_v_t(net764[0:15]),
     .sp4_v_b(net1104[0:15]));
io_col4_BOT I_IO_31_00 ( .ceb(net01234), .bl({bl_31[5], bl_31[4],
     bl_31[37], bl_31[36], bl_31[35], bl_31[34], bl_31[33], bl_31[32],
     bl_31[14], bl_31[20], bl_31[19], bl_31[18], bl_31[17], bl_31[16],
     bl_31[27], bl_31[26], bl_31[25], bl_31[23]}), .sdo(net1106),
     .sdi(net1038), .spiout(spiout_b[61:60]),
     .cdone_in(end_of_startup_bot_r[30]), .spioeb(spioeb_b[61:60]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[56:55]), .pado(pado_b[56:55]),
     .padeb(padeb_b[56:55]), .sp4_h_l(sp4_v_t_31_00[47:0]),
     .sp12_h_l(sp12_v_t_31_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[61:60]), .tnl_op(lft_op_30_00[7:0]),
     .lft_op(lft_op_31_00[7:0]), .bnl_op(lft_op_32_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[359:336]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_31_00[3:0]), .glb_netwk(glb_net_31[7:0]),
     .hold(hold_b_r), .fabric_out(net1207), .sp4_v_t(net1070[0:15]),
     .sp4_v_b(net1138[0:15]));
io_col4_BOT I_IO_20_00 ( .ceb(net01234), .bl({bl_20[5], bl_20[4],
     bl_20[37], bl_20[36], bl_20[35], bl_20[34], bl_20[33], bl_20[32],
     bl_20[14], bl_20[20], bl_20[19], bl_20[18], bl_20[17], bl_20[16],
     bl_20[27], bl_20[26], bl_20[25], bl_20[23]}), .sdo(net1140),
     .sdi(net1004), .spiout(spiout_b[39:38]),
     .cdone_in(end_of_startup_bot_r[19]), .spioeb(spioeb_b[39:38]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[35:34]), .pado(pado_b[35:34]),
     .padeb(padeb_b[35:34]), .sp4_h_l(sp4_v_t_20_00[47:0]),
     .sp12_h_l(sp12_v_t_20_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[39:38]), .tnl_op(lft_op_19_00[7:0]),
     .lft_op(lft_op_20_00[7:0]), .bnl_op(lft_op_21_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[95:72]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_20_00[3:0]), .glb_netwk(glb_net_20[7:0]),
     .hold(hold_b_r), .fabric_out(net1170), .sp4_v_t(net1036[0:15]),
     .sp4_v_b(net1172[0:15]));
io_col4_BOT I_IO_26_00 ( .ceb(net01234), .bl({bl_26[5], bl_26[4],
     bl_26[37], bl_26[36], bl_26[35], bl_26[34], bl_26[33], bl_26[32],
     bl_26[14], bl_26[20], bl_26[19], bl_26[18], bl_26[17], bl_26[16],
     bl_26[27], bl_26[26], bl_26[25], bl_26[23]}), .sdo(net1174),
     .sdi(net664), .spiout(spiout_b[51:50]),
     .cdone_in(end_of_startup_bot_r[25]), .spioeb(spioeb_b[51:50]),
     .mode(net1232), .shift(net1230), .hiz_b(net1236), .r(net1226),
     .bs_en(net1228), .tclk(endtck), .update(net1238),
     .padin(padin_b[47:46]), .pado(pado_b[47:46]),
     .padeb(padeb_b[47:46]), .sp4_h_l(sp4_v_t_26_00[47:0]),
     .sp12_h_l(sp12_v_t_26_00[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[51:50]), .tnl_op(lft_op_25_00[7:0]),
     .lft_op(lft_op_26_00[7:0]), .bnl_op(lft_op_27_00[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_b[239:216]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_26_00[3:0]), .glb_netwk(glb_net_26[7:0]),
     .hold(hold_b_r), .fabric_out(net1249), .sp4_v_t(net696[0:15]),
     .sp4_v_b(net1206[0:15]));
bram_bufferx4 I291 ( .in(ceb_i), .out(net01234));
bram_bufferx4 I892 ( .in(r_i), .out(net1226));
bram_bufferx4 I893 ( .in(bs_en_i), .out(net1228));
bram_bufferx4 I890 ( .in(shift_i), .out(net1230));
bram_bufferx4 I887 ( .in(mode_i), .out(net1232));
bram_bufferx4 I891 ( .in(hiz_b_i), .out(net1236));
bram_bufferx4 I889 ( .in(update_i), .out(net1238));

endmodule
// Library - io, Cell - io_col4_RGT, View - schematic
// LAST TIME SAVED: Feb  5 08:40:49 2008
// NETLIST TIME: Nov 14 16:17:17 2008
`timescale 1ns / 1ns 

module io_col4_RGT ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  pado;
output [23:0]  cf;
output [1:0]  padeb;
output [3:0]  slf_op;
output [1:0]  spi_ss_in_b;

inout [17:0]  bl;
inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_t;

input [1:0]  spioeb;
input [1:0]  spiout;
input [15:0]  pgate;
input [15:0]  vdd_cntl;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [1:0]  padin;
input [7:0]  lft_op;
input [15:0]  reset;
input [15:0]  wl;
input [7:0]  glb_netwk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net262));
rm7  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm7  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm7  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm7  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm7  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm7  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm7  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm7  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm7  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm7  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm7  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm7  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm7  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm7  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm7  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm7  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net262, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(net262),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net262));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net262), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));

endmodule
// Library - leafcell, Cell - array_RGT_IO_1x16, View - schematic
// LAST TIME SAVED: Jan 31 11:19:46 2008
// NETLIST TIME: Nov 14 16:17:17 2008
`timescale 1ns / 1ns 

module array_RGT_IO_1x16 ( cf_r, fabric_out_01, fabric_out_02,
     fabric_out_03, fabric_out_04, fabric_out_05, fabric_out_06,
     fabric_out_07, fabric_out_08, fabric_out_09, fabric_out_10,
     fabric_out_11, fabric_out_12, fabric_out_13, fabric_out_14,
     fabric_out_15, fabric_out_16, padeb, pado, sdo, slf_op_01,
     slf_op_02, slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07,
     slf_op_08, slf_op_09, slf_op_10, slf_op_11, slf_op_12, slf_op_13,
     slf_op_14, slf_op_15, slf_op_16, spi_ss_in_b, SP4_h_l_01,
     SP4_h_l_02, SP4_h_l_03, SP4_h_l_04, SP4_h_l_05, SP4_h_l_06,
     SP4_h_l_07, SP4_h_l_08, SP4_h_l_09, SP4_h_l_10, SP4_h_l_11,
     SP4_h_l_12, SP4_h_l_13, SP4_h_l_14, SP4_h_l_15, SP4_h_l_16,
     SP12_h_l_01, SP12_h_l_02, SP12_h_l_03, SP12_h_l_04, SP12_h_l_05,
     SP12_h_l_06, SP12_h_l_07, SP12_h_l_08, SP12_h_l_09, SP12_h_l_10,
     SP12_h_l_11, SP12_h_l_12, SP12_h_l_13, SP12_h_l_14, SP12_h_l_15,
     SP12_h_l_16, bl, pgate, reset_b, sp4_v_b_01, sp4_v_t_16, vdd_cntl,
     wl, bnl_op_01, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     lft_op_01, lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06,
     lft_op_07, lft_op_08, lft_op_09, lft_op_10, lft_op_11, lft_op_12,
     lft_op_13, lft_op_14, lft_op_15, lft_op_16, mode, padin, prog, r,
     sdi, shift, spioeb, spiout, tclk, tnl_op_16, update );
output  fabric_out_01, fabric_out_02, fabric_out_03, fabric_out_04,
     fabric_out_05, fabric_out_06, fabric_out_07, fabric_out_08,
     fabric_out_09, fabric_out_10, fabric_out_11, fabric_out_12,
     fabric_out_13, fabric_out_14, fabric_out_15, fabric_out_16, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_15;
output [3:0]  slf_op_04;
output [3:0]  slf_op_02;
output [3:0]  slf_op_12;
output [3:0]  slf_op_03;
output [3:0]  slf_op_07;
output [3:0]  slf_op_05;
output [3:0]  slf_op_14;
output [3:0]  slf_op_06;
output [3:0]  slf_op_11;
output [3:0]  slf_op_13;
output [3:0]  slf_op_09;
output [31:0]  spi_ss_in_b;
output [3:0]  slf_op_10;
output [3:0]  slf_op_16;
output [3:0]  slf_op_01;
output [27:0]  padeb;
output [383:0]  cf_r;
output [27:0]  pado;
output [3:0]  slf_op_08;

inout [23:0]  SP12_h_l_12;
inout [23:0]  SP12_h_l_05;
inout [47:0]  SP4_h_l_07;
inout [47:0]  SP4_h_l_12;
inout [23:0]  SP12_h_l_08;
inout [23:0]  SP12_h_l_02;
inout [23:0]  SP12_h_l_16;
inout [23:0]  SP12_h_l_07;
inout [47:0]  SP4_h_l_06;
inout [23:0]  SP12_h_l_03;
inout [47:0]  SP4_h_l_01;
inout [15:0]  sp4_v_b_01;
inout [23:0]  SP12_h_l_15;
inout [47:0]  SP4_h_l_05;
inout [15:0]  sp4_v_t_16;
inout [23:0]  SP12_h_l_11;
inout [47:0]  SP4_h_l_10;
inout [23:0]  SP12_h_l_13;
inout [47:0]  SP4_h_l_14;
inout [47:0]  SP4_h_l_16;
inout [47:0]  SP4_h_l_04;
inout [47:0]  SP4_h_l_09;
inout [47:0]  SP4_h_l_15;
inout [23:0]  SP12_h_l_09;
inout [47:0]  SP4_h_l_08;
inout [47:0]  SP4_h_l_03;
inout [23:0]  SP12_h_l_01;
inout [23:0]  SP12_h_l_04;
inout [47:0]  SP4_h_l_11;
inout [17:0]  bl;
inout [47:0]  SP4_h_l_13;
inout [255:0]  pgate;
inout [23:0]  SP12_h_l_10;
inout [255:0]  vdd_cntl;
inout [255:0]  reset_b;
inout [47:0]  SP4_h_l_02;
inout [23:0]  SP12_h_l_14;
inout [255:0]  wl;
inout [23:0]  SP12_h_l_06;

input [7:0]  glb_netwk_col;
input [7:0]  bnl_op_01;
input [7:0]  lft_op_16;
input [7:0]  lft_op_05;
input [7:0]  lft_op_15;
input [7:0]  lft_op_06;
input [7:0]  lft_op_02;
input [7:0]  lft_op_10;
input [7:0]  lft_op_01;
input [7:0]  lft_op_12;
input [7:0]  lft_op_14;
input [7:0]  lft_op_13;
input [7:0]  lft_op_11;
input [7:0]  lft_op_08;
input [7:0]  lft_op_03;
input [7:0]  lft_op_07;
input [7:0]  lft_op_04;
input [7:0]  tnl_op_16;
input [27:0]  padin;
input [7:0]  lft_op_09;
input [31:0]  spiout;
input [15:0]  cdone_in;
input [31:0]  spioeb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net1138;

wire  [0:15]  net798;

wire  [0:15]  net764;

wire  [0:1]  net1035;

wire  [0:15]  net1172;

wire  [0:1]  net1034;

wire  [0:15]  net832;

wire  [0:15]  net1002;

wire  [0:1]  net1001;

wire  [0:15]  net730;

wire  [0:1]  net1000;

wire  [0:15]  net934;

wire  [0:15]  net696;

wire  [0:15]  net1036;

wire  [0:15]  net662;

wire  [0:15]  net1070;

wire  [7:0]  glb_netwk;

wire  [0:15]  net1104;

wire  [0:15]  net866;

wire  [0:15]  net968;



clk_colbuf8kx8 I105 ( .clko(glb_netwk[7:0]),
     .clki(glb_netwk_col[7:0]));
io_col4_RGT I_io_00_09 ( .ceb(ceb), .sdo(net647), .sdi(net681),
     .spiout(spiout[17:16]), .cdone_in(cdone_in[8]),
     .spioeb(spioeb[17:16]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[13:12]), .pado(pado[13:12]), .padeb(padeb[13:12]),
     .sp4_v_t(net662[0:15]), .spi_ss_in_b(spi_ss_in_b[17:16]),
     .reset(reset_b[143:128]), .sp4_v_b(net696[0:15]),
     .cf(cf_r[215:192]), .bl(bl[17:0]), .slf_op(slf_op_09[3:0]),
     .hold(hold), .fabric_out(fabric_out_09), .prog(prog),
     .lft_op(lft_op_09[7:0]), .sp12_h_l(SP12_h_l_09[23:0]),
     .sp4_h_l(SP4_h_l_09[47:0]), .wl(wl[143:128]),
     .vdd_cntl(vdd_cntl[143:128]), .glb_netwk(glb_netwk[7:0]),
     .pgate(pgate[143:128]), .bnl_op(lft_op_08[7:0]),
     .tnl_op(lft_op_10[7:0]));
io_col4_RGT I_io_00_08 ( .ceb(ceb), .sdo(net681), .sdi(net715),
     .spiout(spiout[15:14]), .cdone_in(cdone_in[7]),
     .spioeb(spioeb[15:14]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[11:10]), .pado(pado[11:10]), .padeb(padeb[11:10]),
     .sp4_v_t(net696[0:15]), .sp4_h_l(SP4_h_l_08[47:0]),
     .sp12_h_l(SP12_h_l_08[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[15:14]), .tnl_op(lft_op_09[7:0]),
     .lft_op(lft_op_08[7:0]), .bnl_op(lft_op_07[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net730[0:15]), .wl(wl[127:112]), .cf(cf_r[191:168]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_08[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_08));
io_col4_RGT I_io_00_07 ( .ceb(ceb), .sdo(net715), .sdi(net953),
     .spiout(spiout[13:12]), .cdone_in(cdone_in[6]),
     .spioeb(spioeb[13:12]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[9:8]), .pado(pado[9:8]), .padeb(padeb[9:8]),
     .sp4_v_t(net730[0:15]), .sp4_h_l(SP4_h_l_07[47:0]),
     .sp12_h_l(SP12_h_l_07[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[13:12]), .tnl_op(lft_op_08[7:0]),
     .lft_op(lft_op_07[7:0]), .bnl_op(lft_op_06[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net968[0:15]), .wl(wl[111:96]), .cf(cf_r[167:144]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_07[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_07));
io_col4_RGT I_io_00_15 ( .ceb(ceb), .sdo(net749), .sdi(net783),
     .spiout(spiout[29:28]), .cdone_in(cdone_in[14]),
     .spioeb(spioeb[29:28]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[25:24]), .pado(pado[25:24]), .padeb(padeb[25:24]),
     .sp4_v_t(net764[0:15]), .sp4_h_l(SP4_h_l_15[47:0]),
     .sp12_h_l(SP12_h_l_15[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[29:28]), .tnl_op(lft_op_16[7:0]),
     .lft_op(lft_op_15[7:0]), .bnl_op(lft_op_14[7:0]),
     .pgate(pgate[239:224]), .reset(reset_b[239:224]),
     .sp4_v_b(net798[0:15]), .wl(wl[239:224]), .cf(cf_r[359:336]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[239:224]),
     .slf_op(slf_op_15[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_15));
io_col4_RGT I_io_00_14 ( .ceb(ceb), .sdo(net783), .sdi(net817),
     .spiout(spiout[27:26]), .cdone_in(cdone_in[13]),
     .spioeb(spioeb[27:26]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[23:22]), .pado(pado[23:22]), .padeb(padeb[23:22]),
     .sp4_v_t(net798[0:15]), .sp4_h_l(SP4_h_l_14[47:0]),
     .sp12_h_l(SP12_h_l_14[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[27:26]), .tnl_op(lft_op_15[7:0]),
     .lft_op(lft_op_14[7:0]), .bnl_op(lft_op_13[7:0]),
     .pgate(pgate[223:208]), .reset(reset_b[223:208]),
     .sp4_v_b(net832[0:15]), .wl(wl[223:208]), .cf(cf_r[335:312]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[223:208]),
     .slf_op(slf_op_14[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_14));
io_col4_RGT I_io_00_13 ( .ceb(ceb), .sdo(net817), .sdi(net851),
     .spiout(spiout[25:24]), .cdone_in(cdone_in[12]),
     .spioeb(spioeb[25:24]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[21:20]), .pado(pado[21:20]), .padeb(padeb[21:20]),
     .sp4_v_t(net832[0:15]), .sp4_h_l(SP4_h_l_13[47:0]),
     .sp12_h_l(SP12_h_l_13[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[25:24]), .tnl_op(lft_op_14[7:0]),
     .lft_op(lft_op_13[7:0]), .bnl_op(lft_op_12[7:0]),
     .pgate(pgate[207:192]), .reset(reset_b[207:192]),
     .sp4_v_b(net866[0:15]), .wl(wl[207:192]), .cf(cf_r[311:288]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[207:192]),
     .slf_op(slf_op_13[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_13));
io_col4_RGT I_io_00_12 ( .ceb(ceb), .sdo(net851), .sdi(net1157),
     .spiout(spiout[23:22]), .cdone_in(cdone_in[11]),
     .spioeb(spioeb[23:22]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[19:18]), .pado(pado[19:18]), .padeb(padeb[19:18]),
     .sp4_v_t(net866[0:15]), .sp4_h_l(SP4_h_l_12[47:0]),
     .sp12_h_l(SP12_h_l_12[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[23:22]), .tnl_op(lft_op_13[7:0]),
     .lft_op(lft_op_12[7:0]), .bnl_op(lft_op_11[7:0]),
     .pgate(pgate[191:176]), .reset(reset_b[191:176]),
     .sp4_v_b(net1172[0:15]), .wl(wl[191:176]), .cf(cf_r[287:264]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[191:176]),
     .slf_op(slf_op_12[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_12));
io_col4_RGT I_io_00_16 ( .ceb(ceb), .sdo(sdo), .sdi(net749),
     .spiout(spiout[31:30]), .cdone_in(cdone_in[15]),
     .spioeb(spioeb[31:30]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[27:26]), .pado(pado[27:26]), .padeb(padeb[27:26]),
     .sp4_v_t(sp4_v_t_16[15:0]), .sp4_h_l(SP4_h_l_16[47:0]),
     .sp12_h_l(SP12_h_l_16[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[31:30]), .tnl_op(tnl_op_16[7:0]),
     .lft_op(lft_op_16[7:0]), .bnl_op(lft_op_15[7:0]),
     .pgate(pgate[255:240]), .reset(reset_b[255:240]),
     .sp4_v_b(net764[0:15]), .wl(wl[255:240]), .cf(cf_r[383:360]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[255:240]),
     .slf_op(slf_op_16[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_16));
io_col4_RGT I_io_00_05 ( .ceb(ceb), .sdo(net919), .sdi(net1089),
     .spiout(spiout[9:8]), .cdone_in(cdone_in[4]),
     .spioeb(spioeb[9:8]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[5:4]), .pado(pado[5:4]), .padeb(padeb[5:4]),
     .sp4_v_t(net934[0:15]), .sp4_h_l(SP4_h_l_05[47:0]),
     .sp12_h_l(SP12_h_l_05[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[9:8]), .tnl_op(lft_op_06[7:0]),
     .lft_op(lft_op_05[7:0]), .bnl_op(lft_op_04[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net1104[0:15]), .wl(wl[79:64]), .cf(cf_r[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_05[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_05));
io_col4_RGT I_io_00_06 ( .ceb(ceb), .sdo(net953), .sdi(net919),
     .spiout(spiout[11:10]), .cdone_in(cdone_in[5]),
     .spioeb(spioeb[11:10]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[7:6]), .pado(pado[7:6]), .padeb(padeb[7:6]),
     .sp4_v_t(net968[0:15]), .sp4_h_l(SP4_h_l_06[47:0]),
     .sp12_h_l(SP12_h_l_06[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[11:10]), .tnl_op(lft_op_07[7:0]),
     .lft_op(lft_op_06[7:0]), .bnl_op(lft_op_05[7:0]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net934[0:15]), .wl(wl[95:80]), .cf(cf_r[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_06[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_06));
io_col4_RGT I_io_00_02 ( .ceb(ceb), .sdo(net987), .sdi(net1021),
     .spiout(spiout[3:2]), .cdone_in(cdone_in[1]),
     .spioeb(spioeb[3:2]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net1000[0:1]), .pado(net1000[0:1]), .padeb(net1001[0:1]),
     .sp4_v_t(net1002[0:15]), .sp4_h_l(SP4_h_l_02[47:0]),
     .sp12_h_l(SP12_h_l_02[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[3:2]), .tnl_op(lft_op_03[7:0]),
     .lft_op(lft_op_02[7:0]), .bnl_op(lft_op_01[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(net1036[0:15]), .wl(wl[31:16]), .cf(cf_r[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_02[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_02));
io_col4_RGT I_io_00_01 ( .ceb(ceb), .sdo(net1021), .sdi(sdi),
     .spiout(spiout[1:0]), .cdone_in(cdone_in[0]),
     .spioeb(spioeb[1:0]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net1034[0:1]), .pado(net1034[0:1]), .padeb(net1035[0:1]),
     .sp4_v_t(net1036[0:15]), .sp4_h_l(SP4_h_l_01[47:0]),
     .sp12_h_l(SP12_h_l_01[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .tnl_op(lft_op_02[7:0]),
     .lft_op(lft_op_01[7:0]), .bnl_op(bnl_op_01[7:0]),
     .pgate(pgate[15:0]), .reset(reset_b[15:0]),
     .sp4_v_b(sp4_v_b_01[15:0]), .wl(wl[15:0]), .cf(cf_r[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[15:0]), .slf_op(slf_op_01[3:0]),
     .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_01));
io_col4_RGT I_io_00_03 ( .ceb(ceb), .sdo(net1055), .sdi(net987),
     .spiout(spiout[5:4]), .cdone_in(cdone_in[2]),
     .spioeb(spioeb[5:4]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[1:0]), .pado(pado[1:0]), .padeb(padeb[1:0]),
     .sp4_v_t(net1070[0:15]), .sp4_h_l(SP4_h_l_03[47:0]),
     .sp12_h_l(SP12_h_l_03[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[5:4]), .tnl_op(lft_op_04[7:0]),
     .lft_op(lft_op_03[7:0]), .bnl_op(lft_op_02[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net1002[0:15]), .wl(wl[47:32]), .cf(cf_r[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_03[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_03));
io_col4_RGT I_io_00_04 ( .ceb(ceb), .sdo(net1089), .sdi(net1055),
     .spiout(spiout[7:6]), .cdone_in(cdone_in[3]),
     .spioeb(spioeb[7:6]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[3:2]), .pado(pado[3:2]), .padeb(padeb[3:2]),
     .sp4_v_t(net1104[0:15]), .sp4_h_l(SP4_h_l_04[47:0]),
     .sp12_h_l(SP12_h_l_04[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[7:6]), .tnl_op(lft_op_05[7:0]),
     .lft_op(lft_op_04[7:0]), .bnl_op(lft_op_03[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net1070[0:15]), .wl(wl[63:48]), .cf(cf_r[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_04[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_04));
io_col4_RGT I_io_00_10 ( .ceb(ceb), .sdo(net1123), .sdi(net647),
     .spiout(spiout[19:18]), .cdone_in(cdone_in[9]),
     .spioeb(spioeb[19:18]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[15:14]), .pado(pado[15:14]), .padeb(padeb[15:14]),
     .sp4_v_t(net1138[0:15]), .sp4_h_l(SP4_h_l_10[47:0]),
     .sp12_h_l(SP12_h_l_10[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[19:18]), .tnl_op(lft_op_11[7:0]),
     .lft_op(lft_op_10[7:0]), .bnl_op(lft_op_09[7:0]),
     .pgate(pgate[159:144]), .reset(reset_b[159:144]),
     .sp4_v_b(net662[0:15]), .wl(wl[159:144]), .cf(cf_r[239:216]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[159:144]),
     .slf_op(slf_op_10[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_10));
io_col4_RGT I_io_00_11 ( .ceb(ceb), .sdo(net1157), .sdi(net1123),
     .spiout(spiout[21:20]), .cdone_in(cdone_in[10]),
     .spioeb(spioeb[21:20]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[17:16]), .pado(pado[17:16]), .padeb(padeb[17:16]),
     .sp4_v_t(net1172[0:15]), .sp4_h_l(SP4_h_l_11[47:0]),
     .sp12_h_l(SP12_h_l_11[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[21:20]), .tnl_op(lft_op_12[7:0]),
     .lft_op(lft_op_11[7:0]), .bnl_op(lft_op_10[7:0]),
     .pgate(pgate[175:160]), .reset(reset_b[175:160]),
     .sp4_v_b(net1138[0:15]), .wl(wl[175:160]), .cf(cf_r[263:240]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[175:160]),
     .slf_op(slf_op_11[3:0]), .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_11));

endmodule
// Library - misc, Cell - ml_osc_stage, View - schematic
// LAST TIME SAVED: Sep  8 19:15:04 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_osc_stage ( out, clkin, oscen_b, pbias, sel_trim );
output  out;

input  clkin, oscen_b, pbias;

input [3:0]  sel_trim;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_mux3_hvt Iml_mux3_hvt_bot ( .in1(loadbot_1), .in0(loadbot_0),
     .out(in_bot), .sel(sel_trim[3:0]), .in2(loadbot_2));
nor2_hvt I228 ( .A(clkin), .B(oscen_b), .Y(net403));
inv_hvt I229 ( .A(net403), .Y(net419));
nch_hvt  MN41 ( .D(loadbot_0), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN39 ( .D(loadbot_2), .B(gnd_), .G(net419), .S(gnd_));
nch_hvt  MN29 ( .D(out), .B(gnd_), .G(in_bot), .S(gnd_));
nch_hvt  MN42 ( .D(loadbot_1), .B(gnd_), .G(net419), .S(gnd_));
pch_hvt  M82 ( .D(vdd_), .B(vdd_), .G(loadbot_1), .S(vdd_));
pch_hvt  M83 ( .D(vdd_), .B(vdd_), .G(loadbot_0), .S(vdd_));
pch_hvt  M85 ( .D(vdd_), .B(vdd_), .G(loadbot_2), .S(vdd_));
pch_hvt  M84 ( .D(vdd_), .B(vdd_), .G(loadbot_1), .S(vdd_));
pch_hvt  M81 ( .D(vdd_), .B(vdd_), .G(loadbot_2), .S(vdd_));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(loadbot_0), .S(vdd_));
pch_hvt  MP73 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net456));
pch_hvt  MP30 ( .D(net452), .B(vdd_), .G(oscen_b), .S(vdd_));
pch_hvt  MP72 ( .D(net456), .B(vdd_), .G(sel_trim[2]), .S(net452));
pch_hvt  MP33 ( .D(out), .B(vdd_), .G(in_bot), .S(vdd_));
pch_hvt  MP74 ( .D(in_bot), .B(vdd_), .G(pbias), .S(net452));

endmodule
// Library - leafcell, Cell - quad_br_ice8, View - schematic
// LAST TIME SAVED: Sep 18 15:35:51 2008
// NETLIST TIME: Nov 14 16:17:17 2008
`timescale 1ns / 1ns 

module quad_br_ice8 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_17_16, carry_out_18_16,
     carry_out_19_16, carry_out_20_16, carry_out_21_16,
     carry_out_22_16, carry_out_23_16, carry_out_24_16,
     carry_out_26_16, carry_out_27_16, carry_out_28_16,
     carry_out_29_16, carry_out_30_16, carry_out_31_16,
     carry_out_32_16, ceb_o, cf_b, cf_r, fabric_out_17_00,
     fabric_out_18_00, fabric_out_32_00, fabric_out_33_01,
     fabric_out_33_02, fabric_out_33_16, hiz_b_o, mode_o, padeb_b,
     padeb_r, padin_81, padin_135, pado_b, pado_r, r_o, sdo, sdo_pad,
     shift_o, slf_op_17_00, slf_op_17_01, slf_op_17_02, slf_op_17_03,
     slf_op_17_04, slf_op_17_05, slf_op_17_06, slf_op_17_07,
     slf_op_17_08, slf_op_17_09, slf_op_17_10, slf_op_17_11,
     slf_op_17_12, slf_op_17_13, slf_op_17_14, slf_op_17_15,
     slf_op_17_16, slf_op_18_16, slf_op_19_16, slf_op_20_16,
     slf_op_21_16, slf_op_22_16, slf_op_23_16, slf_op_24_16,
     slf_op_25_16, slf_op_26_16, slf_op_27_16, slf_op_28_16,
     slf_op_29_16, slf_op_30_16, slf_op_31_16, slf_op_32_16,
     slf_op_33_16, spi_ss_in_b, spi_ss_in_r, tclk_o, update_o, bl,
     pgate_r, reset_r, sp4_h_l_17_00, sp4_h_l_17_01, sp4_h_l_17_02,
     sp4_h_l_17_03, sp4_h_l_17_04, sp4_h_l_17_05, sp4_h_l_17_06,
     sp4_h_l_17_07, sp4_h_l_17_08, sp4_h_l_17_09, sp4_h_l_17_10,
     sp4_h_l_17_11, sp4_h_l_17_12, sp4_h_l_17_13, sp4_h_l_17_14,
     sp4_h_l_17_15, sp4_h_l_17_16, sp4_v_b_17_01, sp4_v_b_17_02,
     sp4_v_b_17_03, sp4_v_b_17_04, sp4_v_b_17_05, sp4_v_b_17_06,
     sp4_v_b_17_07, sp4_v_b_17_08, sp4_v_b_17_09, sp4_v_b_17_10,
     sp4_v_b_17_11, sp4_v_b_17_12, sp4_v_b_17_13, sp4_v_b_17_14,
     sp4_v_b_17_15, sp4_v_b_17_16, sp4_v_t_17_16, sp4_v_t_18_16,
     sp4_v_t_19_16, sp4_v_t_20_16, sp4_v_t_21_16, sp4_v_t_22_16,
     sp4_v_t_23_16, sp4_v_t_24_16, sp4_v_t_25_16, sp4_v_t_26_16,
     sp4_v_t_27_16, sp4_v_t_28_16, sp4_v_t_29_16, sp4_v_t_30_16,
     sp4_v_t_31_16, sp4_v_t_32_16, sp4_v_t_33_16, sp12_h_l_17_01,
     sp12_h_l_17_02, sp12_h_l_17_03, sp12_h_l_17_04, sp12_h_l_17_05,
     sp12_h_l_17_06, sp12_h_l_17_07, sp12_h_l_17_08, sp12_h_l_17_09,
     sp12_h_l_17_10, sp12_h_l_17_11, sp12_h_l_17_12, sp12_h_l_17_13,
     sp12_h_l_17_14, sp12_h_l_17_15, sp12_h_l_17_16, sp12_v_t_17_16,
     sp12_v_t_18_16, sp12_v_t_19_16, sp12_v_t_20_16, sp12_v_t_21_16,
     sp12_v_t_22_16, sp12_v_t_23_16, sp12_v_t_24_16, sp12_v_t_25_16,
     sp12_v_t_26_16, sp12_v_t_27_16, sp12_v_t_28_16, sp12_v_t_29_16,
     sp12_v_t_30_16, sp12_v_t_31_16, sp12_v_t_32_16, vdd_cntl_r, wl_r,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i,
     bnl_op_17_01, bs_en_i, bs_en_mi, ceb_i, ceb_mi,
     end_of_startup_bot_r, end_of_startup_rgt_b, glb_in, hiz_b_i,
     hiz_b_mi, hold_b_r, hold_r_b, lft_op_17_01, lft_op_17_02,
     lft_op_17_03, lft_op_17_04, lft_op_17_05, lft_op_17_06,
     lft_op_17_07, lft_op_17_08, lft_op_17_09, lft_op_17_10,
     lft_op_17_11, lft_op_17_12, lft_op_17_13, lft_op_17_14,
     lft_op_17_15, lft_op_17_16, mode_i, mode_mi, padin_b, padin_r,
     prog, purst, r_i, r_mi, sdi, sdi_pad, shift_i, shift_mi, spioeb_b,
     spioeb_r, spiout_b, spiout_r, tclk_i, tclk_mi, tiegnd,
     tnl_op_17_16, tnl_op_18_16, tnl_op_19_16, tnl_op_20_16,
     tnl_op_21_16, tnl_op_22_16, tnl_op_23_16, tnl_op_24_16,
     tnl_op_25_16, tnl_op_26_16, tnl_op_27_16, tnl_op_28_16,
     tnl_op_29_16, tnl_op_30_16, tnl_op_31_16, tnl_op_32_16,
     tnl_op_33_16, tnr_op_17_16, tnr_op_18_16, tnr_op_19_16,
     tnr_op_20_16, tnr_op_21_16, tnr_op_22_16, tnr_op_23_16,
     tnr_op_24_16, tnr_op_25_16, tnr_op_26_16, tnr_op_27_16,
     tnr_op_28_16, tnr_op_29_16, tnr_op_30_16, tnr_op_31_16,
     tnr_op_32_16, top_op_17_16, top_op_18_16, top_op_19_16,
     top_op_20_16, top_op_21_16, top_op_22_16, top_op_23_16,
     top_op_24_16, top_op_25_16, top_op_26_16, top_op_27_16,
     top_op_28_16, top_op_29_16, top_op_30_16, top_op_31_16,
     top_op_32_16, update_i, update_mi );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sreb_o,
     bm_wdummymux_en_o, bs_en_o, carry_out_17_16, carry_out_18_16,
     carry_out_19_16, carry_out_20_16, carry_out_21_16,
     carry_out_22_16, carry_out_23_16, carry_out_24_16,
     carry_out_26_16, carry_out_27_16, carry_out_28_16,
     carry_out_29_16, carry_out_30_16, carry_out_31_16,
     carry_out_32_16, ceb_o, fabric_out_17_00, fabric_out_18_00,
     fabric_out_32_00, fabric_out_33_01, fabric_out_33_02,
     fabric_out_33_16, hiz_b_o, mode_o, padin_81, padin_135, r_o, sdo,
     sdo_pad, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sreb_i,
     bm_wdummymux_en_i, bs_en_i, bs_en_mi, ceb_i, ceb_mi, hiz_b_i,
     hiz_b_mi, hold_b_r, hold_r_b, mode_i, mode_mi, prog, purst, r_i,
     r_mi, sdi, sdi_pad, shift_i, shift_mi, tclk_i, tclk_mi, tiegnd,
     update_i, update_mi;

output [383:0]  cf_r;
output [7:0]  slf_op_17_08;
output [1:0]  bm_sweb_o;
output [1:0]  bm_sdi_o;
output [56:30]  pado_b;
output [56:30]  padeb_b;
output [7:0]  slf_op_17_13;
output [7:0]  slf_op_24_16;
output [7:0]  slf_op_17_12;
output [7:0]  slf_op_25_16;
output [7:0]  slf_op_17_04;
output [7:0]  slf_op_17_16;
output [7:0]  slf_op_17_06;
output [7:0]  slf_op_26_16;
output [7:0]  slf_op_32_16;
output [7:0]  slf_op_17_07;
output [7:0]  slf_op_31_16;
output [7:0]  slf_op_17_15;
output [3:0]  slf_op_33_16;
output [1:0]  bm_sdo_o;
output [7:0]  slf_op_19_16;
output [1:0]  bm_sclkrw_o;
output [7:0]  slf_op_27_16;
output [31:0]  spi_ss_in_r;
output [7:0]  slf_op_21_16;
output [7:0]  slf_op_17_03;
output [7:0]  slf_op_20_16;
output [7:0]  slf_op_28_16;
output [7:0]  slf_op_18_16;
output [7:0]  slf_op_17_05;
output [27:0]  pado_r;
output [7:0]  slf_op_17_02;
output [7:0]  slf_op_17_14;
output [7:0]  slf_op_17_10;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_17_09;
output [3:0]  slf_op_17_00;
output [7:0]  slf_op_30_16;
output [7:0]  slf_op_17_11;
output [63:32]  spi_ss_in_b;
output [383:0]  cf_b;
output [7:0]  slf_op_29_16;
output [7:0]  slf_op_17_01;
output [7:0]  slf_op_23_16;
output [27:0]  padeb_r;
output [7:0]  slf_op_22_16;

inout [47:0]  sp4_v_t_26_16;
inout [47:0]  sp4_v_b_17_03;
inout [47:0]  sp4_v_b_17_16;
inout [23:0]  sp12_h_l_17_07;
inout [47:0]  sp4_v_t_22_16;
inout [23:0]  sp12_v_t_21_16;
inout [23:0]  sp12_v_t_23_16;
inout [23:0]  sp12_h_l_17_16;
inout [23:0]  sp12_v_t_26_16;
inout [23:0]  sp12_h_l_17_01;
inout [47:0]  sp4_h_l_17_09;
inout [23:0]  sp12_h_l_17_13;
inout [15:0]  sp4_h_l_17_00;
inout [23:0]  sp12_h_l_17_12;
inout [23:0]  sp12_h_l_17_14;
inout [47:0]  sp4_v_t_32_16;
inout [47:0]  sp4_h_l_17_12;
inout [47:0]  sp4_v_t_19_16;
inout [47:0]  sp4_h_l_17_14;
inout [47:0]  sp4_v_b_17_12;
inout [47:0]  sp4_v_t_30_16;
inout [23:0]  sp12_v_t_17_16;
inout [23:0]  sp12_h_l_17_04;
inout [47:0]  sp4_v_b_17_04;
inout [23:0]  sp12_v_t_24_16;
inout [47:0]  sp4_h_l_17_07;
inout [23:0]  sp12_v_t_29_16;
inout [47:0]  sp4_v_t_21_16;
inout [23:0]  sp12_v_t_28_16;
inout [47:0]  sp4_h_l_17_08;
inout [23:0]  sp12_h_l_17_06;
inout [47:0]  sp4_v_t_20_16;
inout [47:0]  sp4_v_t_28_16;
inout [47:0]  sp4_h_l_17_06;
inout [23:0]  sp12_h_l_17_05;
inout [47:0]  sp4_h_l_17_02;
inout [271:0]  reset_r;
inout [23:0]  sp12_h_l_17_15;
inout [15:0]  sp4_v_t_33_16;
inout [23:0]  sp12_h_l_17_02;
inout [23:0]  sp12_v_t_27_16;
inout [47:0]  sp4_h_l_17_11;
inout [23:0]  sp12_h_l_17_09;
inout [47:0]  sp4_v_t_31_16;
inout [47:0]  sp4_v_b_17_09;
inout [47:0]  sp4_v_b_17_06;
inout [23:0]  sp12_v_t_18_16;
inout [47:0]  sp4_v_t_25_16;
inout [47:0]  sp4_v_b_17_10;
inout [47:0]  sp4_v_b_17_13;
inout [23:0]  sp12_v_t_22_16;
inout [47:0]  sp4_v_b_17_14;
inout [23:0]  sp12_v_t_20_16;
inout [47:0]  sp4_v_b_17_01;
inout [47:0]  sp4_v_t_24_16;
inout [47:0]  sp4_v_b_17_11;
inout [23:0]  sp12_v_t_25_16;
inout [47:0]  sp4_v_t_27_16;
inout [47:0]  sp4_h_l_17_04;
inout [47:0]  sp4_h_l_17_15;
inout [47:0]  sp4_v_b_17_08;
inout [47:0]  sp4_v_t_23_16;
inout [47:0]  sp4_h_l_17_03;
inout [47:0]  sp4_v_b_17_02;
inout [47:0]  sp4_v_t_29_16;
inout [47:0]  sp4_v_b_17_05;
inout [23:0]  sp12_v_t_30_16;
inout [23:0]  sp12_h_l_17_11;
inout [23:0]  sp12_h_l_17_03;
inout [271:0]  vdd_cntl_r;
inout [47:0]  sp4_h_l_17_13;
inout [47:0]  sp4_v_t_17_16;
inout [47:0]  sp4_v_t_18_16;
inout [47:0]  sp4_h_l_17_01;
inout [47:0]  sp4_v_b_17_15;
inout [47:0]  sp4_h_l_17_10;
inout [271:0]  pgate_r;
inout [271:0]  wl_r;
inout [1743:874]  bl;
inout [23:0]  sp12_h_l_17_10;
inout [47:0]  sp4_h_l_17_16;
inout [23:0]  sp12_v_t_31_16;
inout [47:0]  sp4_h_l_17_05;
inout [23:0]  sp12_v_t_19_16;
inout [47:0]  sp4_v_b_17_07;
inout [23:0]  sp12_h_l_17_08;
inout [23:0]  sp12_v_t_32_16;

input [7:0]  lft_op_17_16;
input [7:0]  tnl_op_33_16;
input [7:0]  top_op_29_16;
input [7:0]  lft_op_17_13;
input [7:0]  lft_op_17_08;
input [31:0]  spiout_r;
input [7:0]  tnl_op_19_16;
input [7:0]  lft_op_17_02;
input [31:16]  end_of_startup_bot_r;
input [7:0]  tnr_op_30_16;
input [7:0]  lft_op_17_06;
input [7:0]  tnl_op_28_16;
input [7:0]  tnr_op_26_16;
input [7:0]  lft_op_17_07;
input [7:0]  tnr_op_25_16;
input [7:0]  tnr_op_17_16;
input [31:0]  spioeb_r;
input [7:0]  tnr_op_27_16;
input [1:0]  bm_sclkrw_i;
input [7:0]  tnr_op_23_16;
input [7:0]  tnl_op_26_16;
input [7:0]  tnl_op_30_16;
input [7:0]  glb_in;
input [7:0]  tnr_op_24_16;
input [7:0]  tnr_op_28_16;
input [7:0]  top_op_32_16;
input [7:0]  lft_op_17_12;
input [7:0]  bm_sa_i;
input [7:0]  tnl_op_20_16;
input [7:0]  lft_op_17_01;
input [1:0]  bm_sdo_i;
input [1:0]  bm_sweb_i;
input [7:0]  top_op_22_16;
input [7:0]  top_op_25_16;
input [7:0]  lft_op_17_05;
input [3:0]  bnl_op_17_01;
input [7:0]  lft_op_17_14;
input [63:32]  spioeb_b;
input [7:0]  lft_op_17_04;
input [7:0]  top_op_18_16;
input [27:0]  padin_r;
input [7:0]  tnl_op_21_16;
input [7:0]  tnr_op_20_16;
input [7:0]  lft_op_17_10;
input [63:32]  spiout_b;
input [7:0]  lft_op_17_15;
input [7:0]  tnr_op_29_16;
input [7:0]  tnr_op_31_16;
input [7:0]  lft_op_17_09;
input [7:0]  tnr_op_21_16;
input [7:0]  tnl_op_27_16;
input [7:0]  tnr_op_18_16;
input [7:0]  lft_op_17_11;
input [7:0]  top_op_26_16;
input [7:0]  top_op_28_16;
input [7:0]  tnl_op_32_16;
input [7:0]  tnl_op_18_16;
input [7:0]  tnr_op_22_16;
input [1:0]  bm_sdi_i;
input [7:0]  top_op_17_16;
input [7:0]  tnl_op_22_16;
input [7:0]  top_op_24_16;
input [7:0]  tnl_op_25_16;
input [7:0]  top_op_21_16;
input [7:0]  tnr_op_32_16;
input [7:0]  top_op_27_16;
input [56:30]  padin_b;
input [7:0]  top_op_23_16;
input [7:0]  lft_op_17_03;
input [7:0]  tnl_op_29_16;
input [7:0]  tnl_op_31_16;
input [16:1]  end_of_startup_rgt_b;
input [7:0]  top_op_31_16;
input [7:0]  tnl_op_24_16;
input [7:0]  tnl_op_23_16;
input [7:0]  tnr_op_19_16;
input [7:0]  top_op_20_16;
input [7:0]  tnl_op_17_16;
input [7:0]  top_op_30_16;
input [7:0]  top_op_19_16;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net4618;

wire  [0:23]  net3883;

wire  [0:47]  net4932;

wire  [0:47]  net4439;

wire  [0:7]  net4451;

wire  [0:47]  net4256;

wire  [0:47]  net4154;

wire  [0:7]  net3533;

wire  [0:23]  net4045;

wire  [0:7]  net4839;

wire  [0:7]  net2592;

wire  [0:7]  net4837;

wire  [0:23]  net4470;

wire  [0:23]  net3071;

wire  [0:47]  net4853;

wire  [0:47]  net4440;

wire  [0:23]  net4960;

wire  [0:47]  net2585;

wire  [0:7]  net4291;

wire  [0:23]  net4209;

wire  [0:7]  net2718;

wire  [0:23]  net4632;

wire  [0:47]  net4316;

wire  [0:23]  net3980;

wire  [0:7]  net2659;

wire  [0:47]  net3501;

wire  [0:23]  net2678;

wire  [0:47]  net4606;

wire  [0:47]  net2546;

wire  [0:47]  net4092;

wire  [0:47]  net4003;

wire  [0:47]  net2892;

wire  [0:23]  net3721;

wire  [0:47]  net4965;

wire  [0:7]  net4674;

wire  [0:23]  net3560;

wire  [0:23]  net3494;

wire  [0:47]  net4983;

wire  [0:47]  net3336;

wire  [0:7]  net2722;

wire  [0:47]  net4416;

wire  [0:23]  net4860;

wire  [0:7]  net2824;

wire  [0:47]  net3843;

wire  [0:7]  net4711;

wire  [0:23]  net3398;

wire  [0:47]  net2896;

wire  [0:47]  net4280;

wire  [0:47]  net2682;

wire  [0:47]  net4276;

wire  [0:23]  net2401;

wire  [0:47]  net2626;

wire  [0:23]  net2939;

wire  [0:7]  net3473;

wire  [0:47]  net2787;

wire  [0:47]  net4037;

wire  [0:47]  net2110;

wire  [0:7]  net2757;

wire  [0:47]  net3924;

wire  [0:47]  net5013;

wire  [0:7]  net2109;

wire  [0:47]  net4603;

wire  [0:47]  net2189;

wire  [0:47]  net3545;

wire  [0:47]  net2104;

wire  [0:23]  net3397;

wire  [0:23]  net3983;

wire  [0:7]  net3048;

wire  [0:7]  net4558;

wire  [0:7]  net4838;

wire  [0:47]  net3013;

wire  [0:47]  net3026;

wire  [0:23]  net4864;

wire  [0:7]  net5001;

wire  [0:47]  net3989;

wire  [0:23]  net2843;

wire  [0:7]  net2821;

wire  [0:47]  net3441;

wire  [0:7]  net2147;

wire  [0:47]  net3842;

wire  [0:47]  net4277;

wire  [0:7]  net4779;

wire  [0:7]  net4515;

wire  [0:7]  net2434;

wire  [0:47]  net3010;

wire  [0:23]  net3486;

wire  [0:47]  net2945;

wire  [0:47]  net4332;

wire  [0:47]  net3708;

wire  [0:7]  net3407;

wire  [0:7]  net4292;

wire  [0:47]  net3352;

wire  [0:47]  net2458;

wire  [0:7]  net3246;

wire  [0:23]  net2746;

wire  [0:47]  net2540;

wire  [0:47]  net3512;

wire  [0:47]  net4769;

wire  [0:47]  net4522;

wire  [0:47]  net4197;

wire  [0:47]  net4848;

wire  [0:47]  net2352;

wire  [0:47]  net2542;

wire  [0:47]  net2619;

wire  [0:47]  net4819;

wire  [0:47]  net3712;

wire  [0:47]  net3339;

wire  [0:23]  net2389;

wire  [0:47]  net2730;

wire  [0:7]  net2881;

wire  [0:47]  net4442;

wire  [0:47]  net3011;

wire  [0:47]  net4816;

wire  [0:47]  net4980;

wire  [0:47]  net3986;

wire  [0:23]  net3819;

wire  [0:23]  net3396;

wire  [0:47]  net2537;

wire  [0:7]  net3570;

wire  [0:23]  net2393;

wire  [0:7]  net3699;

wire  [0:47]  net3826;

wire  [0:47]  net2732;

wire  [0:7]  net3537;

wire  [0:47]  net3115;

wire  [0:7]  net2436;

wire  [0:47]  net4638;

wire  [0:47]  net2583;

wire  [0:47]  net4805;

wire  [0:47]  net2848;

wire  [0:47]  net2623;

wire  [0:47]  net4850;

wire  [0:47]  net4250;

wire  [0:47]  net4253;

wire  [0:23]  net3975;

wire  [0:23]  net3593;

wire  [0:7]  net2721;

wire  [0:7]  net4513;

wire  [0:47]  net4417;

wire  [0:15]  net2191;

wire  [0:47]  net4443;

wire  [0:47]  net2541;

wire  [0:47]  net4151;

wire  [0:23]  net3722;

wire  [0:47]  net4004;

wire  [0:47]  net4090;

wire  [0:47]  net3953;

wire  [0:47]  net4418;

wire  [0:47]  net4279;

wire  [0:7]  net4511;

wire  [0:7]  net2986;

wire  [0:7]  net3370;

wire  [0:47]  net3438;

wire  [0:23]  net4537;

wire  [0:47]  net2701;

wire  [0:47]  net4093;

wire  [0:47]  net4412;

wire  [0:47]  net4413;

wire  [0:23]  net4538;

wire  [0:7]  net3966;

wire  [0:47]  net4164;

wire  [0:7]  net4454;

wire  [0:23]  net3323;

wire  [0:7]  net2122;

wire  [0:7]  net4942;

wire  [0:47]  net4150;

wire  [0:7]  net3047;

wire  [0:23]  net3918;

wire  [0:47]  net2539;

wire  [0:23]  net3493;

wire  [0:7]  net2108;

wire  [0:7]  net3962;

wire  [0:23]  net4894;

wire  [0:23]  net5028;

wire  [0:23]  net3724;

wire  [0:23]  net4050;

wire  [0:7]  net4780;

wire  [0:7]  net2928;

wire  [0:47]  net4906;

wire  [0:7]  net2441;

wire  [0:47]  net3136;

wire  [0:23]  net2841;

wire  [0:47]  net3790;

wire  [0:23]  net3070;

wire  [0:47]  net2348;

wire  [0:47]  net3060;

wire  [0:47]  net2620;

wire  [0:23]  net2103;

wire  [0:47]  net4005;

wire  [0:23]  net4308;

wire  [0:7]  net3963;

wire  [0:23]  net3657;

wire  [0:23]  net2132;

wire  [0:47]  net2548;

wire  [0:23]  net4080;

wire  [0:23]  net3590;

wire  [0:7]  net4677;

wire  [0:23]  net2940;

wire  [0:23]  net2840;

wire  [0:47]  net2811;

wire  [0:47]  net4818;

wire  [0:47]  net2354;

wire  [0:23]  net4636;

wire  [0:47]  net2450;

wire  [0:23]  net3753;

wire  [0:47]  net3383;

wire  [0:23]  net3492;

wire  [0:23]  net4242;

wire  [0:7]  net2123;

wire  [0:47]  net4153;

wire  [0:23]  net2156;

wire  [0:47]  net3138;

wire  [0:23]  net2677;

wire  [0:47]  net3988;

wire  [0:47]  net4249;

wire  [0:47]  net2782;

wire  [0:47]  net2684;

wire  [0:23]  net4635;

wire  [0:47]  net3827;

wire  [0:7]  net3310;

wire  [0:47]  net3597;

wire  [0:7]  net2138;

wire  [0:7]  net4232;

wire  [0:23]  net4408;

wire  [0:47]  net4492;

wire  [0:23]  net2089;

wire  [0:47]  net3839;

wire  [0:23]  net3329;

wire  [0:7]  net3244;

wire  [0:7]  net3906;

wire  [0:23]  net2615;

wire  [0:47]  net3351;

wire  [0:23]  net2090;

wire  [0:7]  net2884;

wire  [0:23]  net4212;

wire  [0:47]  net2686;

wire  [0:7]  net3640;

wire  [0:47]  net4801;

wire  [0:47]  net3276;

wire  [0:7]  net2184;

wire  [0:47]  net3462;

wire  [0:23]  net3820;

wire  [0:7]  net5003;

wire  [0:23]  net4081;

wire  [0:23]  net4536;

wire  [0:7]  net4189;

wire  [0:47]  net3008;

wire  [0:23]  net2399;

wire  [0:47]  net3990;

wire  [0:47]  net2050;

wire  [0:23]  net2408;

wire  [0:23]  net2743;

wire  [0:47]  net3950;

wire  [0:7]  net4129;

wire  [0:47]  net3354;

wire  [0:47]  net3463;

wire  [0:47]  net3925;

wire  [0:47]  net4149;

wire  [0:7]  net4349;

wire  [0:7]  net2075;

wire  [0:47]  net4685;

wire  [0:7]  net4348;

wire  [0:47]  net4577;

wire  [0:47]  net2646;

wire  [0:47]  net4313;

wire  [0:47]  net4928;

wire  [0:23]  net3101;

wire  [0:23]  net2741;

wire  [0:47]  net3952;

wire  [0:23]  net2680;

wire  [0:47]  net2538;

wire  [0:7]  net2431;

wire  [0:47]  net3871;

wire  [0:47]  net3823;

wire  [0:47]  net3824;

wire  [0:47]  net4653;

wire  [0:7]  net3735;

wire  [0:47]  net2536;

wire  [0:47]  net3497;

wire  [0:7]  net2062;

wire  [0:47]  net2683;

wire  [0:7]  net2661;

wire  [0:47]  net2351;

wire  [0:47]  net2650;

wire  [0:47]  net2621;

wire  [0:23]  net3430;

wire  [0:23]  net4732;

wire  [0:47]  net4523;

wire  [0:7]  net4185;

wire  [0:7]  net4351;

wire  [0:47]  net3057;

wire  [0:47]  net4738;

wire  [0:47]  net2733;

wire  [0:23]  net4144;

wire  [0:47]  net3298;

wire  [0:7]  net2765;

wire  [0:23]  net5026;

wire  [0:23]  net4079;

wire  [0:47]  net4742;

wire  [0:7]  net2074;

wire  [0:7]  net5000;

wire  [0:47]  net2117;

wire  [0:23]  net3655;

wire  [0:23]  net3754;

wire  [0:47]  net4656;

wire  [0:47]  net2125;

wire  [0:23]  net4244;

wire  [0:47]  net4331;

wire  [0:47]  net4576;

wire  [0:47]  net4768;

wire  [0:47]  net2344;

wire  [0:47]  net4330;

wire  [0:23]  net2679;

wire  [0:23]  net4211;

wire  [0:7]  net4024;

wire  [0:7]  net4025;

wire  [0:47]  net2625;

wire  [0:47]  net3278;

wire  [0:47]  net2947;

wire  [0:23]  net4702;

wire  [0:23]  net4568;

wire  [0:47]  net3665;

wire  [0:47]  net3277;

wire  [0:7]  net4876;

wire  [0:47]  net4639;

wire  [0:47]  net2849;

wire  [0:47]  net4251;

wire  [0:23]  net2941;

wire  [0:7]  net4778;

wire  [0:47]  net4686;

wire  [0:47]  net3664;

wire  [0:47]  net3055;

wire  [0:47]  net3923;

wire  [0:47]  net3381;

wire  [0:47]  net4929;

wire  [0:7]  net2102;

wire  [0:47]  net4739;

wire  [0:47]  net3928;

wire  [0:47]  net4168;

wire  [0:23]  net4697;

wire  [0:23]  net4301;

wire  [0:47]  net4118;

wire  [0:47]  net4820;

wire  [0:47]  net3461;

wire  [0:23]  net4627;

wire  [0:7]  net2823;

wire  [0:23]  net3723;

wire  [0:47]  net4765;

wire  [0:47]  net4905;

wire  [0:47]  net4364;

wire  [0:47]  net4902;

wire  [0:7]  net3733;

wire  [0:47]  net2535;

wire  [0:47]  net2729;

wire  [0:7]  net2984;

wire  [0:23]  net2613;

wire  [0:47]  net4479;

wire  [0:7]  net4550;

wire  [0:23]  net3495;

wire  [0:47]  net3709;

wire  [0:47]  net3680;

wire  [0:23]  net3264;

wire  [0:23]  net4861;

wire  [0:23]  net4863;

wire  [0:23]  net4143;

wire  [0:47]  net3302;

wire  [0:47]  net2543;

wire  [0:7]  net3046;

wire  [0:7]  net4395;

wire  [0:23]  net2164;

wire  [0:23]  net3491;

wire  [0:47]  net2894;

wire  [0:23]  net4307;

wire  [0:47]  net2462;

wire  [0:47]  net2972;

wire  [0:47]  net3766;

wire  [0:7]  net3639;

wire  [0:7]  net2885;

wire  [0:23]  net4309;

wire  [0:47]  net2455;

wire  [0:47]  net4802;

wire  [0:23]  net2390;

wire  [0:7]  net4615;

wire  [0:23]  net3428;

wire  [0:47]  net3663;

wire  [0:23]  net2778;

wire  [0:47]  net4196;

wire  [0:47]  net3660;

wire  [0:7]  net2826;

wire  [3:0]  slf_op_29_00;

wire  [3:0]  slf_op_31_00;

wire  [3:0]  slf_op_21_00;

wire  [3:0]  slf_op_19_00;

wire  [3:0]  slf_op_22_00;

wire  [3:0]  slf_op_30_00;

wire  [0:23]  net4047;

wire  [0:23]  net3265;

wire  [0:7]  net4713;

wire  [0:23]  net4699;

wire  [0:23]  net4405;

wire  [0:23]  net3002;

wire  [7:0]  clk_tree_drv;

wire  [0:7]  net3535;

wire  [3:0]  slf_op_26_00;

wire  [3:0]  slf_op_18_00;

wire  [0:7]  net2663;

wire  [0:23]  net2402;

wire  [0:47]  net4767;

wire  [0:7]  net4616;

wire  [0:47]  net2065;

wire  [0:23]  net3395;

wire  [0:23]  net2744;

wire  [0:47]  net3762;

wire  [0:7]  net3896;

wire  [0:7]  net4777;

wire  [0:23]  net4138;

wire  [47:0]  sp4_h_r_17_18;

wire  [47:0]  sp4_h_r_18_19;

wire  [47:0]  sp4_h_r_19_20;

wire  [47:0]  sp4_h_r_20_21;

wire  [3:0]  slf_op_28_00;

wire  [3:0]  slf_op_27_00;

wire  [3:0]  slf_op_25_00;

wire  [3:0]  slf_op_20_00;

wire  [3:0]  slf_op_24_00;

wire  [3:0]  slf_op_32_00;

wire  [0:7]  net2660;

wire  [0:47]  net2687;

wire  [0:7]  net3311;

wire  [0:47]  net3599;

wire  [0:47]  net3337;

wire  [0:47]  net3678;

wire  [0:47]  net4602;

wire  [0:23]  net2906;

wire  [0:47]  net2545;

wire  [0:7]  net2442;

wire  [0:47]  net2341;

wire  [0:47]  net2977;

wire  [0:23]  net2140;

wire  [0:7]  net3700;

wire  [0:47]  net4361;

wire  [0:47]  net2698;

wire  [0:7]  net2435;

wire  [0:7]  net4940;

wire  [0:7]  net2985;

wire  [0:7]  net2594;

wire  [0:47]  net3440;

wire  [0:47]  net2814;

wire  [0:47]  net4038;

wire  [0:47]  net3764;

wire  [0:47]  net2863;

wire  [0:23]  net4310;

wire  [0:47]  net3954;

wire  [0:7]  net2719;

wire  [0:47]  net3675;

wire  [0:47]  net2452;

wire  [0:7]  net2130;

wire  [0:23]  net3169;

wire  [0:7]  net2918;

wire  [0:47]  net4087;

wire  [0:47]  net3930;

wire  [0:23]  net2908;

wire  [0:47]  net3140;

wire  [0:7]  net2882;

wire  [0:47]  net2149;

wire  [0:47]  net5016;

wire  [0:47]  net2449;

wire  [0:47]  net3271;

wire  [0:47]  net2783;

wire  [0:47]  net5011;

wire  [0:23]  net2742;

wire  [0:47]  net3765;

wire  [0:47]  net3951;

wire  [0:47]  net4033;

wire  [0:23]  net3004;

wire  [0:47]  net2353;

wire  [0:7]  net4352;

wire  [0:23]  net3984;

wire  [0:47]  net4817;

wire  [0:7]  net4781;

wire  [0:47]  net4086;

wire  [0:7]  net4059;

wire  [0:47]  net4640;

wire  [0:7]  net3475;

wire  [0:23]  net4406;

wire  [0:23]  net3005;

wire  [0:23]  net3393;

wire  [0:47]  net2456;

wire  [0:47]  net3466;

wire  [0:7]  net4512;

wire  [0:47]  net2459;

wire  [0:47]  net3435;

wire  [0:23]  net4959;

wire  [0:23]  net3230;

wire  [0:7]  net2155;

wire  [0:7]  net3044;

wire  [0:47]  net4278;

wire  [0:23]  net5025;

wire  [0:47]  net3334;

wire  [0:23]  net4796;

wire  [0:23]  net3658;

wire  [0:47]  net4493;

wire  [0:47]  net2648;

wire  [0:23]  net4862;

wire  [0:47]  net2951;

wire  [0:7]  net4455;

wire  [0:7]  net2440;

wire  [0:23]  net3556;

wire  [0:47]  net2451;

wire  [0:23]  net4700;

wire  [0:47]  net4006;

wire  [0:23]  net4958;

wire  [0:23]  net3427;

wire  [0:47]  net3299;

wire  [0:23]  net3394;

wire  [0:47]  net4687;

wire  [0:47]  net2165;

wire  [0:47]  net4444;

wire  [0:7]  net3409;

wire  [0:47]  net2092;

wire  [0:47]  net3338;

wire  [0:47]  net4654;

wire  [0:47]  net3058;

wire  [0:47]  net3059;

wire  [0:7]  net4188;

wire  [0:7]  net4514;

wire  [0:47]  net4931;

wire  [0:7]  net4617;

wire  [0:23]  net3168;

wire  [0:23]  net4147;

wire  [0:7]  net4288;

wire  [0:47]  net4981;

wire  [0:23]  net3068;

wire  [0:47]  net4088;

wire  [0:23]  net2394;

wire  [0:47]  net3661;

wire  [0:7]  net4186;

wire  [0:47]  net2846;

wire  [0:47]  net4964;

wire  [0:23]  net4372;

wire  [0:7]  net2116;

wire  [0:7]  net2087;

wire  [0:47]  net3838;

wire  [0:23]  net3006;

wire  [0:47]  net4933;

wire  [0:23]  net3330;

wire  [0:47]  net4363;

wire  [0:47]  net3135;

wire  [0:23]  net2180;

wire  [0:23]  net3266;

wire  [0:23]  net2671;

wire  [0:23]  net5024;

wire  [0:7]  net4069;

wire  [0:47]  net2952;

wire  [0:23]  net3981;

wire  [0:23]  net2409;

wire  [0:23]  net3558;

wire  [0:47]  net4035;

wire  [0:23]  net4701;

wire  [0:47]  net3549;

wire  [0:23]  net3982;

wire  [0:23]  net2406;

wire  [0:47]  net2463;

wire  [0:7]  net2178;

wire  [0:47]  net2784;

wire  [0:47]  net4312;

wire  [0:23]  net4048;

wire  [0:23]  net3235;

wire  [0:47]  net4091;

wire  [0:7]  net3314;

wire  [0:47]  net2356;

wire  [0:47]  net4117;

wire  [0:7]  net3478;

wire  [0:47]  net2550;

wire  [0:47]  net3547;

wire  [0:47]  net2893;

wire  [0:47]  net4476;

wire  [0:47]  net3788;

wire  [0:47]  net4744;

wire  [0:7]  net3965;

wire  [0:47]  net2624;

wire  [0:23]  net2049;

wire  [0:23]  net2834;

wire  [0:47]  net4655;

wire  [0:23]  net3160;

wire  [0:7]  net4222;

wire  [0:7]  net4452;

wire  [0:23]  net4472;

wire  [0:7]  net2171;

wire  [0:23]  net2997;

wire  [0:23]  net4534;

wire  [0:23]  net4210;

wire  [0:23]  net4798;

wire  [0:23]  net4797;

wire  [0:47]  net3502;

wire  [0:47]  net4360;

wire  [0:23]  net3917;

wire  [0:7]  net4676;

wire  [0:7]  net3313;

wire  [0:47]  net4803;

wire  [0:47]  net2697;

wire  [0:23]  net2612;

wire  [0:23]  net3328;

wire  [0:47]  net3028;

wire  [0:7]  net3799;

wire  [0:47]  net4255;

wire  [0:23]  net3069;

wire  [0:47]  net3603;

wire  [0:7]  net2987;

wire  [0:47]  net4657;

wire  [0:47]  net3870;

wire  [0:23]  net4145;

wire  [0:23]  net3919;

wire  [0:7]  net3967;

wire  [0:7]  net2662;

wire  [0:23]  net4535;

wire  [0:47]  net2133;

wire  [0:47]  net3761;

wire  [0:47]  net4642;

wire  [0:23]  net4897;

wire  [0:23]  net4570;

wire  [0:47]  net3513;

wire  [0:47]  net2549;

wire  [0:47]  net2812;

wire  [0:47]  net2786;

wire  [0:7]  net2443;

wire  [0:23]  net3559;

wire  [0:47]  net4849;

wire  [0:47]  net2734;

wire  [0:47]  net4328;

wire  [0:47]  net3275;

wire  [0:47]  net4582;

wire  [0:23]  net4733;

wire  [0:7]  net4945;

wire  [0:47]  net3927;

wire  [0:7]  net2139;

wire  [0:23]  net4471;

wire  [0:7]  net3580;

wire  [0:47]  net3272;

wire  [0:47]  net4579;

wire  [0:47]  net4851;

wire  [0:47]  net4477;

wire  [0:7]  net4675;

wire  [0:47]  net2685;

wire  [0:47]  net3386;

wire  [0:47]  net4001;

wire  [0:47]  net4525;

wire  [0:47]  net3499;

wire  [0:47]  net4740;

wire  [0:7]  net2720;

wire  [0:7]  net2047;

wire  [0:47]  net4116;

wire  [0:47]  net3139;

wire  [0:7]  net2658;

wire  [0:47]  net3624;

wire  [0:47]  net3188;

wire  [0:23]  net3165;

wire  [0:7]  net3803;

wire  [0:7]  net2177;

wire  [0:47]  net3991;

wire  [0:7]  net4874;

wire  [0:23]  net3656;

wire  [0:47]  net3710;

wire  [0:7]  net2088;

wire  [0:47]  net4908;

wire  [0:23]  net4539;

wire  [0:47]  net4968;

wire  [0:47]  net2789;

wire  [0:47]  net4152;

wire  [0:7]  net3801;

wire  [0:47]  net2349;

wire  [0:47]  net2864;

wire  [0:7]  net3859;

wire  [0:23]  net2091;

wire  [0:23]  net4243;

wire  [0:47]  net3056;

wire  [0:47]  net4524;

wire  [0:23]  net4375;

wire  [0:7]  net3861;

wire  [0:47]  net2454;

wire  [0:7]  net4944;

wire  [0:47]  net4969;

wire  [0:23]  net4634;

wire  [0:7]  net2437;

wire  [0:23]  net2842;

wire  [0:7]  net3862;

wire  [0:7]  net2602;

wire  [0:47]  net4166;

wire  [0:47]  net4327;

wire  [0:23]  net3067;

wire  [0:47]  net4979;

wire  [0:23]  net3561;

wire  [0:47]  net4982;

wire  [0:7]  net3698;

wire  [0:7]  net3696;

wire  [0:7]  net2188;

wire  [0:47]  net2861;

wire  [0:47]  net4581;

wire  [0:7]  net2163;

wire  [0:47]  net2946;

wire  [0:23]  net3232;

wire  [0:47]  net2850;

wire  [0:23]  net4731;

wire  [0:47]  net4907;

wire  [0:7]  net4548;

wire  [0:7]  net2433;

wire  [0:47]  net4478;

wire  [0:47]  net4034;

wire  [0:7]  net3373;

wire  [0:47]  net2731;

wire  [0:47]  net2651;

wire  [0:47]  net2544;

wire  [0:23]  net4734;

wire  [0:47]  net3987;

wire  [0:23]  net2938;

wire  [0:47]  net2845;

wire  [0:47]  net4852;

wire  [0:47]  net3190;

wire  [0:47]  net3349;

wire  [0:47]  net2865;

wire  [0:47]  net3025;

wire  [0:7]  net2988;

wire  [0:7]  net3637;

wire  [0:7]  net2444;

wire  [0:23]  net4146;

wire  [0:23]  net3719;

wire  [0:23]  net2124;

wire  [0:7]  net3536;

wire  [0:47]  net3187;

wire  [0:23]  net3234;

wire  [0:47]  net3929;

wire  [0:23]  net3755;

wire  [0:47]  net2862;

wire  [0:7]  net4022;

wire  [0:23]  net2081;

wire  [0:23]  net3231;

wire  [0:47]  net2457;

wire  [0:47]  net2700;

wire  [0:7]  net2185;

wire  [0:23]  net3591;

wire  [0:47]  net4165;

wire  [0:47]  net4002;

wire  [0:47]  net4169;

wire  [0:7]  net3697;

wire  [0:47]  net2975;

wire  [0:7]  net5002;

wire  [0:23]  net4464;

wire  [0:47]  net4198;

wire  [0:47]  net3353;

wire  [0:47]  net4607;

wire  [0:23]  net3817;

wire  [0:47]  net2813;

wire  [0:7]  net4127;

wire  [0:47]  net3626;

wire  [0:47]  net2346;

wire  [0:23]  net2777;

wire  [0:47]  net2453;

wire  [0:47]  net4115;

wire  [0:7]  net2146;

wire  [0:47]  net3498;

wire  [0:23]  net2905;

wire  [0:47]  net3027;

wire  [0:47]  net3436;

wire  [0:47]  net4441;

wire  [0:7]  net4941;

wire  [0:23]  net3102;

wire  [0:47]  net3303;

wire  [0:7]  net2822;

wire  [0:47]  net4643;

wire  [0:47]  net2809;

wire  [0:7]  net4453;

wire  [0:7]  net3638;

wire  [0:47]  net3548;

wire  [0:7]  net2920;

wire  [0:47]  net3767;

wire  [0:47]  net4575;

wire  [0:23]  net4571;

wire  [0:47]  net3629;

wire  [0:47]  net4641;

wire  [0:7]  net4128;

wire  [0:23]  net4961;

wire  [0:23]  net4082;

wire  [0:47]  net3301;

wire  [0:23]  net3331;

wire  [0:23]  net3003;

wire  [0:47]  net2096;

wire  [0:47]  net2547;

wire  [0:47]  net4604;

wire  [0:47]  net5014;

wire  [0:47]  net3872;

wire  [0:7]  net4782;

wire  [0:47]  net3677;

wire  [0:47]  net4580;

wire  [0:7]  net2154;

wire  [0:23]  net3166;

wire  [0:47]  net4689;

wire  [0:7]  net3477;

wire  [0:7]  net2883;

wire  [0:47]  net2788;

wire  [0:23]  net2676;

wire  [0:47]  net3191;

wire  [0:47]  net3791;

wire  [0:47]  net2357;

wire  [0:23]  net3916;

wire  [0:7]  net4840;

wire  [0:23]  net3267;

wire  [0:7]  net4125;

wire  [0:23]  net3885;

wire  [0:47]  net3828;

wire  [0:47]  net3009;

wire  [0:47]  net4281;

wire  [0:47]  net5012;

wire  [0:47]  net4414;

wire  [0:47]  net4494;

wire  [0:47]  net4903;

wire  [0:47]  net3273;

wire  [0:47]  net2141;

wire  [0:47]  net3384;

wire  [0:23]  net4306;

wire  [0:47]  net4114;

wire  [0:47]  net3189;

wire  [0:7]  net2989;

wire  [0:7]  net4130;

wire  [0:23]  net4962;

wire  [0:7]  net4943;

wire  [0:47]  net2702;

wire  [0:23]  net2404;

wire  [0:47]  net3382;

wire  [0:23]  net3887;

wire  [0:7]  net3254;

wire  [0:47]  net3012;

wire  [0:23]  net2909;

wire  [0:47]  net3707;

wire  [0:7]  net3743;

wire  [0:7]  net3312;

wire  [0:47]  net3464;

wire  [0:23]  net4049;

wire  [0:47]  net3679;

wire  [0:7]  net3636;

wire  [0:23]  net4208;

wire  [0:47]  net3841;

wire  [0:23]  net3756;

wire  [0:23]  net3167;

wire  [0:23]  net3654;

wire  [0:47]  net4254;

wire  [0:7]  net4023;

wire  [0:23]  net2775;

wire  [0:7]  net3045;

wire  [0:23]  net3882;

wire  [0:23]  net4633;

wire  [0:23]  net3818;

wire  [0:47]  net3514;

wire  [0:23]  net2407;

wire  [0:47]  net3350;

wire  [0:7]  net2439;

wire  [0:7]  net4187;

wire  [0:47]  net3787;

wire  [0:47]  net5015;

wire  [0:7]  net4293;

wire  [0:7]  net3534;

wire  [0:23]  net3649;

wire  [0:47]  net3825;

wire  [0:47]  net4527;

wire  [0:47]  net4766;

wire  [0:47]  net2345;

wire  [0:7]  net4456;

wire  [0:47]  net3789;

wire  [0:47]  net4770;

wire  [0:7]  net4026;

wire  [0:23]  net2329;

wire  [0:7]  net3372;

wire  [0:47]  net4490;

wire  [0:47]  net3601;

wire  [0:7]  net3860;

wire  [0:47]  net2182;

wire  [0:47]  net4475;

wire  [0:7]  net4721;

wire  [0:23]  net4865;

wire  [0:7]  net4841;

wire  [0:47]  net2949;

wire  [0:7]  net3802;

wire  [0:47]  net2976;

wire  [0:47]  net4743;

wire  [0:23]  net2904;

wire  [0:47]  net3335;

wire  [0:23]  net4407;

wire  [0:23]  net4245;

wire  [0:47]  net2973;

wire  [0:7]  net4061;

wire  [0:47]  net3604;

wire  [0:47]  net4314;

wire  [0:23]  net3821;

wire  [0:47]  net3137;

wire  [0:23]  net4795;

wire  [0:47]  net3874;

wire  [0:7]  net2825;

wire  [0:47]  net3500;

wire  [0:7]  net2048;

wire  [0:47]  net3515;

wire  [0:23]  net2400;

wire  [0:23]  net4046;

wire  [0:47]  net4317;

wire  [0:47]  net4967;

wire  [0:23]  net2839;

wire  [0:7]  net4678;

wire  [0:23]  net4953;

wire  [0:23]  net2614;

wire  [0:23]  net2148;

wire  [0:47]  net3625;

wire  [0:23]  net4374;

wire  [0:47]  net4199;

wire  [0:47]  net3598;

wire  [0:47]  net4806;

wire  [0:7]  net3898;

wire  [0:23]  net4213;

wire  [0:23]  net4799;

wire  [0:47]  net4804;

wire  [0:47]  net3300;

wire  [0:47]  net2699;

wire  [0:47]  net4605;

wire  [0:47]  net3516;

wire  [0:23]  net2776;

wire  [0:47]  net3873;

wire  [0:7]  net4385;

wire  [0:47]  net2460;

wire  [0:47]  net4359;

wire  [0:47]  net3628;

wire  [0:7]  net3804;

wire  [0:47]  net3186;

wire  [0:23]  net3557;

wire  [0:47]  net3465;

wire  [0:47]  net2950;

wire  [0:23]  net4473;

wire  [0:47]  net4480;

wire  [0:47]  net4526;

wire  [0:47]  net2810;

wire  [0:23]  net3884;

wire  [0:47]  net4690;

wire  [0:47]  net4329;

wire  [0:47]  net2461;

wire  [0:23]  net4376;

wire  [0:23]  net5023;

wire  [0:23]  net3886;

wire  [0:47]  net2350;

wire  [0:47]  net3875;

wire  [0:23]  net3104;

wire  [0:7]  net3800;

wire  [0:7]  net3572;

wire  [0:7]  net2438;

wire  [0:47]  net3023;

wire  [0:7]  net3315;

wire  [0:47]  net3602;

wire  [0:23]  net3720;

wire  [0:47]  net4419;

wire  [0:7]  net2432;

wire  [0:7]  net4350;

wire  [0:7]  net4387;

wire  [0:23]  net2064;

wire  [0:47]  net2347;

wire  [0:7]  net3863;

wire  [0:7]  net3374;

wire  [0:47]  net3439;

wire  [0:47]  net4966;

wire  [0:47]  net2974;

wire  [0:23]  net3072;

wire  [0:7]  net2755;

wire  [0:47]  net4362;

wire  [0:23]  net2745;

wire  [0:7]  net5004;

wire  [0:7]  net3964;

wire  [0:47]  net3792;

wire  [0:23]  net2183;

wire  [0:7]  net4289;

wire  [3:0]  slf_op_33_06;

wire  [3:0]  slf_op_33_05;

wire  [3:0]  slf_op_33_01;

wire  [0:7]  net2063;

wire  [3:0]  slf_op_33_02;

wire  [0:7]  net2101;

wire  [0:23]  net4895;

wire  [0:47]  net2647;

wire  [0:47]  net3955;

wire  [0:47]  net2355;

wire  [0:23]  net4698;

wire  [0:47]  net3024;

wire  [0:7]  net4224;

wire  [0:47]  net3676;

wire  [0:7]  net4290;

wire  [0:23]  net3812;

wire  [0:47]  net3627;

wire  [0:7]  net4614;

wire  [0:47]  net4315;

wire  [0:7]  net4126;

wire  [0:47]  net3544;

wire  [0:47]  net3385;

wire  [0:7]  net3476;

wire  [3:0]  slf_op_33_08;

wire  [3:0]  slf_op_33_12;

wire  [0:47]  net3840;

wire  [3:0]  slf_op_33_13;

wire  [0:23]  net3233;

wire  [0:23]  net3429;

wire  [0:47]  net3662;

wire  [0:47]  net4113;

wire  [0:7]  net2115;

wire  [0:23]  net3103;

wire  [0:23]  net3592;

wire  [3:0]  slf_op_33_03;

wire  [0:23]  net4371;

wire  [3:0]  slf_op_33_14;

wire  [3:0]  slf_op_33_07;

wire  [3:0]  slf_op_33_09;

wire  [3:0]  slf_op_33_10;

wire  [3:0]  slf_op_33_11;

wire  [3:0]  slf_op_33_04;

wire  [3:0]  slf_op_23_00;

wire  [3:0]  slf_op_33_15;

wire  [0:47]  net3546;

wire  [0:47]  net3760;

wire  [0:23]  net3332;

wire  [0:47]  net4036;

wire  [0:47]  net4491;

wire  [0:47]  net2895;

wire  [0:47]  net3711;

wire  [0:23]  net4469;

wire  [0:47]  net4167;

wire  [0:23]  net2907;

wire  [0:47]  net3114;

wire  [0:7]  net3417;

wire  [0:47]  net2358;

wire  [0:23]  net4790;

wire  [0:23]  net2405;

wire  [0:23]  net5027;

wire  [0:23]  net2403;

wire  [0:7]  net4619;

wire  [0:47]  net2860;

wire  [0:23]  net4373;

wire  [0:47]  net2082;

wire  [0:7]  net2131;

wire  [0:47]  net2649;

wire  [0:47]  net4745;

wire  [0:47]  net4901;

wire  [0:7]  net3641;

wire  [0:7]  net3371;

wire  [0:47]  net4200;

wire  [0:23]  net4569;

wire  [0:47]  net4495;

wire  [0:7]  net4884;

wire  [0:47]  net4201;

wire  [0:47]  net2897;

wire  [0:23]  net2172;

wire  [0:7]  net3474;

wire  [0:47]  net2847;

wire  [0:47]  net4688;

wire  [0:47]  net3434;

wire  [0:23]  net4896;

wire  [0:47]  net4930;



lowla_modified I308 ( .clk(tclk_mi), .min(net02093), .lao(net2304));
bram_bufferx4x6 I310 ( .in(sdi_pad), .out(net02093));
tckbufx16 I255 ( .in(tclk_mi), .out(tclk_o));
clk_colbuf8kx8 I346 ( .clko(clk_tree_drv[7:0]), .clki(glb_in[7:0]));
fabric_buf8k I303 ( .f_in(padin_r[27]), .f_out(padin_135));
fabric_buf8k I304 ( .f_in(net2230), .f_out(fabric_out_33_16));
fabric_buf8k I305 ( .f_in(net2237), .f_out(fabric_out_33_02));
fabric_buf8k I306 ( .f_in(net2236), .f_out(fabric_out_33_01));
preio_bot_r I_preio_bot_r ( .ceb_i(ceb_i),
     .tnr_op_32_00({slf_op_33_01[3], slf_op_33_01[2], slf_op_33_01[1],
     slf_op_33_01[0], slf_op_33_01[3], slf_op_33_01[2],
     slf_op_33_01[1], slf_op_33_01[0]}),
     .sp4_h_l_17_00(sp4_h_l_17_00[15:0]),
     .sp4_v_t_17_00(sp4_v_b_17_01[47:0]),
     .sp4_v_t_18_00(net2165[0:47]), .sp4_v_t_19_00(net2149[0:47]),
     .sp4_v_t_20_00(net2141[0:47]), .sp4_v_t_21_00(net2133[0:47]),
     .sp4_v_t_22_00(net2125[0:47]), .sp4_v_t_23_00(net2117[0:47]),
     .sp4_v_t_24_00(net2110[0:47]), .sp4_v_t_25_00(net2104[0:47]),
     .sp4_v_t_26_00(net2096[0:47]), .sp4_v_t_27_00(net2092[0:47]),
     .sp4_v_t_28_00(net2082[0:47]), .sp4_v_t_29_00(net2065[0:47]),
     .sp4_v_t_30_00(net2050[0:47]), .sp4_v_t_31_00(net2182[0:47]),
     .sp4_v_t_32_00(net2189[0:47]), .sp12_v_t_17_00(net2164[0:23]),
     .sp12_v_t_18_00(net2172[0:23]), .sp12_v_t_19_00(net2156[0:23]),
     .sp12_v_t_20_00(net2148[0:23]), .sp12_v_t_21_00(net2140[0:23]),
     .sp12_v_t_22_00(net2132[0:23]), .sp12_v_t_23_00(net2124[0:23]),
     .sp12_v_t_24_00(net2090[0:23]), .sp12_v_t_25_00(net2180[0:23]),
     .sp12_v_t_26_00(net2103[0:23]), .sp12_v_t_27_00(net2091[0:23]),
     .sp12_v_t_28_00(net2089[0:23]), .sp12_v_t_29_00(net2081[0:23]),
     .sp12_v_t_30_00(net2064[0:23]), .sp12_v_t_31_00(net2049[0:23]),
     .sp12_v_t_32_00(net2183[0:23]), .update_i(update_i),
     .lft_op_31_00(net2185[0:7]), .bl_31(bl[1671:1618]),
     .tclk_i(tclk_i), .spiout_b(spiout_b[63:32]),
     .spioeb_b(spioeb_b[63:32]), .shift_i(shift_i), .sdi(sdi),
     .r_i(r_i), .padin_b(padin_b[56:30]), .mode_i(mode_i),
     .slf_op_31_00(slf_op_31_00[3:0]), .glb_net_31(net2048[0:7]),
     .lft_op_30_00(net2047[0:7]), .bl_30(bl[1617:1564]),
     .hold_b_r(hold_b_r), .hiz_b_i(hiz_b_i),
     .end_of_startup_bot_r(end_of_startup_bot_r[31:16]),
     .bs_en_i(bs_en_i), .spi_ss_in_b(spi_ss_in_b[63:32]),
     .slf_op_32_00(slf_op_32_00[3:0]),
     .slf_op_30_00(slf_op_30_00[3:0]), .glb_net_30(net2063[0:7]),
     .lft_op_29_00(net2062[0:7]), .bl_29(bl[1563:1510]),
     .sdo_pad(sdo_pad), .pado_b(pado_b[56:30]), .padin_81(padin_81),
     .padeb_b(padeb_b[56:30]), .slf_op_29_00(slf_op_29_00[3:0]),
     .glb_net_29(net2075[0:7]), .fabric_out_32_00(fabric_out_32_00),
     .fabric_out_18_00(fabric_out_18_00),
     .fabric_out_17_00(fabric_out_17_00), .cf_b(cf_b[383:0]),
     .pgate_r({pgate_r[1], pgate_r[0], pgate_r[2], pgate_r[3],
     pgate_r[5], pgate_r[4], pgate_r[6], pgate_r[7], pgate_r[9],
     pgate_r[8], pgate_r[10], pgate_r[11], pgate_r[13], pgate_r[12],
     pgate_r[14], pgate_r[15]}), .lft_op_28_00(net2074[0:7]),
     .bl_28(bl[1509:1456]), .slf_op_28_00(slf_op_28_00[3:0]),
     .glb_net_28(net2088[0:7]), .lft_op_27_00(net2087[0:7]),
     .bl_27(bl[1455:1402]), .lft_op_26_00(net2177[0:7]),
     .bl_26(bl[1401:1348]), .slf_op_26_00(slf_op_26_00[3:0]),
     .glb_net_26(net2102[0:7]), .lft_op_25_00(net2101[0:7]),
     .slf_op_25_00(slf_op_25_00[3:0]), .glb_net_25(net2109[0:7]),
     .lft_op_24_00(net2108[0:7]), .bl_24(bl[1305:1252]),
     .slf_op_24_00(slf_op_24_00[3:0]), .glb_net_24(net2116[0:7]),
     .lft_op_23_00(net2115[0:7]), .bl_23(bl[1251:1198]),
     .slf_op_23_00(slf_op_23_00[3:0]), .glb_net_23(net2123[0:7]),
     .lft_op_22_00(net2122[0:7]), .bl_22(bl[1197:1144]),
     .slf_op_22_00(slf_op_22_00[3:0]), .glb_net_22(net2131[0:7]),
     .lft_op_21_00(net2130[0:7]), .bl_21(bl[1143:1090]),
     .slf_op_21_00(slf_op_21_00[3:0]), .glb_net_21(net2139[0:7]),
     .lft_op_20_00(net2138[0:7]), .bl_20(bl[1089:1036]),
     .slf_op_20_00(slf_op_20_00[3:0]), .glb_net_20(net2147[0:7]),
     .lft_op_19_00(net2146[0:7]), .bl_19(bl[1035:982]),
     .slf_op_19_00(slf_op_19_00[3:0]), .glb_net_19(net2155[0:7]),
     .lft_op_17_00(slf_op_17_01[7:0]), .bl_17(bl[927:874]),
     .slf_op_17_00(slf_op_17_00[3:0]),
     .tnl_op_17_00(lft_op_17_01[7:0]), .glb_net_17(net2163[0:7]),
     .prog(prog), .lft_op_18_00(net2154[0:7]),
     .slf_op_18_00(slf_op_18_00[3:0]), .glb_net_18(net2171[0:7]),
     .bl_18(bl[981:928]), .wl_r({wl_r[1], wl_r[0], wl_r[2], wl_r[3],
     wl_r[5], wl_r[4], wl_r[6], wl_r[7], wl_r[9], wl_r[8], wl_r[10],
     wl_r[11], wl_r[13], wl_r[12], wl_r[14], wl_r[15]}),
     .slf_op_27_00(slf_op_27_00[3:0]), .glb_net_27(net2178[0:7]),
     .vdd_cntl_r({vdd_cntl_r[1], vdd_cntl_r[0], vdd_cntl_r[2],
     vdd_cntl_r[3], vdd_cntl_r[5], vdd_cntl_r[4], vdd_cntl_r[6],
     vdd_cntl_r[7], vdd_cntl_r[9], vdd_cntl_r[8], vdd_cntl_r[10],
     vdd_cntl_r[11], vdd_cntl_r[13], vdd_cntl_r[12], vdd_cntl_r[14],
     vdd_cntl_r[15]}), .reset_r({reset_r[1], reset_r[0], reset_r[2],
     reset_r[3], reset_r[5], reset_r[4], reset_r[6], reset_r[7],
     reset_r[9], reset_r[8], reset_r[10], reset_r[11], reset_r[13],
     reset_r[12], reset_r[14], reset_r[15]}),
     .glb_net_32(net2184[0:7]), .bl_32(bl[1725:1672]),
     .lft_op_32_00(net2188[0:7]), .bl_25(bl[1347:1306]),
     .sp4_h_r_32_00(net2191[0:15]));
array_RGT_IO_1x16 I_io_33bot ( .ceb(ceb_o), .padin(padin_r[27:0]),
     .padeb(padeb_r[27:0]), .pado(pado_r[27:0]), .cf_r(cf_r[383:0]),
     .bnl_op_01({slf_op_32_00[3], slf_op_32_00[2], slf_op_32_00[1],
     slf_op_32_00[0], slf_op_32_00[3], slf_op_32_00[2],
     slf_op_32_00[1], slf_op_32_00[0]}), .tnl_op_16(tnl_op_33_16[7:0]),
     .lft_op_16(slf_op_32_16[7:0]), .lft_op_15(net3860[0:7]),
     .lft_op_14(net3859[0:7]), .lft_op_13(net3862[0:7]),
     .lft_op_12(net3861[0:7]), .lft_op_11(net3863[0:7]),
     .lft_op_09(net3800[0:7]), .lft_op_10(net3799[0:7]),
     .lft_op_08(net3801[0:7]), .lft_op_07(net3802[0:7]),
     .lft_op_06(net3803[0:7]), .lft_op_04(net3743[0:7]),
     .lft_op_05(net3804[0:7]), .lft_op_01(net2188[0:7]),
     .lft_op_02(net3735[0:7]), .lft_op_03(net3733[0:7]),
     .fabric_out_16(net2230), .fabric_out_15(net2527),
     .fabric_out_14(net2523), .fabric_out_13(net2525),
     .fabric_out_12(net2522), .fabric_out_11(net2571),
     .fabric_out_01(net2236), .fabric_out_02(net2237),
     .fabric_out_03(net2521), .fabric_out_04(net2581),
     .fabric_out_05(net2524), .fabric_out_06(net2526),
     .fabric_out_07(net2558), .fabric_out_08(net2520),
     .fabric_out_09(net2570), .fabric_out_10(net2582),
     .slf_op_16(slf_op_33_16[3:0]), .slf_op_12(slf_op_33_12[3:0]),
     .sp4_v_t_16(sp4_v_t_33_16[15:0]), .reset_b(reset_r[271:16]),
     .slf_op_11(slf_op_33_11[3:0]), .slf_op_09(slf_op_33_09[3:0]),
     .slf_op_08(slf_op_33_08[3:0]), .slf_op_06(slf_op_33_06[3:0]),
     .slf_op_05(slf_op_33_05[3:0]), .SP12_h_l_01(net3104[0:23]),
     .slf_op_10(slf_op_33_10[3:0]), .slf_op_07(slf_op_33_07[3:0]),
     .slf_op_04(slf_op_33_04[3:0]), .wl(wl_r[271:16]),
     .SP4_h_l_06(net3139[0:47]), .SP4_h_l_07(net3138[0:47]),
     .SP4_h_l_04(net2585[0:47]), .SP4_h_l_05(net3140[0:47]),
     .SP4_h_l_02(net3114[0:47]), .SP4_h_l_03(net2583[0:47]),
     .sp4_v_b_01(net2191[0:15]), .slf_op_02(slf_op_33_02[3:0]),
     .slf_op_03(slf_op_33_03[3:0]), .pgate(pgate_r[271:16]),
     .SP12_h_l_16(net3230[0:23]), .SP12_h_l_15(net3232[0:23]),
     .SP12_h_l_14(net3231[0:23]), .SP12_h_l_13(net3234[0:23]),
     .SP12_h_l_12(net3233[0:23]), .SP12_h_l_11(net3235[0:23]),
     .SP12_h_l_10(net3160[0:23]), .SP12_h_l_09(net3169[0:23]),
     .SP12_h_l_08(net3168[0:23]), .SP12_h_l_07(net3167[0:23]),
     .SP12_h_l_06(net3166[0:23]), .SP12_h_l_05(net3165[0:23]),
     .SP12_h_l_04(net3101[0:23]), .SP12_h_l_03(net3102[0:23]),
     .SP12_h_l_02(net3103[0:23]), .slf_op_01(slf_op_33_01[3:0]),
     .SP4_h_l_16(net3191[0:47]), .cdone_in(end_of_startup_rgt_b[16:1]),
     .slf_op_13(slf_op_33_13[3:0]), .slf_op_14(slf_op_33_14[3:0]),
     .slf_op_15(slf_op_33_15[3:0]), .SP4_h_l_15(net3190[0:47]),
     .SP4_h_l_14(net3189[0:47]), .SP4_h_l_13(net3188[0:47]),
     .SP4_h_l_12(net3187[0:47]), .SP4_h_l_11(net3186[0:47]),
     .SP4_h_l_10(net3135[0:47]), .SP4_h_l_09(net3136[0:47]),
     .SP4_h_l_08(net3137[0:47]), .SP4_h_l_01(net3115[0:47]),
     .vdd_cntl(vdd_cntl_r[271:16]), .shift(shift_o), .bs_en(bs_en_o),
     .mode(mode_o), .sdi(net2304), .hiz_b(hiz_b_o), .prog(prog),
     .hold(hold_r_b), .update(update_o),
     .glb_netwk_col(clk_tree_drv[7:0]), .r(r_o),
     .spi_ss_in_b(spi_ss_in_r[31:0]), .sdo(sdo), .bl(bl[1743:1726]),
     .tclk(tclk_o), .spioeb(spioeb_r[31:0]), .spiout(spiout_r[31:0]));
array_BRAM_1x8bot I_bram_25_bot ( .glb_netwk(net2109[0:7]),
     .wl(wl_r[271:16]), .pgate(pgate_r[271:16]),
     .vdd_cntl(vdd_cntl_r[271:16]), .reset_b(reset_r[271:16]),
     .bm_sclkrw_i(bm_sclkrw_i[1:0]), .bm_sdi_i(bm_sdi_i[1:0]),
     .bm_sweb_i(bm_sweb_i[1:0]), .bm_sdo_o(bm_sdo_o[1:0]),
     .bm_sweb_o(bm_sweb_o[1:0]), .bm_sdi_o(bm_sdi_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_o[1:0]), .bm_sdo_i(bm_sdo_i[1:0]),
     .sp12_h_r_01(net2329[0:23]), .lft_op_10(net4125[0:7]),
     .sp4_h_l_04(net3601[0:47]), .sp4_h_l_06(net3628[0:47]),
     .lft_op_09(net4126[0:7]), .lft_op_08(net4127[0:7]),
     .lft_op_06(net4129[0:7]), .lft_op_07(net4128[0:7]),
     .lft_op_05(net4130[0:7]), .lft_op_03(net4059[0:7]),
     .lft_op_04(net4069[0:7]), .lft_op_02(net4061[0:7]),
     .sp4_h_r_09(net2341[0:47]), .bnr_op_01({slf_op_26_00[3],
     slf_op_26_00[2], slf_op_26_00[1], slf_op_26_00[0],
     slf_op_26_00[3], slf_op_26_00[2], slf_op_26_00[1],
     slf_op_26_00[0]}), .sp4_r_v_b_01(net2096[0:47]),
     .sp4_r_v_b_02(net2344[0:47]), .sp4_r_v_b_03(net2345[0:47]),
     .sp4_r_v_b_04(net2346[0:47]), .sp4_r_v_b_05(net2347[0:47]),
     .sp4_r_v_b_06(net2348[0:47]), .sp4_r_v_b_07(net2349[0:47]),
     .sp4_r_v_b_08(net2350[0:47]), .sp4_r_v_b_09(net2351[0:47]),
     .sp4_r_v_b_10(net2352[0:47]), .sp4_r_v_b_11(net2353[0:47]),
     .sp4_r_v_b_12(net2354[0:47]), .sp4_r_v_b_13(net2355[0:47]),
     .sp4_r_v_b_14(net2356[0:47]), .sp4_r_v_b_16(net2357[0:47]),
     .sp4_r_v_b_15(net2358[0:47]), .bnl_op_01({slf_op_24_00[3],
     slf_op_24_00[2], slf_op_24_00[1], slf_op_24_00[0],
     slf_op_24_00[3], slf_op_24_00[2], slf_op_24_00[1],
     slf_op_24_00[0]}), .lft_op_01(net2108[0:7]),
     .bot_op_01({slf_op_25_00[3], slf_op_25_00[2], slf_op_25_00[1],
     slf_op_25_00[0], slf_op_25_00[3], slf_op_25_00[2],
     slf_op_25_00[1], slf_op_25_00[0]}), .sp12_v_b_01(net2180[0:23]),
     .sp4_v_b_16(net3707[0:47]), .sp4_v_b_15(net3708[0:47]),
     .sp4_v_b_14(net3710[0:47]), .sp4_v_b_13(net3709[0:47]),
     .sp4_v_b_12(net3711[0:47]), .sp4_v_b_11(net3712[0:47]),
     .sp4_v_b_10(net3665[0:47]), .sp4_v_b_09(net3664[0:47]),
     .sp4_v_b_08(net3663[0:47]), .sp4_v_b_07(net3662[0:47]),
     .sp4_v_b_06(net3661[0:47]), .sp4_v_b_05(net3660[0:47]),
     .sp4_v_b_04(net3597[0:47]), .sp4_v_b_03(net3598[0:47]),
     .sp4_v_b_02(net3599[0:47]), .sp4_v_b_01(net2104[0:47]),
     .sp12_h_l_10(net3649[0:23]), .sp12_h_l_09(net3658[0:23]),
     .sp12_h_l_08(net3657[0:23]), .sp12_h_l_07(net3656[0:23]),
     .sp12_h_l_06(net3655[0:23]), .sp12_h_l_05(net3654[0:23]),
     .sp12_h_l_04(net3590[0:23]), .sp12_h_l_03(net3591[0:23]),
     .sp12_h_l_02(net3592[0:23]), .sp12_h_l_01(net3593[0:23]),
     .sp12_h_r_10(net2389[0:23]), .sp12_h_r_15(net2390[0:23]),
     .sp12_h_l_15(net3721[0:23]), .sp12_h_l_14(net3720[0:23]),
     .sp12_h_r_14(net2393[0:23]), .sp12_h_r_16(net2394[0:23]),
     .sp12_h_l_16(net3719[0:23]), .sp12_h_l_13(net3723[0:23]),
     .sp12_h_l_12(net3722[0:23]), .sp12_h_l_11(net3724[0:23]),
     .sp12_h_r_13(net2399[0:23]), .sp12_h_r_12(net2400[0:23]),
     .sp12_h_r_11(net2401[0:23]), .sp12_h_r_09(net2402[0:23]),
     .sp12_h_r_08(net2403[0:23]), .sp12_h_r_07(net2404[0:23]),
     .sp12_h_r_06(net2405[0:23]), .sp12_h_r_05(net2406[0:23]),
     .sp12_h_r_04(net2407[0:23]), .sp12_h_r_03(net2408[0:23]),
     .sp12_h_r_02(net2409[0:23]), .lft_op_14(net4185[0:7]),
     .lft_op_13(net4188[0:7]), .lft_op_12(net4187[0:7]),
     .lft_op_11(net4189[0:7]), .lft_op_15(net4186[0:7]),
     .slf_op_15(net3697[0:7]), .slf_op_14(net3696[0:7]),
     .slf_op_13(net3699[0:7]), .slf_op_12(net3698[0:7]),
     .slf_op_11(net3700[0:7]), .slf_op_10(net3636[0:7]),
     .slf_op_09(net3637[0:7]), .slf_op_08(net3638[0:7]),
     .slf_op_07(net3639[0:7]), .slf_op_06(net3640[0:7]),
     .slf_op_05(net3641[0:7]), .slf_op_04(net3580[0:7]),
     .slf_op_03(net3570[0:7]), .slf_op_01(net2101[0:7]),
     .slf_op_02(net3572[0:7]), .rgt_op_01(net2177[0:7]),
     .rgt_op_02(net2431[0:7]), .rgt_op_03(net2432[0:7]),
     .rgt_op_04(net2433[0:7]), .rgt_op_05(net2434[0:7]),
     .rgt_op_06(net2435[0:7]), .rgt_op_07(net2436[0:7]),
     .rgt_op_08(net2437[0:7]), .rgt_op_09(net2438[0:7]),
     .rgt_op_10(net2439[0:7]), .rgt_op_11(net2440[0:7]),
     .rgt_op_12(net2441[0:7]), .rgt_op_13(net2442[0:7]),
     .rgt_op_14(net2443[0:7]), .rgt_op_15(net2444[0:7]),
     .sp4_h_l_05(net3629[0:47]), .sp4_h_l_02(net3603[0:47]),
     .sp4_h_l_03(net3602[0:47]), .sp4_h_l_01(net3604[0:47]),
     .sp4_h_r_01(net2449[0:47]), .sp4_h_r_02(net2450[0:47]),
     .sp4_h_r_03(net2451[0:47]), .sp4_h_r_04(net2452[0:47]),
     .sp4_h_r_05(net2453[0:47]), .sp4_h_r_06(net2454[0:47]),
     .sp4_h_r_07(net2455[0:47]), .sp4_h_r_08(net2456[0:47]),
     .sp4_h_r_10(net2457[0:47]), .sp4_h_r_11(net2458[0:47]),
     .sp4_h_r_12(net2459[0:47]), .sp4_h_r_13(net2460[0:47]),
     .sp4_h_r_14(net2461[0:47]), .sp4_h_r_15(net2462[0:47]),
     .sp4_h_r_16(net2463[0:47]), .lft_op_16(slf_op_24_16[7:0]),
     .tnl_op_16(tnl_op_25_16[7:0]), .sp4_v_t_16(sp4_v_t_25_16[47:0]),
     .top_op_16(top_op_25_16[7:0]), .slf_op_16(slf_op_25_16[7:0]),
     .tnr_op_16(tnr_op_25_16[7:0]), .sp12_v_t_16(sp12_v_t_25_16[23:0]),
     .rgt_op_16(slf_op_26_16[7:0]), .sp4_h_l_16(net3680[0:47]),
     .sp4_h_l_14(net3678[0:47]), .sp4_h_l_15(net3679[0:47]),
     .sp4_h_l_13(net3677[0:47]), .sp4_h_l_12(net3676[0:47]),
     .sp4_h_l_11(net3675[0:47]), .sp4_h_l_10(net3624[0:47]),
     .sp4_h_l_09(net3625[0:47]), .sp4_h_l_08(net3626[0:47]),
     .sp4_h_l_07(net3627[0:47]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_sreb_o(bm_sreb_o), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .bl(bl[1347:1306]), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]));
array_LT1x16 I_lt_21_bot ( .sp12_v_b_01(net2140[0:23]),
     .glb_netwk(net2139[0:7]), .sp12_v_t_16(sp12_v_t_21_16[23:0]),
     .rgt_op_16(slf_op_22_16[7:0]), .top_op_16(top_op_21_16[7:0]),
     .rgt_op_03(net2592[0:7]), .slf_op_02(net4876[0:7]),
     .rgt_op_02(net2594[0:7]), .rgt_op_01(net2122[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3417[0:7]), .lft_op_03(net3407[0:7]),
     .lft_op_02(net3409[0:7]), .lft_op_01(net2138[0:7]),
     .rgt_op_04(net2602[0:7]), .carry_in(net2519),
     .bnl_op_01({slf_op_20_00[3], slf_op_20_00[2], slf_op_20_00[1],
     slf_op_20_00[0], slf_op_20_00[3], slf_op_20_00[2],
     slf_op_20_00[1], slf_op_20_00[0]}), .slf_op_04(net4884[0:7]),
     .slf_op_03(net4874[0:7]), .slf_op_01(net2130[0:7]),
     .sp4_h_l_04(net4905[0:47]), .carry_out(carry_out_21_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net2612[0:23]),
     .sp12_h_r_03(net2613[0:23]), .sp12_h_r_02(net2614[0:23]),
     .sp12_h_r_01(net2615[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_21_16[7:0]), .sp4_v_b_01(net2133[0:47]),
     .sp4_r_v_b_04(net2619[0:47]), .sp4_r_v_b_03(net2620[0:47]),
     .sp4_r_v_b_02(net2621[0:47]), .sp4_r_v_b_01(net2125[0:47]),
     .sp4_h_r_04(net2623[0:47]), .sp4_h_r_03(net2624[0:47]),
     .sp4_h_r_02(net2625[0:47]), .sp4_h_r_01(net2626[0:47]),
     .sp4_h_l_03(net4906[0:47]), .sp4_h_l_02(net4907[0:47]),
     .sp4_h_l_01(net4908[0:47]), .bl(bl[1143:1090]),
     .bot_op_01({slf_op_21_00[3], slf_op_21_00[2], slf_op_21_00[1],
     slf_op_21_00[0], slf_op_21_00[3], slf_op_21_00[2],
     slf_op_21_00[1], slf_op_21_00[0]}), .sp12_h_l_01(net4897[0:23]),
     .sp12_h_l_02(net4896[0:23]), .sp12_h_l_03(net4895[0:23]),
     .sp12_h_l_04(net4894[0:23]), .sp4_v_b_04(net4901[0:47]),
     .sp4_v_b_03(net4902[0:47]), .sp4_v_b_02(net4903[0:47]),
     .bnr_op_01({slf_op_22_00[3], slf_op_22_00[2], slf_op_22_00[1],
     slf_op_22_00[0], slf_op_22_00[3], slf_op_22_00[2],
     slf_op_22_00[1], slf_op_22_00[0]}), .sp4_h_l_05(net4933[0:47]),
     .sp4_h_l_06(net4932[0:47]), .sp4_h_l_07(net4931[0:47]),
     .sp4_h_l_08(net4930[0:47]), .sp4_h_l_09(net4929[0:47]),
     .sp4_h_l_10(net4928[0:47]), .sp4_h_r_10(net2646[0:47]),
     .sp4_h_r_09(net2647[0:47]), .sp4_h_r_08(net2648[0:47]),
     .sp4_h_r_07(net2649[0:47]), .sp4_h_r_06(net2650[0:47]),
     .sp4_h_r_05(net2651[0:47]), .slf_op_05(net4945[0:7]),
     .slf_op_06(net4944[0:7]), .slf_op_07(net4943[0:7]),
     .slf_op_08(net4942[0:7]), .slf_op_09(net4941[0:7]),
     .slf_op_10(net4940[0:7]), .rgt_op_10(net2658[0:7]),
     .rgt_op_09(net2659[0:7]), .rgt_op_08(net2660[0:7]),
     .rgt_op_07(net2661[0:7]), .rgt_op_06(net2662[0:7]),
     .rgt_op_05(net2663[0:7]), .lft_op_10(net3473[0:7]),
     .lft_op_09(net3474[0:7]), .lft_op_08(net3475[0:7]),
     .lft_op_07(net3476[0:7]), .lft_op_06(net3477[0:7]),
     .lft_op_05(net3478[0:7]), .sp12_h_l_10(net4953[0:23]),
     .sp12_h_r_10(net2671[0:23]), .sp12_h_l_09(net4962[0:23]),
     .sp12_h_l_08(net4961[0:23]), .sp12_h_l_07(net4960[0:23]),
     .sp12_h_l_06(net4959[0:23]), .sp12_h_r_05(net2676[0:23]),
     .sp12_h_r_06(net2677[0:23]), .sp12_h_r_07(net2678[0:23]),
     .sp12_h_r_08(net2679[0:23]), .sp12_h_r_09(net2680[0:23]),
     .sp12_h_l_05(net4958[0:23]), .sp4_r_v_b_05(net2682[0:47]),
     .sp4_r_v_b_06(net2683[0:47]), .sp4_r_v_b_07(net2684[0:47]),
     .sp4_r_v_b_08(net2685[0:47]), .sp4_r_v_b_09(net2686[0:47]),
     .sp4_r_v_b_10(net2687[0:47]), .sp4_v_b_10(net4969[0:47]),
     .sp4_v_b_09(net4968[0:47]), .sp4_v_b_08(net4967[0:47]),
     .sp4_v_b_07(net4966[0:47]), .sp4_v_b_06(net4965[0:47]),
     .sp4_v_b_05(net4964[0:47]), .sp4_v_t_16(sp4_v_t_21_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net2697[0:47]), .sp4_h_r_12(net2698[0:47]),
     .sp4_h_r_13(net2699[0:47]), .sp4_h_r_14(net2700[0:47]),
     .sp4_h_r_15(net2701[0:47]), .sp4_h_r_16(net2702[0:47]),
     .sp4_h_l_16(sp4_h_r_20_21[47:0]), .sp4_h_l_15(net4983[0:47]),
     .sp4_h_l_14(net4982[0:47]), .sp4_h_l_13(net4981[0:47]),
     .sp4_h_l_12(net4980[0:47]), .sp4_h_l_11(net4979[0:47]),
     .tnr_op_16(tnr_op_21_16[7:0]), .tnl_op_16(tnl_op_21_16[7:0]),
     .lft_op_16(slf_op_20_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net5001[0:7]), .slf_op_14(net5000[0:7]),
     .slf_op_13(net5003[0:7]), .slf_op_12(net5002[0:7]),
     .slf_op_11(net5004[0:7]), .rgt_op_14(net2718[0:7]),
     .rgt_op_15(net2719[0:7]), .rgt_op_12(net2720[0:7]),
     .rgt_op_13(net2721[0:7]), .rgt_op_11(net2722[0:7]),
     .sp4_v_b_16(net5011[0:47]), .sp4_v_b_14(net5014[0:47]),
     .sp4_v_b_15(net5012[0:47]), .sp4_v_b_13(net5013[0:47]),
     .sp4_v_b_11(net5016[0:47]), .sp4_v_b_12(net5015[0:47]),
     .sp4_r_v_b_16(net2729[0:47]), .sp4_r_v_b_15(net2730[0:47]),
     .sp4_r_v_b_13(net2731[0:47]), .sp4_r_v_b_14(net2732[0:47]),
     .sp4_r_v_b_12(net2733[0:47]), .sp4_r_v_b_11(net2734[0:47]),
     .sp12_h_l_16(net5023[0:23]), .sp12_h_l_15(net5025[0:23]),
     .sp12_h_l_14(net5024[0:23]), .sp12_h_l_13(net5027[0:23]),
     .sp12_h_l_12(net5026[0:23]), .sp12_h_l_11(net5028[0:23]),
     .sp12_h_r_16(net2741[0:23]), .sp12_h_r_14(net2742[0:23]),
     .sp12_h_r_15(net2743[0:23]), .sp12_h_r_12(net2744[0:23]),
     .sp12_h_r_13(net2745[0:23]), .sp12_h_r_11(net2746[0:23]),
     .lft_op_14(net3533[0:7]), .lft_op_15(net3534[0:7]),
     .lft_op_12(net3535[0:7]), .lft_op_11(net3537[0:7]),
     .lft_op_13(net3536[0:7]));
array_LT1x16 I_lt_28_bot ( .sp12_v_b_01(net2089[0:23]),
     .glb_netwk(net2088[0:7]), .sp12_v_t_16(sp12_v_t_28_16[23:0]),
     .rgt_op_16(slf_op_29_16[7:0]), .top_op_16(top_op_28_16[7:0]),
     .rgt_op_03(net2755[0:7]), .slf_op_02(net2920[0:7]),
     .rgt_op_02(net2757[0:7]), .rgt_op_01(net2062[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4395[0:7]), .lft_op_03(net4385[0:7]),
     .lft_op_02(net4387[0:7]), .lft_op_01(net2087[0:7]),
     .rgt_op_04(net2765[0:7]), .carry_in(net2555),
     .bnl_op_01({slf_op_27_00[3], slf_op_27_00[2], slf_op_27_00[1],
     slf_op_27_00[0], slf_op_27_00[3], slf_op_27_00[2],
     slf_op_27_00[1], slf_op_27_00[0]}), .slf_op_04(net2928[0:7]),
     .slf_op_03(net2918[0:7]), .slf_op_01(net2074[0:7]),
     .sp4_h_l_04(net2949[0:47]), .carry_out(carry_out_28_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net2775[0:23]),
     .sp12_h_r_03(net2776[0:23]), .sp12_h_r_02(net2777[0:23]),
     .sp12_h_r_01(net2778[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_28_16[7:0]), .sp4_v_b_01(net2082[0:47]),
     .sp4_r_v_b_04(net2782[0:47]), .sp4_r_v_b_03(net2783[0:47]),
     .sp4_r_v_b_02(net2784[0:47]), .sp4_r_v_b_01(net2065[0:47]),
     .sp4_h_r_04(net2786[0:47]), .sp4_h_r_03(net2787[0:47]),
     .sp4_h_r_02(net2788[0:47]), .sp4_h_r_01(net2789[0:47]),
     .sp4_h_l_03(net2950[0:47]), .sp4_h_l_02(net2951[0:47]),
     .sp4_h_l_01(net2952[0:47]), .bl(bl[1509:1456]),
     .bot_op_01({slf_op_28_00[3], slf_op_28_00[2], slf_op_28_00[1],
     slf_op_28_00[0], slf_op_28_00[3], slf_op_28_00[2],
     slf_op_28_00[1], slf_op_28_00[0]}), .sp12_h_l_01(net2941[0:23]),
     .sp12_h_l_02(net2940[0:23]), .sp12_h_l_03(net2939[0:23]),
     .sp12_h_l_04(net2938[0:23]), .sp4_v_b_04(net2945[0:47]),
     .sp4_v_b_03(net2946[0:47]), .sp4_v_b_02(net2947[0:47]),
     .bnr_op_01({slf_op_29_00[3], slf_op_29_00[2], slf_op_29_00[1],
     slf_op_29_00[0], slf_op_29_00[3], slf_op_29_00[2],
     slf_op_29_00[1], slf_op_29_00[0]}), .sp4_h_l_05(net2977[0:47]),
     .sp4_h_l_06(net2976[0:47]), .sp4_h_l_07(net2975[0:47]),
     .sp4_h_l_08(net2974[0:47]), .sp4_h_l_09(net2973[0:47]),
     .sp4_h_l_10(net2972[0:47]), .sp4_h_r_10(net2809[0:47]),
     .sp4_h_r_09(net2810[0:47]), .sp4_h_r_08(net2811[0:47]),
     .sp4_h_r_07(net2812[0:47]), .sp4_h_r_06(net2813[0:47]),
     .sp4_h_r_05(net2814[0:47]), .slf_op_05(net2989[0:7]),
     .slf_op_06(net2988[0:7]), .slf_op_07(net2987[0:7]),
     .slf_op_08(net2986[0:7]), .slf_op_09(net2985[0:7]),
     .slf_op_10(net2984[0:7]), .rgt_op_10(net2821[0:7]),
     .rgt_op_09(net2822[0:7]), .rgt_op_08(net2823[0:7]),
     .rgt_op_07(net2824[0:7]), .rgt_op_06(net2825[0:7]),
     .rgt_op_05(net2826[0:7]), .lft_op_10(net4451[0:7]),
     .lft_op_09(net4452[0:7]), .lft_op_08(net4453[0:7]),
     .lft_op_07(net4454[0:7]), .lft_op_06(net4455[0:7]),
     .lft_op_05(net4456[0:7]), .sp12_h_l_10(net2997[0:23]),
     .sp12_h_r_10(net2834[0:23]), .sp12_h_l_09(net3006[0:23]),
     .sp12_h_l_08(net3005[0:23]), .sp12_h_l_07(net3004[0:23]),
     .sp12_h_l_06(net3003[0:23]), .sp12_h_r_05(net2839[0:23]),
     .sp12_h_r_06(net2840[0:23]), .sp12_h_r_07(net2841[0:23]),
     .sp12_h_r_08(net2842[0:23]), .sp12_h_r_09(net2843[0:23]),
     .sp12_h_l_05(net3002[0:23]), .sp4_r_v_b_05(net2845[0:47]),
     .sp4_r_v_b_06(net2846[0:47]), .sp4_r_v_b_07(net2847[0:47]),
     .sp4_r_v_b_08(net2848[0:47]), .sp4_r_v_b_09(net2849[0:47]),
     .sp4_r_v_b_10(net2850[0:47]), .sp4_v_b_10(net3013[0:47]),
     .sp4_v_b_09(net3012[0:47]), .sp4_v_b_08(net3011[0:47]),
     .sp4_v_b_07(net3010[0:47]), .sp4_v_b_06(net3009[0:47]),
     .sp4_v_b_05(net3008[0:47]), .sp4_v_t_16(sp4_v_t_28_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net2860[0:47]), .sp4_h_r_12(net2861[0:47]),
     .sp4_h_r_13(net2862[0:47]), .sp4_h_r_14(net2863[0:47]),
     .sp4_h_r_15(net2864[0:47]), .sp4_h_r_16(net2865[0:47]),
     .sp4_h_l_16(net3028[0:47]), .sp4_h_l_15(net3027[0:47]),
     .sp4_h_l_14(net3026[0:47]), .sp4_h_l_13(net3025[0:47]),
     .sp4_h_l_12(net3024[0:47]), .sp4_h_l_11(net3023[0:47]),
     .tnr_op_16(tnr_op_28_16[7:0]), .tnl_op_16(tnl_op_28_16[7:0]),
     .lft_op_16(slf_op_27_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net3045[0:7]), .slf_op_14(net3044[0:7]),
     .slf_op_13(net3047[0:7]), .slf_op_12(net3046[0:7]),
     .slf_op_11(net3048[0:7]), .rgt_op_14(net2881[0:7]),
     .rgt_op_15(net2882[0:7]), .rgt_op_12(net2883[0:7]),
     .rgt_op_13(net2884[0:7]), .rgt_op_11(net2885[0:7]),
     .sp4_v_b_16(net3055[0:47]), .sp4_v_b_14(net3058[0:47]),
     .sp4_v_b_15(net3056[0:47]), .sp4_v_b_13(net3057[0:47]),
     .sp4_v_b_11(net3060[0:47]), .sp4_v_b_12(net3059[0:47]),
     .sp4_r_v_b_16(net2892[0:47]), .sp4_r_v_b_15(net2893[0:47]),
     .sp4_r_v_b_13(net2894[0:47]), .sp4_r_v_b_14(net2895[0:47]),
     .sp4_r_v_b_12(net2896[0:47]), .sp4_r_v_b_11(net2897[0:47]),
     .sp12_h_l_16(net3067[0:23]), .sp12_h_l_15(net3069[0:23]),
     .sp12_h_l_14(net3068[0:23]), .sp12_h_l_13(net3071[0:23]),
     .sp12_h_l_12(net3070[0:23]), .sp12_h_l_11(net3072[0:23]),
     .sp12_h_r_16(net2904[0:23]), .sp12_h_r_14(net2905[0:23]),
     .sp12_h_r_15(net2906[0:23]), .sp12_h_r_12(net2907[0:23]),
     .sp12_h_r_13(net2908[0:23]), .sp12_h_r_11(net2909[0:23]),
     .lft_op_14(net4511[0:7]), .lft_op_15(net4512[0:7]),
     .lft_op_12(net4513[0:7]), .lft_op_11(net4515[0:7]),
     .lft_op_13(net4514[0:7]));
array_LT1x16 I_lt_27_bot ( .sp12_v_b_01(net2091[0:23]),
     .glb_netwk(net2178[0:7]), .sp12_v_t_16(sp12_v_t_27_16[23:0]),
     .rgt_op_16(slf_op_28_16[7:0]), .top_op_16(top_op_27_16[7:0]),
     .rgt_op_03(net2918[0:7]), .slf_op_02(net4387[0:7]),
     .rgt_op_02(net2920[0:7]), .rgt_op_01(net2074[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2433[0:7]), .lft_op_03(net2432[0:7]),
     .lft_op_02(net2431[0:7]), .lft_op_01(net2177[0:7]),
     .rgt_op_04(net2928[0:7]), .carry_in(net2517),
     .bnl_op_01({slf_op_26_00[3], slf_op_26_00[2], slf_op_26_00[1],
     slf_op_26_00[0], slf_op_26_00[3], slf_op_26_00[2],
     slf_op_26_00[1], slf_op_26_00[0]}), .slf_op_04(net4395[0:7]),
     .slf_op_03(net4385[0:7]), .slf_op_01(net2087[0:7]),
     .sp4_h_l_04(net4416[0:47]), .carry_out(carry_out_27_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net2938[0:23]),
     .sp12_h_r_03(net2939[0:23]), .sp12_h_r_02(net2940[0:23]),
     .sp12_h_r_01(net2941[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_27_16[7:0]), .sp4_v_b_01(net2092[0:47]),
     .sp4_r_v_b_04(net2945[0:47]), .sp4_r_v_b_03(net2946[0:47]),
     .sp4_r_v_b_02(net2947[0:47]), .sp4_r_v_b_01(net2082[0:47]),
     .sp4_h_r_04(net2949[0:47]), .sp4_h_r_03(net2950[0:47]),
     .sp4_h_r_02(net2951[0:47]), .sp4_h_r_01(net2952[0:47]),
     .sp4_h_l_03(net4417[0:47]), .sp4_h_l_02(net4418[0:47]),
     .sp4_h_l_01(net4419[0:47]), .bl(bl[1455:1402]),
     .bot_op_01({slf_op_27_00[3], slf_op_27_00[2], slf_op_27_00[1],
     slf_op_27_00[0], slf_op_27_00[3], slf_op_27_00[2],
     slf_op_27_00[1], slf_op_27_00[0]}), .sp12_h_l_01(net4408[0:23]),
     .sp12_h_l_02(net4407[0:23]), .sp12_h_l_03(net4406[0:23]),
     .sp12_h_l_04(net4405[0:23]), .sp4_v_b_04(net4412[0:47]),
     .sp4_v_b_03(net4413[0:47]), .sp4_v_b_02(net4414[0:47]),
     .bnr_op_01({slf_op_28_00[3], slf_op_28_00[2], slf_op_28_00[1],
     slf_op_28_00[0], slf_op_28_00[3], slf_op_28_00[2],
     slf_op_28_00[1], slf_op_28_00[0]}), .sp4_h_l_05(net4444[0:47]),
     .sp4_h_l_06(net4443[0:47]), .sp4_h_l_07(net4442[0:47]),
     .sp4_h_l_08(net4441[0:47]), .sp4_h_l_09(net4440[0:47]),
     .sp4_h_l_10(net4439[0:47]), .sp4_h_r_10(net2972[0:47]),
     .sp4_h_r_09(net2973[0:47]), .sp4_h_r_08(net2974[0:47]),
     .sp4_h_r_07(net2975[0:47]), .sp4_h_r_06(net2976[0:47]),
     .sp4_h_r_05(net2977[0:47]), .slf_op_05(net4456[0:7]),
     .slf_op_06(net4455[0:7]), .slf_op_07(net4454[0:7]),
     .slf_op_08(net4453[0:7]), .slf_op_09(net4452[0:7]),
     .slf_op_10(net4451[0:7]), .rgt_op_10(net2984[0:7]),
     .rgt_op_09(net2985[0:7]), .rgt_op_08(net2986[0:7]),
     .rgt_op_07(net2987[0:7]), .rgt_op_06(net2988[0:7]),
     .rgt_op_05(net2989[0:7]), .lft_op_10(net2439[0:7]),
     .lft_op_09(net2438[0:7]), .lft_op_08(net2437[0:7]),
     .lft_op_07(net2436[0:7]), .lft_op_06(net2435[0:7]),
     .lft_op_05(net2434[0:7]), .sp12_h_l_10(net4464[0:23]),
     .sp12_h_r_10(net2997[0:23]), .sp12_h_l_09(net4473[0:23]),
     .sp12_h_l_08(net4472[0:23]), .sp12_h_l_07(net4471[0:23]),
     .sp12_h_l_06(net4470[0:23]), .sp12_h_r_05(net3002[0:23]),
     .sp12_h_r_06(net3003[0:23]), .sp12_h_r_07(net3004[0:23]),
     .sp12_h_r_08(net3005[0:23]), .sp12_h_r_09(net3006[0:23]),
     .sp12_h_l_05(net4469[0:23]), .sp4_r_v_b_05(net3008[0:47]),
     .sp4_r_v_b_06(net3009[0:47]), .sp4_r_v_b_07(net3010[0:47]),
     .sp4_r_v_b_08(net3011[0:47]), .sp4_r_v_b_09(net3012[0:47]),
     .sp4_r_v_b_10(net3013[0:47]), .sp4_v_b_10(net4480[0:47]),
     .sp4_v_b_09(net4479[0:47]), .sp4_v_b_08(net4478[0:47]),
     .sp4_v_b_07(net4477[0:47]), .sp4_v_b_06(net4476[0:47]),
     .sp4_v_b_05(net4475[0:47]), .sp4_v_t_16(sp4_v_t_27_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net3023[0:47]), .sp4_h_r_12(net3024[0:47]),
     .sp4_h_r_13(net3025[0:47]), .sp4_h_r_14(net3026[0:47]),
     .sp4_h_r_15(net3027[0:47]), .sp4_h_r_16(net3028[0:47]),
     .sp4_h_l_16(net4495[0:47]), .sp4_h_l_15(net4494[0:47]),
     .sp4_h_l_14(net4493[0:47]), .sp4_h_l_13(net4492[0:47]),
     .sp4_h_l_12(net4491[0:47]), .sp4_h_l_11(net4490[0:47]),
     .tnr_op_16(tnr_op_27_16[7:0]), .tnl_op_16(tnl_op_27_16[7:0]),
     .lft_op_16(slf_op_26_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net4512[0:7]), .slf_op_14(net4511[0:7]),
     .slf_op_13(net4514[0:7]), .slf_op_12(net4513[0:7]),
     .slf_op_11(net4515[0:7]), .rgt_op_14(net3044[0:7]),
     .rgt_op_15(net3045[0:7]), .rgt_op_12(net3046[0:7]),
     .rgt_op_13(net3047[0:7]), .rgt_op_11(net3048[0:7]),
     .sp4_v_b_16(net4522[0:47]), .sp4_v_b_14(net4525[0:47]),
     .sp4_v_b_15(net4523[0:47]), .sp4_v_b_13(net4524[0:47]),
     .sp4_v_b_11(net4527[0:47]), .sp4_v_b_12(net4526[0:47]),
     .sp4_r_v_b_16(net3055[0:47]), .sp4_r_v_b_15(net3056[0:47]),
     .sp4_r_v_b_13(net3057[0:47]), .sp4_r_v_b_14(net3058[0:47]),
     .sp4_r_v_b_12(net3059[0:47]), .sp4_r_v_b_11(net3060[0:47]),
     .sp12_h_l_16(net4534[0:23]), .sp12_h_l_15(net4536[0:23]),
     .sp12_h_l_14(net4535[0:23]), .sp12_h_l_13(net4538[0:23]),
     .sp12_h_l_12(net4537[0:23]), .sp12_h_l_11(net4539[0:23]),
     .sp12_h_r_16(net3067[0:23]), .sp12_h_r_14(net3068[0:23]),
     .sp12_h_r_15(net3069[0:23]), .sp12_h_r_12(net3070[0:23]),
     .sp12_h_r_13(net3071[0:23]), .sp12_h_r_11(net3072[0:23]),
     .lft_op_14(net2443[0:7]), .lft_op_15(net2444[0:7]),
     .lft_op_12(net2441[0:7]), .lft_op_11(net2440[0:7]),
     .lft_op_13(net2442[0:7]));
array_LT1x16 I_lt_32_bot ( .sp12_v_b_01(net2183[0:23]),
     .glb_netwk(net2184[0:7]), .sp12_v_t_16(sp12_v_t_32_16[23:0]),
     .rgt_op_16({slf_op_33_16[3], slf_op_33_16[2], slf_op_33_16[1],
     slf_op_33_16[0], slf_op_33_16[3], slf_op_33_16[2],
     slf_op_33_16[1], slf_op_33_16[0]}), .top_op_16(top_op_32_16[7:0]),
     .rgt_op_03({slf_op_33_03[3], slf_op_33_03[2], slf_op_33_03[1],
     slf_op_33_03[0], slf_op_33_03[3], slf_op_33_03[2],
     slf_op_33_03[1], slf_op_33_03[0]}), .slf_op_02(net3735[0:7]),
     .rgt_op_02({slf_op_33_02[3], slf_op_33_02[2], slf_op_33_02[1],
     slf_op_33_02[0], slf_op_33_02[3], slf_op_33_02[2],
     slf_op_33_02[1], slf_op_33_02[0]}), .rgt_op_01({slf_op_33_01[3],
     slf_op_33_01[2], slf_op_33_01[1], slf_op_33_01[0],
     slf_op_33_01[3], slf_op_33_01[2], slf_op_33_01[1],
     slf_op_33_01[0]}), .purst(purst), .prog(prog),
     .lft_op_04(net4232[0:7]), .lft_op_03(net4222[0:7]),
     .lft_op_02(net4224[0:7]), .lft_op_01(net2185[0:7]),
     .rgt_op_04({slf_op_33_04[3], slf_op_33_04[2], slf_op_33_04[1],
     slf_op_33_04[0], slf_op_33_04[3], slf_op_33_04[2],
     slf_op_33_04[1], slf_op_33_04[0]}), .carry_in(net2530),
     .bnl_op_01({slf_op_31_00[3], slf_op_31_00[2], slf_op_31_00[1],
     slf_op_31_00[0], slf_op_31_00[3], slf_op_31_00[2],
     slf_op_31_00[1], slf_op_31_00[0]}), .slf_op_04(net3743[0:7]),
     .slf_op_03(net3733[0:7]), .slf_op_01(net2188[0:7]),
     .sp4_h_l_04(net3764[0:47]), .carry_out(carry_out_32_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net3101[0:23]),
     .sp12_h_r_03(net3102[0:23]), .sp12_h_r_02(net3103[0:23]),
     .sp12_h_r_01(net3104[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_32_16[7:0]), .sp4_v_b_01(net2189[0:47]),
     .sp4_r_v_b_04(net2542[0:47]), .sp4_r_v_b_03(net2541[0:47]),
     .sp4_r_v_b_02(net2539[0:47]), .sp4_r_v_b_01(net2540[0:47]),
     .sp4_h_r_04(net2585[0:47]), .sp4_h_r_03(net2583[0:47]),
     .sp4_h_r_02(net3114[0:47]), .sp4_h_r_01(net3115[0:47]),
     .sp4_h_l_03(net3765[0:47]), .sp4_h_l_02(net3766[0:47]),
     .sp4_h_l_01(net3767[0:47]), .bl(bl[1725:1672]),
     .bot_op_01({slf_op_32_00[3], slf_op_32_00[2], slf_op_32_00[1],
     slf_op_32_00[0], slf_op_32_00[3], slf_op_32_00[2],
     slf_op_32_00[1], slf_op_32_00[0]}), .sp12_h_l_01(net3756[0:23]),
     .sp12_h_l_02(net3755[0:23]), .sp12_h_l_03(net3754[0:23]),
     .sp12_h_l_04(net3753[0:23]), .sp4_v_b_04(net3760[0:47]),
     .sp4_v_b_03(net3761[0:47]), .sp4_v_b_02(net3762[0:47]),
     .bnr_op_01({tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd}), .sp4_h_l_05(net3792[0:47]),
     .sp4_h_l_06(net3791[0:47]), .sp4_h_l_07(net3790[0:47]),
     .sp4_h_l_08(net3789[0:47]), .sp4_h_l_09(net3788[0:47]),
     .sp4_h_l_10(net3787[0:47]), .sp4_h_r_10(net3135[0:47]),
     .sp4_h_r_09(net3136[0:47]), .sp4_h_r_08(net3137[0:47]),
     .sp4_h_r_07(net3138[0:47]), .sp4_h_r_06(net3139[0:47]),
     .sp4_h_r_05(net3140[0:47]), .slf_op_05(net3804[0:7]),
     .slf_op_06(net3803[0:7]), .slf_op_07(net3802[0:7]),
     .slf_op_08(net3801[0:7]), .slf_op_09(net3800[0:7]),
     .slf_op_10(net3799[0:7]), .rgt_op_10({slf_op_33_10[3],
     slf_op_33_10[2], slf_op_33_10[1], slf_op_33_10[0],
     slf_op_33_10[3], slf_op_33_10[2], slf_op_33_10[1],
     slf_op_33_10[0]}), .rgt_op_09({slf_op_33_09[3], slf_op_33_09[2],
     slf_op_33_09[1], slf_op_33_09[0], slf_op_33_09[3],
     slf_op_33_09[2], slf_op_33_09[1], slf_op_33_09[0]}),
     .rgt_op_08({slf_op_33_08[3], slf_op_33_08[2], slf_op_33_08[1],
     slf_op_33_08[0], slf_op_33_08[3], slf_op_33_08[2],
     slf_op_33_08[1], slf_op_33_08[0]}), .rgt_op_07({slf_op_33_07[3],
     slf_op_33_07[2], slf_op_33_07[1], slf_op_33_07[0],
     slf_op_33_07[3], slf_op_33_07[2], slf_op_33_07[1],
     slf_op_33_07[0]}), .rgt_op_06({slf_op_33_06[3], slf_op_33_06[2],
     slf_op_33_06[1], slf_op_33_06[0], slf_op_33_06[3],
     slf_op_33_06[2], slf_op_33_06[1], slf_op_33_06[0]}),
     .rgt_op_05({slf_op_33_05[3], slf_op_33_05[2], slf_op_33_05[1],
     slf_op_33_05[0], slf_op_33_05[3], slf_op_33_05[2],
     slf_op_33_05[1], slf_op_33_05[0]}), .lft_op_10(net4288[0:7]),
     .lft_op_09(net4289[0:7]), .lft_op_08(net4290[0:7]),
     .lft_op_07(net4291[0:7]), .lft_op_06(net4292[0:7]),
     .lft_op_05(net4293[0:7]), .sp12_h_l_10(net3812[0:23]),
     .sp12_h_r_10(net3160[0:23]), .sp12_h_l_09(net3821[0:23]),
     .sp12_h_l_08(net3820[0:23]), .sp12_h_l_07(net3819[0:23]),
     .sp12_h_l_06(net3818[0:23]), .sp12_h_r_05(net3165[0:23]),
     .sp12_h_r_06(net3166[0:23]), .sp12_h_r_07(net3167[0:23]),
     .sp12_h_r_08(net3168[0:23]), .sp12_h_r_09(net3169[0:23]),
     .sp12_h_l_05(net3817[0:23]), .sp4_r_v_b_05(net2537[0:47]),
     .sp4_r_v_b_06(net2538[0:47]), .sp4_r_v_b_07(net2536[0:47]),
     .sp4_r_v_b_08(net2535[0:47]), .sp4_r_v_b_09(net2545[0:47]),
     .sp4_r_v_b_10(net2546[0:47]), .sp4_v_b_10(net3828[0:47]),
     .sp4_v_b_09(net3827[0:47]), .sp4_v_b_08(net3826[0:47]),
     .sp4_v_b_07(net3825[0:47]), .sp4_v_b_06(net3824[0:47]),
     .sp4_v_b_05(net3823[0:47]), .sp4_v_t_16(sp4_v_t_32_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net3186[0:47]), .sp4_h_r_12(net3187[0:47]),
     .sp4_h_r_13(net3188[0:47]), .sp4_h_r_14(net3189[0:47]),
     .sp4_h_r_15(net3190[0:47]), .sp4_h_r_16(net3191[0:47]),
     .sp4_h_l_16(net3843[0:47]), .sp4_h_l_15(net3842[0:47]),
     .sp4_h_l_14(net3841[0:47]), .sp4_h_l_13(net3840[0:47]),
     .sp4_h_l_12(net3839[0:47]), .sp4_h_l_11(net3838[0:47]),
     .tnr_op_16(tnr_op_32_16[7:0]), .tnl_op_16(tnl_op_32_16[7:0]),
     .lft_op_16(slf_op_31_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net3860[0:7]), .slf_op_14(net3859[0:7]),
     .slf_op_13(net3862[0:7]), .slf_op_12(net3861[0:7]),
     .slf_op_11(net3863[0:7]), .rgt_op_14({slf_op_33_14[3],
     slf_op_33_14[2], slf_op_33_14[1], slf_op_33_14[0],
     slf_op_33_14[3], slf_op_33_14[2], slf_op_33_14[1],
     slf_op_33_14[0]}), .rgt_op_15({slf_op_33_15[3], slf_op_33_15[2],
     slf_op_33_15[1], slf_op_33_15[0], slf_op_33_15[3],
     slf_op_33_15[2], slf_op_33_15[1], slf_op_33_15[0]}),
     .rgt_op_12({slf_op_33_12[3], slf_op_33_12[2], slf_op_33_12[1],
     slf_op_33_12[0], slf_op_33_12[3], slf_op_33_12[2],
     slf_op_33_12[1], slf_op_33_12[0]}), .rgt_op_13({slf_op_33_13[3],
     slf_op_33_13[2], slf_op_33_13[1], slf_op_33_13[0],
     slf_op_33_13[3], slf_op_33_13[2], slf_op_33_13[1],
     slf_op_33_13[0]}), .rgt_op_11({slf_op_33_11[3], slf_op_33_11[2],
     slf_op_33_11[1], slf_op_33_11[0], slf_op_33_11[3],
     slf_op_33_11[2], slf_op_33_11[1], slf_op_33_11[0]}),
     .sp4_v_b_16(net3870[0:47]), .sp4_v_b_14(net3873[0:47]),
     .sp4_v_b_15(net3871[0:47]), .sp4_v_b_13(net3872[0:47]),
     .sp4_v_b_11(net3875[0:47]), .sp4_v_b_12(net3874[0:47]),
     .sp4_r_v_b_16(net2550[0:47]), .sp4_r_v_b_15(net2549[0:47]),
     .sp4_r_v_b_13(net2548[0:47]), .sp4_r_v_b_14(net2547[0:47]),
     .sp4_r_v_b_12(net2543[0:47]), .sp4_r_v_b_11(net2544[0:47]),
     .sp12_h_l_16(net3882[0:23]), .sp12_h_l_15(net3884[0:23]),
     .sp12_h_l_14(net3883[0:23]), .sp12_h_l_13(net3886[0:23]),
     .sp12_h_l_12(net3885[0:23]), .sp12_h_l_11(net3887[0:23]),
     .sp12_h_r_16(net3230[0:23]), .sp12_h_r_14(net3231[0:23]),
     .sp12_h_r_15(net3232[0:23]), .sp12_h_r_12(net3233[0:23]),
     .sp12_h_r_13(net3234[0:23]), .sp12_h_r_11(net3235[0:23]),
     .lft_op_14(net4348[0:7]), .lft_op_15(net4349[0:7]),
     .lft_op_12(net4350[0:7]), .lft_op_11(net4352[0:7]),
     .lft_op_13(net4351[0:7]));
array_LT1x16 I_lt_22_bot ( .sp12_v_b_01(net2132[0:23]),
     .glb_netwk(net2131[0:7]), .sp12_v_t_16(sp12_v_t_22_16[23:0]),
     .rgt_op_16(slf_op_23_16[7:0]), .top_op_16(top_op_22_16[7:0]),
     .rgt_op_03(net3244[0:7]), .slf_op_02(net2594[0:7]),
     .rgt_op_02(net3246[0:7]), .rgt_op_01(net2115[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4884[0:7]), .lft_op_03(net4874[0:7]),
     .lft_op_02(net4876[0:7]), .lft_op_01(net2130[0:7]),
     .rgt_op_04(net3254[0:7]), .carry_in(net2518),
     .bnl_op_01({slf_op_21_00[3], slf_op_21_00[2], slf_op_21_00[1],
     slf_op_21_00[0], slf_op_21_00[3], slf_op_21_00[2],
     slf_op_21_00[1], slf_op_21_00[0]}), .slf_op_04(net2602[0:7]),
     .slf_op_03(net2592[0:7]), .slf_op_01(net2122[0:7]),
     .sp4_h_l_04(net2623[0:47]), .carry_out(carry_out_22_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net3264[0:23]),
     .sp12_h_r_03(net3265[0:23]), .sp12_h_r_02(net3266[0:23]),
     .sp12_h_r_01(net3267[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_22_16[7:0]), .sp4_v_b_01(net2125[0:47]),
     .sp4_r_v_b_04(net3271[0:47]), .sp4_r_v_b_03(net3272[0:47]),
     .sp4_r_v_b_02(net3273[0:47]), .sp4_r_v_b_01(net2117[0:47]),
     .sp4_h_r_04(net3275[0:47]), .sp4_h_r_03(net3276[0:47]),
     .sp4_h_r_02(net3277[0:47]), .sp4_h_r_01(net3278[0:47]),
     .sp4_h_l_03(net2624[0:47]), .sp4_h_l_02(net2625[0:47]),
     .sp4_h_l_01(net2626[0:47]), .bl(bl[1197:1144]),
     .bot_op_01({slf_op_22_00[3], slf_op_22_00[2], slf_op_22_00[1],
     slf_op_22_00[0], slf_op_22_00[3], slf_op_22_00[2],
     slf_op_22_00[1], slf_op_22_00[0]}), .sp12_h_l_01(net2615[0:23]),
     .sp12_h_l_02(net2614[0:23]), .sp12_h_l_03(net2613[0:23]),
     .sp12_h_l_04(net2612[0:23]), .sp4_v_b_04(net2619[0:47]),
     .sp4_v_b_03(net2620[0:47]), .sp4_v_b_02(net2621[0:47]),
     .bnr_op_01({slf_op_23_00[3], slf_op_23_00[2], slf_op_23_00[1],
     slf_op_23_00[0], slf_op_23_00[3], slf_op_23_00[2],
     slf_op_23_00[1], slf_op_23_00[0]}), .sp4_h_l_05(net2651[0:47]),
     .sp4_h_l_06(net2650[0:47]), .sp4_h_l_07(net2649[0:47]),
     .sp4_h_l_08(net2648[0:47]), .sp4_h_l_09(net2647[0:47]),
     .sp4_h_l_10(net2646[0:47]), .sp4_h_r_10(net3298[0:47]),
     .sp4_h_r_09(net3299[0:47]), .sp4_h_r_08(net3300[0:47]),
     .sp4_h_r_07(net3301[0:47]), .sp4_h_r_06(net3302[0:47]),
     .sp4_h_r_05(net3303[0:47]), .slf_op_05(net2663[0:7]),
     .slf_op_06(net2662[0:7]), .slf_op_07(net2661[0:7]),
     .slf_op_08(net2660[0:7]), .slf_op_09(net2659[0:7]),
     .slf_op_10(net2658[0:7]), .rgt_op_10(net3310[0:7]),
     .rgt_op_09(net3311[0:7]), .rgt_op_08(net3312[0:7]),
     .rgt_op_07(net3313[0:7]), .rgt_op_06(net3314[0:7]),
     .rgt_op_05(net3315[0:7]), .lft_op_10(net4940[0:7]),
     .lft_op_09(net4941[0:7]), .lft_op_08(net4942[0:7]),
     .lft_op_07(net4943[0:7]), .lft_op_06(net4944[0:7]),
     .lft_op_05(net4945[0:7]), .sp12_h_l_10(net2671[0:23]),
     .sp12_h_r_10(net3323[0:23]), .sp12_h_l_09(net2680[0:23]),
     .sp12_h_l_08(net2679[0:23]), .sp12_h_l_07(net2678[0:23]),
     .sp12_h_l_06(net2677[0:23]), .sp12_h_r_05(net3328[0:23]),
     .sp12_h_r_06(net3329[0:23]), .sp12_h_r_07(net3330[0:23]),
     .sp12_h_r_08(net3331[0:23]), .sp12_h_r_09(net3332[0:23]),
     .sp12_h_l_05(net2676[0:23]), .sp4_r_v_b_05(net3334[0:47]),
     .sp4_r_v_b_06(net3335[0:47]), .sp4_r_v_b_07(net3336[0:47]),
     .sp4_r_v_b_08(net3337[0:47]), .sp4_r_v_b_09(net3338[0:47]),
     .sp4_r_v_b_10(net3339[0:47]), .sp4_v_b_10(net2687[0:47]),
     .sp4_v_b_09(net2686[0:47]), .sp4_v_b_08(net2685[0:47]),
     .sp4_v_b_07(net2684[0:47]), .sp4_v_b_06(net2683[0:47]),
     .sp4_v_b_05(net2682[0:47]), .sp4_v_t_16(sp4_v_t_22_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net3349[0:47]), .sp4_h_r_12(net3350[0:47]),
     .sp4_h_r_13(net3351[0:47]), .sp4_h_r_14(net3352[0:47]),
     .sp4_h_r_15(net3353[0:47]), .sp4_h_r_16(net3354[0:47]),
     .sp4_h_l_16(net2702[0:47]), .sp4_h_l_15(net2701[0:47]),
     .sp4_h_l_14(net2700[0:47]), .sp4_h_l_13(net2699[0:47]),
     .sp4_h_l_12(net2698[0:47]), .sp4_h_l_11(net2697[0:47]),
     .tnr_op_16(tnr_op_22_16[7:0]), .tnl_op_16(tnl_op_22_16[7:0]),
     .lft_op_16(slf_op_21_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net2719[0:7]), .slf_op_14(net2718[0:7]),
     .slf_op_13(net2721[0:7]), .slf_op_12(net2720[0:7]),
     .slf_op_11(net2722[0:7]), .rgt_op_14(net3370[0:7]),
     .rgt_op_15(net3371[0:7]), .rgt_op_12(net3372[0:7]),
     .rgt_op_13(net3373[0:7]), .rgt_op_11(net3374[0:7]),
     .sp4_v_b_16(net2729[0:47]), .sp4_v_b_14(net2732[0:47]),
     .sp4_v_b_15(net2730[0:47]), .sp4_v_b_13(net2731[0:47]),
     .sp4_v_b_11(net2734[0:47]), .sp4_v_b_12(net2733[0:47]),
     .sp4_r_v_b_16(net3381[0:47]), .sp4_r_v_b_15(net3382[0:47]),
     .sp4_r_v_b_13(net3383[0:47]), .sp4_r_v_b_14(net3384[0:47]),
     .sp4_r_v_b_12(net3385[0:47]), .sp4_r_v_b_11(net3386[0:47]),
     .sp12_h_l_16(net2741[0:23]), .sp12_h_l_15(net2743[0:23]),
     .sp12_h_l_14(net2742[0:23]), .sp12_h_l_13(net2745[0:23]),
     .sp12_h_l_12(net2744[0:23]), .sp12_h_l_11(net2746[0:23]),
     .sp12_h_r_16(net3393[0:23]), .sp12_h_r_14(net3394[0:23]),
     .sp12_h_r_15(net3395[0:23]), .sp12_h_r_12(net3396[0:23]),
     .sp12_h_r_13(net3397[0:23]), .sp12_h_r_11(net3398[0:23]),
     .lft_op_14(net5000[0:7]), .lft_op_15(net5001[0:7]),
     .lft_op_12(net5002[0:7]), .lft_op_11(net5004[0:7]),
     .lft_op_13(net5003[0:7]));
array_LT1x16 I_lt_19_bot ( .sp12_v_b_01(net2156[0:23]),
     .glb_netwk(net2155[0:7]), .sp12_v_t_16(sp12_v_t_19_16[23:0]),
     .rgt_op_16(slf_op_20_16[7:0]), .top_op_16(top_op_19_16[7:0]),
     .rgt_op_03(net3407[0:7]), .slf_op_02(net4550[0:7]),
     .rgt_op_02(net3409[0:7]), .rgt_op_01(net2138[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4721[0:7]), .lft_op_03(net4711[0:7]),
     .lft_op_02(net4713[0:7]), .lft_op_01(net2154[0:7]),
     .rgt_op_04(net3417[0:7]), .carry_in(net2533),
     .bnl_op_01({slf_op_18_00[3], slf_op_18_00[2], slf_op_18_00[1],
     slf_op_18_00[0], slf_op_18_00[3], slf_op_18_00[2],
     slf_op_18_00[1], slf_op_18_00[0]}), .slf_op_04(net4558[0:7]),
     .slf_op_03(net4548[0:7]), .slf_op_01(net2146[0:7]),
     .sp4_h_l_04(net4579[0:47]), .carry_out(carry_out_19_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net3427[0:23]),
     .sp12_h_r_03(net3428[0:23]), .sp12_h_r_02(net3429[0:23]),
     .sp12_h_r_01(net3430[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_19_16[7:0]), .sp4_v_b_01(net2149[0:47]),
     .sp4_r_v_b_04(net3434[0:47]), .sp4_r_v_b_03(net3435[0:47]),
     .sp4_r_v_b_02(net3436[0:47]), .sp4_r_v_b_01(net2141[0:47]),
     .sp4_h_r_04(net3438[0:47]), .sp4_h_r_03(net3439[0:47]),
     .sp4_h_r_02(net3440[0:47]), .sp4_h_r_01(net3441[0:47]),
     .sp4_h_l_03(net4580[0:47]), .sp4_h_l_02(net4581[0:47]),
     .sp4_h_l_01(net4582[0:47]), .bl(bl[1035:982]),
     .bot_op_01({slf_op_19_00[3], slf_op_19_00[2], slf_op_19_00[1],
     slf_op_19_00[0], slf_op_19_00[3], slf_op_19_00[2],
     slf_op_19_00[1], slf_op_19_00[0]}), .sp12_h_l_01(net4571[0:23]),
     .sp12_h_l_02(net4570[0:23]), .sp12_h_l_03(net4569[0:23]),
     .sp12_h_l_04(net4568[0:23]), .sp4_v_b_04(net4575[0:47]),
     .sp4_v_b_03(net4576[0:47]), .sp4_v_b_02(net4577[0:47]),
     .bnr_op_01({slf_op_20_00[3], slf_op_20_00[2], slf_op_20_00[1],
     slf_op_20_00[0], slf_op_20_00[3], slf_op_20_00[2],
     slf_op_20_00[1], slf_op_20_00[0]}), .sp4_h_l_05(net4607[0:47]),
     .sp4_h_l_06(net4606[0:47]), .sp4_h_l_07(net4605[0:47]),
     .sp4_h_l_08(net4604[0:47]), .sp4_h_l_09(net4603[0:47]),
     .sp4_h_l_10(net4602[0:47]), .sp4_h_r_10(net3461[0:47]),
     .sp4_h_r_09(net3462[0:47]), .sp4_h_r_08(net3463[0:47]),
     .sp4_h_r_07(net3464[0:47]), .sp4_h_r_06(net3465[0:47]),
     .sp4_h_r_05(net3466[0:47]), .slf_op_05(net4619[0:7]),
     .slf_op_06(net4618[0:7]), .slf_op_07(net4617[0:7]),
     .slf_op_08(net4616[0:7]), .slf_op_09(net4615[0:7]),
     .slf_op_10(net4614[0:7]), .rgt_op_10(net3473[0:7]),
     .rgt_op_09(net3474[0:7]), .rgt_op_08(net3475[0:7]),
     .rgt_op_07(net3476[0:7]), .rgt_op_06(net3477[0:7]),
     .rgt_op_05(net3478[0:7]), .lft_op_10(net4777[0:7]),
     .lft_op_09(net4778[0:7]), .lft_op_08(net4779[0:7]),
     .lft_op_07(net4780[0:7]), .lft_op_06(net4781[0:7]),
     .lft_op_05(net4782[0:7]), .sp12_h_l_10(net4627[0:23]),
     .sp12_h_r_10(net3486[0:23]), .sp12_h_l_09(net4636[0:23]),
     .sp12_h_l_08(net4635[0:23]), .sp12_h_l_07(net4634[0:23]),
     .sp12_h_l_06(net4633[0:23]), .sp12_h_r_05(net3491[0:23]),
     .sp12_h_r_06(net3492[0:23]), .sp12_h_r_07(net3493[0:23]),
     .sp12_h_r_08(net3494[0:23]), .sp12_h_r_09(net3495[0:23]),
     .sp12_h_l_05(net4632[0:23]), .sp4_r_v_b_05(net3497[0:47]),
     .sp4_r_v_b_06(net3498[0:47]), .sp4_r_v_b_07(net3499[0:47]),
     .sp4_r_v_b_08(net3500[0:47]), .sp4_r_v_b_09(net3501[0:47]),
     .sp4_r_v_b_10(net3502[0:47]), .sp4_v_b_10(net4643[0:47]),
     .sp4_v_b_09(net4642[0:47]), .sp4_v_b_08(net4641[0:47]),
     .sp4_v_b_07(net4640[0:47]), .sp4_v_b_06(net4639[0:47]),
     .sp4_v_b_05(net4638[0:47]), .sp4_v_t_16(sp4_v_t_19_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net3512[0:47]), .sp4_h_r_12(net3513[0:47]),
     .sp4_h_r_13(net3514[0:47]), .sp4_h_r_14(net3515[0:47]),
     .sp4_h_r_15(net3516[0:47]), .sp4_h_r_16(sp4_h_r_19_20[47:0]),
     .sp4_h_l_16(sp4_h_r_18_19[47:0]), .sp4_h_l_15(net4657[0:47]),
     .sp4_h_l_14(net4656[0:47]), .sp4_h_l_13(net4655[0:47]),
     .sp4_h_l_12(net4654[0:47]), .sp4_h_l_11(net4653[0:47]),
     .tnr_op_16(tnr_op_19_16[7:0]), .tnl_op_16(tnl_op_19_16[7:0]),
     .lft_op_16(slf_op_18_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net4675[0:7]), .slf_op_14(net4674[0:7]),
     .slf_op_13(net4677[0:7]), .slf_op_12(net4676[0:7]),
     .slf_op_11(net4678[0:7]), .rgt_op_14(net3533[0:7]),
     .rgt_op_15(net3534[0:7]), .rgt_op_12(net3535[0:7]),
     .rgt_op_13(net3536[0:7]), .rgt_op_11(net3537[0:7]),
     .sp4_v_b_16(net4685[0:47]), .sp4_v_b_14(net4688[0:47]),
     .sp4_v_b_15(net4686[0:47]), .sp4_v_b_13(net4687[0:47]),
     .sp4_v_b_11(net4690[0:47]), .sp4_v_b_12(net4689[0:47]),
     .sp4_r_v_b_16(net3544[0:47]), .sp4_r_v_b_15(net3545[0:47]),
     .sp4_r_v_b_13(net3546[0:47]), .sp4_r_v_b_14(net3547[0:47]),
     .sp4_r_v_b_12(net3548[0:47]), .sp4_r_v_b_11(net3549[0:47]),
     .sp12_h_l_16(net4697[0:23]), .sp12_h_l_15(net4699[0:23]),
     .sp12_h_l_14(net4698[0:23]), .sp12_h_l_13(net4701[0:23]),
     .sp12_h_l_12(net4700[0:23]), .sp12_h_l_11(net4702[0:23]),
     .sp12_h_r_16(net3556[0:23]), .sp12_h_r_14(net3557[0:23]),
     .sp12_h_r_15(net3558[0:23]), .sp12_h_r_12(net3559[0:23]),
     .sp12_h_r_13(net3560[0:23]), .sp12_h_r_11(net3561[0:23]),
     .lft_op_14(net4837[0:7]), .lft_op_15(net4838[0:7]),
     .lft_op_12(net4839[0:7]), .lft_op_11(net4841[0:7]),
     .lft_op_13(net4840[0:7]));
array_LT1x16 I_lt_24_bot ( .sp12_v_b_01(net2090[0:23]),
     .glb_netwk(net2116[0:7]), .sp12_v_t_16(sp12_v_t_24_16[23:0]),
     .rgt_op_16(slf_op_25_16[7:0]), .top_op_16(top_op_24_16[7:0]),
     .rgt_op_03(net3570[0:7]), .slf_op_02(net4061[0:7]),
     .rgt_op_02(net3572[0:7]), .rgt_op_01(net2101[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3254[0:7]), .lft_op_03(net3244[0:7]),
     .lft_op_02(net3246[0:7]), .lft_op_01(net2115[0:7]),
     .rgt_op_04(net3580[0:7]), .carry_in(net2513),
     .bnl_op_01({slf_op_23_00[3], slf_op_23_00[2], slf_op_23_00[1],
     slf_op_23_00[0], slf_op_23_00[3], slf_op_23_00[2],
     slf_op_23_00[1], slf_op_23_00[0]}), .slf_op_04(net4069[0:7]),
     .slf_op_03(net4059[0:7]), .slf_op_01(net2108[0:7]),
     .sp4_h_l_04(net4090[0:47]), .carry_out(carry_out_24_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net3590[0:23]),
     .sp12_h_r_03(net3591[0:23]), .sp12_h_r_02(net3592[0:23]),
     .sp12_h_r_01(net3593[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_24_16[7:0]), .sp4_v_b_01(net2110[0:47]),
     .sp4_r_v_b_04(net3597[0:47]), .sp4_r_v_b_03(net3598[0:47]),
     .sp4_r_v_b_02(net3599[0:47]), .sp4_r_v_b_01(net2104[0:47]),
     .sp4_h_r_04(net3601[0:47]), .sp4_h_r_03(net3602[0:47]),
     .sp4_h_r_02(net3603[0:47]), .sp4_h_r_01(net3604[0:47]),
     .sp4_h_l_03(net4091[0:47]), .sp4_h_l_02(net4092[0:47]),
     .sp4_h_l_01(net4093[0:47]), .bl(bl[1305:1252]),
     .bot_op_01({slf_op_24_00[3], slf_op_24_00[2], slf_op_24_00[1],
     slf_op_24_00[0], slf_op_24_00[3], slf_op_24_00[2],
     slf_op_24_00[1], slf_op_24_00[0]}), .sp12_h_l_01(net4082[0:23]),
     .sp12_h_l_02(net4081[0:23]), .sp12_h_l_03(net4080[0:23]),
     .sp12_h_l_04(net4079[0:23]), .sp4_v_b_04(net4086[0:47]),
     .sp4_v_b_03(net4087[0:47]), .sp4_v_b_02(net4088[0:47]),
     .bnr_op_01({slf_op_25_00[3], slf_op_25_00[2], slf_op_25_00[1],
     slf_op_25_00[0], slf_op_25_00[3], slf_op_25_00[2],
     slf_op_25_00[1], slf_op_25_00[0]}), .sp4_h_l_05(net4118[0:47]),
     .sp4_h_l_06(net4117[0:47]), .sp4_h_l_07(net4116[0:47]),
     .sp4_h_l_08(net4115[0:47]), .sp4_h_l_09(net4114[0:47]),
     .sp4_h_l_10(net4113[0:47]), .sp4_h_r_10(net3624[0:47]),
     .sp4_h_r_09(net3625[0:47]), .sp4_h_r_08(net3626[0:47]),
     .sp4_h_r_07(net3627[0:47]), .sp4_h_r_06(net3628[0:47]),
     .sp4_h_r_05(net3629[0:47]), .slf_op_05(net4130[0:7]),
     .slf_op_06(net4129[0:7]), .slf_op_07(net4128[0:7]),
     .slf_op_08(net4127[0:7]), .slf_op_09(net4126[0:7]),
     .slf_op_10(net4125[0:7]), .rgt_op_10(net3636[0:7]),
     .rgt_op_09(net3637[0:7]), .rgt_op_08(net3638[0:7]),
     .rgt_op_07(net3639[0:7]), .rgt_op_06(net3640[0:7]),
     .rgt_op_05(net3641[0:7]), .lft_op_10(net3310[0:7]),
     .lft_op_09(net3311[0:7]), .lft_op_08(net3312[0:7]),
     .lft_op_07(net3313[0:7]), .lft_op_06(net3314[0:7]),
     .lft_op_05(net3315[0:7]), .sp12_h_l_10(net4138[0:23]),
     .sp12_h_r_10(net3649[0:23]), .sp12_h_l_09(net4147[0:23]),
     .sp12_h_l_08(net4146[0:23]), .sp12_h_l_07(net4145[0:23]),
     .sp12_h_l_06(net4144[0:23]), .sp12_h_r_05(net3654[0:23]),
     .sp12_h_r_06(net3655[0:23]), .sp12_h_r_07(net3656[0:23]),
     .sp12_h_r_08(net3657[0:23]), .sp12_h_r_09(net3658[0:23]),
     .sp12_h_l_05(net4143[0:23]), .sp4_r_v_b_05(net3660[0:47]),
     .sp4_r_v_b_06(net3661[0:47]), .sp4_r_v_b_07(net3662[0:47]),
     .sp4_r_v_b_08(net3663[0:47]), .sp4_r_v_b_09(net3664[0:47]),
     .sp4_r_v_b_10(net3665[0:47]), .sp4_v_b_10(net4154[0:47]),
     .sp4_v_b_09(net4153[0:47]), .sp4_v_b_08(net4152[0:47]),
     .sp4_v_b_07(net4151[0:47]), .sp4_v_b_06(net4150[0:47]),
     .sp4_v_b_05(net4149[0:47]), .sp4_v_t_16(sp4_v_t_24_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net3675[0:47]), .sp4_h_r_12(net3676[0:47]),
     .sp4_h_r_13(net3677[0:47]), .sp4_h_r_14(net3678[0:47]),
     .sp4_h_r_15(net3679[0:47]), .sp4_h_r_16(net3680[0:47]),
     .sp4_h_l_16(net4169[0:47]), .sp4_h_l_15(net4168[0:47]),
     .sp4_h_l_14(net4167[0:47]), .sp4_h_l_13(net4166[0:47]),
     .sp4_h_l_12(net4165[0:47]), .sp4_h_l_11(net4164[0:47]),
     .tnr_op_16(tnr_op_24_16[7:0]), .tnl_op_16(tnl_op_24_16[7:0]),
     .lft_op_16(slf_op_23_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net4186[0:7]), .slf_op_14(net4185[0:7]),
     .slf_op_13(net4188[0:7]), .slf_op_12(net4187[0:7]),
     .slf_op_11(net4189[0:7]), .rgt_op_14(net3696[0:7]),
     .rgt_op_15(net3697[0:7]), .rgt_op_12(net3698[0:7]),
     .rgt_op_13(net3699[0:7]), .rgt_op_11(net3700[0:7]),
     .sp4_v_b_16(net4196[0:47]), .sp4_v_b_14(net4199[0:47]),
     .sp4_v_b_15(net4197[0:47]), .sp4_v_b_13(net4198[0:47]),
     .sp4_v_b_11(net4201[0:47]), .sp4_v_b_12(net4200[0:47]),
     .sp4_r_v_b_16(net3707[0:47]), .sp4_r_v_b_15(net3708[0:47]),
     .sp4_r_v_b_13(net3709[0:47]), .sp4_r_v_b_14(net3710[0:47]),
     .sp4_r_v_b_12(net3711[0:47]), .sp4_r_v_b_11(net3712[0:47]),
     .sp12_h_l_16(net4208[0:23]), .sp12_h_l_15(net4210[0:23]),
     .sp12_h_l_14(net4209[0:23]), .sp12_h_l_13(net4212[0:23]),
     .sp12_h_l_12(net4211[0:23]), .sp12_h_l_11(net4213[0:23]),
     .sp12_h_r_16(net3719[0:23]), .sp12_h_r_14(net3720[0:23]),
     .sp12_h_r_15(net3721[0:23]), .sp12_h_r_12(net3722[0:23]),
     .sp12_h_r_13(net3723[0:23]), .sp12_h_r_11(net3724[0:23]),
     .lft_op_14(net3370[0:7]), .lft_op_15(net3371[0:7]),
     .lft_op_12(net3372[0:7]), .lft_op_11(net3374[0:7]),
     .lft_op_13(net3373[0:7]));
array_LT1x16 I_lt_31_bot ( .sp12_v_b_01(net2049[0:23]),
     .glb_netwk(net2048[0:7]), .sp12_v_t_16(sp12_v_t_31_16[23:0]),
     .rgt_op_16(slf_op_32_16[7:0]), .top_op_16(top_op_31_16[7:0]),
     .rgt_op_03(net3733[0:7]), .slf_op_02(net4224[0:7]),
     .rgt_op_02(net3735[0:7]), .rgt_op_01(net2188[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3906[0:7]), .lft_op_03(net3896[0:7]),
     .lft_op_02(net3898[0:7]), .lft_op_01(net2047[0:7]),
     .rgt_op_04(net3743[0:7]), .carry_in(net2528),
     .bnl_op_01({slf_op_30_00[3], slf_op_30_00[2], slf_op_30_00[1],
     slf_op_30_00[0], slf_op_30_00[3], slf_op_30_00[2],
     slf_op_30_00[1], slf_op_30_00[0]}), .slf_op_04(net4232[0:7]),
     .slf_op_03(net4222[0:7]), .slf_op_01(net2185[0:7]),
     .sp4_h_l_04(net4253[0:47]), .carry_out(carry_out_31_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net3753[0:23]),
     .sp12_h_r_03(net3754[0:23]), .sp12_h_r_02(net3755[0:23]),
     .sp12_h_r_01(net3756[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_31_16[7:0]), .sp4_v_b_01(net2182[0:47]),
     .sp4_r_v_b_04(net3760[0:47]), .sp4_r_v_b_03(net3761[0:47]),
     .sp4_r_v_b_02(net3762[0:47]), .sp4_r_v_b_01(net2189[0:47]),
     .sp4_h_r_04(net3764[0:47]), .sp4_h_r_03(net3765[0:47]),
     .sp4_h_r_02(net3766[0:47]), .sp4_h_r_01(net3767[0:47]),
     .sp4_h_l_03(net4254[0:47]), .sp4_h_l_02(net4255[0:47]),
     .sp4_h_l_01(net4256[0:47]), .bl(bl[1671:1618]),
     .bot_op_01({slf_op_31_00[3], slf_op_31_00[2], slf_op_31_00[1],
     slf_op_31_00[0], slf_op_31_00[3], slf_op_31_00[2],
     slf_op_31_00[1], slf_op_31_00[0]}), .sp12_h_l_01(net4245[0:23]),
     .sp12_h_l_02(net4244[0:23]), .sp12_h_l_03(net4243[0:23]),
     .sp12_h_l_04(net4242[0:23]), .sp4_v_b_04(net4249[0:47]),
     .sp4_v_b_03(net4250[0:47]), .sp4_v_b_02(net4251[0:47]),
     .bnr_op_01({slf_op_32_00[3], slf_op_32_00[2], slf_op_32_00[1],
     slf_op_32_00[0], slf_op_32_00[3], slf_op_32_00[2],
     slf_op_32_00[1], slf_op_32_00[0]}), .sp4_h_l_05(net4281[0:47]),
     .sp4_h_l_06(net4280[0:47]), .sp4_h_l_07(net4279[0:47]),
     .sp4_h_l_08(net4278[0:47]), .sp4_h_l_09(net4277[0:47]),
     .sp4_h_l_10(net4276[0:47]), .sp4_h_r_10(net3787[0:47]),
     .sp4_h_r_09(net3788[0:47]), .sp4_h_r_08(net3789[0:47]),
     .sp4_h_r_07(net3790[0:47]), .sp4_h_r_06(net3791[0:47]),
     .sp4_h_r_05(net3792[0:47]), .slf_op_05(net4293[0:7]),
     .slf_op_06(net4292[0:7]), .slf_op_07(net4291[0:7]),
     .slf_op_08(net4290[0:7]), .slf_op_09(net4289[0:7]),
     .slf_op_10(net4288[0:7]), .rgt_op_10(net3799[0:7]),
     .rgt_op_09(net3800[0:7]), .rgt_op_08(net3801[0:7]),
     .rgt_op_07(net3802[0:7]), .rgt_op_06(net3803[0:7]),
     .rgt_op_05(net3804[0:7]), .lft_op_10(net3962[0:7]),
     .lft_op_09(net3963[0:7]), .lft_op_08(net3964[0:7]),
     .lft_op_07(net3965[0:7]), .lft_op_06(net3966[0:7]),
     .lft_op_05(net3967[0:7]), .sp12_h_l_10(net4301[0:23]),
     .sp12_h_r_10(net3812[0:23]), .sp12_h_l_09(net4310[0:23]),
     .sp12_h_l_08(net4309[0:23]), .sp12_h_l_07(net4308[0:23]),
     .sp12_h_l_06(net4307[0:23]), .sp12_h_r_05(net3817[0:23]),
     .sp12_h_r_06(net3818[0:23]), .sp12_h_r_07(net3819[0:23]),
     .sp12_h_r_08(net3820[0:23]), .sp12_h_r_09(net3821[0:23]),
     .sp12_h_l_05(net4306[0:23]), .sp4_r_v_b_05(net3823[0:47]),
     .sp4_r_v_b_06(net3824[0:47]), .sp4_r_v_b_07(net3825[0:47]),
     .sp4_r_v_b_08(net3826[0:47]), .sp4_r_v_b_09(net3827[0:47]),
     .sp4_r_v_b_10(net3828[0:47]), .sp4_v_b_10(net4317[0:47]),
     .sp4_v_b_09(net4316[0:47]), .sp4_v_b_08(net4315[0:47]),
     .sp4_v_b_07(net4314[0:47]), .sp4_v_b_06(net4313[0:47]),
     .sp4_v_b_05(net4312[0:47]), .sp4_v_t_16(sp4_v_t_31_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net3838[0:47]), .sp4_h_r_12(net3839[0:47]),
     .sp4_h_r_13(net3840[0:47]), .sp4_h_r_14(net3841[0:47]),
     .sp4_h_r_15(net3842[0:47]), .sp4_h_r_16(net3843[0:47]),
     .sp4_h_l_16(net4332[0:47]), .sp4_h_l_15(net4331[0:47]),
     .sp4_h_l_14(net4330[0:47]), .sp4_h_l_13(net4329[0:47]),
     .sp4_h_l_12(net4328[0:47]), .sp4_h_l_11(net4327[0:47]),
     .tnr_op_16(tnr_op_31_16[7:0]), .tnl_op_16(tnl_op_31_16[7:0]),
     .lft_op_16(slf_op_30_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net4349[0:7]), .slf_op_14(net4348[0:7]),
     .slf_op_13(net4351[0:7]), .slf_op_12(net4350[0:7]),
     .slf_op_11(net4352[0:7]), .rgt_op_14(net3859[0:7]),
     .rgt_op_15(net3860[0:7]), .rgt_op_12(net3861[0:7]),
     .rgt_op_13(net3862[0:7]), .rgt_op_11(net3863[0:7]),
     .sp4_v_b_16(net4359[0:47]), .sp4_v_b_14(net4362[0:47]),
     .sp4_v_b_15(net4360[0:47]), .sp4_v_b_13(net4361[0:47]),
     .sp4_v_b_11(net4364[0:47]), .sp4_v_b_12(net4363[0:47]),
     .sp4_r_v_b_16(net3870[0:47]), .sp4_r_v_b_15(net3871[0:47]),
     .sp4_r_v_b_13(net3872[0:47]), .sp4_r_v_b_14(net3873[0:47]),
     .sp4_r_v_b_12(net3874[0:47]), .sp4_r_v_b_11(net3875[0:47]),
     .sp12_h_l_16(net4371[0:23]), .sp12_h_l_15(net4373[0:23]),
     .sp12_h_l_14(net4372[0:23]), .sp12_h_l_13(net4375[0:23]),
     .sp12_h_l_12(net4374[0:23]), .sp12_h_l_11(net4376[0:23]),
     .sp12_h_r_16(net3882[0:23]), .sp12_h_r_14(net3883[0:23]),
     .sp12_h_r_15(net3884[0:23]), .sp12_h_r_12(net3885[0:23]),
     .sp12_h_r_13(net3886[0:23]), .sp12_h_r_11(net3887[0:23]),
     .lft_op_14(net4022[0:7]), .lft_op_15(net4023[0:7]),
     .lft_op_12(net4024[0:7]), .lft_op_11(net4026[0:7]),
     .lft_op_13(net4025[0:7]));
array_LT1x16 I_lt_29_bot ( .sp12_v_b_01(net2081[0:23]),
     .glb_netwk(net2075[0:7]), .sp12_v_t_16(sp12_v_t_29_16[23:0]),
     .rgt_op_16(slf_op_30_16[7:0]), .top_op_16(top_op_29_16[7:0]),
     .rgt_op_03(net3896[0:7]), .slf_op_02(net2757[0:7]),
     .rgt_op_02(net3898[0:7]), .rgt_op_01(net2047[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2928[0:7]), .lft_op_03(net2918[0:7]),
     .lft_op_02(net2920[0:7]), .lft_op_01(net2074[0:7]),
     .rgt_op_04(net3906[0:7]), .carry_in(net2553),
     .bnl_op_01({slf_op_28_00[3], slf_op_28_00[2], slf_op_28_00[1],
     slf_op_28_00[0], slf_op_28_00[3], slf_op_28_00[2],
     slf_op_28_00[1], slf_op_28_00[0]}), .slf_op_04(net2765[0:7]),
     .slf_op_03(net2755[0:7]), .slf_op_01(net2062[0:7]),
     .sp4_h_l_04(net2786[0:47]), .carry_out(carry_out_29_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net3916[0:23]),
     .sp12_h_r_03(net3917[0:23]), .sp12_h_r_02(net3918[0:23]),
     .sp12_h_r_01(net3919[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_29_16[7:0]), .sp4_v_b_01(net2065[0:47]),
     .sp4_r_v_b_04(net3923[0:47]), .sp4_r_v_b_03(net3924[0:47]),
     .sp4_r_v_b_02(net3925[0:47]), .sp4_r_v_b_01(net2050[0:47]),
     .sp4_h_r_04(net3927[0:47]), .sp4_h_r_03(net3928[0:47]),
     .sp4_h_r_02(net3929[0:47]), .sp4_h_r_01(net3930[0:47]),
     .sp4_h_l_03(net2787[0:47]), .sp4_h_l_02(net2788[0:47]),
     .sp4_h_l_01(net2789[0:47]), .bl(bl[1563:1510]),
     .bot_op_01({slf_op_29_00[3], slf_op_29_00[2], slf_op_29_00[1],
     slf_op_29_00[0], slf_op_29_00[3], slf_op_29_00[2],
     slf_op_29_00[1], slf_op_29_00[0]}), .sp12_h_l_01(net2778[0:23]),
     .sp12_h_l_02(net2777[0:23]), .sp12_h_l_03(net2776[0:23]),
     .sp12_h_l_04(net2775[0:23]), .sp4_v_b_04(net2782[0:47]),
     .sp4_v_b_03(net2783[0:47]), .sp4_v_b_02(net2784[0:47]),
     .bnr_op_01({slf_op_30_00[3], slf_op_30_00[2], slf_op_30_00[1],
     slf_op_30_00[0], slf_op_30_00[3], slf_op_30_00[2],
     slf_op_30_00[1], slf_op_30_00[0]}), .sp4_h_l_05(net2814[0:47]),
     .sp4_h_l_06(net2813[0:47]), .sp4_h_l_07(net2812[0:47]),
     .sp4_h_l_08(net2811[0:47]), .sp4_h_l_09(net2810[0:47]),
     .sp4_h_l_10(net2809[0:47]), .sp4_h_r_10(net3950[0:47]),
     .sp4_h_r_09(net3951[0:47]), .sp4_h_r_08(net3952[0:47]),
     .sp4_h_r_07(net3953[0:47]), .sp4_h_r_06(net3954[0:47]),
     .sp4_h_r_05(net3955[0:47]), .slf_op_05(net2826[0:7]),
     .slf_op_06(net2825[0:7]), .slf_op_07(net2824[0:7]),
     .slf_op_08(net2823[0:7]), .slf_op_09(net2822[0:7]),
     .slf_op_10(net2821[0:7]), .rgt_op_10(net3962[0:7]),
     .rgt_op_09(net3963[0:7]), .rgt_op_08(net3964[0:7]),
     .rgt_op_07(net3965[0:7]), .rgt_op_06(net3966[0:7]),
     .rgt_op_05(net3967[0:7]), .lft_op_10(net2984[0:7]),
     .lft_op_09(net2985[0:7]), .lft_op_08(net2986[0:7]),
     .lft_op_07(net2987[0:7]), .lft_op_06(net2988[0:7]),
     .lft_op_05(net2989[0:7]), .sp12_h_l_10(net2834[0:23]),
     .sp12_h_r_10(net3975[0:23]), .sp12_h_l_09(net2843[0:23]),
     .sp12_h_l_08(net2842[0:23]), .sp12_h_l_07(net2841[0:23]),
     .sp12_h_l_06(net2840[0:23]), .sp12_h_r_05(net3980[0:23]),
     .sp12_h_r_06(net3981[0:23]), .sp12_h_r_07(net3982[0:23]),
     .sp12_h_r_08(net3983[0:23]), .sp12_h_r_09(net3984[0:23]),
     .sp12_h_l_05(net2839[0:23]), .sp4_r_v_b_05(net3986[0:47]),
     .sp4_r_v_b_06(net3987[0:47]), .sp4_r_v_b_07(net3988[0:47]),
     .sp4_r_v_b_08(net3989[0:47]), .sp4_r_v_b_09(net3990[0:47]),
     .sp4_r_v_b_10(net3991[0:47]), .sp4_v_b_10(net2850[0:47]),
     .sp4_v_b_09(net2849[0:47]), .sp4_v_b_08(net2848[0:47]),
     .sp4_v_b_07(net2847[0:47]), .sp4_v_b_06(net2846[0:47]),
     .sp4_v_b_05(net2845[0:47]), .sp4_v_t_16(sp4_v_t_29_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net4001[0:47]), .sp4_h_r_12(net4002[0:47]),
     .sp4_h_r_13(net4003[0:47]), .sp4_h_r_14(net4004[0:47]),
     .sp4_h_r_15(net4005[0:47]), .sp4_h_r_16(net4006[0:47]),
     .sp4_h_l_16(net2865[0:47]), .sp4_h_l_15(net2864[0:47]),
     .sp4_h_l_14(net2863[0:47]), .sp4_h_l_13(net2862[0:47]),
     .sp4_h_l_12(net2861[0:47]), .sp4_h_l_11(net2860[0:47]),
     .tnr_op_16(tnr_op_29_16[7:0]), .tnl_op_16(tnl_op_29_16[7:0]),
     .lft_op_16(slf_op_28_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net2882[0:7]), .slf_op_14(net2881[0:7]),
     .slf_op_13(net2884[0:7]), .slf_op_12(net2883[0:7]),
     .slf_op_11(net2885[0:7]), .rgt_op_14(net4022[0:7]),
     .rgt_op_15(net4023[0:7]), .rgt_op_12(net4024[0:7]),
     .rgt_op_13(net4025[0:7]), .rgt_op_11(net4026[0:7]),
     .sp4_v_b_16(net2892[0:47]), .sp4_v_b_14(net2895[0:47]),
     .sp4_v_b_15(net2893[0:47]), .sp4_v_b_13(net2894[0:47]),
     .sp4_v_b_11(net2897[0:47]), .sp4_v_b_12(net2896[0:47]),
     .sp4_r_v_b_16(net4033[0:47]), .sp4_r_v_b_15(net4034[0:47]),
     .sp4_r_v_b_13(net4035[0:47]), .sp4_r_v_b_14(net4036[0:47]),
     .sp4_r_v_b_12(net4037[0:47]), .sp4_r_v_b_11(net4038[0:47]),
     .sp12_h_l_16(net2904[0:23]), .sp12_h_l_15(net2906[0:23]),
     .sp12_h_l_14(net2905[0:23]), .sp12_h_l_13(net2908[0:23]),
     .sp12_h_l_12(net2907[0:23]), .sp12_h_l_11(net2909[0:23]),
     .sp12_h_r_16(net4045[0:23]), .sp12_h_r_14(net4046[0:23]),
     .sp12_h_r_15(net4047[0:23]), .sp12_h_r_12(net4048[0:23]),
     .sp12_h_r_13(net4049[0:23]), .sp12_h_r_11(net4050[0:23]),
     .lft_op_14(net3044[0:7]), .lft_op_15(net3045[0:7]),
     .lft_op_12(net3046[0:7]), .lft_op_11(net3048[0:7]),
     .lft_op_13(net3047[0:7]));
array_LT1x16 I_lt_23_bot ( .sp12_v_b_01(net2124[0:23]),
     .glb_netwk(net2123[0:7]), .sp12_v_t_16(sp12_v_t_23_16[23:0]),
     .rgt_op_16(slf_op_24_16[7:0]), .top_op_16(top_op_23_16[7:0]),
     .rgt_op_03(net4059[0:7]), .slf_op_02(net3246[0:7]),
     .rgt_op_02(net4061[0:7]), .rgt_op_01(net2108[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2602[0:7]), .lft_op_03(net2592[0:7]),
     .lft_op_02(net2594[0:7]), .lft_op_01(net2122[0:7]),
     .rgt_op_04(net4069[0:7]), .carry_in(net2515),
     .bnl_op_01({slf_op_22_00[3], slf_op_22_00[2], slf_op_22_00[1],
     slf_op_22_00[0], slf_op_22_00[3], slf_op_22_00[2],
     slf_op_22_00[1], slf_op_22_00[0]}), .slf_op_04(net3254[0:7]),
     .slf_op_03(net3244[0:7]), .slf_op_01(net2115[0:7]),
     .sp4_h_l_04(net3275[0:47]), .carry_out(carry_out_23_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net4079[0:23]),
     .sp12_h_r_03(net4080[0:23]), .sp12_h_r_02(net4081[0:23]),
     .sp12_h_r_01(net4082[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_23_16[7:0]), .sp4_v_b_01(net2117[0:47]),
     .sp4_r_v_b_04(net4086[0:47]), .sp4_r_v_b_03(net4087[0:47]),
     .sp4_r_v_b_02(net4088[0:47]), .sp4_r_v_b_01(net2110[0:47]),
     .sp4_h_r_04(net4090[0:47]), .sp4_h_r_03(net4091[0:47]),
     .sp4_h_r_02(net4092[0:47]), .sp4_h_r_01(net4093[0:47]),
     .sp4_h_l_03(net3276[0:47]), .sp4_h_l_02(net3277[0:47]),
     .sp4_h_l_01(net3278[0:47]), .bl(bl[1251:1198]),
     .bot_op_01({slf_op_23_00[3], slf_op_23_00[2], slf_op_23_00[1],
     slf_op_23_00[0], slf_op_23_00[3], slf_op_23_00[2],
     slf_op_23_00[1], slf_op_23_00[0]}), .sp12_h_l_01(net3267[0:23]),
     .sp12_h_l_02(net3266[0:23]), .sp12_h_l_03(net3265[0:23]),
     .sp12_h_l_04(net3264[0:23]), .sp4_v_b_04(net3271[0:47]),
     .sp4_v_b_03(net3272[0:47]), .sp4_v_b_02(net3273[0:47]),
     .bnr_op_01({slf_op_24_00[3], slf_op_24_00[2], slf_op_24_00[1],
     slf_op_24_00[0], slf_op_24_00[3], slf_op_24_00[2],
     slf_op_24_00[1], slf_op_24_00[0]}), .sp4_h_l_05(net3303[0:47]),
     .sp4_h_l_06(net3302[0:47]), .sp4_h_l_07(net3301[0:47]),
     .sp4_h_l_08(net3300[0:47]), .sp4_h_l_09(net3299[0:47]),
     .sp4_h_l_10(net3298[0:47]), .sp4_h_r_10(net4113[0:47]),
     .sp4_h_r_09(net4114[0:47]), .sp4_h_r_08(net4115[0:47]),
     .sp4_h_r_07(net4116[0:47]), .sp4_h_r_06(net4117[0:47]),
     .sp4_h_r_05(net4118[0:47]), .slf_op_05(net3315[0:7]),
     .slf_op_06(net3314[0:7]), .slf_op_07(net3313[0:7]),
     .slf_op_08(net3312[0:7]), .slf_op_09(net3311[0:7]),
     .slf_op_10(net3310[0:7]), .rgt_op_10(net4125[0:7]),
     .rgt_op_09(net4126[0:7]), .rgt_op_08(net4127[0:7]),
     .rgt_op_07(net4128[0:7]), .rgt_op_06(net4129[0:7]),
     .rgt_op_05(net4130[0:7]), .lft_op_10(net2658[0:7]),
     .lft_op_09(net2659[0:7]), .lft_op_08(net2660[0:7]),
     .lft_op_07(net2661[0:7]), .lft_op_06(net2662[0:7]),
     .lft_op_05(net2663[0:7]), .sp12_h_l_10(net3323[0:23]),
     .sp12_h_r_10(net4138[0:23]), .sp12_h_l_09(net3332[0:23]),
     .sp12_h_l_08(net3331[0:23]), .sp12_h_l_07(net3330[0:23]),
     .sp12_h_l_06(net3329[0:23]), .sp12_h_r_05(net4143[0:23]),
     .sp12_h_r_06(net4144[0:23]), .sp12_h_r_07(net4145[0:23]),
     .sp12_h_r_08(net4146[0:23]), .sp12_h_r_09(net4147[0:23]),
     .sp12_h_l_05(net3328[0:23]), .sp4_r_v_b_05(net4149[0:47]),
     .sp4_r_v_b_06(net4150[0:47]), .sp4_r_v_b_07(net4151[0:47]),
     .sp4_r_v_b_08(net4152[0:47]), .sp4_r_v_b_09(net4153[0:47]),
     .sp4_r_v_b_10(net4154[0:47]), .sp4_v_b_10(net3339[0:47]),
     .sp4_v_b_09(net3338[0:47]), .sp4_v_b_08(net3337[0:47]),
     .sp4_v_b_07(net3336[0:47]), .sp4_v_b_06(net3335[0:47]),
     .sp4_v_b_05(net3334[0:47]), .sp4_v_t_16(sp4_v_t_23_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net4164[0:47]), .sp4_h_r_12(net4165[0:47]),
     .sp4_h_r_13(net4166[0:47]), .sp4_h_r_14(net4167[0:47]),
     .sp4_h_r_15(net4168[0:47]), .sp4_h_r_16(net4169[0:47]),
     .sp4_h_l_16(net3354[0:47]), .sp4_h_l_15(net3353[0:47]),
     .sp4_h_l_14(net3352[0:47]), .sp4_h_l_13(net3351[0:47]),
     .sp4_h_l_12(net3350[0:47]), .sp4_h_l_11(net3349[0:47]),
     .tnr_op_16(tnr_op_23_16[7:0]), .tnl_op_16(tnl_op_23_16[7:0]),
     .lft_op_16(slf_op_22_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net3371[0:7]), .slf_op_14(net3370[0:7]),
     .slf_op_13(net3373[0:7]), .slf_op_12(net3372[0:7]),
     .slf_op_11(net3374[0:7]), .rgt_op_14(net4185[0:7]),
     .rgt_op_15(net4186[0:7]), .rgt_op_12(net4187[0:7]),
     .rgt_op_13(net4188[0:7]), .rgt_op_11(net4189[0:7]),
     .sp4_v_b_16(net3381[0:47]), .sp4_v_b_14(net3384[0:47]),
     .sp4_v_b_15(net3382[0:47]), .sp4_v_b_13(net3383[0:47]),
     .sp4_v_b_11(net3386[0:47]), .sp4_v_b_12(net3385[0:47]),
     .sp4_r_v_b_16(net4196[0:47]), .sp4_r_v_b_15(net4197[0:47]),
     .sp4_r_v_b_13(net4198[0:47]), .sp4_r_v_b_14(net4199[0:47]),
     .sp4_r_v_b_12(net4200[0:47]), .sp4_r_v_b_11(net4201[0:47]),
     .sp12_h_l_16(net3393[0:23]), .sp12_h_l_15(net3395[0:23]),
     .sp12_h_l_14(net3394[0:23]), .sp12_h_l_13(net3397[0:23]),
     .sp12_h_l_12(net3396[0:23]), .sp12_h_l_11(net3398[0:23]),
     .sp12_h_r_16(net4208[0:23]), .sp12_h_r_14(net4209[0:23]),
     .sp12_h_r_15(net4210[0:23]), .sp12_h_r_12(net4211[0:23]),
     .sp12_h_r_13(net4212[0:23]), .sp12_h_r_11(net4213[0:23]),
     .lft_op_14(net2718[0:7]), .lft_op_15(net2719[0:7]),
     .lft_op_12(net2720[0:7]), .lft_op_11(net2722[0:7]),
     .lft_op_13(net2721[0:7]));
array_LT1x16 I_lt_30_bot ( .sp12_v_b_01(net2064[0:23]),
     .glb_netwk(net2063[0:7]), .sp12_v_t_16(sp12_v_t_30_16[23:0]),
     .rgt_op_16(slf_op_31_16[7:0]), .top_op_16(top_op_30_16[7:0]),
     .rgt_op_03(net4222[0:7]), .slf_op_02(net3898[0:7]),
     .rgt_op_02(net4224[0:7]), .rgt_op_01(net2185[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net2765[0:7]), .lft_op_03(net2755[0:7]),
     .lft_op_02(net2757[0:7]), .lft_op_01(net2062[0:7]),
     .rgt_op_04(net4232[0:7]), .carry_in(net2529),
     .bnl_op_01({slf_op_29_00[3], slf_op_29_00[2], slf_op_29_00[1],
     slf_op_29_00[0], slf_op_29_00[3], slf_op_29_00[2],
     slf_op_29_00[1], slf_op_29_00[0]}), .slf_op_04(net3906[0:7]),
     .slf_op_03(net3896[0:7]), .slf_op_01(net2047[0:7]),
     .sp4_h_l_04(net3927[0:47]), .carry_out(carry_out_30_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net4242[0:23]),
     .sp12_h_r_03(net4243[0:23]), .sp12_h_r_02(net4244[0:23]),
     .sp12_h_r_01(net4245[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_30_16[7:0]), .sp4_v_b_01(net2050[0:47]),
     .sp4_r_v_b_04(net4249[0:47]), .sp4_r_v_b_03(net4250[0:47]),
     .sp4_r_v_b_02(net4251[0:47]), .sp4_r_v_b_01(net2182[0:47]),
     .sp4_h_r_04(net4253[0:47]), .sp4_h_r_03(net4254[0:47]),
     .sp4_h_r_02(net4255[0:47]), .sp4_h_r_01(net4256[0:47]),
     .sp4_h_l_03(net3928[0:47]), .sp4_h_l_02(net3929[0:47]),
     .sp4_h_l_01(net3930[0:47]), .bl(bl[1617:1564]),
     .bot_op_01({slf_op_30_00[3], slf_op_30_00[2], slf_op_30_00[1],
     slf_op_30_00[0], slf_op_30_00[3], slf_op_30_00[2],
     slf_op_30_00[1], slf_op_30_00[0]}), .sp12_h_l_01(net3919[0:23]),
     .sp12_h_l_02(net3918[0:23]), .sp12_h_l_03(net3917[0:23]),
     .sp12_h_l_04(net3916[0:23]), .sp4_v_b_04(net3923[0:47]),
     .sp4_v_b_03(net3924[0:47]), .sp4_v_b_02(net3925[0:47]),
     .bnr_op_01({slf_op_31_00[3], slf_op_31_00[2], slf_op_31_00[1],
     slf_op_31_00[0], slf_op_31_00[3], slf_op_31_00[2],
     slf_op_31_00[1], slf_op_31_00[0]}), .sp4_h_l_05(net3955[0:47]),
     .sp4_h_l_06(net3954[0:47]), .sp4_h_l_07(net3953[0:47]),
     .sp4_h_l_08(net3952[0:47]), .sp4_h_l_09(net3951[0:47]),
     .sp4_h_l_10(net3950[0:47]), .sp4_h_r_10(net4276[0:47]),
     .sp4_h_r_09(net4277[0:47]), .sp4_h_r_08(net4278[0:47]),
     .sp4_h_r_07(net4279[0:47]), .sp4_h_r_06(net4280[0:47]),
     .sp4_h_r_05(net4281[0:47]), .slf_op_05(net3967[0:7]),
     .slf_op_06(net3966[0:7]), .slf_op_07(net3965[0:7]),
     .slf_op_08(net3964[0:7]), .slf_op_09(net3963[0:7]),
     .slf_op_10(net3962[0:7]), .rgt_op_10(net4288[0:7]),
     .rgt_op_09(net4289[0:7]), .rgt_op_08(net4290[0:7]),
     .rgt_op_07(net4291[0:7]), .rgt_op_06(net4292[0:7]),
     .rgt_op_05(net4293[0:7]), .lft_op_10(net2821[0:7]),
     .lft_op_09(net2822[0:7]), .lft_op_08(net2823[0:7]),
     .lft_op_07(net2824[0:7]), .lft_op_06(net2825[0:7]),
     .lft_op_05(net2826[0:7]), .sp12_h_l_10(net3975[0:23]),
     .sp12_h_r_10(net4301[0:23]), .sp12_h_l_09(net3984[0:23]),
     .sp12_h_l_08(net3983[0:23]), .sp12_h_l_07(net3982[0:23]),
     .sp12_h_l_06(net3981[0:23]), .sp12_h_r_05(net4306[0:23]),
     .sp12_h_r_06(net4307[0:23]), .sp12_h_r_07(net4308[0:23]),
     .sp12_h_r_08(net4309[0:23]), .sp12_h_r_09(net4310[0:23]),
     .sp12_h_l_05(net3980[0:23]), .sp4_r_v_b_05(net4312[0:47]),
     .sp4_r_v_b_06(net4313[0:47]), .sp4_r_v_b_07(net4314[0:47]),
     .sp4_r_v_b_08(net4315[0:47]), .sp4_r_v_b_09(net4316[0:47]),
     .sp4_r_v_b_10(net4317[0:47]), .sp4_v_b_10(net3991[0:47]),
     .sp4_v_b_09(net3990[0:47]), .sp4_v_b_08(net3989[0:47]),
     .sp4_v_b_07(net3988[0:47]), .sp4_v_b_06(net3987[0:47]),
     .sp4_v_b_05(net3986[0:47]), .sp4_v_t_16(sp4_v_t_30_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net4327[0:47]), .sp4_h_r_12(net4328[0:47]),
     .sp4_h_r_13(net4329[0:47]), .sp4_h_r_14(net4330[0:47]),
     .sp4_h_r_15(net4331[0:47]), .sp4_h_r_16(net4332[0:47]),
     .sp4_h_l_16(net4006[0:47]), .sp4_h_l_15(net4005[0:47]),
     .sp4_h_l_14(net4004[0:47]), .sp4_h_l_13(net4003[0:47]),
     .sp4_h_l_12(net4002[0:47]), .sp4_h_l_11(net4001[0:47]),
     .tnr_op_16(tnr_op_30_16[7:0]), .tnl_op_16(tnl_op_30_16[7:0]),
     .lft_op_16(slf_op_29_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net4023[0:7]), .slf_op_14(net4022[0:7]),
     .slf_op_13(net4025[0:7]), .slf_op_12(net4024[0:7]),
     .slf_op_11(net4026[0:7]), .rgt_op_14(net4348[0:7]),
     .rgt_op_15(net4349[0:7]), .rgt_op_12(net4350[0:7]),
     .rgt_op_13(net4351[0:7]), .rgt_op_11(net4352[0:7]),
     .sp4_v_b_16(net4033[0:47]), .sp4_v_b_14(net4036[0:47]),
     .sp4_v_b_15(net4034[0:47]), .sp4_v_b_13(net4035[0:47]),
     .sp4_v_b_11(net4038[0:47]), .sp4_v_b_12(net4037[0:47]),
     .sp4_r_v_b_16(net4359[0:47]), .sp4_r_v_b_15(net4360[0:47]),
     .sp4_r_v_b_13(net4361[0:47]), .sp4_r_v_b_14(net4362[0:47]),
     .sp4_r_v_b_12(net4363[0:47]), .sp4_r_v_b_11(net4364[0:47]),
     .sp12_h_l_16(net4045[0:23]), .sp12_h_l_15(net4047[0:23]),
     .sp12_h_l_14(net4046[0:23]), .sp12_h_l_13(net4049[0:23]),
     .sp12_h_l_12(net4048[0:23]), .sp12_h_l_11(net4050[0:23]),
     .sp12_h_r_16(net4371[0:23]), .sp12_h_r_14(net4372[0:23]),
     .sp12_h_r_15(net4373[0:23]), .sp12_h_r_12(net4374[0:23]),
     .sp12_h_r_13(net4375[0:23]), .sp12_h_r_11(net4376[0:23]),
     .lft_op_14(net2881[0:7]), .lft_op_15(net2882[0:7]),
     .lft_op_12(net2883[0:7]), .lft_op_11(net2885[0:7]),
     .lft_op_13(net2884[0:7]));
array_LT1x16 I_lt_26_bot ( .sp12_v_b_01(net2103[0:23]),
     .glb_netwk(net2102[0:7]), .sp12_v_t_16(sp12_v_t_26_16[23:0]),
     .rgt_op_16(slf_op_27_16[7:0]), .top_op_16(top_op_26_16[7:0]),
     .rgt_op_03(net4385[0:7]), .slf_op_02(net2431[0:7]),
     .rgt_op_02(net4387[0:7]), .rgt_op_01(net2087[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net3580[0:7]), .lft_op_03(net3570[0:7]),
     .lft_op_02(net3572[0:7]), .lft_op_01(net2101[0:7]),
     .rgt_op_04(net4395[0:7]), .carry_in(net2516),
     .bnl_op_01({slf_op_25_00[3], slf_op_25_00[2], slf_op_25_00[1],
     slf_op_25_00[0], slf_op_25_00[3], slf_op_25_00[2],
     slf_op_25_00[1], slf_op_25_00[0]}), .slf_op_04(net2433[0:7]),
     .slf_op_03(net2432[0:7]), .slf_op_01(net2177[0:7]),
     .sp4_h_l_04(net2452[0:47]), .carry_out(carry_out_26_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net4405[0:23]),
     .sp12_h_r_03(net4406[0:23]), .sp12_h_r_02(net4407[0:23]),
     .sp12_h_r_01(net4408[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_26_16[7:0]), .sp4_v_b_01(net2096[0:47]),
     .sp4_r_v_b_04(net4412[0:47]), .sp4_r_v_b_03(net4413[0:47]),
     .sp4_r_v_b_02(net4414[0:47]), .sp4_r_v_b_01(net2092[0:47]),
     .sp4_h_r_04(net4416[0:47]), .sp4_h_r_03(net4417[0:47]),
     .sp4_h_r_02(net4418[0:47]), .sp4_h_r_01(net4419[0:47]),
     .sp4_h_l_03(net2451[0:47]), .sp4_h_l_02(net2450[0:47]),
     .sp4_h_l_01(net2449[0:47]), .bl(bl[1401:1348]),
     .bot_op_01({slf_op_26_00[3], slf_op_26_00[2], slf_op_26_00[1],
     slf_op_26_00[0], slf_op_26_00[3], slf_op_26_00[2],
     slf_op_26_00[1], slf_op_26_00[0]}), .sp12_h_l_01(net2329[0:23]),
     .sp12_h_l_02(net2409[0:23]), .sp12_h_l_03(net2408[0:23]),
     .sp12_h_l_04(net2407[0:23]), .sp4_v_b_04(net2346[0:47]),
     .sp4_v_b_03(net2345[0:47]), .sp4_v_b_02(net2344[0:47]),
     .bnr_op_01({slf_op_27_00[3], slf_op_27_00[2], slf_op_27_00[1],
     slf_op_27_00[0], slf_op_27_00[3], slf_op_27_00[2],
     slf_op_27_00[1], slf_op_27_00[0]}), .sp4_h_l_05(net2453[0:47]),
     .sp4_h_l_06(net2454[0:47]), .sp4_h_l_07(net2455[0:47]),
     .sp4_h_l_08(net2456[0:47]), .sp4_h_l_09(net2341[0:47]),
     .sp4_h_l_10(net2457[0:47]), .sp4_h_r_10(net4439[0:47]),
     .sp4_h_r_09(net4440[0:47]), .sp4_h_r_08(net4441[0:47]),
     .sp4_h_r_07(net4442[0:47]), .sp4_h_r_06(net4443[0:47]),
     .sp4_h_r_05(net4444[0:47]), .slf_op_05(net2434[0:7]),
     .slf_op_06(net2435[0:7]), .slf_op_07(net2436[0:7]),
     .slf_op_08(net2437[0:7]), .slf_op_09(net2438[0:7]),
     .slf_op_10(net2439[0:7]), .rgt_op_10(net4451[0:7]),
     .rgt_op_09(net4452[0:7]), .rgt_op_08(net4453[0:7]),
     .rgt_op_07(net4454[0:7]), .rgt_op_06(net4455[0:7]),
     .rgt_op_05(net4456[0:7]), .lft_op_10(net3636[0:7]),
     .lft_op_09(net3637[0:7]), .lft_op_08(net3638[0:7]),
     .lft_op_07(net3639[0:7]), .lft_op_06(net3640[0:7]),
     .lft_op_05(net3641[0:7]), .sp12_h_l_10(net2389[0:23]),
     .sp12_h_r_10(net4464[0:23]), .sp12_h_l_09(net2402[0:23]),
     .sp12_h_l_08(net2403[0:23]), .sp12_h_l_07(net2404[0:23]),
     .sp12_h_l_06(net2405[0:23]), .sp12_h_r_05(net4469[0:23]),
     .sp12_h_r_06(net4470[0:23]), .sp12_h_r_07(net4471[0:23]),
     .sp12_h_r_08(net4472[0:23]), .sp12_h_r_09(net4473[0:23]),
     .sp12_h_l_05(net2406[0:23]), .sp4_r_v_b_05(net4475[0:47]),
     .sp4_r_v_b_06(net4476[0:47]), .sp4_r_v_b_07(net4477[0:47]),
     .sp4_r_v_b_08(net4478[0:47]), .sp4_r_v_b_09(net4479[0:47]),
     .sp4_r_v_b_10(net4480[0:47]), .sp4_v_b_10(net2352[0:47]),
     .sp4_v_b_09(net2351[0:47]), .sp4_v_b_08(net2350[0:47]),
     .sp4_v_b_07(net2349[0:47]), .sp4_v_b_06(net2348[0:47]),
     .sp4_v_b_05(net2347[0:47]), .sp4_v_t_16(sp4_v_t_26_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net4490[0:47]), .sp4_h_r_12(net4491[0:47]),
     .sp4_h_r_13(net4492[0:47]), .sp4_h_r_14(net4493[0:47]),
     .sp4_h_r_15(net4494[0:47]), .sp4_h_r_16(net4495[0:47]),
     .sp4_h_l_16(net2463[0:47]), .sp4_h_l_15(net2462[0:47]),
     .sp4_h_l_14(net2461[0:47]), .sp4_h_l_13(net2460[0:47]),
     .sp4_h_l_12(net2459[0:47]), .sp4_h_l_11(net2458[0:47]),
     .tnr_op_16(tnr_op_26_16[7:0]), .tnl_op_16(tnl_op_26_16[7:0]),
     .lft_op_16(slf_op_25_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net2444[0:7]), .slf_op_14(net2443[0:7]),
     .slf_op_13(net2442[0:7]), .slf_op_12(net2441[0:7]),
     .slf_op_11(net2440[0:7]), .rgt_op_14(net4511[0:7]),
     .rgt_op_15(net4512[0:7]), .rgt_op_12(net4513[0:7]),
     .rgt_op_13(net4514[0:7]), .rgt_op_11(net4515[0:7]),
     .sp4_v_b_16(net2357[0:47]), .sp4_v_b_14(net2356[0:47]),
     .sp4_v_b_15(net2358[0:47]), .sp4_v_b_13(net2355[0:47]),
     .sp4_v_b_11(net2353[0:47]), .sp4_v_b_12(net2354[0:47]),
     .sp4_r_v_b_16(net4522[0:47]), .sp4_r_v_b_15(net4523[0:47]),
     .sp4_r_v_b_13(net4524[0:47]), .sp4_r_v_b_14(net4525[0:47]),
     .sp4_r_v_b_12(net4526[0:47]), .sp4_r_v_b_11(net4527[0:47]),
     .sp12_h_l_16(net2394[0:23]), .sp12_h_l_15(net2390[0:23]),
     .sp12_h_l_14(net2393[0:23]), .sp12_h_l_13(net2399[0:23]),
     .sp12_h_l_12(net2400[0:23]), .sp12_h_l_11(net2401[0:23]),
     .sp12_h_r_16(net4534[0:23]), .sp12_h_r_14(net4535[0:23]),
     .sp12_h_r_15(net4536[0:23]), .sp12_h_r_12(net4537[0:23]),
     .sp12_h_r_13(net4538[0:23]), .sp12_h_r_11(net4539[0:23]),
     .lft_op_14(net3696[0:7]), .lft_op_15(net3697[0:7]),
     .lft_op_12(net3698[0:7]), .lft_op_11(net3700[0:7]),
     .lft_op_13(net3699[0:7]));
array_LT1x16 I_lt_18_bot ( .sp12_v_b_01(net2172[0:23]),
     .glb_netwk(net2171[0:7]), .sp12_v_t_16(sp12_v_t_18_16[23:0]),
     .rgt_op_16(slf_op_19_16[7:0]), .top_op_16(top_op_18_16[7:0]),
     .rgt_op_03(net4548[0:7]), .slf_op_02(net4713[0:7]),
     .rgt_op_02(net4550[0:7]), .rgt_op_01(net2146[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(slf_op_17_04[7:0]),
     .lft_op_03(slf_op_17_03[7:0]), .lft_op_02(slf_op_17_02[7:0]),
     .lft_op_01(slf_op_17_01[7:0]), .rgt_op_04(net4558[0:7]),
     .carry_in(net2532), .bnl_op_01({slf_op_17_00[3], slf_op_17_00[2],
     slf_op_17_00[1], slf_op_17_00[0], slf_op_17_00[3],
     slf_op_17_00[2], slf_op_17_00[1], slf_op_17_00[0]}),
     .slf_op_04(net4721[0:7]), .slf_op_03(net4711[0:7]),
     .slf_op_01(net2154[0:7]), .sp4_h_l_04(net4742[0:47]),
     .carry_out(carry_out_18_16), .vdd_cntl(vdd_cntl_r[271:16]),
     .sp12_h_r_04(net4568[0:23]), .sp12_h_r_03(net4569[0:23]),
     .sp12_h_r_02(net4570[0:23]), .sp12_h_r_01(net4571[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(slf_op_18_16[7:0]),
     .sp4_v_b_01(net2165[0:47]), .sp4_r_v_b_04(net4575[0:47]),
     .sp4_r_v_b_03(net4576[0:47]), .sp4_r_v_b_02(net4577[0:47]),
     .sp4_r_v_b_01(net2149[0:47]), .sp4_h_r_04(net4579[0:47]),
     .sp4_h_r_03(net4580[0:47]), .sp4_h_r_02(net4581[0:47]),
     .sp4_h_r_01(net4582[0:47]), .sp4_h_l_03(net4743[0:47]),
     .sp4_h_l_02(net4744[0:47]), .sp4_h_l_01(net4745[0:47]),
     .bl(bl[981:928]), .bot_op_01({slf_op_18_00[3], slf_op_18_00[2],
     slf_op_18_00[1], slf_op_18_00[0], slf_op_18_00[3],
     slf_op_18_00[2], slf_op_18_00[1], slf_op_18_00[0]}),
     .sp12_h_l_01(net4734[0:23]), .sp12_h_l_02(net4733[0:23]),
     .sp12_h_l_03(net4732[0:23]), .sp12_h_l_04(net4731[0:23]),
     .sp4_v_b_04(net4738[0:47]), .sp4_v_b_03(net4739[0:47]),
     .sp4_v_b_02(net4740[0:47]), .bnr_op_01({slf_op_19_00[3],
     slf_op_19_00[2], slf_op_19_00[1], slf_op_19_00[0],
     slf_op_19_00[3], slf_op_19_00[2], slf_op_19_00[1],
     slf_op_19_00[0]}), .sp4_h_l_05(net4770[0:47]),
     .sp4_h_l_06(net4769[0:47]), .sp4_h_l_07(net4768[0:47]),
     .sp4_h_l_08(net4767[0:47]), .sp4_h_l_09(net4766[0:47]),
     .sp4_h_l_10(net4765[0:47]), .sp4_h_r_10(net4602[0:47]),
     .sp4_h_r_09(net4603[0:47]), .sp4_h_r_08(net4604[0:47]),
     .sp4_h_r_07(net4605[0:47]), .sp4_h_r_06(net4606[0:47]),
     .sp4_h_r_05(net4607[0:47]), .slf_op_05(net4782[0:7]),
     .slf_op_06(net4781[0:7]), .slf_op_07(net4780[0:7]),
     .slf_op_08(net4779[0:7]), .slf_op_09(net4778[0:7]),
     .slf_op_10(net4777[0:7]), .rgt_op_10(net4614[0:7]),
     .rgt_op_09(net4615[0:7]), .rgt_op_08(net4616[0:7]),
     .rgt_op_07(net4617[0:7]), .rgt_op_06(net4618[0:7]),
     .rgt_op_05(net4619[0:7]), .lft_op_10(slf_op_17_10[7:0]),
     .lft_op_09(slf_op_17_09[7:0]), .lft_op_08(slf_op_17_08[7:0]),
     .lft_op_07(slf_op_17_07[7:0]), .lft_op_06(slf_op_17_06[7:0]),
     .lft_op_05(slf_op_17_05[7:0]), .sp12_h_l_10(net4790[0:23]),
     .sp12_h_r_10(net4627[0:23]), .sp12_h_l_09(net4799[0:23]),
     .sp12_h_l_08(net4798[0:23]), .sp12_h_l_07(net4797[0:23]),
     .sp12_h_l_06(net4796[0:23]), .sp12_h_r_05(net4632[0:23]),
     .sp12_h_r_06(net4633[0:23]), .sp12_h_r_07(net4634[0:23]),
     .sp12_h_r_08(net4635[0:23]), .sp12_h_r_09(net4636[0:23]),
     .sp12_h_l_05(net4795[0:23]), .sp4_r_v_b_05(net4638[0:47]),
     .sp4_r_v_b_06(net4639[0:47]), .sp4_r_v_b_07(net4640[0:47]),
     .sp4_r_v_b_08(net4641[0:47]), .sp4_r_v_b_09(net4642[0:47]),
     .sp4_r_v_b_10(net4643[0:47]), .sp4_v_b_10(net4806[0:47]),
     .sp4_v_b_09(net4805[0:47]), .sp4_v_b_08(net4804[0:47]),
     .sp4_v_b_07(net4803[0:47]), .sp4_v_b_06(net4802[0:47]),
     .sp4_v_b_05(net4801[0:47]), .sp4_v_t_16(sp4_v_t_18_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net4653[0:47]), .sp4_h_r_12(net4654[0:47]),
     .sp4_h_r_13(net4655[0:47]), .sp4_h_r_14(net4656[0:47]),
     .sp4_h_r_15(net4657[0:47]), .sp4_h_r_16(sp4_h_r_18_19[47:0]),
     .sp4_h_l_16(sp4_h_r_17_18[47:0]), .sp4_h_l_15(net4820[0:47]),
     .sp4_h_l_14(net4819[0:47]), .sp4_h_l_13(net4818[0:47]),
     .sp4_h_l_12(net4817[0:47]), .sp4_h_l_11(net4816[0:47]),
     .tnr_op_16(tnr_op_18_16[7:0]), .tnl_op_16(tnl_op_18_16[7:0]),
     .lft_op_16(slf_op_17_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net4838[0:7]), .slf_op_14(net4837[0:7]),
     .slf_op_13(net4840[0:7]), .slf_op_12(net4839[0:7]),
     .slf_op_11(net4841[0:7]), .rgt_op_14(net4674[0:7]),
     .rgt_op_15(net4675[0:7]), .rgt_op_12(net4676[0:7]),
     .rgt_op_13(net4677[0:7]), .rgt_op_11(net4678[0:7]),
     .sp4_v_b_16(net4848[0:47]), .sp4_v_b_14(net4851[0:47]),
     .sp4_v_b_15(net4849[0:47]), .sp4_v_b_13(net4850[0:47]),
     .sp4_v_b_11(net4853[0:47]), .sp4_v_b_12(net4852[0:47]),
     .sp4_r_v_b_16(net4685[0:47]), .sp4_r_v_b_15(net4686[0:47]),
     .sp4_r_v_b_13(net4687[0:47]), .sp4_r_v_b_14(net4688[0:47]),
     .sp4_r_v_b_12(net4689[0:47]), .sp4_r_v_b_11(net4690[0:47]),
     .sp12_h_l_16(net4860[0:23]), .sp12_h_l_15(net4862[0:23]),
     .sp12_h_l_14(net4861[0:23]), .sp12_h_l_13(net4864[0:23]),
     .sp12_h_l_12(net4863[0:23]), .sp12_h_l_11(net4865[0:23]),
     .sp12_h_r_16(net4697[0:23]), .sp12_h_r_14(net4698[0:23]),
     .sp12_h_r_15(net4699[0:23]), .sp12_h_r_12(net4700[0:23]),
     .sp12_h_r_13(net4701[0:23]), .sp12_h_r_11(net4702[0:23]),
     .lft_op_14(slf_op_17_14[7:0]), .lft_op_15(slf_op_17_15[7:0]),
     .lft_op_12(slf_op_17_12[7:0]), .lft_op_11(slf_op_17_11[7:0]),
     .lft_op_13(slf_op_17_13[7:0]));
array_LT1x16 I_lt_17_bot ( .sp12_v_b_01(net2164[0:23]),
     .glb_netwk(net2163[0:7]), .sp12_v_t_16(sp12_v_t_17_16[23:0]),
     .rgt_op_16(slf_op_18_16[7:0]), .top_op_16(top_op_17_16[7:0]),
     .rgt_op_03(net4711[0:7]), .slf_op_02(slf_op_17_02[7:0]),
     .rgt_op_02(net4713[0:7]), .rgt_op_01(net2154[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(lft_op_17_04[7:0]),
     .lft_op_03(lft_op_17_03[7:0]), .lft_op_02(lft_op_17_02[7:0]),
     .lft_op_01(lft_op_17_01[7:0]), .rgt_op_04(net4721[0:7]),
     .carry_in(net2534), .bnl_op_01({bnl_op_17_01[3], bnl_op_17_01[2],
     bnl_op_17_01[1], bnl_op_17_01[0], bnl_op_17_01[3],
     bnl_op_17_01[2], bnl_op_17_01[1], bnl_op_17_01[0]}),
     .slf_op_04(slf_op_17_04[7:0]), .slf_op_03(slf_op_17_03[7:0]),
     .slf_op_01(slf_op_17_01[7:0]), .sp4_h_l_04(sp4_h_l_17_04[47:0]),
     .carry_out(carry_out_17_16), .vdd_cntl(vdd_cntl_r[271:16]),
     .sp12_h_r_04(net4731[0:23]), .sp12_h_r_03(net4732[0:23]),
     .sp12_h_r_02(net4733[0:23]), .sp12_h_r_01(net4734[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(slf_op_17_16[7:0]),
     .sp4_v_b_01(sp4_v_b_17_01[47:0]), .sp4_r_v_b_04(net4738[0:47]),
     .sp4_r_v_b_03(net4739[0:47]), .sp4_r_v_b_02(net4740[0:47]),
     .sp4_r_v_b_01(net2165[0:47]), .sp4_h_r_04(net4742[0:47]),
     .sp4_h_r_03(net4743[0:47]), .sp4_h_r_02(net4744[0:47]),
     .sp4_h_r_01(net4745[0:47]), .sp4_h_l_03(sp4_h_l_17_03[47:0]),
     .sp4_h_l_02(sp4_h_l_17_02[47:0]),
     .sp4_h_l_01(sp4_h_l_17_01[47:0]), .bl(bl[927:874]),
     .bot_op_01({slf_op_17_00[3], slf_op_17_00[2], slf_op_17_00[1],
     slf_op_17_00[0], slf_op_17_00[3], slf_op_17_00[2],
     slf_op_17_00[1], slf_op_17_00[0]}),
     .sp12_h_l_01(sp12_h_l_17_01[23:0]),
     .sp12_h_l_02(sp12_h_l_17_02[23:0]),
     .sp12_h_l_03(sp12_h_l_17_03[23:0]),
     .sp12_h_l_04(sp12_h_l_17_04[23:0]),
     .sp4_v_b_04(sp4_v_b_17_04[47:0]),
     .sp4_v_b_03(sp4_v_b_17_03[47:0]),
     .sp4_v_b_02(sp4_v_b_17_02[47:0]), .bnr_op_01({slf_op_18_00[3],
     slf_op_18_00[2], slf_op_18_00[1], slf_op_18_00[0],
     slf_op_18_00[3], slf_op_18_00[2], slf_op_18_00[1],
     slf_op_18_00[0]}), .sp4_h_l_05(sp4_h_l_17_05[47:0]),
     .sp4_h_l_06(sp4_h_l_17_06[47:0]),
     .sp4_h_l_07(sp4_h_l_17_07[47:0]),
     .sp4_h_l_08(sp4_h_l_17_08[47:0]),
     .sp4_h_l_09(sp4_h_l_17_09[47:0]),
     .sp4_h_l_10(sp4_h_l_17_10[47:0]), .sp4_h_r_10(net4765[0:47]),
     .sp4_h_r_09(net4766[0:47]), .sp4_h_r_08(net4767[0:47]),
     .sp4_h_r_07(net4768[0:47]), .sp4_h_r_06(net4769[0:47]),
     .sp4_h_r_05(net4770[0:47]), .slf_op_05(slf_op_17_05[7:0]),
     .slf_op_06(slf_op_17_06[7:0]), .slf_op_07(slf_op_17_07[7:0]),
     .slf_op_08(slf_op_17_08[7:0]), .slf_op_09(slf_op_17_09[7:0]),
     .slf_op_10(slf_op_17_10[7:0]), .rgt_op_10(net4777[0:7]),
     .rgt_op_09(net4778[0:7]), .rgt_op_08(net4779[0:7]),
     .rgt_op_07(net4780[0:7]), .rgt_op_06(net4781[0:7]),
     .rgt_op_05(net4782[0:7]), .lft_op_10(lft_op_17_10[7:0]),
     .lft_op_09(lft_op_17_09[7:0]), .lft_op_08(lft_op_17_08[7:0]),
     .lft_op_07(lft_op_17_07[7:0]), .lft_op_06(lft_op_17_06[7:0]),
     .lft_op_05(lft_op_17_05[7:0]), .sp12_h_l_10(sp12_h_l_17_10[23:0]),
     .sp12_h_r_10(net4790[0:23]), .sp12_h_l_09(sp12_h_l_17_09[23:0]),
     .sp12_h_l_08(sp12_h_l_17_08[23:0]),
     .sp12_h_l_07(sp12_h_l_17_07[23:0]),
     .sp12_h_l_06(sp12_h_l_17_06[23:0]), .sp12_h_r_05(net4795[0:23]),
     .sp12_h_r_06(net4796[0:23]), .sp12_h_r_07(net4797[0:23]),
     .sp12_h_r_08(net4798[0:23]), .sp12_h_r_09(net4799[0:23]),
     .sp12_h_l_05(sp12_h_l_17_05[23:0]), .sp4_r_v_b_05(net4801[0:47]),
     .sp4_r_v_b_06(net4802[0:47]), .sp4_r_v_b_07(net4803[0:47]),
     .sp4_r_v_b_08(net4804[0:47]), .sp4_r_v_b_09(net4805[0:47]),
     .sp4_r_v_b_10(net4806[0:47]), .sp4_v_b_10(sp4_v_b_17_10[47:0]),
     .sp4_v_b_09(sp4_v_b_17_09[47:0]),
     .sp4_v_b_08(sp4_v_b_17_08[47:0]),
     .sp4_v_b_07(sp4_v_b_17_07[47:0]),
     .sp4_v_b_06(sp4_v_b_17_06[47:0]),
     .sp4_v_b_05(sp4_v_b_17_05[47:0]),
     .sp4_v_t_16(sp4_v_t_17_16[47:0]), .pgate(pgate_r[271:16]),
     .reset_b(reset_r[271:16]), .sp4_h_r_11(net4816[0:47]),
     .sp4_h_r_12(net4817[0:47]), .sp4_h_r_13(net4818[0:47]),
     .sp4_h_r_14(net4819[0:47]), .sp4_h_r_15(net4820[0:47]),
     .sp4_h_r_16(sp4_h_r_17_18[47:0]),
     .sp4_h_l_16(sp4_h_l_17_16[47:0]),
     .sp4_h_l_15(sp4_h_l_17_15[47:0]),
     .sp4_h_l_14(sp4_h_l_17_14[47:0]),
     .sp4_h_l_13(sp4_h_l_17_13[47:0]),
     .sp4_h_l_12(sp4_h_l_17_12[47:0]),
     .sp4_h_l_11(sp4_h_l_17_11[47:0]), .tnr_op_16(tnr_op_17_16[7:0]),
     .tnl_op_16(tnl_op_17_16[7:0]), .lft_op_16(lft_op_17_16[7:0]),
     .wl(wl_r[271:16]), .slf_op_15(slf_op_17_15[7:0]),
     .slf_op_14(slf_op_17_14[7:0]), .slf_op_13(slf_op_17_13[7:0]),
     .slf_op_12(slf_op_17_12[7:0]), .slf_op_11(slf_op_17_11[7:0]),
     .rgt_op_14(net4837[0:7]), .rgt_op_15(net4838[0:7]),
     .rgt_op_12(net4839[0:7]), .rgt_op_13(net4840[0:7]),
     .rgt_op_11(net4841[0:7]), .sp4_v_b_16(sp4_v_b_17_16[47:0]),
     .sp4_v_b_14(sp4_v_b_17_14[47:0]),
     .sp4_v_b_15(sp4_v_b_17_15[47:0]),
     .sp4_v_b_13(sp4_v_b_17_13[47:0]),
     .sp4_v_b_11(sp4_v_b_17_11[47:0]),
     .sp4_v_b_12(sp4_v_b_17_12[47:0]), .sp4_r_v_b_16(net4848[0:47]),
     .sp4_r_v_b_15(net4849[0:47]), .sp4_r_v_b_13(net4850[0:47]),
     .sp4_r_v_b_14(net4851[0:47]), .sp4_r_v_b_12(net4852[0:47]),
     .sp4_r_v_b_11(net4853[0:47]), .sp12_h_l_16(sp12_h_l_17_16[23:0]),
     .sp12_h_l_15(sp12_h_l_17_15[23:0]),
     .sp12_h_l_14(sp12_h_l_17_14[23:0]),
     .sp12_h_l_13(sp12_h_l_17_13[23:0]),
     .sp12_h_l_12(sp12_h_l_17_12[23:0]),
     .sp12_h_l_11(sp12_h_l_17_11[23:0]), .sp12_h_r_16(net4860[0:23]),
     .sp12_h_r_14(net4861[0:23]), .sp12_h_r_15(net4862[0:23]),
     .sp12_h_r_12(net4863[0:23]), .sp12_h_r_13(net4864[0:23]),
     .sp12_h_r_11(net4865[0:23]), .lft_op_14(lft_op_17_14[7:0]),
     .lft_op_15(lft_op_17_15[7:0]), .lft_op_12(lft_op_17_12[7:0]),
     .lft_op_11(lft_op_17_11[7:0]), .lft_op_13(lft_op_17_13[7:0]));
array_LT1x16 I_lt_20_bot ( .sp12_v_b_01(net2148[0:23]),
     .glb_netwk(net2147[0:7]), .sp12_v_t_16(sp12_v_t_20_16[23:0]),
     .rgt_op_16(slf_op_21_16[7:0]), .top_op_16(top_op_20_16[7:0]),
     .rgt_op_03(net4874[0:7]), .slf_op_02(net3409[0:7]),
     .rgt_op_02(net4876[0:7]), .rgt_op_01(net2130[0:7]), .purst(purst),
     .prog(prog), .lft_op_04(net4558[0:7]), .lft_op_03(net4548[0:7]),
     .lft_op_02(net4550[0:7]), .lft_op_01(net2146[0:7]),
     .rgt_op_04(net4884[0:7]), .carry_in(net2514),
     .bnl_op_01({slf_op_19_00[3], slf_op_19_00[2], slf_op_19_00[1],
     slf_op_19_00[0], slf_op_19_00[3], slf_op_19_00[2],
     slf_op_19_00[1], slf_op_19_00[0]}), .slf_op_04(net3417[0:7]),
     .slf_op_03(net3407[0:7]), .slf_op_01(net2138[0:7]),
     .sp4_h_l_04(net3438[0:47]), .carry_out(carry_out_20_16),
     .vdd_cntl(vdd_cntl_r[271:16]), .sp12_h_r_04(net4894[0:23]),
     .sp12_h_r_03(net4895[0:23]), .sp12_h_r_02(net4896[0:23]),
     .sp12_h_r_01(net4897[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(slf_op_20_16[7:0]), .sp4_v_b_01(net2141[0:47]),
     .sp4_r_v_b_04(net4901[0:47]), .sp4_r_v_b_03(net4902[0:47]),
     .sp4_r_v_b_02(net4903[0:47]), .sp4_r_v_b_01(net2133[0:47]),
     .sp4_h_r_04(net4905[0:47]), .sp4_h_r_03(net4906[0:47]),
     .sp4_h_r_02(net4907[0:47]), .sp4_h_r_01(net4908[0:47]),
     .sp4_h_l_03(net3439[0:47]), .sp4_h_l_02(net3440[0:47]),
     .sp4_h_l_01(net3441[0:47]), .bl(bl[1089:1036]),
     .bot_op_01({slf_op_20_00[3], slf_op_20_00[2], slf_op_20_00[1],
     slf_op_20_00[0], slf_op_20_00[3], slf_op_20_00[2],
     slf_op_20_00[1], slf_op_20_00[0]}), .sp12_h_l_01(net3430[0:23]),
     .sp12_h_l_02(net3429[0:23]), .sp12_h_l_03(net3428[0:23]),
     .sp12_h_l_04(net3427[0:23]), .sp4_v_b_04(net3434[0:47]),
     .sp4_v_b_03(net3435[0:47]), .sp4_v_b_02(net3436[0:47]),
     .bnr_op_01({slf_op_21_00[3], slf_op_21_00[2], slf_op_21_00[1],
     slf_op_21_00[0], slf_op_21_00[3], slf_op_21_00[2],
     slf_op_21_00[1], slf_op_21_00[0]}), .sp4_h_l_05(net3466[0:47]),
     .sp4_h_l_06(net3465[0:47]), .sp4_h_l_07(net3464[0:47]),
     .sp4_h_l_08(net3463[0:47]), .sp4_h_l_09(net3462[0:47]),
     .sp4_h_l_10(net3461[0:47]), .sp4_h_r_10(net4928[0:47]),
     .sp4_h_r_09(net4929[0:47]), .sp4_h_r_08(net4930[0:47]),
     .sp4_h_r_07(net4931[0:47]), .sp4_h_r_06(net4932[0:47]),
     .sp4_h_r_05(net4933[0:47]), .slf_op_05(net3478[0:7]),
     .slf_op_06(net3477[0:7]), .slf_op_07(net3476[0:7]),
     .slf_op_08(net3475[0:7]), .slf_op_09(net3474[0:7]),
     .slf_op_10(net3473[0:7]), .rgt_op_10(net4940[0:7]),
     .rgt_op_09(net4941[0:7]), .rgt_op_08(net4942[0:7]),
     .rgt_op_07(net4943[0:7]), .rgt_op_06(net4944[0:7]),
     .rgt_op_05(net4945[0:7]), .lft_op_10(net4614[0:7]),
     .lft_op_09(net4615[0:7]), .lft_op_08(net4616[0:7]),
     .lft_op_07(net4617[0:7]), .lft_op_06(net4618[0:7]),
     .lft_op_05(net4619[0:7]), .sp12_h_l_10(net3486[0:23]),
     .sp12_h_r_10(net4953[0:23]), .sp12_h_l_09(net3495[0:23]),
     .sp12_h_l_08(net3494[0:23]), .sp12_h_l_07(net3493[0:23]),
     .sp12_h_l_06(net3492[0:23]), .sp12_h_r_05(net4958[0:23]),
     .sp12_h_r_06(net4959[0:23]), .sp12_h_r_07(net4960[0:23]),
     .sp12_h_r_08(net4961[0:23]), .sp12_h_r_09(net4962[0:23]),
     .sp12_h_l_05(net3491[0:23]), .sp4_r_v_b_05(net4964[0:47]),
     .sp4_r_v_b_06(net4965[0:47]), .sp4_r_v_b_07(net4966[0:47]),
     .sp4_r_v_b_08(net4967[0:47]), .sp4_r_v_b_09(net4968[0:47]),
     .sp4_r_v_b_10(net4969[0:47]), .sp4_v_b_10(net3502[0:47]),
     .sp4_v_b_09(net3501[0:47]), .sp4_v_b_08(net3500[0:47]),
     .sp4_v_b_07(net3499[0:47]), .sp4_v_b_06(net3498[0:47]),
     .sp4_v_b_05(net3497[0:47]), .sp4_v_t_16(sp4_v_t_20_16[47:0]),
     .pgate(pgate_r[271:16]), .reset_b(reset_r[271:16]),
     .sp4_h_r_11(net4979[0:47]), .sp4_h_r_12(net4980[0:47]),
     .sp4_h_r_13(net4981[0:47]), .sp4_h_r_14(net4982[0:47]),
     .sp4_h_r_15(net4983[0:47]), .sp4_h_r_16(sp4_h_r_20_21[47:0]),
     .sp4_h_l_16(sp4_h_r_19_20[47:0]), .sp4_h_l_15(net3516[0:47]),
     .sp4_h_l_14(net3515[0:47]), .sp4_h_l_13(net3514[0:47]),
     .sp4_h_l_12(net3513[0:47]), .sp4_h_l_11(net3512[0:47]),
     .tnr_op_16(tnr_op_20_16[7:0]), .tnl_op_16(tnl_op_20_16[7:0]),
     .lft_op_16(slf_op_19_16[7:0]), .wl(wl_r[271:16]),
     .slf_op_15(net3534[0:7]), .slf_op_14(net3533[0:7]),
     .slf_op_13(net3536[0:7]), .slf_op_12(net3535[0:7]),
     .slf_op_11(net3537[0:7]), .rgt_op_14(net5000[0:7]),
     .rgt_op_15(net5001[0:7]), .rgt_op_12(net5002[0:7]),
     .rgt_op_13(net5003[0:7]), .rgt_op_11(net5004[0:7]),
     .sp4_v_b_16(net3544[0:47]), .sp4_v_b_14(net3547[0:47]),
     .sp4_v_b_15(net3545[0:47]), .sp4_v_b_13(net3546[0:47]),
     .sp4_v_b_11(net3549[0:47]), .sp4_v_b_12(net3548[0:47]),
     .sp4_r_v_b_16(net5011[0:47]), .sp4_r_v_b_15(net5012[0:47]),
     .sp4_r_v_b_13(net5013[0:47]), .sp4_r_v_b_14(net5014[0:47]),
     .sp4_r_v_b_12(net5015[0:47]), .sp4_r_v_b_11(net5016[0:47]),
     .sp12_h_l_16(net3556[0:23]), .sp12_h_l_15(net3558[0:23]),
     .sp12_h_l_14(net3557[0:23]), .sp12_h_l_13(net3560[0:23]),
     .sp12_h_l_12(net3559[0:23]), .sp12_h_l_11(net3561[0:23]),
     .sp12_h_r_16(net5023[0:23]), .sp12_h_r_14(net5024[0:23]),
     .sp12_h_r_15(net5025[0:23]), .sp12_h_r_12(net5026[0:23]),
     .sp12_h_r_13(net5027[0:23]), .sp12_h_r_11(net5028[0:23]),
     .lft_op_14(net4674[0:7]), .lft_op_15(net4675[0:7]),
     .lft_op_12(net4676[0:7]), .lft_op_11(net4678[0:7]),
     .lft_op_13(net4677[0:7]));
bram_bufferx4 I307 ( .in(ceb_mi), .out(ceb_o));
bram_bufferx4 I254 ( .in(mode_mi), .out(mode_o));
bram_bufferx4 I256 ( .in(r_mi), .out(r_o));
bram_bufferx4 I257 ( .in(update_mi), .out(update_o));
bram_bufferx4 I258 ( .in(shift_mi), .out(shift_o));
bram_bufferx4 I259 ( .in(hiz_b_mi), .out(hiz_b_o));
bram_bufferx4 I260 ( .in(bs_en_mi), .out(bs_en_o));

endmodule
// Library - leafcell, Cell - array_RGT_IO_1x16top, View - schematic
// LAST TIME SAVED: Apr  7 12:04:40 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module array_RGT_IO_1x16top ( cf_l, fabric_out_17, fabric_out_18,
     fabric_out_19, fabric_out_20, fabric_out_21, fabric_out_22,
     fabric_out_23, fabric_out_24, fabric_out_25, fabric_out_26,
     fabric_out_27, fabric_out_28, fabric_out_29, fabric_out_30,
     fabric_out_31, fabric_out_32, padeb, pado, sdo, slf_op_00_17,
     slf_op_00_18, slf_op_00_19, slf_op_00_20, slf_op_00_21,
     slf_op_00_22, slf_op_00_23, slf_op_00_24, slf_op_00_25,
     slf_op_00_26, slf_op_00_27, slf_op_00_28, slf_op_00_29,
     slf_op_00_30, slf_op_00_31, slf_op_00_32, spi_ss_in_b,
     SP4_h_l_00_17, SP4_h_l_00_18, SP4_h_l_00_19, SP4_h_l_00_20,
     SP4_h_l_00_21, SP4_h_l_00_22, SP4_h_l_00_23, SP4_h_l_00_24,
     SP4_h_l_00_25, SP4_h_l_00_26, SP4_h_l_00_27, SP4_h_l_00_28,
     SP4_h_l_00_29, SP4_h_l_00_30, SP4_h_l_00_31, SP4_h_l_00_32,
     SP12_h_l_00_17, SP12_h_l_00_18, SP12_h_l_00_19, SP12_h_l_00_20,
     SP12_h_l_00_21, SP12_h_l_00_22, SP12_h_l_00_23, SP12_h_l_00_24,
     SP12_h_l_00_25, SP12_h_l_00_26, SP12_h_l_00_27, SP12_h_l_00_28,
     SP12_h_l_00_29, SP12_h_l_00_30, SP12_h_l_00_31, SP12_h_l_00_32,
     bl, pgate, reset_b, sp4_v_b_00_17, sp4_v_t_00_32, vdd_cntl, wl,
     bnl_op_00_32, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     lft_op_00_17, lft_op_00_18, lft_op_00_19, lft_op_00_20,
     lft_op_00_21, lft_op_00_22, lft_op_00_23, lft_op_00_24,
     lft_op_00_25, lft_op_00_26, lft_op_00_27, lft_op_00_28,
     lft_op_00_29, lft_op_00_30, lft_op_00_31, lft_op_00_32, mode,
     padin, prog, r, sdi, shift, spioeb, spiout, tclk, tnl_op_00_17,
     update );
output  fabric_out_17, fabric_out_18, fabric_out_19, fabric_out_20,
     fabric_out_21, fabric_out_22, fabric_out_23, fabric_out_24,
     fabric_out_25, fabric_out_26, fabric_out_27, fabric_out_28,
     fabric_out_29, fabric_out_30, fabric_out_31, fabric_out_32, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_00_22;
output [3:0]  slf_op_00_17;
output [3:0]  slf_op_00_30;
output [3:0]  slf_op_00_21;
output [3:0]  slf_op_00_18;
output [3:0]  slf_op_00_27;
output [3:0]  slf_op_00_23;
output [3:0]  slf_op_00_19;
output [3:0]  slf_op_00_29;
output [3:0]  slf_op_00_28;
output [3:0]  slf_op_00_24;
output [54:28]  pado;
output [54:28]  padeb;
output [3:0]  slf_op_00_25;
output [3:0]  slf_op_00_20;
output [383:0]  cf_l;
output [31:0]  spi_ss_in_b;
output [3:0]  slf_op_00_32;
output [3:0]  slf_op_00_31;
output [3:0]  slf_op_00_26;

inout [23:0]  SP12_h_l_00_23;
inout [23:0]  SP12_h_l_00_24;
inout [23:0]  SP12_h_l_00_22;
inout [23:0]  SP12_h_l_00_31;
inout [47:0]  SP4_h_l_00_25;
inout [23:0]  SP12_h_l_00_18;
inout [23:0]  SP12_h_l_00_28;
inout [47:0]  SP4_h_l_00_29;
inout [47:0]  SP4_h_l_00_27;
inout [47:0]  SP4_h_l_00_17;
inout [23:0]  SP12_h_l_00_21;
inout [47:0]  SP4_h_l_00_32;
inout [23:0]  SP12_h_l_00_25;
inout [15:0]  sp4_v_t_00_32;
inout [23:0]  SP12_h_l_00_17;
inout [47:0]  SP4_h_l_00_20;
inout [23:0]  SP12_h_l_00_19;
inout [47:0]  SP4_h_l_00_24;
inout [47:0]  SP4_h_l_00_22;
inout [47:0]  SP4_h_l_00_19;
inout [47:0]  SP4_h_l_00_23;
inout [23:0]  SP12_h_l_00_26;
inout [47:0]  SP4_h_l_00_26;
inout [271:16]  reset_b;
inout [23:0]  SP12_h_l_00_32;
inout [23:0]  SP12_h_l_00_29;
inout [47:0]  SP4_h_l_00_28;
inout [271:16]  pgate;
inout [15:0]  sp4_v_b_00_17;
inout [271:16]  wl;
inout [271:16]  vdd_cntl;
inout [47:0]  SP4_h_l_00_21;
inout [23:0]  SP12_h_l_00_30;
inout [23:0]  SP12_h_l_00_20;
inout [47:0]  SP4_h_l_00_31;
inout [23:0]  SP12_h_l_00_27;
inout [47:0]  SP4_h_l_00_30;
inout [47:0]  SP4_h_l_00_18;
inout [17:0]  bl;

input [7:0]  lft_op_00_21;
input [7:0]  lft_op_00_19;
input [7:0]  lft_op_00_26;
input [7:0]  lft_op_00_31;
input [7:0]  glb_netwk_col;
input [7:0]  lft_op_00_25;
input [7:0]  lft_op_00_24;
input [7:0]  bnl_op_00_32;
input [7:0]  lft_op_00_23;
input [7:0]  lft_op_00_28;
input [7:0]  lft_op_00_20;
input [7:0]  lft_op_00_32;
input [7:0]  lft_op_00_30;
input [32:17]  cdone_in;
input [7:0]  tnl_op_00_17;
input [54:28]  padin;
input [7:0]  lft_op_00_18;
input [7:0]  lft_op_00_29;
input [7:0]  lft_op_00_17;
input [7:0]  lft_op_00_27;
input [31:0]  spiout;
input [7:0]  lft_op_00_22;
input [31:0]  spioeb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net1097;

wire  [0:15]  net1063;

wire  [0:15]  net791;

wire  [0:15]  net961;

wire  [0:15]  net689;

wire  [0:15]  net927;

wire  [0:15]  net655;

wire  [0:15]  net1165;

wire  [7:0]  glb_netwk;

wire  [0:1]  net891;

wire  [0:1]  net01185;

wire  [0:15]  net995;

wire  [0:15]  net723;

wire  [0:1]  net0991;

wire  [0:15]  net757;

wire  [0:15]  net859;

wire  [0:15]  net825;

wire  [0:15]  net1029;

wire  [0:15]  net1131;

wire  [0:1]  net1186;



clk_colbuf8kx8 I107 ( .clko(glb_netwk[7:0]),
     .clki(glb_netwk_col[7:0]));
io_col4_RGT I_io_00_25 ( .ceb(ceb), .sdo(net640), .sdi(net674),
     .spiout(spiout[17:16]), .cdone_in(cdone_in[25]),
     .spioeb(spioeb[17:16]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[43:42]), .pado(pado[43:42]), .padeb(padeb[43:42]),
     .sp4_v_t(net655[0:15]), .spi_ss_in_b(spi_ss_in_b[17:16]),
     .reset(reset_b[159:144]), .sp4_v_b(net689[0:15]),
     .cf(cf_l[215:192]), .bl(bl[17:0]), .slf_op(slf_op_00_25[3:0]),
     .hold(hold), .fabric_out(fabric_out_25), .prog(prog),
     .lft_op(lft_op_00_25[7:0]), .sp12_h_l(SP12_h_l_00_25[23:0]),
     .sp4_h_l(SP4_h_l_00_25[47:0]), .wl(wl[159:144]),
     .vdd_cntl(vdd_cntl[159:144]), .glb_netwk(glb_netwk[7:0]),
     .pgate(pgate[159:144]), .bnl_op(lft_op_00_24[7:0]),
     .tnl_op(lft_op_00_26[7:0]));
io_col4_RGT I_io_00_24 ( .ceb(ceb), .sdo(net674), .sdi(net708),
     .spiout(spiout[15:14]), .cdone_in(cdone_in[24]),
     .spioeb(spioeb[15:14]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[41:40]), .pado(pado[41:40]), .padeb(padeb[41:40]),
     .sp4_v_t(net689[0:15]), .sp4_h_l(SP4_h_l_00_24[47:0]),
     .sp12_h_l(SP12_h_l_00_24[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[15:14]), .tnl_op(lft_op_00_25[7:0]),
     .lft_op(lft_op_00_24[7:0]), .bnl_op(lft_op_00_23[7:0]),
     .pgate(pgate[143:128]), .reset(reset_b[143:128]),
     .sp4_v_b(net723[0:15]), .wl(wl[143:128]), .cf(cf_l[191:168]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[143:128]),
     .slf_op(slf_op_00_24[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_24));
io_col4_RGT I_io_00_23 ( .ceb(ceb), .sdo(net708), .sdi(net946),
     .spiout(spiout[13:12]), .cdone_in(cdone_in[23]),
     .spioeb(spioeb[13:12]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[39:38]), .pado(pado[39:38]), .padeb(padeb[39:38]),
     .sp4_v_t(net723[0:15]), .sp4_h_l(SP4_h_l_00_23[47:0]),
     .sp12_h_l(SP12_h_l_00_23[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[13:12]), .tnl_op(lft_op_00_24[7:0]),
     .lft_op(lft_op_00_23[7:0]), .bnl_op(lft_op_00_22[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net961[0:15]), .wl(wl[127:112]), .cf(cf_l[167:144]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_00_23[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_23));
io_col4_RGT I_io_00_31 ( .ceb(ceb), .sdo(net742), .sdi(net776),
     .spiout(spiout[29:28]), .cdone_in(cdone_in[31]),
     .spioeb(spioeb[29:28]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin({n_short, padin[54]}), .pado({n_short, pado[54]}),
     .padeb({n_idle, padeb[54]}), .sp4_v_t(net757[0:15]),
     .sp4_h_l(SP4_h_l_00_31[47:0]), .sp12_h_l(SP12_h_l_00_31[23:0]),
     .prog(prog), .spi_ss_in_b(spi_ss_in_b[29:28]),
     .tnl_op(lft_op_00_32[7:0]), .lft_op(lft_op_00_31[7:0]),
     .bnl_op(lft_op_00_30[7:0]), .pgate(pgate[255:240]),
     .reset(reset_b[255:240]), .sp4_v_b(net791[0:15]),
     .wl(wl[255:240]), .cf(cf_l[359:336]), .bl(bl[17:0]),
     .vdd_cntl(vdd_cntl[255:240]), .slf_op(slf_op_00_31[3:0]),
     .glb_netwk(glb_netwk[7:0]), .hold(hold),
     .fabric_out(fabric_out_31));
io_col4_RGT I_io_00_30 ( .ceb(ceb), .sdo(net776), .sdi(net810),
     .spiout(spiout[27:26]), .cdone_in(cdone_in[30]),
     .spioeb(spioeb[27:26]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[53:52]), .pado(pado[53:52]), .padeb(padeb[53:52]),
     .sp4_v_t(net791[0:15]), .sp4_h_l(SP4_h_l_00_30[47:0]),
     .sp12_h_l(SP12_h_l_00_30[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[27:26]), .tnl_op(lft_op_00_31[7:0]),
     .lft_op(lft_op_00_30[7:0]), .bnl_op(lft_op_00_29[7:0]),
     .pgate(pgate[239:224]), .reset(reset_b[239:224]),
     .sp4_v_b(net825[0:15]), .wl(wl[239:224]), .cf(cf_l[335:312]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[239:224]),
     .slf_op(slf_op_00_30[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_30));
io_col4_RGT I_io_00_29 ( .ceb(ceb), .sdo(net810), .sdi(net844),
     .spiout(spiout[25:24]), .cdone_in(cdone_in[29]),
     .spioeb(spioeb[25:24]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[51:50]), .pado(pado[51:50]), .padeb(padeb[51:50]),
     .sp4_v_t(net825[0:15]), .sp4_h_l(SP4_h_l_00_29[47:0]),
     .sp12_h_l(SP12_h_l_00_29[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[25:24]), .tnl_op(lft_op_00_30[7:0]),
     .lft_op(lft_op_00_29[7:0]), .bnl_op(lft_op_00_28[7:0]),
     .pgate(pgate[223:208]), .reset(reset_b[223:208]),
     .sp4_v_b(net859[0:15]), .wl(wl[223:208]), .cf(cf_l[311:288]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[223:208]),
     .slf_op(slf_op_00_29[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_29));
io_col4_RGT I_io_00_28 ( .ceb(ceb), .sdo(net844), .sdi(net1150),
     .spiout(spiout[23:22]), .cdone_in(cdone_in[28]),
     .spioeb(spioeb[23:22]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[49:48]), .pado(pado[49:48]), .padeb(padeb[49:48]),
     .sp4_v_t(net859[0:15]), .sp4_h_l(SP4_h_l_00_28[47:0]),
     .sp12_h_l(SP12_h_l_00_28[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[23:22]), .tnl_op(lft_op_00_29[7:0]),
     .lft_op(lft_op_00_28[7:0]), .bnl_op(lft_op_00_27[7:0]),
     .pgate(pgate[207:192]), .reset(reset_b[207:192]),
     .sp4_v_b(net1165[0:15]), .wl(wl[207:192]), .cf(cf_l[287:264]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[207:192]),
     .slf_op(slf_op_00_28[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_28));
io_col4_RGT I_io_00_32 ( .ceb(ceb), .sdo(sdo), .sdi(net742),
     .spiout(spiout[31:30]), .cdone_in(cdone_in[32]),
     .spioeb(spioeb[31:30]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net891[0:1]), .pado(net891[0:1]), .padeb(net1186[0:1]),
     .sp4_v_t(sp4_v_t_00_32[15:0]), .sp4_h_l(SP4_h_l_00_32[47:0]),
     .sp12_h_l(SP12_h_l_00_32[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[31:30]), .tnl_op(tnl_op_00_17[7:0]),
     .lft_op(lft_op_00_32[7:0]), .bnl_op(lft_op_00_31[7:0]),
     .pgate(pgate[271:256]), .reset(reset_b[271:256]),
     .sp4_v_b(net757[0:15]), .wl(wl[271:256]), .cf(cf_l[383:360]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[271:256]),
     .slf_op(slf_op_00_32[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_32));
io_col4_RGT I_io_00_21 ( .ceb(ceb), .sdo(net912), .sdi(net1082),
     .spiout(spiout[9:8]), .cdone_in(cdone_in[21]),
     .spioeb(spioeb[9:8]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[35:34]), .pado(pado[35:34]), .padeb(padeb[35:34]),
     .sp4_v_t(net927[0:15]), .sp4_h_l(SP4_h_l_00_21[47:0]),
     .sp12_h_l(SP12_h_l_00_21[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[9:8]), .tnl_op(lft_op_00_22[7:0]),
     .lft_op(lft_op_00_21[7:0]), .bnl_op(lft_op_00_20[7:0]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net1097[0:15]), .wl(wl[95:80]), .cf(cf_l[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_00_21[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_21));
io_col4_RGT I_io_00_22 ( .ceb(ceb), .sdo(net946), .sdi(net912),
     .spiout(spiout[11:10]), .cdone_in(cdone_in[22]),
     .spioeb(spioeb[11:10]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[37:36]), .pado(pado[37:36]), .padeb(padeb[37:36]),
     .sp4_v_t(net961[0:15]), .sp4_h_l(SP4_h_l_00_22[47:0]),
     .sp12_h_l(SP12_h_l_00_22[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[11:10]), .tnl_op(lft_op_00_23[7:0]),
     .lft_op(lft_op_00_22[7:0]), .bnl_op(lft_op_00_21[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net927[0:15]), .wl(wl[111:96]), .cf(cf_l[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_00_22[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_22));
io_col4_RGT I_io_00_18 ( .ceb(ceb), .sdo(net980), .sdi(net1014),
     .spiout(spiout[3:2]), .cdone_in(cdone_in[18]),
     .spioeb(spioeb[3:2]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net0991[0:1]), .pado(net0991[0:1]), .padeb(net01185[0:1]),
     .sp4_v_t(net995[0:15]), .sp4_h_l(SP4_h_l_00_18[47:0]),
     .sp12_h_l(SP12_h_l_00_18[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[3:2]), .tnl_op(lft_op_00_19[7:0]),
     .lft_op(lft_op_00_18[7:0]), .bnl_op(lft_op_00_17[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net1029[0:15]), .wl(wl[47:32]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_00_18[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_18));
io_col4_RGT I_io_00_17 ( .ceb(ceb), .sdo(net1014), .sdi(sdi),
     .spiout(spiout[1:0]), .cdone_in(cdone_in[17]),
     .spioeb(spioeb[1:0]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[29:28]), .pado(pado[29:28]), .padeb(padeb[29:28]),
     .sp4_v_t(net1029[0:15]), .sp4_h_l(SP4_h_l_00_17[47:0]),
     .sp12_h_l(SP12_h_l_00_17[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .tnl_op(lft_op_00_18[7:0]),
     .lft_op(lft_op_00_17[7:0]), .bnl_op(bnl_op_00_32[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(sp4_v_b_00_17[15:0]), .wl(wl[31:16]), .cf(cf_l[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_00_17[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_17));
io_col4_RGT I_io_00_19 ( .ceb(ceb), .sdo(net1048), .sdi(net980),
     .spiout(spiout[5:4]), .cdone_in(cdone_in[19]),
     .spioeb(spioeb[5:4]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[31:30]), .pado(pado[31:30]), .padeb(padeb[31:30]),
     .sp4_v_t(net1063[0:15]), .sp4_h_l(SP4_h_l_00_19[47:0]),
     .sp12_h_l(SP12_h_l_00_19[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[5:4]), .tnl_op(lft_op_00_20[7:0]),
     .lft_op(lft_op_00_19[7:0]), .bnl_op(lft_op_00_18[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net995[0:15]), .wl(wl[63:48]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_00_19[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_19));
io_col4_RGT I_io_00_20 ( .ceb(ceb), .sdo(net1082), .sdi(net1048),
     .spiout(spiout[7:6]), .cdone_in(cdone_in[20]),
     .spioeb(spioeb[7:6]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[33:32]), .pado(pado[33:32]), .padeb(padeb[33:32]),
     .sp4_v_t(net1097[0:15]), .sp4_h_l(SP4_h_l_00_20[47:0]),
     .sp12_h_l(SP12_h_l_00_20[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[7:6]), .tnl_op(lft_op_00_21[7:0]),
     .lft_op(lft_op_00_20[7:0]), .bnl_op(lft_op_00_19[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net1063[0:15]), .wl(wl[79:64]), .cf(cf_l[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_00_20[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_20));
io_col4_RGT I_io_00_26 ( .ceb(ceb), .sdo(net1116), .sdi(net640),
     .spiout(spiout[19:18]), .cdone_in(cdone_in[26]),
     .spioeb(spioeb[19:18]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[45:44]), .pado(pado[45:44]), .padeb(padeb[45:44]),
     .sp4_v_t(net1131[0:15]), .sp4_h_l(SP4_h_l_00_26[47:0]),
     .sp12_h_l(SP12_h_l_00_26[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[19:18]), .tnl_op(lft_op_00_27[7:0]),
     .lft_op(lft_op_00_26[7:0]), .bnl_op(lft_op_00_25[7:0]),
     .pgate(pgate[175:160]), .reset(reset_b[175:160]),
     .sp4_v_b(net655[0:15]), .wl(wl[175:160]), .cf(cf_l[239:216]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[175:160]),
     .slf_op(slf_op_00_26[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_26));
io_col4_RGT I_io_00_27 ( .ceb(ceb), .sdo(net1150), .sdi(net1116),
     .spiout(spiout[21:20]), .cdone_in(cdone_in[27]),
     .spioeb(spioeb[21:20]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[47:46]), .pado(pado[47:46]), .padeb(padeb[47:46]),
     .sp4_v_t(net1165[0:15]), .sp4_h_l(SP4_h_l_00_27[47:0]),
     .sp12_h_l(SP12_h_l_00_27[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[21:20]), .tnl_op(lft_op_00_28[7:0]),
     .lft_op(lft_op_00_27[7:0]), .bnl_op(lft_op_00_26[7:0]),
     .pgate(pgate[191:176]), .reset(reset_b[191:176]),
     .sp4_v_b(net1131[0:15]), .wl(wl[191:176]), .cf(cf_l[263:240]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[191:176]),
     .slf_op(slf_op_00_27[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_27));

endmodule
// Library - leafcell, Cell - bram_4kbankout_pbuffer_top, View -
//schematic
// LAST TIME SAVED: Aug 24 17:34:59 2007
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module bram_4kbankout_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [15:0]  bm_bweb;
input [15:0]  bm_d;
input [7:0]  bm_aa;
input [7:0]  bm_sa_i;
input [7:0]  bm_ab;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_bankout I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));
bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbankout, View -
//schematic
// LAST TIME SAVED: Mar  6 11:51:24 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module bram_4kprouting_tbankout ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_v_t_top;
inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_v_b_top;
inout [23:0]  sp12_h_r_top;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_bot;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_v_b_bot;

input [7:0]  rgt_op_top;
input [7:0]  bnr_op_top;
input [7:0]  glb_netwk;
input [7:0]  lft_op_bot;
input [7:0]  bnl_op_top;
input [7:0]  top_op_top;
input [7:0]  bm_sa_i;
input [7:0]  tnr_op_bot;
input [7:0]  tnl_op_bot;
input [7:0]  bnl_op_bot;
input [7:0]  lft_op_top;
input [7:0]  bot_op_bot;
input [15:0]  pgate_top;
input [15:0]  reset_b_top;
input [7:0]  tnl_op_top;
input [7:0]  tnr_op_top;
input [7:0]  bnr_op_bot;
input [15:0]  wl_top;
input [7:0]  rgt_op_bot;
input [15:0]  vdd_cntl_top;
input [15:0]  vdd_cntl_bot;
input [15:0]  pgate_bot;
input [15:0]  wl_bot;
input [15:0]  reset_b_bot;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net316;

wire  [0:7]  net243;

wire  [0:7]  net240;

wire  [0:7]  net295;

wire  [0:7]  net211;

wire  [0:7]  net210;

wire  [0:7]  net209;

wire  [0:7]  net208;

wire  [0:7]  net242;

wire  [0:7]  net241;

wire  [7:0]  in2_top;

wire  [15:0]  bm_bweb;

wire  [23:0]  sp12_v_b_top;

wire  [15:0]  bm_d;

wire  [7:0]  in2_bot;



bram_routing_tracks4rev I_bot ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}), .s_r(net213),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(tnr_op_bot[7:0]),
     .tnl_op(tnl_op_bot[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net0227),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev I_top ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}), .s_r(net245),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net0226),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbankout_pbuffer_top I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net245), .bm_wen(net213),
     .bm_d(bm_d[15:0]), .bm_clkr(net244), .bm_clkw(net212),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sdo_i(bm_sdo_i),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(bm_sdi_o),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net295[0:7]),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15],
     vdd_cntl_bot[12], vdd_cntl_bot[13], vdd_cntl_bot[10],
     vdd_cntl_bot[11], vdd_cntl_bot[8], vdd_cntl_bot[9],
     vdd_cntl_bot[6], vdd_cntl_bot[7], vdd_cntl_bot[4],
     vdd_cntl_bot[5], vdd_cntl_bot[2], vdd_cntl_bot[3],
     vdd_cntl_bot[0], vdd_cntl_bot[1]}), .bl(bl[41:26]),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net295[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15],
     vdd_cntl_top[12], vdd_cntl_top[13], vdd_cntl_top[10],
     vdd_cntl_top[11], vdd_cntl_top[8], vdd_cntl_top[9],
     vdd_cntl_top[6], vdd_cntl_top[7], vdd_cntl_top[4],
     vdd_cntl_top[5], vdd_cntl_top[2], vdd_cntl_top[3],
     vdd_cntl_top[0], vdd_cntl_top[1]}), .bl(bl[41:26]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}), .op(slf_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net316[0:7]));
tielo I14 ( .tielo(net0226));
tielo I15 ( .tielo(net0227));

endmodule
// Library - leafcell, Cell - bram_4kbank_pbuffer_top, View - schematic
// LAST TIME SAVED: Aug 24 17:33:08 2007
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module bram_4kbank_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [15:0]  bm_q;
output [7:0]  bm_sa_o;

input [15:0]  bm_bweb;
input [7:0]  bm_aa;
input [7:0]  bm_ab;
input [15:0]  bm_d;
input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbank, View - schematic
// LAST TIME SAVED: Mar  6 11:38:00 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module bram_4kprouting_tbank ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  slf_op_top;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;

inout [23:0]  sp12_h_l_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_h_l_top;
inout [23:0]  sp12_h_r_top;
inout [23:0]  sp12_v_t_top;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [47:0]  sp4_v_t_top;
inout [41:0]  bl;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_v_b_bot;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_l_bot;
inout [47:0]  sp4_v_b_top;
inout [47:0]  sp4_r_v_b_top;
inout [47:0]  sp4_h_r_top;

input [7:0]  bot_op_bot;
input [7:0]  tnr_op_top;
input [7:0]  bm_sa_i;
input [7:0]  tnr_op_bot;
input [7:0]  bnl_op_top;
input [7:0]  glb_netwk;
input [7:0]  rgt_op_bot;
input [7:0]  lft_op_bot;
input [7:0]  bnl_op_bot;
input [7:0]  tnl_op_bot;
input [7:0]  tnl_op_top;
input [15:0]  pgate_bot;
input [7:0]  bnr_op_bot;
input [7:0]  rgt_op_top;
input [15:0]  reset_b_bot;
input [7:0]  top_op_top;
input [7:0]  bnr_op_top;
input [15:0]  vdd_cntl_top;
input [15:0]  pgate_top;
input [15:0]  reset_b_top;
input [15:0]  vdd_cntl_bot;
input [15:0]  wl_bot;
input [15:0]  wl_top;
input [7:0]  lft_op_top;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net211;

wire  [0:7]  net316;

wire  [0:7]  net243;

wire  [0:7]  net240;

wire  [0:7]  net241;

wire  [7:0]  in2_top;

wire  [15:0]  bm_d;

wire  [15:0]  bm_bweb;

wire  [0:7]  net210;

wire  [0:7]  net209;

wire  [0:7]  net208;

wire  [0:7]  net242;

wire  [7:0]  in2_bot;

wire  [0:7]  net295;

wire  [23:0]  sp12_v_b_top;



bram_routing_tracks4rev I_bot ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}), .s_r(net213),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(tnr_op_bot[7:0]),
     .tnl_op(tnl_op_bot[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net0227),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev I_top ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}), .s_r(net245),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net0226),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbank_pbuffer_top I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net245), .bm_wen(net213),
     .bm_d(bm_d[15:0]), .bm_clkr(net244), .bm_clkw(net212),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sdo_i(bm_sdo_i),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(bm_sdi_o),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net295[0:7]),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15],
     vdd_cntl_bot[12], vdd_cntl_bot[13], vdd_cntl_bot[10],
     vdd_cntl_bot[11], vdd_cntl_bot[8], vdd_cntl_bot[9],
     vdd_cntl_bot[6], vdd_cntl_bot[7], vdd_cntl_bot[4],
     vdd_cntl_bot[5], vdd_cntl_bot[2], vdd_cntl_bot[3],
     vdd_cntl_bot[0], vdd_cntl_bot[1]}), .bl(bl[41:26]),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net295[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15],
     vdd_cntl_top[12], vdd_cntl_top[13], vdd_cntl_top[10],
     vdd_cntl_top[11], vdd_cntl_top[8], vdd_cntl_top[9],
     vdd_cntl_top[6], vdd_cntl_top[7], vdd_cntl_top[4],
     vdd_cntl_top[5], vdd_cntl_top[2], vdd_cntl_top[3],
     vdd_cntl_top[0], vdd_cntl_top[1]}), .bl(bl[41:26]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}), .op(slf_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net316[0:7]));
tielo I14 ( .tielo(net0226));
tielo I15 ( .tielo(net0227));

endmodule
// Library - leafcell, Cell - bram_4kbankin_pbuffer_top, View -
//schematic
// LAST TIME SAVED: Aug 24 17:33:59 2007
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module bram_4kbankin_pbuffer_top ( bm_init_o, bm_q, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_aa, bm_ab, bm_bweb, bm_clkr,
     bm_clkw, bm_d, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;

input  bm_clkr, bm_clkw, bm_init_i, bm_rcapmux_en_i, bm_ren, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bm_wen;

output [7:0]  bm_sa_o;
output [15:0]  bm_q;

input [7:0]  bm_sa_i;
input [7:0]  bm_ab;
input [7:0]  bm_aa;
input [15:0]  bm_d;
input [15:0]  bm_bweb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_4k_buffer I13 ( .bm_sdo_o(bm_sdo_o), .bm_sdo_i(net101),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sdi_i(bm_sdi_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_init_i(bm_init_i),
     .bm_sweb_o(bm_sweb_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_init_o(bm_init_o));
bram_4k_bankin I2 ( .bm_q(bm_q[15:0]), .bm_sclk(bm_sclk_o),
     .bm_wdummymux_en(bm_wdummymux_en_o),
     .bm_rcapmux_en(bm_rcapmux_en_o), .bm_bweb(bm_bweb[15:0]),
     .bm_ren(bm_ren), .bm_wen(bm_wen), .bm_clkr(bm_clkr),
     .bm_sweb(bm_sweb_o), .bm_sreb(bm_sreb_o), .bm_sdi(bm_sdo_i),
     .bm_sclkrw(bm_sclkrw_o), .bm_sa(bm_sa_o[7:0]),
     .bm_init(bm_init_o), .bm_d(bm_d[15:0]), .bm_clkw(bm_clkw),
     .bm_ab(bm_ab[7:0]), .bm_aa(bm_aa[7:0]), .bm_sdo(net101));

endmodule
// Library - leafcell, Cell - bram_4kprouting_tbankin, View - schematic
// LAST TIME SAVED: Mar  6 11:48:18 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module bram_4kprouting_tbankin ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, slf_op_bot, slf_op_top, bl, sp4_h_l_bot,
     sp4_h_l_top, sp4_h_r_bot, sp4_h_r_top, sp4_r_v_b_bot,
     sp4_r_v_b_top, sp4_v_b_bot, sp4_v_b_top, sp4_v_t_top,
     sp12_h_l_bot, sp12_h_l_top, sp12_h_r_bot, sp12_h_r_top,
     sp12_v_b_bot, sp12_v_t_top, bm_init_i, bm_rcapmux_en_i, bm_sa_i,
     bm_sclk_i, bm_sclkrw_i, bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i,
     bm_wdummymux_en_i, bnl_op_bot, bnl_op_top, bnr_op_bot, bnr_op_top,
     bot_op_bot, glb_netwk, lft_op_bot, lft_op_top, pgate_bot,
     pgate_top, prog, reset_b_bot, reset_b_top, rgt_op_bot, rgt_op_top,
     tnl_op_bot, tnl_op_top, tnr_op_bot, tnr_op_top, top_op_top,
     vdd_cntl_bot, vdd_cntl_top, wl_bot, wl_top );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  bm_sa_o;
output [7:0]  slf_op_bot;
output [7:0]  slf_op_top;

inout [23:0]  sp12_h_l_bot;
inout [23:0]  sp12_v_t_top;
inout [47:0]  sp4_h_l_top;
inout [47:0]  sp4_h_l_bot;
inout [47:0]  sp4_r_v_b_top;
inout [23:0]  sp12_v_b_bot;
inout [47:0]  sp4_h_r_bot;
inout [47:0]  sp4_r_v_b_bot;
inout [47:0]  sp4_v_t_top;
inout [47:0]  sp4_v_b_bot;
inout [47:0]  sp4_h_r_top;
inout [47:0]  sp4_v_b_top;
inout [23:0]  sp12_h_r_top;
inout [41:0]  bl;
inout [23:0]  sp12_h_r_bot;
inout [23:0]  sp12_h_l_top;

input [7:0]  bnr_op_bot;
input [7:0]  rgt_op_top;
input [7:0]  lft_op_bot;
input [7:0]  tnr_op_bot;
input [7:0]  bnr_op_top;
input [7:0]  tnl_op_top;
input [7:0]  top_op_top;
input [7:0]  tnl_op_bot;
input [7:0]  bnl_op_bot;
input [7:0]  rgt_op_bot;
input [7:0]  lft_op_top;
input [7:0]  bm_sa_i;
input [15:0]  wl_top;
input [15:0]  wl_bot;
input [7:0]  tnr_op_top;
input [7:0]  bot_op_bot;
input [7:0]  glb_netwk;
input [15:0]  pgate_top;
input [15:0]  reset_b_top;
input [15:0]  vdd_cntl_top;
input [15:0]  pgate_bot;
input [15:0]  vdd_cntl_bot;
input [15:0]  reset_b_bot;
input [7:0]  bnl_op_top;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net316;

wire  [0:7]  net243;

wire  [0:7]  net240;

wire  [23:0]  sp12_v_b_top;

wire  [0:7]  net241;

wire  [7:0]  in2_top;

wire  [0:7]  net211;

wire  [0:7]  net242;

wire  [0:7]  net208;

wire  [0:7]  net209;

wire  [0:7]  net210;

wire  [0:7]  net295;

wire  [7:0]  in2_bot;

wire  [15:0]  bm_bweb;

wire  [15:0]  bm_d;



bram_routing_tracks4rev I_bot ( .vdd_cntl({vdd_cntl_bot[14],
     vdd_cntl_bot[15], vdd_cntl_bot[12], vdd_cntl_bot[13],
     vdd_cntl_bot[10], vdd_cntl_bot[11], vdd_cntl_bot[8],
     vdd_cntl_bot[9], vdd_cntl_bot[6], vdd_cntl_bot[7],
     vdd_cntl_bot[4], vdd_cntl_bot[5], vdd_cntl_bot[2],
     vdd_cntl_bot[3], vdd_cntl_bot[0], vdd_cntl_bot[1]}), .s_r(net213),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .top_op(slf_op_top[7:0]), .tnr_op(tnr_op_bot[7:0]),
     .tnl_op(tnl_op_bot[7:0]), .slf_op(slf_op_bot[7:0]),
     .rgt_op(rgt_op_bot[7:0]), .reset_b({reset_b_bot[14],
     reset_b_bot[15], reset_b_bot[12], reset_b_bot[13],
     reset_b_bot[10], reset_b_bot[11], reset_b_bot[8], reset_b_bot[9],
     reset_b_bot[6], reset_b_bot[7], reset_b_bot[4], reset_b_bot[5],
     reset_b_bot[2], reset_b_bot[3], reset_b_bot[0], reset_b_bot[1]}),
     .prog(prog), .pgate({pgate_bot[14], pgate_bot[15], pgate_bot[12],
     pgate_bot[13], pgate_bot[10], pgate_bot[11], pgate_bot[8],
     pgate_bot[9], pgate_bot[6], pgate_bot[7], pgate_bot[4],
     pgate_bot[5], pgate_bot[2], pgate_bot[3], pgate_bot[0],
     pgate_bot[1]}), .lft_op(lft_op_bot[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net0227),
     .bot_op(bot_op_bot[7:0]), .bnr_op(bnr_op_bot[7:0]),
     .bnl_op(bnl_op_bot[7:0]), .lc_trk_g3(net208[0:7]),
     .lc_trk_g2(net209[0:7]), .lc_trk_g1(net210[0:7]),
     .lc_trk_g0(net211[0:7]), .clk(net212),
     .sp12_v_t(sp12_v_b_top[23:0]), .sp12_v_b(sp12_v_b_bot[23:0]),
     .sp12_h_r(sp12_h_r_bot[23:0]), .sp12_h_l(sp12_h_l_bot[23:0]),
     .sp4_v_t(sp4_v_b_top[47:0]), .sp4_v_b(sp4_v_b_bot[47:0]),
     .sp4_r_v_b(sp4_r_v_b_bot[47:0]), .sp4_h_r(sp4_h_r_bot[47:0]),
     .sp4_h_l(sp4_h_l_bot[47:0]), .bl(bl[25:0]));
bram_routing_tracks4rev I_top ( .vdd_cntl({vdd_cntl_top[14],
     vdd_cntl_top[15], vdd_cntl_top[12], vdd_cntl_top[13],
     vdd_cntl_top[10], vdd_cntl_top[11], vdd_cntl_top[8],
     vdd_cntl_top[9], vdd_cntl_top[6], vdd_cntl_top[7],
     vdd_cntl_top[4], vdd_cntl_top[5], vdd_cntl_top[2],
     vdd_cntl_top[3], vdd_cntl_top[0], vdd_cntl_top[1]}), .s_r(net245),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .top_op(top_op_top[7:0]), .tnr_op(tnr_op_top[7:0]),
     .tnl_op(tnl_op_top[7:0]), .slf_op(slf_op_top[7:0]),
     .rgt_op(rgt_op_top[7:0]), .reset_b({reset_b_top[14],
     reset_b_top[15], reset_b_top[12], reset_b_top[13],
     reset_b_top[10], reset_b_top[11], reset_b_top[8], reset_b_top[9],
     reset_b_top[6], reset_b_top[7], reset_b_top[4], reset_b_top[5],
     reset_b_top[2], reset_b_top[3], reset_b_top[0], reset_b_top[1]}),
     .prog(prog), .pgate({pgate_top[14], pgate_top[15], pgate_top[12],
     pgate_top[13], pgate_top[10], pgate_top[11], pgate_top[8],
     pgate_top[9], pgate_top[6], pgate_top[7], pgate_top[4],
     pgate_top[5], pgate_top[2], pgate_top[3], pgate_top[0],
     pgate_top[1]}), .lft_op(lft_op_top[7:0]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net0226),
     .bot_op(slf_op_bot[7:0]), .bnr_op(bnr_op_top[7:0]),
     .bnl_op(bnl_op_top[7:0]), .lc_trk_g3(net240[0:7]),
     .lc_trk_g2(net241[0:7]), .lc_trk_g1(net242[0:7]),
     .lc_trk_g0(net243[0:7]), .clk(net244),
     .sp12_v_t(sp12_v_t_top[23:0]), .sp12_v_b(sp12_v_b_top[23:0]),
     .sp12_h_r(sp12_h_r_top[23:0]), .sp12_h_l(sp12_h_l_top[23:0]),
     .sp4_v_t(sp4_v_t_top[47:0]), .sp4_v_b(sp4_v_b_top[47:0]),
     .sp4_r_v_b(sp4_r_v_b_top[47:0]), .sp4_h_r(sp4_h_r_top[47:0]),
     .sp4_h_l(sp4_h_l_top[47:0]), .bl(bl[25:0]));
bram_4kbankin_pbuffer_top I19 ( .bm_q({slf_op_top[7:0],
     slf_op_bot[7:0]}), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_init_i(bm_init_i), .bm_ren(net245), .bm_wen(net213),
     .bm_d(bm_d[15:0]), .bm_clkr(net244), .bm_clkw(net212),
     .bm_bweb(bm_bweb[15:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_sdo_o(bm_sdo_o), .bm_sdi_i(bm_sdi_i), .bm_ab(net316[0:7]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sdo_i(bm_sdo_i),
     .bm_sreb_i(bm_sreb_i), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(bm_sdi_o),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_aa(net295[0:7]),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_sweb_o(bm_sweb_o),
     .bm_wdummymux_en_o(bm_wdummymux_en_o));
bram_4k_inmux_8x4 I6 ( .vdd_cntl({vdd_cntl_bot[14], vdd_cntl_bot[15],
     vdd_cntl_bot[12], vdd_cntl_bot[13], vdd_cntl_bot[10],
     vdd_cntl_bot[11], vdd_cntl_bot[8], vdd_cntl_bot[9],
     vdd_cntl_bot[6], vdd_cntl_bot[7], vdd_cntl_bot[4],
     vdd_cntl_bot[5], vdd_cntl_bot[2], vdd_cntl_bot[3],
     vdd_cntl_bot[0], vdd_cntl_bot[1]}), .bl(bl[41:26]),
     .wl({wl_bot[14], wl_bot[15], wl_bot[12], wl_bot[13], wl_bot[10],
     wl_bot[11], wl_bot[8], wl_bot[9], wl_bot[6], wl_bot[7], wl_bot[4],
     wl_bot[5], wl_bot[2], wl_bot[3], wl_bot[0], wl_bot[1]}),
     .reset_b({reset_b_bot[14], reset_b_bot[15], reset_b_bot[12],
     reset_b_bot[13], reset_b_bot[10], reset_b_bot[11], reset_b_bot[8],
     reset_b_bot[9], reset_b_bot[6], reset_b_bot[7], reset_b_bot[4],
     reset_b_bot[5], reset_b_bot[2], reset_b_bot[3], reset_b_bot[0],
     reset_b_bot[1]}), .prog(prog), .pgate({pgate_bot[14],
     pgate_bot[15], pgate_bot[12], pgate_bot[13], pgate_bot[10],
     pgate_bot[11], pgate_bot[8], pgate_bot[9], pgate_bot[6],
     pgate_bot[7], pgate_bot[4], pgate_bot[5], pgate_bot[2],
     pgate_bot[3], pgate_bot[0], pgate_bot[1]}), .op(slf_op_bot[7:0]),
     .lc_trk_g3(net208[0:7]), .lc_trk_g2(net209[0:7]),
     .lc_trk_g1(net210[0:7]), .lc_trk_g0(net211[0:7]),
     .sp12_h_r({sp12_h_r_bot[22], sp12_h_r_bot[6], sp12_h_r_bot[20],
     sp12_h_r_bot[4], sp12_h_r_bot[18], sp12_h_r_bot[2],
     sp12_h_r_bot[16], sp12_h_r_bot[0], sp12_h_r_bot[14],
     sp12_h_r_bot[12], sp12_h_r_bot[10], sp12_h_r_bot[8]}),
     .sp4_v_b({sp4_v_b_bot[46], sp4_v_b_bot[30], sp4_v_b_bot[14],
     sp4_v_b_bot[44], sp4_v_b_bot[28], sp4_v_b_bot[12],
     sp4_v_b_bot[42], sp4_v_b_bot[26], sp4_v_b_bot[10],
     sp4_v_b_bot[40], sp4_v_b_bot[24], sp4_v_b_bot[8], sp4_v_b_bot[38],
     sp4_v_b_bot[22], sp4_v_b_bot[6], sp4_v_b_bot[36], sp4_v_b_bot[20],
     sp4_v_b_bot[4], sp4_v_b_bot[34], sp4_v_b_bot[18], sp4_v_b_bot[2],
     sp4_v_b_bot[32], sp4_v_b_bot[16], sp4_v_b_bot[0]}),
     .sp4_r_v_b({sp4_r_v_b_bot[47], sp4_r_v_b_bot[31],
     sp4_r_v_b_bot[15], sp4_r_v_b_bot[45], sp4_r_v_b_bot[29],
     sp4_r_v_b_bot[13], sp4_r_v_b_bot[43], sp4_r_v_b_bot[27],
     sp4_r_v_b_bot[11], sp4_r_v_b_bot[41], sp4_r_v_b_bot[25],
     sp4_r_v_b_bot[9], sp4_r_v_b_bot[39], sp4_r_v_b_bot[23],
     sp4_r_v_b_bot[7], sp4_r_v_b_bot[37], sp4_r_v_b_bot[21],
     sp4_r_v_b_bot[5], sp4_r_v_b_bot[35], sp4_r_v_b_bot[19],
     sp4_r_v_b_bot[3], sp4_r_v_b_bot[33], sp4_r_v_b_bot[17],
     sp4_r_v_b_bot[1]}), .sp4_h_r({sp4_h_r_bot[46], sp4_h_r_bot[30],
     sp4_h_r_bot[14], sp4_h_r_bot[44], sp4_h_r_bot[28],
     sp4_h_r_bot[12], sp4_h_r_bot[42], sp4_h_r_bot[26],
     sp4_h_r_bot[10], sp4_h_r_bot[40], sp4_h_r_bot[24], sp4_h_r_bot[8],
     sp4_h_r_bot[38], sp4_h_r_bot[22], sp4_h_r_bot[6], sp4_h_r_bot[36],
     sp4_h_r_bot[20], sp4_h_r_bot[4], sp4_h_r_bot[34], sp4_h_r_bot[18],
     sp4_h_r_bot[2], sp4_h_r_bot[32], sp4_h_r_bot[16],
     sp4_h_r_bot[0]}), .in3(bm_bweb[7:0]), .in2(in2_bot[7:0]),
     .in1(bm_d[7:0]), .in0(net295[0:7]), .sp12_v_b({sp12_v_b_bot[14],
     sp12_v_b_bot[12], sp12_v_b_bot[10], sp12_v_b_bot[8],
     sp12_v_b_bot[22], sp12_v_b_bot[6], sp12_v_b_bot[20],
     sp12_v_b_bot[4], sp12_v_b_bot[18], sp12_v_b_bot[2],
     sp12_v_b_bot[16], sp12_v_b_bot[0]}));
bram_4k_inmux_8x4 I0 ( .vdd_cntl({vdd_cntl_top[14], vdd_cntl_top[15],
     vdd_cntl_top[12], vdd_cntl_top[13], vdd_cntl_top[10],
     vdd_cntl_top[11], vdd_cntl_top[8], vdd_cntl_top[9],
     vdd_cntl_top[6], vdd_cntl_top[7], vdd_cntl_top[4],
     vdd_cntl_top[5], vdd_cntl_top[2], vdd_cntl_top[3],
     vdd_cntl_top[0], vdd_cntl_top[1]}), .bl(bl[41:26]),
     .sp12_v_b({sp12_v_b_top[14], sp12_v_b_top[12], sp12_v_b_top[10],
     sp12_v_b_top[8], sp12_v_b_top[22], sp12_v_b_top[6],
     sp12_v_b_top[20], sp12_v_b_top[4], sp12_v_b_top[18],
     sp12_v_b_top[2], sp12_v_b_top[16], sp12_v_b_top[0]}),
     .wl({wl_top[14], wl_top[15], wl_top[12], wl_top[13], wl_top[10],
     wl_top[11], wl_top[8], wl_top[9], wl_top[6], wl_top[7], wl_top[4],
     wl_top[5], wl_top[2], wl_top[3], wl_top[0], wl_top[1]}),
     .reset_b({reset_b_top[14], reset_b_top[15], reset_b_top[12],
     reset_b_top[13], reset_b_top[10], reset_b_top[11], reset_b_top[8],
     reset_b_top[9], reset_b_top[6], reset_b_top[7], reset_b_top[4],
     reset_b_top[5], reset_b_top[2], reset_b_top[3], reset_b_top[0],
     reset_b_top[1]}), .prog(prog), .pgate({pgate_top[14],
     pgate_top[15], pgate_top[12], pgate_top[13], pgate_top[10],
     pgate_top[11], pgate_top[8], pgate_top[9], pgate_top[6],
     pgate_top[7], pgate_top[4], pgate_top[5], pgate_top[2],
     pgate_top[3], pgate_top[0], pgate_top[1]}), .op(slf_op_top[7:0]),
     .lc_trk_g3(net240[0:7]), .lc_trk_g2(net241[0:7]),
     .lc_trk_g1(net242[0:7]), .lc_trk_g0(net243[0:7]),
     .sp12_h_r({sp12_h_r_top[22], sp12_h_r_top[6], sp12_h_r_top[20],
     sp12_h_r_top[4], sp12_h_r_top[18], sp12_h_r_top[2],
     sp12_h_r_top[16], sp12_h_r_top[0], sp12_h_r_top[14],
     sp12_h_r_top[12], sp12_h_r_top[10], sp12_h_r_top[8]}),
     .sp4_v_b({sp4_v_b_top[46], sp4_v_b_top[30], sp4_v_b_top[14],
     sp4_v_b_top[44], sp4_v_b_top[28], sp4_v_b_top[12],
     sp4_v_b_top[42], sp4_v_b_top[26], sp4_v_b_top[10],
     sp4_v_b_top[40], sp4_v_b_top[24], sp4_v_b_top[8], sp4_v_b_top[38],
     sp4_v_b_top[22], sp4_v_b_top[6], sp4_v_b_top[36], sp4_v_b_top[20],
     sp4_v_b_top[4], sp4_v_b_top[34], sp4_v_b_top[18], sp4_v_b_top[2],
     sp4_v_b_top[32], sp4_v_b_top[16], sp4_v_b_top[0]}),
     .sp4_r_v_b({sp4_r_v_b_top[47], sp4_r_v_b_top[31],
     sp4_r_v_b_top[15], sp4_r_v_b_top[45], sp4_r_v_b_top[29],
     sp4_r_v_b_top[13], sp4_r_v_b_top[43], sp4_r_v_b_top[27],
     sp4_r_v_b_top[11], sp4_r_v_b_top[41], sp4_r_v_b_top[25],
     sp4_r_v_b_top[9], sp4_r_v_b_top[39], sp4_r_v_b_top[23],
     sp4_r_v_b_top[7], sp4_r_v_b_top[37], sp4_r_v_b_top[21],
     sp4_r_v_b_top[5], sp4_r_v_b_top[35], sp4_r_v_b_top[19],
     sp4_r_v_b_top[3], sp4_r_v_b_top[33], sp4_r_v_b_top[17],
     sp4_r_v_b_top[1]}), .sp4_h_r({sp4_h_r_top[46], sp4_h_r_top[30],
     sp4_h_r_top[14], sp4_h_r_top[44], sp4_h_r_top[28],
     sp4_h_r_top[12], sp4_h_r_top[42], sp4_h_r_top[26],
     sp4_h_r_top[10], sp4_h_r_top[40], sp4_h_r_top[24], sp4_h_r_top[8],
     sp4_h_r_top[38], sp4_h_r_top[22], sp4_h_r_top[6], sp4_h_r_top[36],
     sp4_h_r_top[20], sp4_h_r_top[4], sp4_h_r_top[34], sp4_h_r_top[18],
     sp4_h_r_top[2], sp4_h_r_top[32], sp4_h_r_top[16],
     sp4_h_r_top[0]}), .in3(bm_bweb[15:8]), .in2(in2_top[7:0]),
     .in1(bm_d[15:8]), .in0(net316[0:7]));
tielo I14 ( .tielo(net0226));
tielo I15 ( .tielo(net0227));

endmodule
// Library - leafcell, Cell - array_BRAM_1x8top, View - schematic
// LAST TIME SAVED: Feb 28 14:10:09 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module array_BRAM_1x8top ( bm_init_o, bm_rcapmux_en_o, bm_sa_o,
     bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, glb_netwk, slf_op_01, slf_op_02, slf_op_03,
     slf_op_04, slf_op_05, slf_op_06, slf_op_07, slf_op_08, slf_op_09,
     slf_op_10, slf_op_11, slf_op_12, slf_op_13, slf_op_14, slf_op_15,
     slf_op_16, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02, sp4_h_l_03,
     sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07, sp4_h_l_08,
     sp4_h_l_09, sp4_h_l_10, sp4_h_l_11, sp4_h_l_12, sp4_h_l_13,
     sp4_h_l_14, sp4_h_l_15, sp4_h_l_16, sp4_h_r_01, sp4_h_r_02,
     sp4_h_r_03, sp4_h_r_04, sp4_h_r_05, sp4_h_r_06, sp4_h_r_07,
     sp4_h_r_08, sp4_h_r_09, sp4_h_r_10, sp4_h_r_11, sp4_h_r_12,
     sp4_h_r_13, sp4_h_r_14, sp4_h_r_15, sp4_h_r_16, sp4_r_v_b_01,
     sp4_r_v_b_02, sp4_r_v_b_03, sp4_r_v_b_04, sp4_r_v_b_05,
     sp4_r_v_b_06, sp4_r_v_b_07, sp4_r_v_b_08, sp4_r_v_b_09,
     sp4_r_v_b_10, sp4_r_v_b_11, sp4_r_v_b_12, sp4_r_v_b_13,
     sp4_r_v_b_14, sp4_r_v_b_15, sp4_r_v_b_16, sp4_v_b_01, sp4_v_b_02,
     sp4_v_b_03, sp4_v_b_04, sp4_v_b_05, sp4_v_b_06, sp4_v_b_07,
     sp4_v_b_08, sp4_v_b_09, sp4_v_b_10, sp4_v_b_11, sp4_v_b_12,
     sp4_v_b_13, sp4_v_b_14, sp4_v_b_15, sp4_v_b_16, sp4_v_t_16,
     sp12_h_l_01, sp12_h_l_02, sp12_h_l_03, sp12_h_l_04, sp12_h_l_05,
     sp12_h_l_06, sp12_h_l_07, sp12_h_l_08, sp12_h_l_09, sp12_h_l_10,
     sp12_h_l_11, sp12_h_l_12, sp12_h_l_13, sp12_h_l_14, sp12_h_l_15,
     sp12_h_l_16, sp12_h_r_01, sp12_h_r_02, sp12_h_r_03, sp12_h_r_04,
     sp12_h_r_05, sp12_h_r_06, sp12_h_r_07, sp12_h_r_08, sp12_h_r_09,
     sp12_h_r_10, sp12_h_r_11, sp12_h_r_12, sp12_h_r_13, sp12_h_r_14,
     sp12_h_r_15, sp12_h_r_16, sp12_v_b_01, sp12_v_t_16, vdd_cntl, wl,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i,
     bnl_op_01, bnr_op_01, bot_op_01, glb_netwk_col, lft_op_01,
     lft_op_02, lft_op_03, lft_op_04, lft_op_05, lft_op_06, lft_op_07,
     lft_op_08, lft_op_09, lft_op_10, lft_op_11, lft_op_12, lft_op_13,
     lft_op_14, lft_op_15, lft_op_16, prog, rgt_op_01, rgt_op_02,
     rgt_op_03, rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08,
     rgt_op_09, rgt_op_10, rgt_op_11, rgt_op_12, rgt_op_13, rgt_op_14,
     rgt_op_15, rgt_op_16, tnl_op_16, tnr_op_16, top_op_16 );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, prog;

output [7:0]  slf_op_03;
output [7:0]  slf_op_08;
output [7:0]  slf_op_01;
output [7:0]  slf_op_15;
output [7:0]  slf_op_02;
output [7:0]  slf_op_09;
output [7:0]  slf_op_10;
output [7:0]  slf_op_06;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_11;
output [7:0]  slf_op_12;
output [7:0]  slf_op_14;
output [7:0]  slf_op_05;
output [7:0]  slf_op_07;
output [7:0]  slf_op_16;
output [7:0]  slf_op_13;
output [7:0]  slf_op_04;
output [7:0]  glb_netwk;

inout [23:0]  sp12_h_r_03;
inout [23:0]  sp12_h_r_09;
inout [47:0]  sp4_h_l_15;
inout [47:0]  sp4_v_b_15;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_r_15;
inout [47:0]  sp4_h_r_14;
inout [47:0]  sp4_v_b_09;
inout [23:0]  sp12_h_r_14;
inout [23:0]  sp12_h_l_14;
inout [47:0]  sp4_r_v_b_10;
inout [23:0]  sp12_h_r_12;
inout [23:0]  sp12_h_r_10;
inout [47:0]  sp4_v_b_10;
inout [47:0]  sp4_h_r_02;
inout [47:0]  sp4_v_b_06;
inout [23:0]  sp12_h_l_10;
inout [41:0]  bl;
inout [47:0]  sp4_h_r_10;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_r_v_b_14;
inout [47:0]  sp4_h_r_04;
inout [47:0]  sp4_h_r_09;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_h_l_12;
inout [23:0]  sp12_h_l_12;
inout [47:0]  sp4_h_l_09;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_r_v_b_13;
inout [47:0]  sp4_h_r_08;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_r_v_b_11;
inout [23:0]  sp12_v_t_16;
inout [47:0]  sp4_r_v_b_01;
inout [23:0]  sp12_h_l_13;
inout [47:0]  sp4_r_v_b_02;
inout [47:0]  sp4_r_v_b_09;
inout [47:0]  sp4_h_l_07;
inout [23:0]  sp12_h_l_04;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_r_v_b_05;
inout [23:0]  sp12_h_r_13;
inout [47:0]  sp4_h_r_07;
inout [23:0]  sp12_h_r_07;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_h_l_04;
inout [47:0]  sp4_v_b_05;
inout [23:0]  sp12_v_b_01;
inout [47:0]  sp4_h_l_01;
inout [23:0]  sp12_h_l_05;
inout [23:0]  sp12_h_r_11;
inout [47:0]  sp4_h_r_11;
inout [47:0]  sp4_h_r_06;
inout [23:0]  sp12_h_r_16;
inout [47:0]  sp4_r_v_b_06;
inout [47:0]  sp4_h_l_02;
inout [47:0]  sp4_v_b_16;
inout [47:0]  sp4_r_v_b_12;
inout [23:0]  sp12_h_l_09;
inout [47:0]  sp4_r_v_b_03;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_h_r_16;
inout [23:0]  sp12_h_r_08;
inout [47:0]  sp4_v_b_14;
inout [47:0]  sp4_h_l_11;
inout [23:0]  sp12_h_r_04;
inout [23:0]  sp12_h_r_05;
inout [23:0]  sp12_h_l_16;
inout [47:0]  sp4_v_b_04;
inout [47:0]  sp4_h_r_13;
inout [47:0]  sp4_r_v_b_16;
inout [47:0]  sp4_v_b_12;
inout [23:0]  sp12_h_r_15;
inout [23:0]  sp12_h_l_15;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_h_r_01;
inout [23:0]  sp12_h_l_06;
inout [47:0]  sp4_v_b_03;
inout [47:0]  sp4_v_t_16;
inout [23:0]  sp12_h_l_01;
inout [47:0]  sp4_h_r_12;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_h_l_08;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_h_l_10;
inout [47:0]  sp4_h_l_14;
inout [47:0]  sp4_h_l_03;
inout [47:0]  sp4_v_b_13;
inout [47:0]  sp4_v_b_11;
inout [47:0]  sp4_r_v_b_15;
inout [47:0]  sp4_h_l_16;
inout [23:0]  sp12_h_l_08;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_h_l_13;
inout [271:16]  wl;
inout [271:16]  vdd_cntl;
inout [271:16]  pgate;
inout [271:16]  reset_b;
inout [23:0]  sp12_h_l_11;
inout [47:0]  sp4_v_b_08;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_h_l_06;

input [7:0]  lft_op_06;
input [7:0]  lft_op_01;
input [7:0]  bnr_op_01;
input [7:0]  rgt_op_13;
input [7:0]  rgt_op_09;
input [7:0]  lft_op_14;
input [7:0]  rgt_op_16;
input [7:0]  bot_op_01;
input [7:0]  rgt_op_02;
input [7:0]  tnl_op_16;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_01;
input [7:0]  lft_op_08;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_12;
input [7:0]  lft_op_07;
input [7:0]  lft_op_04;
input [7:0]  bm_sa_i;
input [7:0]  rgt_op_10;
input [7:0]  lft_op_13;
input [7:0]  rgt_op_11;
input [7:0]  lft_op_10;
input [7:0]  lft_op_09;
input [7:0]  top_op_16;
input [7:0]  lft_op_16;
input [7:0]  rgt_op_15;
input [7:0]  glb_netwk_col;
input [7:0]  lft_op_11;
input [7:0]  rgt_op_14;
input [7:0]  lft_op_02;
input [7:0]  rgt_op_05;
input [7:0]  rgt_op_06;
input [7:0]  tnr_op_16;
input [7:0]  lft_op_05;
input [7:0]  bnl_op_01;
input [7:0]  lft_op_15;
input [7:0]  rgt_op_08;
input [7:0]  lft_op_03;
input [7:0]  lft_op_12;
input [7:0]  rgt_op_04;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:23]  net970;

wire  [0:23]  net908;

wire  [0:23]  net787;

wire  [0:7]  net686;

wire  [0:7]  net873;

wire  [0:7]  net997;

wire  [0:7]  net935;

wire  [0:23]  net663;

wire  [0:7]  net813;

wire  [0:23]  net725;

wire  [0:23]  net846;

wire  [0:7]  net1061;

wire  [0:23]  net1035;

wire  [0:7]  net751;



clk_colbuf8kx8 I107 ( .clko(glb_netwk[7:0]),
     .clki(glb_netwk_col[7:0]));
bram_4kprouting_tbankout I_bram_out_0825_18 ( .bm_sdo_o(bm_sdo_o),
     .bm_sdi_i(bm_sdi_i), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sdo_i(net1008), .bm_sweb_i(bm_sweb_i), .bm_sdi_o(net1010),
     .bm_sclkrw_o(net1011), .bm_sweb_o(net1012),
     .slf_op_top(slf_op_02[7:0]), .slf_op_bot(slf_op_01[7:0]),
     .wl_top(wl[47:32]), .wl_bot(wl[31:16]),
     .top_op_top(slf_op_03[7:0]), .tnl_op_top(lft_op_03[7:0]),
     .tnl_op_bot(lft_op_02[7:0]), .reset_b_top(reset_b[47:32]),
     .reset_b_bot(reset_b[31:16]), .prog(prog),
     .pgate_top(pgate[47:32]), .pgate_bot(pgate[31:16]),
     .lft_op_top(lft_op_02[7:0]), .lft_op_bot(lft_op_01[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bot_op_bot(bot_op_01[7:0]), .sp4_h_r_top(sp4_h_r_02[47:0]),
     .bnl_op_top(lft_op_01[7:0]), .bnl_op_bot(bnl_op_01[7:0]),
     .bnr_op_bot(bnr_op_01[7:0]), .sp4_h_r_bot(sp4_h_r_01[47:0]),
     .sp12_v_t_top(net1035[0:23]), .sp12_v_b_bot(sp12_v_b_01[23:0]),
     .bm_init_i(bm_init_i), .sp12_h_l_top(sp12_h_l_02[23:0]),
     .sp12_h_r_bot(sp12_h_r_01[23:0]),
     .sp12_h_l_bot(sp12_h_l_01[23:0]),
     .sp12_h_r_top(sp12_h_r_02[23:0]), .sp4_v_t_top(sp4_v_b_03[47:0]),
     .sp4_v_b_top(sp4_v_b_02[47:0]), .sp4_v_b_bot(sp4_v_b_01[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_01[47:0]),
     .sp4_h_l_top(sp4_h_l_02[47:0]), .tnr_op_top(rgt_op_03[7:0]),
     .sp4_h_l_bot(sp4_h_l_01[47:0]), .tnr_op_bot(rgt_op_02[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .sp4_r_v_b_top(sp4_r_v_b_02[47:0]), .rgt_op_bot(rgt_op_01[7:0]),
     .rgt_op_top(rgt_op_02[7:0]), .bnr_op_top(rgt_op_01[7:0]),
     .bm_sa_i(bm_sa_i[7:0]), .bm_sclk_i(bm_sclk_i),
     .bm_sreb_i(bm_sreb_i), .bm_rcapmux_en_o(net1059),
     .bm_init_o(net1060), .bm_sa_o(net1061[0:7]), .bm_sclk_o(net1062),
     .bm_sreb_o(net1063), .bm_wdummymux_en_o(net1064),
     .vdd_cntl_top(vdd_cntl[47:32]), .vdd_cntl_bot(vdd_cntl[31:16]));
bram_4kprouting_tbank I_bram_0825_24 ( .bm_sdo_o(net698),
     .bm_sdi_i(net700), .bm_sclkrw_i(net701), .bm_sdo_i(net636),
     .bm_sweb_i(net702), .bm_sdi_o(net638), .bm_sclkrw_o(net639),
     .bm_sweb_o(net640), .slf_op_top(slf_op_08[7:0]),
     .slf_op_bot(slf_op_07[7:0]), .wl_bot(wl[127:112]),
     .top_op_top(slf_op_09[7:0]), .sp12_h_l_bot(sp12_h_l_07[23:0]),
     .sp4_h_l_bot(sp4_h_l_07[47:0]), .tnl_op_top(lft_op_09[7:0]),
     .tnl_op_bot(lft_op_08[7:0]), .reset_b_top(reset_b[143:128]),
     .reset_b_bot(reset_b[127:112]), .vdd_cntl_top(vdd_cntl[143:128]),
     .prog(prog), .pgate_top(pgate[143:128]),
     .pgate_bot(pgate[127:112]), .lft_op_bot(lft_op_07[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(net754),
     .bot_op_bot(slf_op_06[7:0]), .rgt_op_bot(rgt_op_07[7:0]),
     .bnl_op_top(lft_op_07[7:0]), .bnl_op_bot(lft_op_06[7:0]),
     .sp4_h_r_top(sp4_h_r_08[47:0]), .sp12_v_t_top(net663[0:23]),
     .sp12_v_b_bot(net725[0:23]), .bm_init_i(net750),
     .sp4_h_r_bot(sp4_h_r_07[47:0]), .sp12_h_r_bot(sp12_h_r_07[23:0]),
     .sp4_v_t_top(sp4_v_b_09[47:0]), .sp4_v_b_bot(sp4_v_b_07[47:0]),
     .sp12_h_r_top(sp12_h_r_08[23:0]), .tnr_op_bot(rgt_op_08[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net749),
     .sp4_h_l_top(sp4_h_l_08[47:0]), .lft_op_top(lft_op_08[7:0]),
     .wl_top(wl[143:128]), .sp12_h_l_top(sp12_h_l_08[23:0]),
     .sp4_v_b_top(sp4_v_b_08[47:0]), .tnr_op_top(rgt_op_09[7:0]),
     .rgt_op_top(rgt_op_08[7:0]), .bm_sa_i(net751[0:7]),
     .bm_sclk_i(net752), .bm_sreb_i(net753), .bm_rcapmux_en_o(net684),
     .bm_init_o(net685), .bm_sa_o(net686[0:7]), .bm_sclk_o(net687),
     .bm_sreb_o(net688), .bm_wdummymux_en_o(net689),
     .vdd_cntl_bot(vdd_cntl[127:112]), .bnr_op_bot(rgt_op_06[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_07[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_08[47:0]), .bnr_op_top(rgt_op_07[7:0]));
bram_4kprouting_tbank I_bram_0825_22 ( .bm_sdo_o(net760),
     .bm_sdi_i(net762), .bm_sclkrw_i(net763), .bm_sdo_i(net698),
     .bm_sweb_i(net764), .bm_sdi_o(net700), .bm_sclkrw_o(net701),
     .bm_sweb_o(net702), .slf_op_top(slf_op_06[7:0]),
     .slf_op_bot(slf_op_05[7:0]), .wl_top(wl[111:96]),
     .wl_bot(wl[95:80]), .top_op_top(slf_op_07[7:0]),
     .tnl_op_top(lft_op_07[7:0]), .tnl_op_bot(lft_op_06[7:0]),
     .reset_b_top(reset_b[111:96]), .reset_b_bot(reset_b[95:80]),
     .prog(prog), .pgate_top(pgate[111:96]), .pgate_bot(pgate[95:80]),
     .lft_op_top(lft_op_06[7:0]), .lft_op_bot(lft_op_05[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(net816),
     .bot_op_bot(slf_op_04[7:0]), .sp4_h_r_top(sp4_h_r_06[47:0]),
     .bnl_op_top(lft_op_05[7:0]), .bnl_op_bot(lft_op_04[7:0]),
     .bnr_op_bot(rgt_op_04[7:0]), .sp4_h_r_bot(sp4_h_r_05[47:0]),
     .sp12_v_t_top(net725[0:23]), .sp12_v_b_bot(net787[0:23]),
     .bm_init_i(net812), .sp12_h_l_top(sp12_h_l_06[23:0]),
     .sp12_h_r_bot(sp12_h_r_05[23:0]),
     .sp12_h_l_bot(sp12_h_l_05[23:0]),
     .sp12_h_r_top(sp12_h_r_06[23:0]), .sp4_v_t_top(sp4_v_b_07[47:0]),
     .sp4_v_b_top(sp4_v_b_06[47:0]), .sp4_v_b_bot(sp4_v_b_05[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_05[47:0]),
     .sp4_h_l_top(sp4_h_l_06[47:0]), .tnr_op_top(rgt_op_07[7:0]),
     .sp4_h_l_bot(sp4_h_l_05[47:0]), .tnr_op_bot(rgt_op_06[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net811),
     .sp4_r_v_b_top(sp4_r_v_b_06[47:0]), .rgt_op_bot(rgt_op_05[7:0]),
     .rgt_op_top(rgt_op_06[7:0]), .bnr_op_top(rgt_op_05[7:0]),
     .bm_sa_i(net813[0:7]), .bm_sclk_i(net814), .bm_sreb_i(net815),
     .bm_rcapmux_en_o(net749), .bm_init_o(net750),
     .bm_sa_o(net751[0:7]), .bm_sclk_o(net752), .bm_sreb_o(net753),
     .bm_wdummymux_en_o(net754), .vdd_cntl_top(vdd_cntl[111:96]),
     .vdd_cntl_bot(vdd_cntl[95:80]));
bram_4kprouting_tbank I_bram_0825_20 ( .bm_sdo_o(net1008),
     .bm_sdi_i(net1010), .bm_sclkrw_i(net1011), .bm_sdo_i(net760),
     .bm_sweb_i(net1012), .bm_sdi_o(net762), .bm_sclkrw_o(net763),
     .bm_sweb_o(net764), .slf_op_top(slf_op_04[7:0]),
     .slf_op_bot(slf_op_03[7:0]), .wl_top(wl[79:64]),
     .wl_bot(wl[63:48]), .top_op_top(slf_op_05[7:0]),
     .tnl_op_top(lft_op_05[7:0]), .tnl_op_bot(lft_op_04[7:0]),
     .reset_b_top(reset_b[79:64]), .reset_b_bot(reset_b[63:48]),
     .prog(prog), .pgate_top(pgate[79:64]), .pgate_bot(pgate[63:48]),
     .lft_op_top(lft_op_04[7:0]), .lft_op_bot(lft_op_03[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bm_wdummymux_en_i(net1064),
     .bot_op_bot(slf_op_02[7:0]), .sp4_h_r_top(sp4_h_r_04[47:0]),
     .bnl_op_top(lft_op_03[7:0]), .bnl_op_bot(lft_op_02[7:0]),
     .bnr_op_bot(rgt_op_02[7:0]), .sp4_h_r_bot(sp4_h_r_03[47:0]),
     .sp12_v_t_top(net787[0:23]), .sp12_v_b_bot(net1035[0:23]),
     .bm_init_i(net1060), .sp12_h_l_top(sp12_h_l_04[23:0]),
     .sp12_h_r_bot(sp12_h_r_03[23:0]),
     .sp12_h_l_bot(sp12_h_l_03[23:0]),
     .sp12_h_r_top(sp12_h_r_04[23:0]), .sp4_v_t_top(sp4_v_b_05[47:0]),
     .sp4_v_b_top(sp4_v_b_04[47:0]), .sp4_v_b_bot(sp4_v_b_03[47:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_03[47:0]),
     .sp4_h_l_top(sp4_h_l_04[47:0]), .tnr_op_top(rgt_op_05[7:0]),
     .sp4_h_l_bot(sp4_h_l_03[47:0]), .tnr_op_bot(rgt_op_04[7:0]),
     .bl(bl[41:0]), .bm_rcapmux_en_i(net1059),
     .sp4_r_v_b_top(sp4_r_v_b_04[47:0]), .rgt_op_bot(rgt_op_03[7:0]),
     .rgt_op_top(rgt_op_04[7:0]), .bnr_op_top(rgt_op_03[7:0]),
     .bm_sa_i(net1061[0:7]), .bm_sclk_i(net1062), .bm_sreb_i(net1063),
     .bm_rcapmux_en_o(net811), .bm_init_o(net812),
     .bm_sa_o(net813[0:7]), .bm_sclk_o(net814), .bm_sreb_o(net815),
     .bm_wdummymux_en_o(net816), .vdd_cntl_top(vdd_cntl[79:64]),
     .vdd_cntl_bot(vdd_cntl[63:48]));
bram_4kprouting_tbank I_bram_0825_28 ( .slf_op_top(slf_op_12[7:0]),
     .sp4_h_l_bot(sp4_h_l_11[47:0]), .slf_op_bot(slf_op_11[7:0]),
     .sp4_r_v_b_top(sp4_r_v_b_12[47:0]),
     .reset_b_top(reset_b[207:192]), .tnl_op_top(lft_op_13[7:0]),
     .top_op_top(slf_op_13[7:0]), .rgt_op_bot(rgt_op_11[7:0]),
     .tnl_op_bot(lft_op_12[7:0]), .prog(prog),
     .lft_op_top(lft_op_12[7:0]), .lft_op_bot(lft_op_11[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bnl_op_top(lft_op_11[7:0]),
     .rgt_op_top(rgt_op_12[7:0]), .bnl_op_bot(lft_op_10[7:0]),
     .sp12_h_l_top(sp12_h_l_12[23:0]), .sp4_v_b_top(sp4_v_b_12[47:0]),
     .bl(bl[41:0]), .bm_wdummymux_en_i(net939),
     .bot_op_bot(slf_op_10[7:0]), .tnr_op_bot(rgt_op_12[7:0]),
     .bnr_op_bot(rgt_op_10[7:0]), .sp4_h_l_top(sp4_h_l_12[47:0]),
     .wl_bot(wl[191:176]), .sp4_r_v_b_bot(sp4_r_v_b_11[47:0]),
     .tnr_op_top(rgt_op_13[7:0]), .sp12_v_t_top(net846[0:23]),
     .sp12_v_b_bot(net908[0:23]), .bm_init_i(net934),
     .sp4_h_r_bot(sp4_h_r_11[47:0]), .pgate_top(pgate[207:192]),
     .sp12_h_r_bot(sp12_h_r_11[23:0]), .sp4_v_t_top(sp4_v_b_13[47:0]),
     .sp12_h_r_top(sp12_h_r_12[23:0]), .sp4_v_b_bot(sp4_v_b_11[47:0]),
     .bnr_op_top(rgt_op_11[7:0]), .reset_b_bot(reset_b[191:176]),
     .wl_top(wl[207:192]), .sp4_h_r_top(sp4_h_r_12[47:0]),
     .bm_rcapmux_en_i(net932), .bm_sdo_o(net928), .bm_sdi_i(net931),
     .pgate_bot(pgate[191:176]), .bm_sa_i(net935[0:7]),
     .bm_sclk_i(net936), .bm_sclkrw_i(net933), .bm_sdo_i(net866),
     .bm_sreb_i(net937), .bm_sweb_i(net938), .bm_sdi_o(net869),
     .bm_rcapmux_en_o(net870), .bm_sclkrw_o(net871),
     .bm_init_o(net872), .bm_sa_o(net873[0:7]), .bm_sclk_o(net874),
     .bm_sreb_o(net875), .bm_sweb_o(net876),
     .bm_wdummymux_en_o(net877), .vdd_cntl_bot(vdd_cntl[191:176]),
     .vdd_cntl_top(vdd_cntl[207:192]),
     .sp12_h_l_bot(sp12_h_l_11[23:0]));
bram_4kprouting_tbank I_bram_0825_26 ( .slf_op_top(slf_op_10[7:0]),
     .sp4_h_l_bot(sp4_h_l_09[47:0]), .slf_op_bot(slf_op_09[7:0]),
     .sp4_r_v_b_top(sp4_r_v_b_10[47:0]),
     .reset_b_top(reset_b[175:160]), .tnl_op_top(lft_op_11[7:0]),
     .top_op_top(slf_op_11[7:0]), .rgt_op_bot(rgt_op_09[7:0]),
     .tnl_op_bot(lft_op_10[7:0]), .prog(prog),
     .lft_op_top(lft_op_10[7:0]), .lft_op_bot(lft_op_09[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bnl_op_top(lft_op_09[7:0]),
     .rgt_op_top(rgt_op_10[7:0]), .bnl_op_bot(lft_op_08[7:0]),
     .sp12_h_l_top(sp12_h_l_10[23:0]), .sp4_v_b_top(sp4_v_b_10[47:0]),
     .bl(bl[41:0]), .bm_wdummymux_en_i(net689),
     .bot_op_bot(slf_op_08[7:0]), .tnr_op_bot(rgt_op_10[7:0]),
     .bnr_op_bot(rgt_op_08[7:0]), .sp4_h_l_top(sp4_h_l_10[47:0]),
     .wl_bot(wl[159:144]), .sp4_r_v_b_bot(sp4_r_v_b_09[47:0]),
     .tnr_op_top(rgt_op_11[7:0]), .sp12_v_t_top(net908[0:23]),
     .sp12_v_b_bot(net663[0:23]), .bm_init_i(net685),
     .sp4_h_r_bot(sp4_h_r_09[47:0]), .pgate_top(pgate[175:160]),
     .sp12_h_r_bot(sp12_h_r_09[23:0]), .sp4_v_t_top(sp4_v_b_11[47:0]),
     .sp12_h_r_top(sp12_h_r_10[23:0]), .sp4_v_b_bot(sp4_v_b_09[47:0]),
     .bnr_op_top(rgt_op_09[7:0]), .reset_b_bot(reset_b[159:144]),
     .wl_top(wl[175:160]), .sp4_h_r_top(sp4_h_r_10[47:0]),
     .bm_rcapmux_en_i(net684), .bm_sdo_o(net636), .bm_sdi_i(net638),
     .pgate_bot(pgate[159:144]), .bm_sa_i(net686[0:7]),
     .bm_sclk_i(net687), .bm_sclkrw_i(net639), .bm_sdo_i(net928),
     .bm_sreb_i(net688), .bm_sweb_i(net640), .bm_sdi_o(net931),
     .bm_rcapmux_en_o(net932), .bm_sclkrw_o(net933),
     .bm_init_o(net934), .bm_sa_o(net935[0:7]), .bm_sclk_o(net936),
     .bm_sreb_o(net937), .bm_sweb_o(net938),
     .bm_wdummymux_en_o(net939), .vdd_cntl_bot(vdd_cntl[159:144]),
     .vdd_cntl_top(vdd_cntl[175:160]),
     .sp12_h_l_bot(sp12_h_l_09[23:0]));
bram_4kprouting_tbank I_bram_0825_30 ( .slf_op_top(slf_op_14[7:0]),
     .sp4_h_l_bot(sp4_h_l_13[47:0]), .slf_op_bot(slf_op_13[7:0]),
     .sp4_r_v_b_top(sp4_r_v_b_14[47:0]),
     .reset_b_top(reset_b[239:224]), .tnl_op_top(lft_op_15[7:0]),
     .top_op_top(slf_op_15[7:0]), .rgt_op_bot(rgt_op_13[7:0]),
     .tnl_op_bot(lft_op_14[7:0]), .prog(prog),
     .lft_op_top(lft_op_14[7:0]), .lft_op_bot(lft_op_13[7:0]),
     .glb_netwk(glb_netwk[7:0]), .bnl_op_top(lft_op_13[7:0]),
     .rgt_op_top(rgt_op_14[7:0]), .bnl_op_bot(lft_op_12[7:0]),
     .sp12_h_l_top(sp12_h_l_14[23:0]), .sp4_v_b_top(sp4_v_b_14[47:0]),
     .bl(bl[41:0]), .bm_wdummymux_en_i(net877),
     .bot_op_bot(slf_op_12[7:0]), .tnr_op_bot(rgt_op_14[7:0]),
     .bnr_op_bot(rgt_op_12[7:0]), .sp4_h_l_top(sp4_h_l_14[47:0]),
     .wl_bot(wl[223:208]), .sp4_r_v_b_bot(sp4_r_v_b_13[47:0]),
     .tnr_op_top(rgt_op_15[7:0]), .sp12_v_t_top(net970[0:23]),
     .sp12_v_b_bot(net846[0:23]), .bm_init_i(net872),
     .sp4_h_r_bot(sp4_h_r_13[47:0]), .pgate_top(pgate[239:224]),
     .sp12_h_r_bot(sp12_h_r_13[23:0]), .sp4_v_t_top(sp4_v_b_15[47:0]),
     .sp12_h_r_top(sp12_h_r_14[23:0]), .sp4_v_b_bot(sp4_v_b_13[47:0]),
     .bnr_op_top(rgt_op_13[7:0]), .reset_b_bot(reset_b[223:208]),
     .wl_top(wl[239:224]), .sp4_h_r_top(sp4_h_r_14[47:0]),
     .bm_rcapmux_en_i(net870), .bm_sdo_o(net866), .bm_sdi_i(net869),
     .pgate_bot(pgate[223:208]), .bm_sa_i(net873[0:7]),
     .bm_sclk_i(net874), .bm_sclkrw_i(net871), .bm_sdo_i(net990),
     .bm_sreb_i(net875), .bm_sweb_i(net876), .bm_sdi_o(net993),
     .bm_rcapmux_en_o(net994), .bm_sclkrw_o(net995),
     .bm_init_o(net996), .bm_sa_o(net997[0:7]), .bm_sclk_o(net998),
     .bm_sreb_o(net999), .bm_sweb_o(net1000),
     .bm_wdummymux_en_o(net1001), .vdd_cntl_bot(vdd_cntl[223:208]),
     .vdd_cntl_top(vdd_cntl[239:224]),
     .sp12_h_l_bot(sp12_h_l_13[23:0]));
bram_4kprouting_tbankin I_bram_in_0825_32 ( .bm_sdo_o(net990),
     .bm_sdi_i(net993), .bm_sclkrw_i(net995), .bm_sdo_i(bm_sdo_i),
     .bm_sweb_i(net1000), .bm_sdi_o(bm_sdi_o),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_sweb_o(bm_sweb_o),
     .slf_op_top(slf_op_16[7:0]), .slf_op_bot(slf_op_15[7:0]),
     .wl_bot(wl[255:240]), .top_op_top(top_op_16[7:0]),
     .sp12_h_l_bot(sp12_h_l_15[23:0]), .sp4_h_l_bot(sp4_h_l_15[47:0]),
     .tnl_op_top(tnl_op_16[7:0]), .tnl_op_bot(lft_op_16[7:0]),
     .reset_b_top(reset_b[271:256]), .reset_b_bot(reset_b[255:240]),
     .vdd_cntl_top(vdd_cntl[271:256]), .prog(prog),
     .pgate_top(pgate[271:256]), .pgate_bot(pgate[255:240]),
     .lft_op_bot(lft_op_15[7:0]), .glb_netwk(glb_netwk[7:0]),
     .bm_wdummymux_en_i(net1001), .bot_op_bot(slf_op_14[7:0]),
     .rgt_op_bot(rgt_op_15[7:0]), .bnl_op_top(lft_op_15[7:0]),
     .bnl_op_bot(lft_op_14[7:0]), .sp4_h_r_top(sp4_h_r_16[47:0]),
     .sp12_v_t_top(sp12_v_t_16[23:0]), .sp12_v_b_bot(net970[0:23]),
     .bm_init_i(net996), .sp4_h_r_bot(sp4_h_r_15[47:0]),
     .sp12_h_r_bot(sp12_h_r_15[23:0]), .sp4_v_t_top(sp4_v_t_16[47:0]),
     .sp4_v_b_bot(sp4_v_b_15[47:0]), .sp12_h_r_top(sp12_h_r_16[23:0]),
     .tnr_op_bot(rgt_op_16[7:0]), .bl(bl[41:0]),
     .bm_rcapmux_en_i(net994), .sp4_h_l_top(sp4_h_l_16[47:0]),
     .lft_op_top(lft_op_16[7:0]), .wl_top(wl[271:256]),
     .sp12_h_l_top(sp12_h_l_16[23:0]), .sp4_v_b_top(sp4_v_b_16[47:0]),
     .tnr_op_top(tnr_op_16[7:0]), .rgt_op_top(rgt_op_16[7:0]),
     .bm_sa_i(net997[0:7]), .bm_sclk_i(net998), .bm_sreb_i(net999),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_sclk_o(bm_sclk_o),
     .bm_sreb_o(bm_sreb_o), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .vdd_cntl_bot(vdd_cntl[255:240]), .bnr_op_bot(rgt_op_14[7:0]),
     .sp4_r_v_b_bot(sp4_r_v_b_15[47:0]),
     .sp4_r_v_b_top(sp4_r_v_b_16[47:0]), .bnr_op_top(rgt_op_15[7:0]));

endmodule
// Library - leafcell, Cell - array_LT1x16top, View - schematic
// LAST TIME SAVED: Jun 12 09:54:14 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module array_LT1x16top ( carry_out, glb_netwk, slf_op_01, slf_op_02,
     slf_op_03, slf_op_04, slf_op_05, slf_op_06, slf_op_07, slf_op_08,
     slf_op_09, slf_op_10, slf_op_11, slf_op_12, slf_op_13, slf_op_14,
     slf_op_15, slf_op_16, bl, pgate, reset_b, sp4_h_l_01, sp4_h_l_02,
     sp4_h_l_03, sp4_h_l_04, sp4_h_l_05, sp4_h_l_06, sp4_h_l_07,
     sp4_h_l_08, sp4_h_l_09, sp4_h_l_10, sp4_h_l_11, sp4_h_l_12,
     sp4_h_l_13, sp4_h_l_14, sp4_h_l_15, sp4_h_l_16, sp4_h_r_01,
     sp4_h_r_02, sp4_h_r_03, sp4_h_r_04, sp4_h_r_05, sp4_h_r_06,
     sp4_h_r_07, sp4_h_r_08, sp4_h_r_09, sp4_h_r_10, sp4_h_r_11,
     sp4_h_r_12, sp4_h_r_13, sp4_h_r_14, sp4_h_r_15, sp4_h_r_16,
     sp4_r_v_b_01, sp4_r_v_b_02, sp4_r_v_b_03, sp4_r_v_b_04,
     sp4_r_v_b_05, sp4_r_v_b_06, sp4_r_v_b_07, sp4_r_v_b_08,
     sp4_r_v_b_09, sp4_r_v_b_10, sp4_r_v_b_11, sp4_r_v_b_12,
     sp4_r_v_b_13, sp4_r_v_b_14, sp4_r_v_b_15, sp4_r_v_b_16,
     sp4_v_b_01, sp4_v_b_02, sp4_v_b_03, sp4_v_b_04, sp4_v_b_05,
     sp4_v_b_06, sp4_v_b_07, sp4_v_b_08, sp4_v_b_09, sp4_v_b_10,
     sp4_v_b_11, sp4_v_b_12, sp4_v_b_13, sp4_v_b_14, sp4_v_b_15,
     sp4_v_b_16, sp4_v_t_16, sp12_h_l_01, sp12_h_l_02, sp12_h_l_03,
     sp12_h_l_04, sp12_h_l_05, sp12_h_l_06, sp12_h_l_07, sp12_h_l_08,
     sp12_h_l_09, sp12_h_l_10, sp12_h_l_11, sp12_h_l_12, sp12_h_l_13,
     sp12_h_l_14, sp12_h_l_15, sp12_h_l_16, sp12_h_r_01, sp12_h_r_02,
     sp12_h_r_03, sp12_h_r_04, sp12_h_r_05, sp12_h_r_06, sp12_h_r_07,
     sp12_h_r_08, sp12_h_r_09, sp12_h_r_10, sp12_h_r_11, sp12_h_r_12,
     sp12_h_r_13, sp12_h_r_14, sp12_h_r_15, sp12_h_r_16, sp12_v_b__01,
     sp12_v_t_16, vdd_cntl, wl, bnl_op_01, bnr_op_01, bot_op_01,
     carry_in, glb_netwk_col, lft_op_01, lft_op_02, lft_op_03,
     lft_op_04, lft_op_05, lft_op_06, lft_op_07, lft_op_08, lft_op_09,
     lft_op_10, lft_op_11, lft_op_12, lft_op_13, lft_op_14, lft_op_15,
     lft_op_16, prog, purst, rgt_op_01, rgt_op_02, rgt_op_03,
     rgt_op_04, rgt_op_05, rgt_op_06, rgt_op_07, rgt_op_08, rgt_op_09,
     rgt_op_10, rgt_op_11, rgt_op_12, rgt_op_13, rgt_op_14, rgt_op_15,
     rgt_op_16, tnl_op_16, tnr_op_16, top_op_16 );
output  carry_out;


input  carry_in, prog, purst;

output [7:0]  slf_op_16;
output [7:0]  slf_op_01;
output [7:0]  slf_op_10;
output [7:0]  slf_op_08;
output [7:0]  slf_op_07;
output [7:0]  slf_op_11;
output [7:0]  slf_op_02;
output [7:0]  slf_op_12;
output [7:0]  glb_netwk;
output [7:0]  slf_op_06;
output [7:0]  slf_op_03;
output [7:0]  slf_op_09;
output [7:0]  slf_op_13;
output [7:0]  slf_op_15;
output [7:0]  slf_op_04;
output [7:0]  slf_op_05;
output [7:0]  slf_op_14;

inout [47:0]  sp4_r_v_b_15;
inout [47:0]  sp4_h_l_10;
inout [23:0]  sp12_h_l_16;
inout [47:0]  sp4_h_r_16;
inout [23:0]  sp12_h_l_04;
inout [23:0]  sp12_h_l_02;
inout [47:0]  sp4_v_b_05;
inout [47:0]  sp4_v_b_16;
inout [47:0]  sp4_h_l_07;
inout [47:0]  sp4_r_v_b_16;
inout [23:0]  sp12_h_r_13;
inout [47:0]  sp4_r_v_b_01;
inout [47:0]  sp4_v_b_15;
inout [47:0]  sp4_v_b_06;
inout [47:0]  sp4_v_b_13;
inout [47:0]  sp4_h_l_12;
inout [47:0]  sp4_h_l_16;
inout [47:0]  sp4_h_r_13;
inout [47:0]  sp4_v_b_12;
inout [47:0]  sp4_v_b_09;
inout [47:0]  sp4_r_v_b_11;
inout [23:0]  sp12_h_r_11;
inout [47:0]  sp4_v_b_14;
inout [47:0]  sp4_h_r_11;
inout [23:0]  sp12_h_r_06;
inout [47:0]  sp4_r_v_b_04;
inout [47:0]  sp4_h_r_08;
inout [23:0]  sp12_h_l_05;
inout [47:0]  sp4_r_v_b_07;
inout [47:0]  sp4_v_t_16;
inout [23:0]  sp12_h_r_01;
inout [47:0]  sp4_h_l_11;
inout [47:0]  sp4_r_v_b_14;
inout [23:0]  sp12_h_l_12;
inout [23:0]  sp12_h_l_06;
inout [23:0]  sp12_h_r_02;
inout [47:0]  sp4_v_b_02;
inout [47:0]  sp4_h_l_05;
inout [47:0]  sp4_h_l_13;
inout [47:0]  sp4_r_v_b_10;
inout [23:0]  sp12_h_l_11;
inout [23:0]  sp12_h_r_15;
inout [47:0]  sp4_h_l_14;
inout [47:0]  sp4_h_l_06;
inout [255:0]  wl;
inout [47:0]  sp4_h_r_03;
inout [47:0]  sp4_r_v_b_06;
inout [255:0]  reset_b;
inout [47:0]  sp4_h_r_06;
inout [47:0]  sp4_r_v_b_03;
inout [23:0]  sp12_h_r_08;
inout [47:0]  sp4_h_r_01;
inout [47:0]  sp4_h_l_02;
inout [23:0]  sp12_h_l_09;
inout [23:0]  sp12_h_r_10;
inout [47:0]  sp4_h_l_09;
inout [47:0]  sp4_h_r_05;
inout [47:0]  sp4_h_r_12;
inout [47:0]  sp4_h_l_08;
inout [23:0]  sp12_h_r_12;
inout [255:0]  pgate;
inout [47:0]  sp4_v_b_07;
inout [47:0]  sp4_v_b_10;
inout [23:0]  sp12_h_r_16;
inout [47:0]  sp4_h_r_02;
inout [23:0]  sp12_h_l_08;
inout [23:0]  sp12_h_l_03;
inout [47:0]  sp4_h_l_01;
inout [23:0]  sp12_h_r_14;
inout [47:0]  sp4_r_v_b_02;
inout [255:0]  vdd_cntl;
inout [23:0]  sp12_v_t_16;
inout [47:0]  sp4_r_v_b_12;
inout [47:0]  sp4_h_r_04;
inout [23:0]  sp12_h_l_10;
inout [47:0]  sp4_h_l_15;
inout [23:0]  sp12_h_l_15;
inout [23:0]  sp12_h_r_03;
inout [47:0]  sp4_h_r_15;
inout [23:0]  sp12_h_l_07;
inout [47:0]  sp4_h_r_07;
inout [47:0]  sp4_r_v_b_08;
inout [47:0]  sp4_v_b_01;
inout [47:0]  sp4_h_l_04;
inout [23:0]  sp12_h_r_07;
inout [23:0]  sp12_h_l_13;
inout [23:0]  sp12_h_r_04;
inout [47:0]  sp4_v_b_08;
inout [47:0]  sp4_r_v_b_13;
inout [47:0]  sp4_v_b_04;
inout [23:0]  sp12_h_r_05;
inout [47:0]  sp4_r_v_b_05;
inout [47:0]  sp4_h_r_14;
inout [53:0]  bl;
inout [47:0]  sp4_h_r_10;
inout [47:0]  sp4_v_b_11;
inout [23:0]  sp12_v_b__01;
inout [47:0]  sp4_h_l_03;
inout [47:0]  sp4_v_b_03;
inout [47:0]  sp4_h_r_09;
inout [47:0]  sp4_r_v_b_09;
inout [23:0]  sp12_h_l_01;
inout [23:0]  sp12_h_l_14;
inout [23:0]  sp12_h_r_09;

input [7:0]  rgt_op_15;
input [7:0]  rgt_op_04;
input [7:0]  lft_op_04;
input [7:0]  lft_op_03;
input [7:0]  lft_op_08;
input [7:0]  rgt_op_06;
input [7:0]  tnr_op_16;
input [7:0]  lft_op_06;
input [7:0]  lft_op_15;
input [7:0]  rgt_op_10;
input [7:0]  tnl_op_16;
input [7:0]  rgt_op_12;
input [7:0]  lft_op_05;
input [7:0]  bot_op_01;
input [7:0]  bnl_op_01;
input [7:0]  bnr_op_01;
input [7:0]  lft_op_16;
input [7:0]  rgt_op_14;
input [7:0]  rgt_op_07;
input [7:0]  rgt_op_09;
input [7:0]  rgt_op_13;
input [7:0]  lft_op_11;
input [7:0]  lft_op_10;
input [7:0]  rgt_op_03;
input [7:0]  rgt_op_16;
input [7:0]  lft_op_12;
input [7:0]  lft_op_02;
input [7:0]  rgt_op_08;
input [7:0]  rgt_op_05;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_11;
input [7:0]  lft_op_09;
input [7:0]  lft_op_14;
input [7:0]  top_op_16;
input [7:0]  lft_op_13;
input [7:0]  lft_op_01;
input [7:0]  rgt_op_02;
input [7:0]  rgt_op_01;
input [7:0]  lft_op_07;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:23]  net983;

wire  [0:23]  net1039;

wire  [0:23]  net675;

wire  [0:23]  net899;

wire  [0:23]  net787;

wire  [0:23]  net843;

wire  [0:23]  net731;

wire  [0:23]  net871;

wire  [0:23]  net815;

wire  [0:23]  net1011;

wire  [0:23]  net647;

wire  [0:23]  net619;

wire  [0:23]  net759;

wire  [0:23]  net927;

wire  [0:23]  net955;



ltile4rev0 I_LT06 ( .prog(prog), .carry_out(net779),
     .lft_op(lft_op_06[7:0]), .sp12_h_l(sp12_h_l_06[23:0]),
     .sp4_h_l(sp4_h_l_06[47:0]), .sp4_v_b(sp4_v_b_06[47:0]),
     .sp12_v_b(net871[0:23]), .sp12_h_r(sp12_h_r_06[23:0]),
     .sp4_h_r(sp4_h_r_06[47:0]), .sp12_v_t(net787[0:23]),
     .sp4_v_t(sp4_v_b_07[47:0]), .sp4_r_v_b(sp4_r_v_b_06[47:0]),
     .wl(wl[95:80]), .top_op(slf_op_07[7:0]), .rgt_op(rgt_op_06[7:0]),
     .bot_op(slf_op_05[7:0]), .bl(bl[53:0]), .reset_b(reset_b[95:80]),
     .vdd_cntl(vdd_cntl[95:80]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net863), .purst(purst), .slf_op(slf_op_06[7:0]),
     .pgate(pgate[95:80]), .bnr_op(rgt_op_05[7:0]),
     .bnl_op(lft_op_05[7:0]), .tnr_op(rgt_op_07[7:0]),
     .tnl_op(lft_op_07[7:0]));
ltile4rev0 I_LT03 ( .prog(prog), .carry_out(net807),
     .lft_op(lft_op_03[7:0]), .sp12_h_l(sp12_h_l_03[23:0]),
     .sp4_h_l(sp4_h_l_03[47:0]), .sp4_v_b(sp4_v_b_03[47:0]),
     .sp12_v_b(net927[0:23]), .sp12_h_r(sp12_h_r_03[23:0]),
     .sp4_h_r(sp4_h_r_03[47:0]), .sp12_v_t(net815[0:23]),
     .sp4_v_t(sp4_v_b_04[47:0]), .sp4_r_v_b(sp4_r_v_b_03[47:0]),
     .wl(wl[47:32]), .top_op(slf_op_04[7:0]), .rgt_op(rgt_op_03[7:0]),
     .bot_op(slf_op_02[7:0]), .bl(bl[53:0]), .reset_b(reset_b[47:32]),
     .vdd_cntl(vdd_cntl[47:32]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net919), .purst(purst), .slf_op(slf_op_03[7:0]),
     .pgate(pgate[47:32]), .bnr_op(rgt_op_02[7:0]),
     .bnl_op(lft_op_02[7:0]), .tnr_op(rgt_op_04[7:0]),
     .tnl_op(lft_op_04[7:0]));
ltile4rev0 I_LT04 ( .prog(prog), .carry_out(net835),
     .lft_op(lft_op_04[7:0]), .sp12_h_l(sp12_h_l_04[23:0]),
     .sp4_h_l(sp4_h_l_04[47:0]), .sp4_v_b(sp4_v_b_04[47:0]),
     .sp12_v_b(net815[0:23]), .sp12_h_r(sp12_h_r_04[23:0]),
     .sp4_h_r(sp4_h_r_04[47:0]), .sp12_v_t(net843[0:23]),
     .sp4_v_t(sp4_v_b_05[47:0]), .sp4_r_v_b(sp4_r_v_b_04[47:0]),
     .wl(wl[63:48]), .top_op(slf_op_05[7:0]), .rgt_op(rgt_op_04[7:0]),
     .bot_op(slf_op_03[7:0]), .bl(bl[53:0]), .reset_b(reset_b[63:48]),
     .vdd_cntl(vdd_cntl[63:48]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net807), .purst(purst), .slf_op(slf_op_04[7:0]),
     .pgate(pgate[63:48]), .bnr_op(rgt_op_03[7:0]),
     .bnl_op(lft_op_03[7:0]), .tnr_op(rgt_op_05[7:0]),
     .tnl_op(lft_op_05[7:0]));
ltile4rev0 I_LT05 ( .prog(prog), .carry_out(net863),
     .lft_op(lft_op_05[7:0]), .sp12_h_l(sp12_h_l_05[23:0]),
     .sp4_h_l(sp4_h_l_05[47:0]), .sp4_v_b(sp4_v_b_05[47:0]),
     .sp12_v_b(net843[0:23]), .sp12_h_r(sp12_h_r_05[23:0]),
     .sp4_h_r(sp4_h_r_05[47:0]), .sp12_v_t(net871[0:23]),
     .sp4_v_t(sp4_v_b_06[47:0]), .sp4_r_v_b(sp4_r_v_b_05[47:0]),
     .wl(wl[79:64]), .top_op(slf_op_06[7:0]), .rgt_op(rgt_op_05[7:0]),
     .bot_op(slf_op_04[7:0]), .bl(bl[53:0]), .reset_b(reset_b[79:64]),
     .vdd_cntl(vdd_cntl[79:64]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net835), .purst(purst), .slf_op(slf_op_05[7:0]),
     .pgate(pgate[79:64]), .bnr_op(rgt_op_04[7:0]),
     .bnl_op(lft_op_04[7:0]), .tnr_op(rgt_op_06[7:0]),
     .tnl_op(lft_op_06[7:0]));
ltile4rev0 I_LT12 ( .prog(prog), .carry_out(net751),
     .lft_op(lft_op_12[7:0]), .sp12_h_l(sp12_h_l_12[23:0]),
     .sp4_h_l(sp4_h_l_12[47:0]), .sp4_v_b(sp4_v_b_12[47:0]),
     .sp12_v_b(net731[0:23]), .sp12_h_r(sp12_h_r_12[23:0]),
     .sp4_h_r(sp4_h_r_12[47:0]), .sp12_v_t(net759[0:23]),
     .sp4_v_t(sp4_v_b_13[47:0]), .sp4_r_v_b(sp4_r_v_b_12[47:0]),
     .wl(wl[191:176]), .top_op(slf_op_13[7:0]),
     .rgt_op(rgt_op_12[7:0]), .bot_op(slf_op_11[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[191:176]), .vdd_cntl(vdd_cntl[191:176]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net723), .purst(purst),
     .slf_op(slf_op_12[7:0]), .pgate(pgate[191:176]),
     .bnr_op(rgt_op_11[7:0]), .bnl_op(lft_op_11[7:0]),
     .tnr_op(rgt_op_13[7:0]), .tnl_op(lft_op_13[7:0]));
ltile4rev0 I_LT11 ( .prog(prog), .carry_out(net723),
     .lft_op(lft_op_11[7:0]), .sp12_h_l(sp12_h_l_11[23:0]),
     .sp4_h_l(sp4_h_l_11[47:0]), .sp4_v_b(sp4_v_b_11[47:0]),
     .sp12_v_b(net955[0:23]), .sp12_h_r(sp12_h_r_11[23:0]),
     .sp4_h_r(sp4_h_r_11[47:0]), .sp12_v_t(net731[0:23]),
     .sp4_v_t(sp4_v_b_12[47:0]), .sp4_r_v_b(sp4_r_v_b_11[47:0]),
     .wl(wl[175:160]), .top_op(slf_op_12[7:0]),
     .rgt_op(rgt_op_11[7:0]), .bot_op(slf_op_10[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[175:160]), .vdd_cntl(vdd_cntl[175:160]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net947), .purst(purst),
     .slf_op(slf_op_11[7:0]), .pgate(pgate[175:160]),
     .bnr_op(rgt_op_10[7:0]), .bnl_op(lft_op_10[7:0]),
     .tnr_op(rgt_op_12[7:0]), .tnl_op(lft_op_12[7:0]));
ltile4rev0 I_LT16 ( .prog(prog), .carry_out(carry_out),
     .lft_op(lft_op_16[7:0]), .sp12_h_l(sp12_h_l_16[23:0]),
     .sp4_h_l(sp4_h_l_16[47:0]), .sp4_v_b(sp4_v_b_16[47:0]),
     .sp12_v_b(net619[0:23]), .sp12_h_r(sp12_h_r_16[23:0]),
     .sp4_h_r(sp4_h_r_16[47:0]), .sp12_v_t(sp12_v_t_16[23:0]),
     .sp4_v_t(sp4_v_t_16[47:0]), .sp4_r_v_b(sp4_r_v_b_16[47:0]),
     .wl(wl[255:240]), .top_op(top_op_16[7:0]),
     .rgt_op(rgt_op_16[7:0]), .bot_op(slf_op_15[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[255:240]), .vdd_cntl(vdd_cntl[255:240]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net611), .purst(purst),
     .slf_op(slf_op_16[7:0]), .pgate(pgate[255:240]),
     .bnr_op(rgt_op_15[7:0]), .bnl_op(lft_op_15[7:0]),
     .tnr_op(tnr_op_16[7:0]), .tnl_op(tnl_op_16[7:0]));
ltile4rev0 I_LT14 ( .prog(prog), .carry_out(net667),
     .lft_op(lft_op_14[7:0]), .sp12_h_l(sp12_h_l_14[23:0]),
     .sp4_h_l(sp4_h_l_14[47:0]), .sp4_v_b(sp4_v_b_14[47:0]),
     .sp12_v_b(net647[0:23]), .sp12_h_r(sp12_h_r_14[23:0]),
     .sp4_h_r(sp4_h_r_14[47:0]), .sp12_v_t(net675[0:23]),
     .sp4_v_t(sp4_v_b_15[47:0]), .sp4_r_v_b(sp4_r_v_b_14[47:0]),
     .wl(wl[223:208]), .top_op(slf_op_15[7:0]),
     .rgt_op(rgt_op_14[7:0]), .bot_op(slf_op_13[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[223:208]), .vdd_cntl(vdd_cntl[223:208]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net639), .purst(purst),
     .slf_op(slf_op_14[7:0]), .pgate(pgate[223:208]),
     .bnr_op(rgt_op_13[7:0]), .bnl_op(lft_op_13[7:0]),
     .tnr_op(rgt_op_15[7:0]), .tnl_op(lft_op_15[7:0]));
ltile4rev0 I_LT13 ( .prog(prog), .carry_out(net639),
     .lft_op(lft_op_13[7:0]), .sp12_h_l(sp12_h_l_13[23:0]),
     .sp4_h_l(sp4_h_l_13[47:0]), .sp4_v_b(sp4_v_b_13[47:0]),
     .sp12_v_b(net759[0:23]), .sp12_h_r(sp12_h_r_13[23:0]),
     .sp4_h_r(sp4_h_r_13[47:0]), .sp12_v_t(net647[0:23]),
     .sp4_v_t(sp4_v_b_14[47:0]), .sp4_r_v_b(sp4_r_v_b_13[47:0]),
     .wl(wl[207:192]), .top_op(slf_op_14[7:0]),
     .rgt_op(rgt_op_13[7:0]), .bot_op(slf_op_12[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[207:192]), .vdd_cntl(vdd_cntl[207:192]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net751), .purst(purst),
     .slf_op(slf_op_13[7:0]), .pgate(pgate[207:192]),
     .bnr_op(rgt_op_12[7:0]), .bnl_op(lft_op_12[7:0]),
     .tnr_op(rgt_op_14[7:0]), .tnl_op(lft_op_14[7:0]));
ltile4rev0 I_LT15 ( .prog(prog), .carry_out(net611),
     .lft_op(lft_op_15[7:0]), .sp12_h_l(sp12_h_l_15[23:0]),
     .sp4_h_l(sp4_h_l_15[47:0]), .sp4_v_b(sp4_v_b_15[47:0]),
     .sp12_v_b(net675[0:23]), .sp12_h_r(sp12_h_r_15[23:0]),
     .sp4_h_r(sp4_h_r_15[47:0]), .sp12_v_t(net619[0:23]),
     .sp4_v_t(sp4_v_b_16[47:0]), .sp4_r_v_b(sp4_r_v_b_15[47:0]),
     .wl(wl[239:224]), .top_op(slf_op_16[7:0]),
     .rgt_op(rgt_op_15[7:0]), .bot_op(slf_op_14[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[239:224]), .vdd_cntl(vdd_cntl[239:224]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net667), .purst(purst),
     .slf_op(slf_op_15[7:0]), .pgate(pgate[239:224]),
     .bnr_op(rgt_op_14[7:0]), .bnl_op(lft_op_14[7:0]),
     .tnr_op(rgt_op_16[7:0]), .tnl_op(lft_op_16[7:0]));
ltile4rev0 I_LT01 ( .prog(prog), .carry_out(net891),
     .lft_op(lft_op_01[7:0]), .sp12_h_l(sp12_h_l_01[23:0]),
     .sp4_h_l(sp4_h_l_01[47:0]), .sp4_v_b(sp4_v_b_01[47:0]),
     .sp12_v_b(sp12_v_b__01[23:0]), .sp12_h_r(sp12_h_r_01[23:0]),
     .sp4_h_r(sp4_h_r_01[47:0]), .sp12_v_t(net899[0:23]),
     .sp4_v_t(sp4_v_b_02[47:0]), .sp4_r_v_b(sp4_r_v_b_01[47:0]),
     .wl(wl[15:0]), .top_op(slf_op_02[7:0]), .rgt_op(rgt_op_01[7:0]),
     .bot_op(bot_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[15:0]),
     .vdd_cntl(vdd_cntl[15:0]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(carry_in), .purst(purst), .slf_op(slf_op_01[7:0]),
     .pgate(pgate[15:0]), .bnr_op(bnr_op_01[7:0]),
     .bnl_op(bnl_op_01[7:0]), .tnr_op(rgt_op_02[7:0]),
     .tnl_op(lft_op_02[7:0]));
ltile4rev0 I_LT02 ( .prog(prog), .carry_out(net919),
     .lft_op(lft_op_02[7:0]), .sp12_h_l(sp12_h_l_02[23:0]),
     .sp4_h_l(sp4_h_l_02[47:0]), .sp4_v_b(sp4_v_b_02[47:0]),
     .sp12_v_b(net899[0:23]), .sp12_h_r(sp12_h_r_02[23:0]),
     .sp4_h_r(sp4_h_r_02[47:0]), .sp12_v_t(net927[0:23]),
     .sp4_v_t(sp4_v_b_03[47:0]), .sp4_r_v_b(sp4_r_v_b_02[47:0]),
     .wl(wl[31:16]), .top_op(slf_op_03[7:0]), .rgt_op(rgt_op_02[7:0]),
     .bot_op(slf_op_01[7:0]), .bl(bl[53:0]), .reset_b(reset_b[31:16]),
     .vdd_cntl(vdd_cntl[31:16]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net891), .purst(purst), .slf_op(slf_op_02[7:0]),
     .pgate(pgate[31:16]), .bnr_op(rgt_op_01[7:0]),
     .bnl_op(lft_op_01[7:0]), .tnr_op(rgt_op_03[7:0]),
     .tnl_op(lft_op_03[7:0]));
ltile4rev0 I_LT10 ( .prog(prog), .carry_out(net947),
     .lft_op(lft_op_10[7:0]), .sp12_h_l(sp12_h_l_10[23:0]),
     .sp4_h_l(sp4_h_l_10[47:0]), .sp4_v_b(sp4_v_b_10[47:0]),
     .sp12_v_b(net1039[0:23]), .sp12_h_r(sp12_h_r_10[23:0]),
     .sp4_h_r(sp4_h_r_10[47:0]), .sp12_v_t(net955[0:23]),
     .sp4_v_t(sp4_v_b_11[47:0]), .sp4_r_v_b(sp4_r_v_b_10[47:0]),
     .wl(wl[159:144]), .top_op(slf_op_11[7:0]),
     .rgt_op(rgt_op_10[7:0]), .bot_op(slf_op_09[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[159:144]), .vdd_cntl(vdd_cntl[159:144]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net1031), .purst(purst),
     .slf_op(slf_op_10[7:0]), .pgate(pgate[159:144]),
     .bnr_op(rgt_op_09[7:0]), .bnl_op(lft_op_09[7:0]),
     .tnr_op(rgt_op_11[7:0]), .tnl_op(lft_op_11[7:0]));
ltile4rev0 I_LT08 ( .prog(prog), .carry_out(net975),
     .lft_op(lft_op_08[7:0]), .sp12_h_l(sp12_h_l_08[23:0]),
     .sp4_h_l(sp4_h_l_08[47:0]), .sp4_v_b(sp4_v_b_08[47:0]),
     .sp12_v_b(net1011[0:23]), .sp12_h_r(sp12_h_r_08[23:0]),
     .sp4_h_r(sp4_h_r_08[47:0]), .sp12_v_t(net983[0:23]),
     .sp4_v_t(sp4_v_b_09[47:0]), .sp4_r_v_b(sp4_r_v_b_08[47:0]),
     .wl(wl[127:112]), .top_op(slf_op_09[7:0]),
     .rgt_op(rgt_op_08[7:0]), .bot_op(slf_op_07[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[127:112]), .vdd_cntl(vdd_cntl[127:112]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net1003), .purst(purst),
     .slf_op(slf_op_08[7:0]), .pgate(pgate[127:112]),
     .bnr_op(rgt_op_07[7:0]), .bnl_op(lft_op_07[7:0]),
     .tnr_op(rgt_op_09[7:0]), .tnl_op(lft_op_09[7:0]));
ltile4rev0 I_LT07 ( .prog(prog), .carry_out(net1003),
     .lft_op(lft_op_07[7:0]), .sp12_h_l(sp12_h_l_07[23:0]),
     .sp4_h_l(sp4_h_l_07[47:0]), .sp4_v_b(sp4_v_b_07[47:0]),
     .sp12_v_b(net787[0:23]), .sp12_h_r(sp12_h_r_07[23:0]),
     .sp4_h_r(sp4_h_r_07[47:0]), .sp12_v_t(net1011[0:23]),
     .sp4_v_t(sp4_v_b_08[47:0]), .sp4_r_v_b(sp4_r_v_b_07[47:0]),
     .wl(wl[111:96]), .top_op(slf_op_08[7:0]), .rgt_op(rgt_op_07[7:0]),
     .bot_op(slf_op_06[7:0]), .bl(bl[53:0]), .reset_b(reset_b[111:96]),
     .vdd_cntl(vdd_cntl[111:96]), .glb_netwk(glb_netwk[7:0]),
     .carry_in(net779), .purst(purst), .slf_op(slf_op_07[7:0]),
     .pgate(pgate[111:96]), .bnr_op(rgt_op_06[7:0]),
     .bnl_op(lft_op_06[7:0]), .tnr_op(rgt_op_08[7:0]),
     .tnl_op(lft_op_08[7:0]));
ltile4rev0 I_LT09 ( .prog(prog), .carry_out(net1031),
     .lft_op(lft_op_09[7:0]), .sp12_h_l(sp12_h_l_09[23:0]),
     .sp4_h_l(sp4_h_l_09[47:0]), .sp4_v_b(sp4_v_b_09[47:0]),
     .sp12_v_b(net983[0:23]), .sp12_h_r(sp12_h_r_09[23:0]),
     .sp4_h_r(sp4_h_r_09[47:0]), .sp12_v_t(net1039[0:23]),
     .sp4_v_t(sp4_v_b_10[47:0]), .sp4_r_v_b(sp4_r_v_b_09[47:0]),
     .wl(wl[143:128]), .top_op(slf_op_10[7:0]),
     .rgt_op(rgt_op_09[7:0]), .bot_op(slf_op_08[7:0]), .bl(bl[53:0]),
     .reset_b(reset_b[143:128]), .vdd_cntl(vdd_cntl[143:128]),
     .glb_netwk(glb_netwk[7:0]), .carry_in(net975), .purst(purst),
     .slf_op(slf_op_09[7:0]), .pgate(pgate[143:128]),
     .bnr_op(rgt_op_08[7:0]), .bnl_op(lft_op_08[7:0]),
     .tnr_op(rgt_op_10[7:0]), .tnl_op(lft_op_10[7:0]));
clk_colbuf8kx8 I78 ( .clko(glb_netwk[7:0]), .clki(glb_netwk_col[7:0]));

endmodule
// Library - misc, Cell - ml_mux2_hvt, View - schematic
// LAST TIME SAVED: Apr  5 16:31:59 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_mux2_hvt ( out, in0, in1, sel );
output  out;

input  in0, in1, sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



txgate_hvt I31 ( .in(in1), .out(out), .pp(net25), .nn(sel));
txgate_hvt I32 ( .in(in0), .out(out), .pp(sel), .nn(net25));
inv_hvt I220 ( .A(sel), .Y(net25));

endmodule
// Library - io, Cell - io_col4_BRAM_TOP, View - schematic
// LAST TIME SAVED: Feb  5 08:39:17 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module io_col4_BRAM_TOP ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [1:0]  spi_ss_in_b;
output [23:0]  cf;
output [1:0]  padeb;
output [1:0]  pado;
output [3:0]  slf_op;

inout [15:0]  sp4_v_t;
inout [17:0]  bl;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [15:0]  sp4_v_b;

input [1:0]  padin;
input [1:0]  spioeb;
input [15:0]  pgate;
input [15:0]  reset;
input [15:0]  wl;
input [15:0]  vdd_cntl;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [1:0]  spiout;
input [7:0]  lft_op;
input [7:0]  glb_netwk;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net129));
rm6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net129, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(net129),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net129));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net129), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));

endmodule
// Library - io, Cell - io_col4_TOP, View - schematic
// LAST TIME SAVED: Feb  5 08:41:32 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module io_col4_TOP ( cf, fabric_out, padeb, pado, sdo, slf_op,
     spi_ss_in_b, bl, sp4_h_l, sp4_v_b, sp4_v_t, sp12_h_l, bnl_op,
     bs_en, cdone_in, ceb, glb_netwk, hiz_b, hold, lft_op, mode, padin,
     pgate, prog, r, reset, sdi, shift, spioeb, spiout, tclk, tnl_op,
     update, vdd_cntl, wl );
output  fabric_out, sdo;


input  bs_en, cdone_in, ceb, hiz_b, hold, mode, prog, r, sdi, shift,
     tclk, update;

output [23:0]  cf;
output [1:0]  pado;
output [1:0]  padeb;
output [3:0]  slf_op;
output [1:0]  spi_ss_in_b;

inout [15:0]  sp4_v_b;
inout [23:0]  sp12_h_l;
inout [47:0]  sp4_h_l;
inout [17:0]  bl;
inout [15:0]  sp4_v_t;

input [1:0]  padin;
input [1:0]  spioeb;
input [15:0]  vdd_cntl;
input [15:0]  wl;
input [15:0]  pgate;
input [15:0]  reset;
input [1:0]  spiout;
input [7:0]  tnl_op;
input [7:0]  bnl_op;
input [7:0]  glb_netwk;
input [7:0]  lft_op;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:0]  om;

wire  [5:0]  ti;

wire  [1:0]  oenm;

wire  [3:0]  t_mid;

wire  [7:0]  lc_trk_g0;

wire  [7:0]  lc_trk_g1;



inv_hvt I90 ( .A(prog), .Y(progb));
inv_hvt I89 ( .A(progb), .Y(net128));
rm6  R0_15_ ( .MINUS(sp4_v_b[15]), .PLUS(sp4_v_t[11]));
rm6  R0_14_ ( .MINUS(sp4_v_b[14]), .PLUS(sp4_v_t[10]));
rm6  R0_13_ ( .MINUS(sp4_v_b[13]), .PLUS(sp4_v_t[9]));
rm6  R0_12_ ( .MINUS(sp4_v_b[12]), .PLUS(sp4_v_t[8]));
rm6  R0_11_ ( .MINUS(sp4_v_b[11]), .PLUS(sp4_v_t[7]));
rm6  R0_10_ ( .MINUS(sp4_v_b[10]), .PLUS(sp4_v_t[6]));
rm6  R0_9_ ( .MINUS(sp4_v_b[9]), .PLUS(sp4_v_t[5]));
rm6  R0_8_ ( .MINUS(sp4_v_b[8]), .PLUS(sp4_v_t[4]));
rm6  R0_7_ ( .MINUS(sp4_v_b[7]), .PLUS(sp4_v_t[3]));
rm6  R0_6_ ( .MINUS(sp4_v_b[6]), .PLUS(sp4_v_t[2]));
rm6  R0_5_ ( .MINUS(sp4_v_b[5]), .PLUS(sp4_v_t[1]));
rm6  R0_4_ ( .MINUS(sp4_v_b[4]), .PLUS(sp4_v_t[0]));
rm6  R0_3_ ( .MINUS(t_mid[3]), .PLUS(sp4_v_t[15]));
rm6  R0_2_ ( .MINUS(t_mid[2]), .PLUS(sp4_v_t[14]));
rm6  R0_1_ ( .MINUS(t_mid[1]), .PLUS(sp4_v_t[13]));
rm6  R0_0_ ( .MINUS(t_mid[0]), .PLUS(sp4_v_t[12]));
io_col_odrv4_x40bare I_io_odrv4x40 ( cf[23:0], bl[3:0], sp4_h_l[47:0],
     sp4_v_b[15:0], {slf_op[0], slf_op[2]}, {slf_op[1], slf_op[3]},
     {pgate[14], pgate[15], pgate[12], pgate[13], pgate[10], pgate[11],
     pgate[8], pgate[9], pgate[6], pgate[7], pgate[4], pgate[5],
     pgate[2], pgate[3], pgate[0], pgate[1]}, net128, {reset[14],
     reset[15], reset[12], reset[13], reset[10], reset[11], reset[8],
     reset[9], reset[6], reset[7], reset[4], reset[5], reset[2],
     reset[3], reset[0], reset[1]}, {vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]},
     {wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]});
io_gmux_x16bare I_io_gmux_x16 ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .min7({sp4_h_l[47], sp4_h_l[39], sp4_h_l[31], sp4_h_l[23],
     sp4_h_l[15], sp4_h_l[7], sp12_h_l[23], sp12_h_l[15], sp12_h_l[7],
     sp4_v_b[15], sp4_v_b[7], bnl_op[7], lft_op[7], tnl_op[7], gnd_,
     gnd_}), .min6({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30], sp4_h_l[22],
     sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14], sp12_h_l[6],
     sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6], tnl_op[6], gnd_,
     gnd_}), .min5({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min4({sp4_h_l[44], sp4_h_l[36], sp4_h_l[28], sp4_h_l[20],
     sp4_h_l[12], sp4_h_l[4], sp12_h_l[20], sp12_h_l[12], sp12_h_l[4],
     sp4_v_b[12], sp4_v_b[4], bnl_op[4], lft_op[4], tnl_op[4], gnd_,
     gnd_}), .min3({sp4_h_l[43], sp4_h_l[35], sp4_h_l[27], sp4_h_l[19],
     sp4_h_l[11], sp4_h_l[3], sp12_h_l[19], sp12_h_l[11], sp12_h_l[3],
     sp4_v_b[11], sp4_v_b[3], bnl_op[3], lft_op[3], tnl_op[3], gnd_,
     gnd_}), .min2({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26], sp4_h_l[18],
     sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10], sp12_h_l[2],
     sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2], tnl_op[2], gnd_,
     gnd_}), .min1({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min0({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min8({sp4_h_l[40], sp4_h_l[32], sp4_h_l[24], sp4_h_l[16],
     sp4_h_l[8], sp4_h_l[0], sp12_h_l[16], sp12_h_l[8], sp12_h_l[0],
     sp4_v_b[8], sp4_v_b[0], bnl_op[0], lft_op[0], tnl_op[0], gnd_,
     gnd_}), .min9({sp4_h_l[41], sp4_h_l[33], sp4_h_l[25], sp4_h_l[17],
     sp4_h_l[9], sp4_h_l[1], sp12_h_l[17], sp12_h_l[9], sp12_h_l[1],
     sp4_v_b[9], sp4_v_b[1], bnl_op[1], lft_op[1], tnl_op[1], gnd_,
     gnd_}), .min10({sp4_h_l[42], sp4_h_l[34], sp4_h_l[26],
     sp4_h_l[18], sp4_h_l[10], sp4_h_l[2], sp12_h_l[18], sp12_h_l[10],
     sp12_h_l[2], sp4_v_b[10], sp4_v_b[2], bnl_op[2], lft_op[2],
     tnl_op[2], gnd_, gnd_}), .min11({sp4_h_l[43], sp4_h_l[35],
     sp4_h_l[27], sp4_h_l[19], sp4_h_l[11], sp4_h_l[3], sp12_h_l[19],
     sp12_h_l[11], sp12_h_l[3], sp4_v_b[11], sp4_v_b[3], bnl_op[3],
     lft_op[3], tnl_op[3], gnd_, gnd_}), .min12({sp4_h_l[44],
     sp4_h_l[36], sp4_h_l[28], sp4_h_l[20], sp4_h_l[12], sp4_h_l[4],
     sp12_h_l[20], sp12_h_l[12], sp12_h_l[4], sp4_v_b[12], sp4_v_b[4],
     bnl_op[4], lft_op[4], tnl_op[4], gnd_, gnd_}),
     .min13({sp4_h_l[45], sp4_h_l[37], sp4_h_l[29], sp4_h_l[21],
     sp4_h_l[13], sp4_h_l[5], sp12_h_l[21], sp12_h_l[13], sp12_h_l[5],
     sp4_v_b[13], sp4_v_b[5], bnl_op[5], lft_op[5], tnl_op[5], gnd_,
     gnd_}), .min14({sp4_h_l[46], sp4_h_l[38], sp4_h_l[30],
     sp4_h_l[22], sp4_h_l[14], sp4_h_l[6], sp12_h_l[22], sp12_h_l[14],
     sp12_h_l[6], sp4_v_b[14], sp4_v_b[6], bnl_op[6], lft_op[6],
     tnl_op[6], gnd_, gnd_}), .min15({sp4_h_l[47], sp4_h_l[39],
     sp4_h_l[31], sp4_h_l[23], sp4_h_l[15], sp4_h_l[7], sp12_h_l[23],
     sp12_h_l[15], sp12_h_l[7], sp4_v_b[15], sp4_v_b[7], bnl_op[7],
     lft_op[7], tnl_op[7], gnd_, gnd_}), .bl(bl[9:4]), .wl({wl[14],
     wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9], wl[6],
     wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}),
     .lc_trk_g0(lc_trk_g0[7:0]), .prog(net128),
     .lc_trk_g1(lc_trk_g1[7:0]));
sbox1_colbdlc Isbox1_col ( .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .outclk(outclk), .fabric_out(fabric_out), .min6({lc_trk_g1[6],
     lc_trk_g1[4], lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7],
     lc_trk_g0[5], lc_trk_g0[3], lc_trk_g0[1]}),
     .inclk_in({lc_trk_g1[3], lc_trk_g1[0], lc_trk_g0[3], lc_trk_g0[0],
     glb_netwk[7:0]}), .ceb_in({lc_trk_g1[5], lc_trk_g1[2],
     lc_trk_g0[5], lc_trk_g0[2], glb_netwk[7], glb_netwk[5],
     glb_netwk[3], glb_netwk[1]}), .clk_in({lc_trk_g1[4], lc_trk_g1[1],
     lc_trk_g0[4], lc_trk_g0[1], glb_netwk[7:0]}), .update(update),
     .spiout(spiout[1:0]), .spioeb(spioeb[1:0]), .padin(padin[1:0]),
     .out(om[1:0]), .oeb(oenm[1:0]), .min5({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min4({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min3({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min2({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .min1({lc_trk_g1[7], lc_trk_g1[5],
     lc_trk_g1[3], lc_trk_g1[1], lc_trk_g0[6], lc_trk_g0[4],
     lc_trk_g0[2], lc_trk_g0[0]}), .min0({lc_trk_g1[6], lc_trk_g1[4],
     lc_trk_g1[2], lc_trk_g1[0], lc_trk_g0[7], lc_trk_g0[5],
     lc_trk_g0[3], lc_trk_g0[1]}), .cdone_in(cdone_in), .bs_en(bs_en),
     .updt(enable_update), .ti(ti[5:0]),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .pado(pado[1:0]),
     .padeb(padeb[1:0]), .t_mid(t_mid[3:0]), .sp4_v_b(sp4_v_b[3:0]),
     .r({sp4_h_l[19], sp4_h_l[13], sp4_h_l[7], sp4_h_l[1]}),
     .l({sp4_h_l[43], sp4_h_l[37], sp4_h_l[31], sp4_h_l[25]}),
     .bl(bl[15:10]), .inclk(inclk), .wl({wl[14], wl[15], wl[12],
     wl[13], wl[10], wl[11], wl[8], wl[9], wl[6], wl[7], wl[4], wl[5],
     wl[2], wl[3], wl[0], wl[1]}), .reset({reset[14], reset[15],
     reset[12], reset[13], reset[10], reset[11], reset[8], reset[9],
     reset[6], reset[7], reset[4], reset[5], reset[2], reset[3],
     reset[0], reset[1]}), .pgate({pgate[14], pgate[15], pgate[12],
     pgate[13], pgate[10], pgate[11], pgate[8], pgate[9], pgate[6],
     pgate[7], pgate[4], pgate[5], pgate[2], pgate[3], pgate[0],
     pgate[1]}), .prog(net128));
ioe_col2 I_ioe_col2 ( .ceb(ceb), .vdd_cntl({vdd_cntl[14], vdd_cntl[15],
     vdd_cntl[12], vdd_cntl[13], vdd_cntl[10], vdd_cntl[11],
     vdd_cntl[8], vdd_cntl[9], vdd_cntl[6], vdd_cntl[7], vdd_cntl[4],
     vdd_cntl[5], vdd_cntl[2], vdd_cntl[3], vdd_cntl[0], vdd_cntl[1]}),
     .dout(slf_op[3:0]), .outclk(outclk), .hold(hold), .rstio(r),
     .wl({wl[14], wl[15], wl[12], wl[13], wl[10], wl[11], wl[8], wl[9],
     wl[6], wl[7], wl[4], wl[5], wl[2], wl[3], wl[0], wl[1]}),
     .reset({reset[14], reset[15], reset[12], reset[13], reset[10],
     reset[11], reset[8], reset[9], reset[6], reset[7], reset[4],
     reset[5], reset[2], reset[3], reset[0], reset[1]}),
     .pgate({pgate[14], pgate[15], pgate[12], pgate[13], pgate[10],
     pgate[11], pgate[8], pgate[9], pgate[6], pgate[7], pgate[4],
     pgate[5], pgate[2], pgate[3], pgate[0], pgate[1]}), .hiz_b(hiz_b),
     .update(enable_update), .ti(ti[5:0]), .tclk(tclk), .shift(shift),
     .sdi(sdi), .prog(net128), .padin(padin[1:0]), .mode(mode),
     .inclk(inclk), .bs_en(bs_en), .sp12_h_l(sp12_h_l[23:0]),
     .sdo(sdo), .pado(om[1:0]), .padeb(oenm[1:0]), .bl(bl[17:16]));

endmodule
// Library - leafcell, Cell - preio_top_r, View - schematic
// LAST TIME SAVED: Sep 18 15:38:10 2008
// NETLIST TIME: Nov 14 16:17:18 2008
`timescale 1ns / 1ns 

module preio_top_r ( bs_en_o, ceb_o, cf_t, fabric_out_17_33, hiz_b_o,
     mode_o, padeb_t, padin_192, pado_t, r_o, sdo, shift_o,
     slf_op_17_33, slf_op_18_33, slf_op_19_33, slf_op_20_33,
     slf_op_21_33, slf_op_22_33, slf_op_23_33, slf_op_24_33,
     slf_op_25_33, slf_op_26_33, slf_op_27_33, slf_op_28_33,
     slf_op_29_33, slf_op_30_33, slf_op_31_33, slf_op_32_33, tclk_o,
     update_o, bl_17, bl_18, bl_19, bl_20, bl_21, bl_22, bl_23, bl_24,
     bl_25, bl_26, bl_27, bl_28, bl_29, bl_30, bl_31, bl_32,
     sp4_h_l_17_33, sp4_h_r_32_33, sp4_v_b_17_33, sp4_v_b_18_33,
     sp4_v_b_19_33, sp4_v_b_20_33, sp4_v_b_21_33, sp4_v_b_22_33,
     sp4_v_b_23_33, sp4_v_b_24_33, sp4_v_b_25_33, sp4_v_b_26_33,
     sp4_v_b_27_33, sp4_v_b_28_33, sp4_v_b_29_33, sp4_v_b_30_33,
     sp4_v_b_31_33, sp4_v_b_32_33, sp12_v_b_17_33, sp12_v_b_18_33,
     sp12_v_b_19_33, sp12_v_b_20_33, sp12_v_b_21_33, sp12_v_b_22_33,
     sp12_v_b_23_33, sp12_v_b_24_33, sp12_v_b_25_33, sp12_v_b_26_33,
     sp12_v_b_27_33, sp12_v_b_28_33, sp12_v_b_29_33, sp12_v_b_30_33,
     sp12_v_b_31_33, sp12_v_b_32_33, bnl_op_17_33, bnr_op_32_33,
     bs_en_i, ceb_i, end_of_startup_top_r, glb_net_17, glb_net_18,
     glb_net_19, glb_net_20, glb_net_21, glb_net_22, glb_net_23,
     glb_net_24, glb_net_25, glb_net_26, glb_net_27, glb_net_28,
     glb_net_29, glb_net_30, glb_net_31, glb_net_32, hiz_b_i, hold_t_r,
     lft_op_17_33, lft_op_18_33, lft_op_19_33, lft_op_20_33,
     lft_op_21_33, lft_op_22_33, lft_op_23_33, lft_op_24_33,
     lft_op_25_33, lft_op_26_33, lft_op_27_33, lft_op_28_33,
     lft_op_29_33, lft_op_30_33, lft_op_31_33, lft_op_32_33, mode_i,
     padin_t, pgate_r, prog, r_i, reset_r, sdi, shift_i, tclk_i,
     tiegnd, tievdd, update_i, vdd_cntl_r, wl_r );
output  bs_en_o, ceb_o, fabric_out_17_33, hiz_b_o, mode_o, padin_192,
     r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_r, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, tiegnd, tievdd, update_i;

output [3:0]  slf_op_28_33;
output [3:0]  slf_op_24_33;
output [3:0]  slf_op_22_33;
output [3:0]  slf_op_18_33;
output [3:0]  slf_op_29_33;
output [3:0]  slf_op_21_33;
output [3:0]  slf_op_20_33;
output [3:0]  slf_op_23_33;
output [3:0]  slf_op_17_33;
output [3:0]  slf_op_19_33;
output [3:0]  slf_op_31_33;
output [3:0]  slf_op_25_33;
output [59:30]  padeb_t;
output [59:30]  pado_t;
output [383:0]  cf_t;
output [3:0]  slf_op_30_33;
output [3:0]  slf_op_26_33;
output [3:0]  slf_op_32_33;
output [3:0]  slf_op_27_33;

inout [23:0]  sp12_v_b_17_33;
inout [47:0]  sp4_v_b_23_33;
inout [47:0]  sp4_v_b_27_33;
inout [47:0]  sp4_v_b_26_33;
inout [47:0]  sp4_v_b_31_33;
inout [47:0]  sp4_v_b_29_33;
inout [47:0]  sp4_v_b_21_33;
inout [23:0]  sp12_v_b_32_33;
inout [23:0]  sp12_v_b_25_33;
inout [47:0]  sp4_v_b_30_33;
inout [23:0]  sp12_v_b_24_33;
inout [53:0]  bl_29;
inout [53:0]  bl_28;
inout [23:0]  sp12_v_b_22_33;
inout [53:0]  bl_27;
inout [23:0]  sp12_v_b_28_33;
inout [23:0]  sp12_v_b_31_33;
inout [47:0]  sp4_v_b_19_33;
inout [23:0]  sp12_v_b_21_33;
inout [47:0]  sp4_v_b_22_33;
inout [15:0]  sp4_h_r_32_33;
inout [23:0]  sp12_v_b_19_33;
inout [53:0]  bl_30;
inout [47:0]  sp4_v_b_24_33;
inout [47:0]  sp4_v_b_18_33;
inout [15:0]  sp4_h_l_17_33;
inout [23:0]  sp12_v_b_26_33;
inout [53:0]  bl_26;
inout [47:0]  sp4_v_b_25_33;
inout [23:0]  sp12_v_b_23_33;
inout [23:0]  sp12_v_b_18_33;
inout [47:0]  sp4_v_b_28_33;
inout [53:0]  bl_23;
inout [53:0]  bl_19;
inout [53:0]  bl_20;
inout [53:0]  bl_21;
inout [53:0]  bl_22;
inout [41:0]  bl_25;
inout [53:0]  bl_32;
inout [53:0]  bl_18;
inout [53:0]  bl_17;
inout [23:0]  sp12_v_b_29_33;
inout [23:0]  sp12_v_b_30_33;
inout [23:0]  sp12_v_b_20_33;
inout [53:0]  bl_24;
inout [53:0]  bl_31;
inout [47:0]  sp4_v_b_32_33;
inout [47:0]  sp4_v_b_20_33;
inout [47:0]  sp4_v_b_17_33;
inout [23:0]  sp12_v_b_27_33;

input [7:0]  lft_op_22_33;
input [7:0]  glb_net_32;
input [7:0]  lft_op_24_33;
input [7:0]  lft_op_31_33;
input [7:0]  bnl_op_17_33;
input [7:0]  glb_net_28;
input [15:0]  wl_r;
input [7:0]  glb_net_24;
input [7:0]  lft_op_26_33;
input [7:0]  lft_op_17_33;
input [7:0]  glb_net_18;
input [7:0]  glb_net_29;
input [7:0]  lft_op_18_33;
input [7:0]  glb_net_30;
input [7:0]  glb_net_20;
input [7:0]  lft_op_32_33;
input [7:0]  lft_op_20_33;
input [7:0]  glb_net_26;
input [7:0]  bnr_op_32_33;
input [7:0]  lft_op_23_33;
input [7:0]  glb_net_25;
input [7:0]  glb_net_21;
input [7:0]  lft_op_28_33;
input [7:0]  lft_op_30_33;
input [15:0]  vdd_cntl_r;
input [7:0]  glb_net_31;
input [7:0]  lft_op_25_33;
input [7:0]  lft_op_27_33;
input [7:0]  glb_net_17;
input [59:30]  padin_t;
input [32:17]  end_of_startup_top_r;
input [7:0]  glb_net_22;
input [7:0]  glb_net_23;
input [7:0]  glb_net_27;
input [7:0]  glb_net_19;
input [7:0]  lft_op_21_33;
input [7:0]  lft_op_29_33;
input [15:0]  reset_r;
input [7:0]  lft_op_19_33;
input [15:0]  pgate_r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net842;

wire  [0:1]  net813;

wire  [0:1]  net1246;

wire  [0:1]  net1255;

wire  [0:1]  net1237;

wire  [0:15]  net757;

wire  [0:15]  net792;

wire  [0:15]  net827;

wire  [0:15]  net967;

wire  [0:1]  net1128;

wire  [0:1]  net1244;

wire  [0:1]  net848;

wire  [0:1]  net1235;

wire  [0:1]  net1257;

wire  [0:15]  net1107;

wire  [0:1]  net1243;

wire  [0:15]  net1212;

wire  [0:15]  net890;

wire  [0:15]  net722;

wire  [0:15]  net932;

wire  [0:15]  net687;

wire  [0:15]  net1177;

wire  [0:15]  net1002;

wire  [0:1]  net778;

wire  [0:1]  net844;

wire  [0:15]  net1072;

wire  [0:1]  net1163;

wire  [0:15]  net1142;

wire  [0:15]  net1037;

wire  [0:1]  net1198;

wire  [0:1]  net918;

wire  [0:1]  net1245;

wire  [0:1]  net953;



lowla_modified I342 ( .clk(tclk_i), .min(net0615), .lao(net831));
bram_bufferx4x6 I345 ( .in(sdi), .out(net0615));
fabric_buf8k I343 ( .f_in(net790), .f_out(fabric_out_17_33));
fabric_buf8k I344 ( .f_in(padin_t[30]), .f_out(padin_192));
tckbufx16 I339 ( .in(tclk_i), .out(tclk_o));
io_col4_BRAM_TOP I_IO_25_33bram ( .ceb(ceb_o), .bl({bl_25[5], bl_25[4],
     bl_25[37], bl_25[36], bl_25[35], bl_25[34], bl_25[33], bl_25[32],
     bl_25[14], bl_25[20], bl_25[19], bl_25[18], bl_25[17], bl_25[16],
     bl_25[27], bl_25[26], bl_25[25], bl_25[23]}), .sdo(net866),
     .sdi(net656), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[25]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[47:46]), .pado(pado_t[47:46]),
     .padeb(padeb_t[47:46]), .sp4_h_l(sp4_v_b_25_33[47:0]),
     .sp12_h_l(sp12_v_b_25_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1244[0:1]), .tnl_op(lft_op_24_33[7:0]),
     .lft_op(lft_op_25_33[7:0]), .bnl_op(lft_op_26_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[215:192]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_25_33[3:0]), .glb_netwk(glb_net_25[7:0]),
     .hold(hold_t_r), .fabric_out(net1236), .sp4_v_t(net890[0:15]),
     .sp4_v_b(net687[0:15]));
io_col4_TOP I_IO_18_33 ( .ceb(ceb_o), .bl({bl_18[5], bl_18[4],
     bl_18[37], bl_18[36], bl_18[35], bl_18[34], bl_18[33], bl_18[32],
     bl_18[14], bl_18[20], bl_18[19], bl_18[18], bl_18[17], bl_18[16],
     bl_18[27], bl_18[26], bl_18[25], bl_18[23]}), .sdo(net761),
     .sdi(net691), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[18]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[33:32]), .pado(pado_t[33:32]),
     .padeb(padeb_t[33:32]), .sp4_h_l(sp4_v_b_18_33[47:0]),
     .sp12_h_l(sp12_v_b_18_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1235[0:1]), .tnl_op(lft_op_17_33[7:0]),
     .lft_op(lft_op_18_33[7:0]), .bnl_op(lft_op_19_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[47:24]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_18_33[3:0]), .glb_netwk(glb_net_18[7:0]),
     .hold(hold_t_r), .fabric_out(net1248), .sp4_v_t(net792[0:15]),
     .sp4_v_b(net722[0:15]));
io_col4_TOP I_IO_28_33 ( .ceb(ceb_o), .bl({bl_28[5], bl_28[4],
     bl_28[37], bl_28[36], bl_28[35], bl_28[34], bl_28[33], bl_28[32],
     bl_28[14], bl_28[20], bl_28[19], bl_28[18], bl_28[17], bl_28[16],
     bl_28[27], bl_28[26], bl_28[25], bl_28[23]}), .sdo(net796),
     .sdi(net726), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[28]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[53:52]), .pado(pado_t[53:52]),
     .padeb(padeb_t[53:52]), .sp4_h_l(sp4_v_b_28_33[47:0]),
     .sp12_h_l(sp12_v_b_28_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1245[0:1]), .tnl_op(lft_op_27_33[7:0]),
     .lft_op(lft_op_28_33[7:0]), .bnl_op(lft_op_29_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[287:264]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_28_33[3:0]), .glb_netwk(glb_net_28[7:0]),
     .hold(hold_t_r), .fabric_out(net1249), .sp4_v_t(net827[0:15]),
     .sp4_v_b(net757[0:15]));
io_col4_TOP I_IO_17_33 ( .ceb(ceb_o), .bl({bl_17[5], bl_17[4],
     bl_17[37], bl_17[36], bl_17[35], bl_17[34], bl_17[33], bl_17[32],
     bl_17[14], bl_17[20], bl_17[19], bl_17[18], bl_17[17], bl_17[16],
     bl_17[27], bl_17[26], bl_17[25], bl_17[23]}), .sdo(sdo),
     .sdi(net761), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[17]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[31:30]), .pado(pado_t[31:30]),
     .padeb(padeb_t[31:30]), .sp4_h_l(sp4_v_b_17_33[47:0]),
     .sp12_h_l(sp12_v_b_17_33[23:0]), .prog(prog),
     .spi_ss_in_b(net778[0:1]), .tnl_op(bnl_op_17_33[7:0]),
     .lft_op(lft_op_17_33[7:0]), .bnl_op(lft_op_18_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[23:0]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_17_33[3:0]), .glb_netwk(glb_net_17[7:0]),
     .hold(hold_t_r), .fabric_out(net790),
     .sp4_v_t(sp4_h_l_17_33[15:0]), .sp4_v_b(net792[0:15]));
io_col4_TOP I_IO_27_33 ( .ceb(ceb_o), .bl({bl_27[5], bl_27[4],
     bl_27[37], bl_27[36], bl_27[35], bl_27[34], bl_27[33], bl_27[32],
     bl_27[14], bl_27[20], bl_27[19], bl_27[18], bl_27[17], bl_27[16],
     bl_27[27], bl_27[26], bl_27[25], bl_27[23]}), .sdo(net1181),
     .sdi(net796), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[27]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[51:50]), .pado(pado_t[51:50]),
     .padeb(padeb_t[51:50]), .sp4_h_l(sp4_v_b_27_33[47:0]),
     .sp12_h_l(sp12_v_b_27_33[23:0]), .prog(prog),
     .spi_ss_in_b(net813[0:1]), .tnl_op(lft_op_26_33[7:0]),
     .lft_op(lft_op_27_33[7:0]), .bnl_op(lft_op_28_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[263:240]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_27_33[3:0]), .glb_netwk(glb_net_27[7:0]),
     .hold(hold_t_r), .fabric_out(net825), .sp4_v_t(net1212[0:15]),
     .sp4_v_b(net827[0:15]));
io_col4_TOP I_IO_32_33 ( .ceb(ceb_o), .bl({bl_32[5], bl_32[4],
     bl_32[37], bl_32[36], bl_32[35], bl_32[34], bl_32[33], bl_32[32],
     bl_32[14], bl_32[20], bl_32[19], bl_32[18], bl_32[17], bl_32[16],
     bl_32[27], bl_32[26], bl_32[25], bl_32[23]}), .sdo(net1111),
     .sdi(net831), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[32]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(net842[0:1]), .pado(net842[0:1]), .padeb(net844[0:1]),
     .sp4_h_l(sp4_v_b_32_33[47:0]), .sp12_h_l(sp12_v_b_32_33[23:0]),
     .prog(prog), .spi_ss_in_b(net848[0:1]),
     .tnl_op(lft_op_31_33[7:0]), .lft_op(lft_op_32_33[7:0]),
     .bnl_op(bnr_op_32_33[7:0]), .pgate(pgate_r[15:0]),
     .reset(reset_r[15:0]), .wl(wl_r[15:0]), .cf(cf_t[383:360]),
     .vdd_cntl(vdd_cntl_r[15:0]), .slf_op(slf_op_32_33[3:0]),
     .glb_netwk(glb_net_32[7:0]), .hold(hold_t_r), .fabric_out(net860),
     .sp4_v_t(net1142[0:15]), .sp4_v_b(sp4_h_r_32_33[15:0]));
io_col4_TOP I_IO_24_33 ( .ceb(ceb_o), .bl({bl_24[5], bl_24[4],
     bl_24[37], bl_24[36], bl_24[35], bl_24[34], bl_24[33], bl_24[32],
     bl_24[14], bl_24[20], bl_24[19], bl_24[18], bl_24[17], bl_24[16],
     bl_24[27], bl_24[26], bl_24[25], bl_24[23]}), .sdo(net936),
     .sdi(net866), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[24]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[45:44]), .pado(pado_t[45:44]),
     .padeb(padeb_t[45:44]), .sp4_v_t(net967[0:15]),
     .sp4_h_l(sp4_v_b_24_33[47:0]), .sp12_h_l(sp12_v_b_24_33[23:0]),
     .prog(prog), .spi_ss_in_b(net1255[0:1]),
     .tnl_op(lft_op_23_33[7:0]), .lft_op(lft_op_24_33[7:0]),
     .bnl_op(lft_op_25_33[7:0]), .pgate(pgate_r[15:0]),
     .reset(reset_r[15:0]), .sp4_v_b(net890[0:15]), .wl(wl_r[15:0]),
     .cf(cf_t[191:168]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_24_33[3:0]), .glb_netwk(glb_net_24[7:0]),
     .hold(hold_t_r), .fabric_out(net1252));
io_col4_TOP I_IO_21_33 ( .ceb(ceb_o), .bl({bl_21[5], bl_21[4],
     bl_21[37], bl_21[36], bl_21[35], bl_21[34], bl_21[33], bl_21[32],
     bl_21[14], bl_21[20], bl_21[19], bl_21[18], bl_21[17], bl_21[16],
     bl_21[27], bl_21[26], bl_21[25], bl_21[23]}), .sdo(net1146),
     .sdi(net901), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[21]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[39:38]), .pado(pado_t[39:38]),
     .padeb(padeb_t[39:38]), .sp4_h_l(sp4_v_b_21_33[47:0]),
     .sp12_h_l(sp12_v_b_21_33[23:0]), .prog(prog),
     .spi_ss_in_b(net918[0:1]), .tnl_op(lft_op_20_33[7:0]),
     .lft_op(lft_op_21_33[7:0]), .bnl_op(lft_op_22_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[119:96]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_21_33[3:0]), .glb_netwk(glb_net_21[7:0]),
     .hold(hold_t_r), .fabric_out(net1240), .sp4_v_t(net1177[0:15]),
     .sp4_v_b(net932[0:15]));
io_col4_TOP I_IO_23_33 ( .ceb(ceb_o), .bl({bl_23[5], bl_23[4],
     bl_23[37], bl_23[36], bl_23[35], bl_23[34], bl_23[33], bl_23[32],
     bl_23[14], bl_23[20], bl_23[19], bl_23[18], bl_23[17], bl_23[16],
     bl_23[27], bl_23[26], bl_23[25], bl_23[23]}), .sdo(net971),
     .sdi(net936), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[23]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[43:42]), .pado(pado_t[43:42]),
     .padeb(padeb_t[43:42]), .sp4_h_l(sp4_v_b_23_33[47:0]),
     .sp12_h_l(sp12_v_b_23_33[23:0]), .prog(prog),
     .spi_ss_in_b(net953[0:1]), .tnl_op(lft_op_22_33[7:0]),
     .lft_op(lft_op_23_33[7:0]), .bnl_op(lft_op_24_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[167:144]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_23_33[3:0]), .glb_netwk(glb_net_23[7:0]),
     .hold(hold_t_r), .fabric_out(net965), .sp4_v_t(net1002[0:15]),
     .sp4_v_b(net967[0:15]));
io_col4_TOP I_IO_22_33 ( .ceb(ceb_o), .bl({bl_22[5], bl_22[4],
     bl_22[37], bl_22[36], bl_22[35], bl_22[34], bl_22[33], bl_22[32],
     bl_22[14], bl_22[20], bl_22[19], bl_22[18], bl_22[17], bl_22[16],
     bl_22[27], bl_22[26], bl_22[25], bl_22[23]}), .sdo(net901),
     .sdi(net971), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[22]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[41:40]), .pado(pado_t[41:40]),
     .padeb(padeb_t[41:40]), .sp4_h_l(sp4_v_b_22_33[47:0]),
     .sp12_h_l(sp12_v_b_22_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1237[0:1]), .tnl_op(lft_op_21_33[7:0]),
     .lft_op(lft_op_22_33[7:0]), .bnl_op(lft_op_23_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[143:120]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_22_33[3:0]), .glb_netwk(glb_net_22[7:0]),
     .hold(hold_t_r), .fabric_out(net1000), .sp4_v_t(net932[0:15]),
     .sp4_v_b(net1002[0:15]));
io_col4_TOP I_IO_19_33 ( .ceb(ceb_o), .bl({bl_19[5], bl_19[4],
     bl_19[37], bl_19[36], bl_19[35], bl_19[34], bl_19[33], bl_19[32],
     bl_19[14], bl_19[20], bl_19[19], bl_19[18], bl_19[17], bl_19[16],
     bl_19[27], bl_19[26], bl_19[25], bl_19[23]}), .sdo(net691),
     .sdi(net1006), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[19]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[35:34]), .pado(pado_t[35:34]),
     .padeb(padeb_t[35:34]), .sp4_h_l(sp4_v_b_19_33[47:0]),
     .sp12_h_l(sp12_v_b_19_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1243[0:1]), .tnl_op(lft_op_18_33[7:0]),
     .lft_op(lft_op_19_33[7:0]), .bnl_op(lft_op_20_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[71:48]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_19_33[3:0]), .glb_netwk(glb_net_19[7:0]),
     .hold(hold_t_r), .fabric_out(net1239), .sp4_v_t(net722[0:15]),
     .sp4_v_b(net1037[0:15]));
io_col4_TOP I_IO_30_33 ( .ceb(ceb_o), .bl({bl_30[5], bl_30[4],
     bl_30[37], bl_30[36], bl_30[35], bl_30[34], bl_30[33], bl_30[32],
     bl_30[14], bl_30[20], bl_30[19], bl_30[18], bl_30[17], bl_30[16],
     bl_30[27], bl_30[26], bl_30[25], bl_30[23]}), .sdo(net1076),
     .sdi(net1041), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[30]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[57:56]), .pado(pado_t[57:56]),
     .padeb(padeb_t[57:56]), .sp4_h_l(sp4_v_b_30_33[47:0]),
     .sp12_h_l(sp12_v_b_30_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1257[0:1]), .tnl_op(lft_op_29_33[7:0]),
     .lft_op(lft_op_30_33[7:0]), .bnl_op(lft_op_31_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[335:312]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_30_33[3:0]), .glb_netwk(glb_net_30[7:0]),
     .hold(hold_t_r), .fabric_out(net1253), .sp4_v_t(net1107[0:15]),
     .sp4_v_b(net1072[0:15]));
io_col4_TOP I_IO_29_33 ( .ceb(ceb_o), .bl({bl_29[5], bl_29[4],
     bl_29[37], bl_29[36], bl_29[35], bl_29[34], bl_29[33], bl_29[32],
     bl_29[14], bl_29[20], bl_29[19], bl_29[18], bl_29[17], bl_29[16],
     bl_29[27], bl_29[26], bl_29[25], bl_29[23]}), .sdo(net726),
     .sdi(net1076), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[29]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[55:54]), .pado(pado_t[55:54]),
     .padeb(padeb_t[55:54]), .sp4_h_l(sp4_v_b_29_33[47:0]),
     .sp12_h_l(sp12_v_b_29_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1246[0:1]), .tnl_op(lft_op_28_33[7:0]),
     .lft_op(lft_op_29_33[7:0]), .bnl_op(lft_op_30_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[311:288]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_29_33[3:0]), .glb_netwk(glb_net_29[7:0]),
     .hold(hold_t_r), .fabric_out(net1258), .sp4_v_t(net757[0:15]),
     .sp4_v_b(net1107[0:15]));
io_col4_TOP I_IO_31_33 ( .ceb(ceb_o), .bl({bl_31[5], bl_31[4],
     bl_31[37], bl_31[36], bl_31[35], bl_31[34], bl_31[33], bl_31[32],
     bl_31[14], bl_31[20], bl_31[19], bl_31[18], bl_31[17], bl_31[16],
     bl_31[27], bl_31[26], bl_31[25], bl_31[23]}), .sdo(net1041),
     .sdi(net1111), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[31]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[59:58]), .pado(pado_t[59:58]),
     .padeb(padeb_t[59:58]), .sp4_h_l(sp4_v_b_31_33[47:0]),
     .sp12_h_l(sp12_v_b_31_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1128[0:1]), .tnl_op(lft_op_30_33[7:0]),
     .lft_op(lft_op_31_33[7:0]), .bnl_op(lft_op_32_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[359:336]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_31_33[3:0]), .glb_netwk(glb_net_31[7:0]),
     .hold(hold_t_r), .fabric_out(net1140), .sp4_v_t(net1072[0:15]),
     .sp4_v_b(net1142[0:15]));
io_col4_TOP I_IO_20_33 ( .ceb(ceb_o), .bl({bl_20[5], bl_20[4],
     bl_20[37], bl_20[36], bl_20[35], bl_20[34], bl_20[33], bl_20[32],
     bl_20[14], bl_20[20], bl_20[19], bl_20[18], bl_20[17], bl_20[16],
     bl_20[27], bl_20[26], bl_20[25], bl_20[23]}), .sdo(net1006),
     .sdi(net1146), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[20]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[37:36]), .pado(pado_t[37:36]),
     .padeb(padeb_t[37:36]), .sp4_h_l(sp4_v_b_20_33[47:0]),
     .sp12_h_l(sp12_v_b_20_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1163[0:1]), .tnl_op(lft_op_19_33[7:0]),
     .lft_op(lft_op_20_33[7:0]), .bnl_op(lft_op_21_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[95:72]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_20_33[3:0]), .glb_netwk(glb_net_20[7:0]),
     .hold(hold_t_r), .fabric_out(net1175), .sp4_v_t(net1037[0:15]),
     .sp4_v_b(net1177[0:15]));
io_col4_TOP I_IO_26_33 ( .ceb(ceb_o), .bl({bl_26[5], bl_26[4],
     bl_26[37], bl_26[36], bl_26[35], bl_26[34], bl_26[33], bl_26[32],
     bl_26[14], bl_26[20], bl_26[19], bl_26[18], bl_26[17], bl_26[16],
     bl_26[27], bl_26[26], bl_26[25], bl_26[23]}), .sdo(net656),
     .sdi(net1181), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_r[26]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t[49:48]), .pado(pado_t[49:48]),
     .padeb(padeb_t[49:48]), .sp4_h_l(sp4_v_b_26_33[47:0]),
     .sp12_h_l(sp12_v_b_26_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1198[0:1]), .tnl_op(lft_op_25_33[7:0]),
     .lft_op(lft_op_26_33[7:0]), .bnl_op(lft_op_27_33[7:0]),
     .pgate(pgate_r[15:0]), .reset(reset_r[15:0]), .wl(wl_r[15:0]),
     .cf(cf_t[239:216]), .vdd_cntl(vdd_cntl_r[15:0]),
     .slf_op(slf_op_26_33[3:0]), .glb_netwk(glb_net_26[7:0]),
     .hold(hold_t_r), .fabric_out(net1210), .sp4_v_t(net687[0:15]),
     .sp4_v_b(net1212[0:15]));
bram_bufferx4 I340 ( .in(ceb_i), .out(ceb_o));
bram_bufferx4 I1079 ( .in(bs_en_i), .out(bs_en_o));
bram_bufferx4 I1082 ( .in(update_i), .out(update_o));
bram_bufferx4 I1076 ( .in(mode_i), .out(mode_o));
bram_bufferx4 I1078 ( .in(shift_i), .out(shift_o));
bram_bufferx4 I1080 ( .in(r_i), .out(r_o));
bram_bufferx4 I1081 ( .in(hiz_b_i), .out(hiz_b_o));

endmodule
// Library - leafcell, Cell - quad_tr_ice8, View - schematic
// LAST TIME SAVED: Sep 18 15:38:25 2008
// NETLIST TIME: Nov 14 16:17:19 2008
`timescale 1ns / 1ns 

module quad_tr_ice8 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, ceb_o, cf_r, cf_t, fabric_out_17_33,
     fabric_out_33_17, fabric_out_33_18, hiz_b_o, mode_o, padeb_r,
     padeb_t, padin_136, padin_192, pado_r, pado_t, r_o, sdo, shift_o,
     slf_op_17_17, slf_op_17_18, slf_op_17_19, slf_op_17_20,
     slf_op_17_21, slf_op_17_22, slf_op_17_23, slf_op_17_24,
     slf_op_17_25, slf_op_17_26, slf_op_17_27, slf_op_17_28,
     slf_op_17_29, slf_op_17_30, slf_op_17_31, slf_op_17_32,
     slf_op_17_33, slf_op_18_17, slf_op_19_17, slf_op_20_17,
     slf_op_21_17, slf_op_22_17, slf_op_23_17, slf_op_24_17,
     slf_op_25_17, slf_op_26_17, slf_op_27_17, slf_op_28_17,
     slf_op_29_17, slf_op_30_17, slf_op_31_17, slf_op_32_17,
     slf_op_33_17, spi_ss_in_b_r, tclk_o, update_o, bl, pgate_r,
     reset_r, sp4_h_l_17_17, sp4_h_l_17_18, sp4_h_l_17_19,
     sp4_h_l_17_20, sp4_h_l_17_21, sp4_h_l_17_22, sp4_h_l_17_23,
     sp4_h_l_17_24, sp4_h_l_17_25, sp4_h_l_17_26, sp4_h_l_17_27,
     sp4_h_l_17_28, sp4_h_l_17_29, sp4_h_l_17_30, sp4_h_l_17_31,
     sp4_h_l_17_32, sp4_h_l_17_33, sp4_v_b_17_17, sp4_v_b_17_18,
     sp4_v_b_17_19, sp4_v_b_17_20, sp4_v_b_17_21, sp4_v_b_17_22,
     sp4_v_b_17_23, sp4_v_b_17_24, sp4_v_b_17_25, sp4_v_b_17_26,
     sp4_v_b_17_27, sp4_v_b_17_28, sp4_v_b_17_29, sp4_v_b_17_30,
     sp4_v_b_17_31, sp4_v_b_17_32, sp4_v_b_18_17, sp4_v_b_19_17,
     sp4_v_b_20_17, sp4_v_b_21_17, sp4_v_b_22_17, sp4_v_b_23_17,
     sp4_v_b_24_17, sp4_v_b_25_17, sp4_v_b_26_17, sp4_v_b_27_17,
     sp4_v_b_28_17, sp4_v_b_29_17, sp4_v_b_30_17, sp4_v_b_31_17,
     sp4_v_b_32_17, sp4_v_b_33_17, sp12_h_l_17_17, sp12_h_l_17_18,
     sp12_h_l_17_19, sp12_h_l_17_20, sp12_h_l_17_21, sp12_h_l_17_22,
     sp12_h_l_17_23, sp12_h_l_17_24, sp12_h_l_17_25, sp12_h_l_17_26,
     sp12_h_l_17_27, sp12_h_l_17_28, sp12_h_l_17_29, sp12_h_l_17_30,
     sp12_h_l_17_31, sp12_h_l_17_32, sp12_v_b_17_17, sp12_v_b_18_17,
     sp12_v_b_19_17, sp12_v_b_20_17, sp12_v_b_21_17, sp12_v_b_22_17,
     sp12_v_b_23_17, sp12_v_b_24_17, sp12_v_b_25_17, sp12_v_b_26_17,
     sp12_v_b_27_17, sp12_v_b_28_17, sp12_v_b_29_17, sp12_v_b_30_17,
     sp12_v_b_31_17, sp12_v_b_32_17, vdd_cntl_r, wl_r, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_17_17,
     bnl_op_18_17, bnl_op_19_17, bnl_op_20_17, bnl_op_21_17,
     bnl_op_22_17, bnl_op_23_17, bnl_op_24_17, bnl_op_25_17,
     bnl_op_26_17, bnl_op_27_17, bnl_op_28_17, bnl_op_29_17,
     bnl_op_30_17, bnl_op_31_17, bnl_op_32_17, bnl_op_33_17,
     bnr_op_17_17, bnr_op_18_17, bnr_op_19_17, bnr_op_20_17,
     bnr_op_21_17, bnr_op_22_17, bnr_op_23_17, bnr_op_24_17,
     bnr_op_25_17, bnr_op_26_17, bnr_op_27_17, bnr_op_28_17,
     bnr_op_29_17, bnr_op_30_17, bnr_op_31_17, bnr_op_32_17,
     bot_op_17_17, bot_op_18_17, bot_op_19_17, bot_op_20_17,
     bot_op_21_17, bot_op_22_17, bot_op_23_17, bot_op_24_17,
     bot_op_25_17, bot_op_26_17, bot_op_27_17, bot_op_28_17,
     bot_op_29_17, bot_op_30_17, bot_op_31_17, bot_op_32_17, bs_en_i,
     carry_in_17_17, carry_in_18_17, carry_in_19_17, carry_in_20_17,
     carry_in_21_17, carry_in_22_17, carry_in_23_17, carry_in_24_17,
     carry_in_26_17, carry_in_27_17, carry_in_28_17, carry_in_29_17,
     carry_in_30_17, carry_in_31_17, carry_in_32_17, ceb_i,
     end_of_startup_lft_b, end_of_startup_top_r, glb_in, hiz_b_i,
     hold_r_t, hold_t_r, lft_op_17_17, lft_op_17_18, lft_op_17_19,
     lft_op_17_20, lft_op_17_21, lft_op_17_22, lft_op_17_23,
     lft_op_17_24, lft_op_17_25, lft_op_17_26, lft_op_17_27,
     lft_op_17_28, lft_op_17_29, lft_op_17_30, lft_op_17_31,
     lft_op_17_32, mode_i, padin_r, padin_t, prog, purst, r_i, sdi,
     shift_i, tclk_i, tiegnd, tievdd, tnl_op_17_32, update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bs_en_o, ceb_o,
     fabric_out_17_33, fabric_out_33_17, fabric_out_33_18, hiz_b_o,
     mode_o, padin_136, padin_192, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en_i,
     carry_in_17_17, carry_in_18_17, carry_in_19_17, carry_in_20_17,
     carry_in_21_17, carry_in_22_17, carry_in_23_17, carry_in_24_17,
     carry_in_26_17, carry_in_27_17, carry_in_28_17, carry_in_29_17,
     carry_in_30_17, carry_in_31_17, carry_in_32_17, ceb_i, hiz_b_i,
     hold_r_t, hold_t_r, mode_i, prog, purst, r_i, sdi, shift_i,
     tclk_i, tiegnd, tievdd, update_i;

output [7:0]  slf_op_17_26;
output [7:0]  slf_op_24_17;
output [7:0]  slf_op_20_17;
output [7:0]  slf_op_17_28;
output [7:0]  slf_op_17_29;
output [54:28]  padeb_r;
output [7:0]  slf_op_26_17;
output [383:0]  cf_t;
output [7:0]  slf_op_21_17;
output [7:0]  slf_op_17_18;
output [7:0]  slf_op_17_19;
output [7:0]  slf_op_17_25;
output [7:0]  slf_op_30_17;
output [7:0]  slf_op_17_20;
output [7:0]  slf_op_27_17;
output [7:0]  slf_op_17_23;
output [7:0]  slf_op_19_17;
output [59:30]  pado_t;
output [7:0]  slf_op_31_17;
output [59:30]  padeb_t;
output [7:0]  slf_op_17_22;
output [383:0]  cf_r;
output [7:0]  slf_op_17_30;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_22_17;
output [7:0]  slf_op_17_31;
output [3:0]  slf_op_17_33;
output [3:0]  slf_op_33_17;
output [7:0]  slf_op_25_17;
output [7:0]  slf_op_18_17;
output [7:0]  slf_op_29_17;
output [7:0]  slf_op_17_24;
output [7:0]  slf_op_17_17;
output [63:32]  spi_ss_in_b_r;
output [7:0]  slf_op_17_27;
output [7:0]  slf_op_32_17;
output [7:0]  slf_op_28_17;
output [7:0]  slf_op_23_17;
output [54:28]  pado_r;
output [7:0]  slf_op_17_32;
output [7:0]  slf_op_17_21;

inout [47:0]  sp4_h_l_17_25;
inout [47:0]  sp4_v_b_18_17;
inout [23:0]  sp12_h_l_17_18;
inout [23:0]  sp12_h_l_17_30;
inout [23:0]  sp12_v_b_32_17;
inout [23:0]  sp12_v_b_22_17;
inout [23:0]  sp12_v_b_27_17;
inout [47:0]  sp4_v_b_17_21;
inout [47:0]  sp4_v_b_17_23;
inout [47:0]  sp4_h_l_17_27;
inout [23:0]  sp12_v_b_26_17;
inout [47:0]  sp4_v_b_32_17;
inout [47:0]  sp4_v_b_17_30;
inout [47:0]  sp4_v_b_20_17;
inout [47:0]  sp4_v_b_17_32;
inout [23:0]  sp12_h_l_17_28;
inout [15:0]  sp4_v_b_33_17;
inout [47:0]  sp4_h_l_17_19;
inout [47:0]  sp4_v_b_19_17;
inout [47:0]  sp4_h_l_17_24;
inout [47:0]  sp4_h_l_17_22;
inout [47:0]  sp4_v_b_28_17;
inout [47:0]  sp4_v_b_24_17;
inout [23:0]  sp12_v_b_23_17;
inout [23:0]  sp12_h_l_17_27;
inout [23:0]  sp12_h_l_17_21;
inout [23:0]  sp12_h_l_17_23;
inout [23:0]  sp12_h_l_17_29;
inout [23:0]  sp12_v_b_28_17;
inout [23:0]  sp12_h_l_17_20;
inout [47:0]  sp4_v_b_17_29;
inout [47:0]  sp4_h_l_17_20;
inout [23:0]  sp12_v_b_29_17;
inout [23:0]  sp12_v_b_30_17;
inout [47:0]  sp4_v_b_17_25;
inout [47:0]  sp4_v_b_17_20;
inout [23:0]  sp12_h_l_17_31;
inout [47:0]  sp4_v_b_17_26;
inout [23:0]  sp12_h_l_17_32;
inout [47:0]  sp4_v_b_17_17;
inout [23:0]  sp12_v_b_19_17;
inout [47:0]  sp4_v_b_29_17;
inout [47:0]  sp4_h_l_17_21;
inout [23:0]  sp12_v_b_17_17;
inout [23:0]  sp12_h_l_17_24;
inout [23:0]  sp12_v_b_31_17;
inout [47:0]  sp4_h_l_17_28;
inout [47:0]  sp4_v_b_21_17;
inout [23:0]  sp12_h_l_17_25;
inout [47:0]  sp4_h_l_17_30;
inout [47:0]  sp4_v_b_23_17;
inout [23:0]  sp12_h_l_17_26;
inout [47:0]  sp4_h_l_17_26;
inout [47:0]  sp4_v_b_17_24;
inout [47:0]  sp4_h_l_17_23;
inout [47:0]  sp4_h_l_17_32;
inout [1743:874]  bl;
inout [271:0]  pgate_r;
inout [271:0]  wl_r;
inout [47:0]  sp4_v_b_25_17;
inout [47:0]  sp4_v_b_31_17;
inout [47:0]  sp4_h_l_17_17;
inout [47:0]  sp4_v_b_26_17;
inout [47:0]  sp4_v_b_17_31;
inout [23:0]  sp12_v_b_25_17;
inout [23:0]  sp12_h_l_17_17;
inout [47:0]  sp4_v_b_27_17;
inout [23:0]  sp12_h_l_17_22;
inout [23:0]  sp12_v_b_20_17;
inout [271:0]  vdd_cntl_r;
inout [271:0]  reset_r;
inout [47:0]  sp4_h_l_17_18;
inout [47:0]  sp4_v_b_17_19;
inout [23:0]  sp12_v_b_24_17;
inout [47:0]  sp4_v_b_17_27;
inout [47:0]  sp4_v_b_30_17;
inout [47:0]  sp4_v_b_22_17;
inout [47:0]  sp4_h_l_17_29;
inout [47:0]  sp4_v_b_17_22;
inout [47:0]  sp4_h_l_17_31;
inout [23:0]  sp12_v_b_21_17;
inout [15:0]  sp4_h_l_17_33;
inout [47:0]  sp4_v_b_17_28;
inout [23:0]  sp12_v_b_18_17;
inout [23:0]  sp12_h_l_17_19;
inout [47:0]  sp4_v_b_17_18;

input [7:0]  bnl_op_25_17;
input [7:0]  lft_op_17_19;
input [7:0]  lft_op_17_22;
input [7:0]  bnl_op_17_17;
input [7:0]  bnr_op_21_17;
input [7:0]  bot_op_28_17;
input [7:0]  bnr_op_28_17;
input [7:0]  bnr_op_17_17;
input [7:0]  bnr_op_20_17;
input [7:0]  bnr_op_23_17;
input [7:0]  bnl_op_22_17;
input [7:0]  lft_op_17_32;
input [7:0]  lft_op_17_18;
input [7:0]  bnl_op_18_17;
input [7:0]  bot_op_21_17;
input [7:0]  bnl_op_23_17;
input [7:0]  lft_op_17_26;
input [7:0]  bnr_op_29_17;
input [7:0]  lft_op_17_29;
input [7:0]  bot_op_19_17;
input [7:0]  bot_op_32_17;
input [7:0]  bot_op_29_17;
input [7:0]  lft_op_17_31;
input [7:0]  lft_op_17_20;
input [7:0]  bot_op_31_17;
input [7:0]  bot_op_27_17;
input [7:0]  bnl_op_24_17;
input [7:0]  bot_op_25_17;
input [16:1]  end_of_startup_lft_b;
input [7:0]  bnr_op_31_17;
input [7:0]  bnl_op_33_17;
input [7:0]  bnl_op_21_17;
input [7:0]  bnr_op_26_17;
input [7:0]  lft_op_17_28;
input [7:0]  bnr_op_24_17;
input [7:0]  lft_op_17_25;
input [7:0]  bot_op_20_17;
input [7:0]  bnr_op_30_17;
input [7:0]  bnl_op_28_17;
input [7:0]  bot_op_22_17;
input [7:0]  lft_op_17_27;
input [7:0]  bnl_op_29_17;
input [7:0]  bot_op_18_17;
input [7:0]  bnr_op_32_17;
input [7:0]  bnr_op_19_17;
input [7:0]  glb_in;
input [7:0]  lft_op_17_21;
input [7:0]  lft_op_17_17;
input [59:30]  padin_t;
input [7:0]  lft_op_17_30;
input [7:0]  bot_op_26_17;
input [7:0]  bot_op_24_17;
input [7:0]  bnl_op_32_17;
input [3:0]  tnl_op_17_32;
input [7:0]  lft_op_17_24;
input [7:0]  bnl_op_30_17;
input [7:0]  bm_sa_i;
input [7:0]  lft_op_17_23;
input [7:0]  bnr_op_18_17;
input [7:0]  bnr_op_25_17;
input [7:0]  bot_op_23_17;
input [7:0]  bnl_op_20_17;
input [7:0]  bnr_op_27_17;
input [54:28]  padin_r;
input [7:0]  bnl_op_26_17;
input [7:0]  bnl_op_31_17;
input [7:0]  bnl_op_19_17;
input [7:0]  bot_op_17_17;
input [7:0]  bnl_op_27_17;
input [7:0]  bot_op_30_17;
input [7:0]  bnr_op_22_17;
input [32:17]  end_of_startup_top_r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:7]  net3935;

wire  [0:23]  net3194;

wire  [0:47]  net2443;

wire  [0:47]  net3755;

wire  [0:47]  net4465;

wire  [0:47]  net3591;

wire  [0:47]  net2658;

wire  [0:23]  net2902;

wire  [0:47]  net4795;

wire  [0:23]  net3686;

wire  [0:23]  net4508;

wire  [0:47]  net3734;

wire  [0:7]  net2621;

wire  [0:7]  net2327;

wire  [0:47]  net2909;

wire  [0:23]  net3396;

wire  [0:7]  net4425;

wire  [0:23]  net3124;

wire  [0:7]  net2787;

wire  [0:23]  net3230;

wire  [0:47]  net3594;

wire  [0:47]  net4794;

wire  [0:47]  net4467;

wire  [0:47]  net4662;

wire  [0:47]  net3956;

wire  [0:47]  net2422;

wire  [0:7]  net2784;

wire  [0:23]  net2539;

wire  [0:23]  net2475;

wire  [0:7]  net3499;

wire  [0:23]  net4682;

wire  [0:7]  net2847;

wire  [0:7]  net4812;

wire  [0:47]  net3564;

wire  [0:23]  net2574;

wire  [0:47]  net2494;

wire  [0:47]  net3898;

wire  [0:47]  net4170;

wire  [0:7]  net4025;

wire  [0:47]  net2235;

wire  [0:23]  net3359;

wire  [0:7]  net3207;

wire  [0:47]  net3631;

wire  [0:7]  net3045;

wire  [0:7]  net4815;

wire  [0:47]  net3074;

wire  [0:47]  net4085;

wire  [0:7]  net4319;

wire  [0:47]  net2745;

wire  [0:47]  net2346;

wire  [0:7]  net3369;

wire  [0:47]  net2351;

wire  [0:7]  net3211;

wire  [0:23]  net4436;

wire  [0:7]  net3666;

wire  [0:47]  net2444;

wire  [0:47]  net2776;

wire  [0:47]  net4495;

wire  [0:23]  net4344;

wire  [0:47]  net2936;

wire  [0:23]  net4836;

wire  [0:47]  net2809;

wire  [0:23]  net4706;

wire  [0:47]  net3757;

wire  [0:47]  net3475;

wire  [0:47]  net4335;

wire  [0:7]  net2359;

wire  [0:47]  net4167;

wire  [0:23]  net4445;

wire  [0:7]  net2713;

wire  [0:7]  net4193;

wire  [0:7]  net3772;

wire  [0:23]  net3953;

wire  [0:23]  net2878;

wire  [0:47]  net4385;

wire  [0:7]  net3994;

wire  [0:23]  net4049;

wire  [0:47]  net3314;

wire  [0:23]  net4115;

wire  [0:7]  net3932;

wire  [0:47]  net3478;

wire  [0:23]  net3031;

wire  [0:47]  net4791;

wire  [0:47]  net3971;

wire  [0:47]  net4411;

wire  [0:47]  net2751;

wire  [0:47]  net3140;

wire  [0:23]  net3133;

wire  [0:47]  net3182;

wire  [0:47]  net2912;

wire  [0:23]  net3131;

wire  [0:47]  net2610;

wire  [0:47]  net3629;

wire  [0:47]  net2240;

wire  [0:7]  net2389;

wire  [0:23]  net4543;

wire  [0:47]  net2823;

wire  [0:7]  net4357;

wire  [0:47]  net4744;

wire  [0:47]  net2349;

wire  [0:47]  net2244;

wire  [0:47]  net3510;

wire  [0:23]  net3197;

wire  [0:47]  net3842;

wire  [0:47]  net3674;

wire  [0:47]  net4168;

wire  [0:47]  net2750;

wire  [0:47]  net3955;

wire  [0:47]  net2690;

wire  [0:7]  net3114;

wire  [0:7]  net3219;

wire  [0:47]  net2229;

wire  [0:47]  net2987;

wire  [0:47]  net3264;

wire  [0:47]  net3839;

wire  [0:7]  net3711;

wire  [0:47]  net3022;

wire  [0:7]  net4191;

wire  [0:47]  net4628;

wire  [0:7]  net2844;

wire  [0:47]  net3020;

wire  [0:23]  net4705;

wire  [0:47]  net3809;

wire  [0:47]  net2495;

wire  [0:47]  net3268;

wire  [0:47]  net3566;

wire  [0:47]  net4659;

wire  [0:23]  net4019;

wire  [0:47]  net2824;

wire  [0:47]  net2855;

wire  [0:47]  net4224;

wire  [0:47]  net2484;

wire  [0:23]  net2386;

wire  [0:23]  net3132;

wire  [0:7]  net4752;

wire  [0:47]  net4494;

wire  [0:47]  net3628;

wire  [0:23]  net3363;

wire  [0:47]  net3184;

wire  [0:47]  net2243;

wire  [0:47]  net3104;

wire  [3:0]  slf_op_32_33;

wire  [0:23]  net3952;

wire  [0:47]  net4332;

wire  [0:47]  net3632;

wire  [0:7]  net3828;

wire  [0:47]  net2986;

wire  [3:0]  slf_op_30_33;

wire  [0:23]  net3130;

wire  [0:47]  net2242;

wire  [3:0]  slf_op_24_33;

wire  [3:0]  slf_op_26_33;

wire  [3:0]  slf_op_27_33;

wire  [3:0]  slf_op_28_33;

wire  [3:0]  slf_op_33_24;

wire  [3:0]  slf_op_33_21;

wire  [3:0]  slf_op_23_33;

wire  [3:0]  slf_op_31_33;

wire  [3:0]  slf_op_22_33;

wire  [3:0]  slf_op_18_33;

wire  [3:0]  slf_op_19_33;

wire  [3:0]  slf_op_33_25;

wire  [3:0]  slf_op_21_33;

wire  [3:0]  slf_op_29_33;

wire  [3:0]  slf_op_33_22;

wire  [3:0]  slf_op_20_33;

wire  [3:0]  slf_op_25_00;

wire  [3:0]  slf_op_33_27;

wire  [3:0]  slf_op_33_32;

wire  [3:0]  slf_op_33_26;

wire  [3:0]  slf_op_33_31;

wire  [3:0]  slf_op_33_19;

wire  [3:0]  slf_op_33_18;

wire  [3:0]  slf_op_33_28;

wire  [3:0]  slf_op_33_30;

wire  [3:0]  slf_op_33_23;

wire  [3:0]  slf_op_33_20;

wire  [3:0]  slf_op_33_29;

wire  [0:7]  net4517;

wire  [7:0]  clk_tree_drv;

wire  [0:23]  net2904;

wire  [0:23]  net3691;

wire  [0:7]  net2456;

wire  [0:47]  net4627;

wire  [0:47]  net3728;

wire  [0:7]  net4264;

wire  [0:47]  net3267;

wire  [0:23]  net4213;

wire  [0:47]  net2350;

wire  [0:7]  net3767;

wire  [0:7]  net3174;

wire  [0:23]  net3457;

wire  [0:47]  net3406;

wire  [0:23]  net3395;

wire  [0:23]  net3853;

wire  [0:47]  net3676;

wire  [0:23]  net3525;

wire  [0:47]  net4631;

wire  [0:7]  net4484;

wire  [0:23]  net2411;

wire  [0:23]  net3788;

wire  [0:7]  net2622;

wire  [0:23]  net2477;

wire  [0:7]  net3827;

wire  [0:47]  net2479;

wire  [0:47]  net3974;

wire  [0:47]  net2587;

wire  [0:23]  net2640;

wire  [0:47]  net2938;

wire  [0:47]  net3183;

wire  [0:23]  net2542;

wire  [0:23]  net4600;

wire  [0:7]  net4751;

wire  [0:47]  net3318;

wire  [0:47]  net3404;

wire  [0:7]  net3991;

wire  [0:47]  net3646;

wire  [0:47]  net4555;

wire  [0:15]  net4847;

wire  [0:23]  net2576;

wire  [0:47]  net3970;

wire  [0:7]  net2719;

wire  [0:47]  net2446;

wire  [0:47]  net4384;

wire  [0:7]  net2328;

wire  [0:47]  net3759;

wire  [0:7]  net2518;

wire  [0:47]  net2911;

wire  [0:47]  net3795;

wire  [0:47]  net4499;

wire  [0:7]  net4321;

wire  [0:47]  net4287;

wire  [0:47]  net3185;

wire  [0:7]  net3173;

wire  [0:47]  net4123;

wire  [0:7]  net3439;

wire  [0:47]  net3465;

wire  [0:7]  net2332;

wire  [0:7]  net4590;

wire  [0:47]  net4718;

wire  [0:7]  net3703;

wire  [0:47]  net4298;

wire  [0:23]  net4116;

wire  [0:47]  net4449;

wire  [0:7]  net2319;

wire  [0:47]  net4388;

wire  [0:7]  net4427;

wire  [0:23]  net4280;

wire  [0:47]  net2746;

wire  [0:23]  net4018;

wire  [0:7]  net2519;

wire  [0:47]  net4777;

wire  [0:23]  net3944;

wire  [0:23]  net4835;

wire  [0:7]  net4811;

wire  [0:47]  net2807;

wire  [0:47]  net4615;

wire  [0:47]  net4252;

wire  [0:7]  net2517;

wire  [0:47]  net2908;

wire  [0:47]  net4249;

wire  [0:7]  net2681;

wire  [0:47]  net4416;

wire  [0:47]  net2825;

wire  [0:23]  net4272;

wire  [0:47]  net4577;

wire  [0:47]  net4169;

wire  [0:47]  net4062;

wire  [0:47]  net3803;

wire  [0:47]  net3021;

wire  [0:47]  net2694;

wire  [0:23]  net2641;

wire  [0:47]  net2748;

wire  [0:47]  net2339;

wire  [0:23]  net2294;

wire  [0:47]  net2937;

wire  [0:47]  net3735;

wire  [0:23]  net4181;

wire  [0:23]  net3690;

wire  [0:47]  net3794;

wire  [0:47]  net4776;

wire  [0:47]  net3511;

wire  [0:7]  net3375;

wire  [0:23]  net3030;

wire  [0:23]  net3623;

wire  [0:23]  net3885;

wire  [0:7]  net4203;

wire  [0:47]  net3514;

wire  [0:7]  net4485;

wire  [0:7]  net3335;

wire  [0:23]  net4182;

wire  [0:23]  net2707;

wire  [0:47]  net4787;

wire  [0:23]  net3066;

wire  [0:7]  net3337;

wire  [0:23]  net2637;

wire  [0:23]  net4108;

wire  [0:23]  net4378;

wire  [0:47]  net2811;

wire  [0:47]  net2659;

wire  [0:23]  net4608;

wire  [0:23]  net3557;

wire  [0:47]  net3919;

wire  [0:47]  net2238;

wire  [0:23]  net2358;

wire  [0:7]  net3699;

wire  [0:47]  net3644;

wire  [0:23]  net3458;

wire  [0:7]  net3608;

wire  [0:47]  net4719;

wire  [0:47]  net2245;

wire  [0:23]  net4379;

wire  [0:23]  net3951;

wire  [0:23]  net2296;

wire  [0:47]  net3569;

wire  [0:47]  net4578;

wire  [0:47]  net3079;

wire  [0:23]  net4541;

wire  [0:47]  net2344;

wire  [0:47]  net4121;

wire  [0:47]  net3808;

wire  [0:23]  net4216;

wire  [0:7]  net4756;

wire  [0:47]  net2655;

wire  [0:47]  net2527;

wire  [0:23]  net3622;

wire  [0:47]  net2644;

wire  [0:7]  net2515;

wire  [0:23]  net4606;

wire  [0:23]  net3358;

wire  [0:47]  net3467;

wire  [0:47]  net3923;

wire  [0:23]  net4113;

wire  [0:7]  net3539;

wire  [0:47]  net3187;

wire  [0:23]  net2805;

wire  [0:47]  net2826;

wire  [0:47]  net3242;

wire  [0:23]  net3689;

wire  [0:23]  net2702;

wire  [0:47]  net2749;

wire  [0:47]  net3136;

wire  [0:7]  net4483;

wire  [0:7]  net4591;

wire  [0:23]  net3722;

wire  [0:23]  net3461;

wire  [0:23]  net2801;

wire  [0:47]  net4496;

wire  [0:7]  net4323;

wire  [0:47]  net3479;

wire  [0:7]  net3209;

wire  [0:23]  net2287;

wire  [0:47]  net4124;

wire  [0:47]  net2423;

wire  [0:23]  net3035;

wire  [0:47]  net3645;

wire  [0:47]  net3350;

wire  [0:7]  net2455;

wire  [0:47]  net4248;

wire  [0:47]  net2771;

wire  [0:47]  net2345;

wire  [0:47]  net2973;

wire  [0:7]  net4521;

wire  [0:7]  net3444;

wire  [0:47]  net4251;

wire  [0:7]  net4259;

wire  [0:47]  net4086;

wire  [0:7]  net4095;

wire  [0:23]  net2282;

wire  [0:23]  net3526;

wire  [0:7]  net4587;

wire  [0:47]  net4823;

wire  [0:47]  net3959;

wire  [0:47]  net3147;

wire  [0:7]  net3665;

wire  [0:47]  net3103;

wire  [0:7]  net3336;

wire  [0:23]  net3862;

wire  [0:23]  net2639;

wire  [0:7]  net4650;

wire  [0:7]  net3697;

wire  [0:47]  net2607;

wire  [0:7]  net3442;

wire  [0:7]  net2323;

wire  [0:47]  net4661;

wire  [0:47]  net3482;

wire  [0:23]  net4342;

wire  [0:7]  net2330;

wire  [0:7]  net3606;

wire  [0:23]  net3360;

wire  [0:7]  net4263;

wire  [0:47]  net3894;

wire  [0:7]  net4359;

wire  [0:47]  net3427;

wire  [0:7]  net2715;

wire  [0:47]  net3240;

wire  [0:7]  net4097;

wire  [0:23]  net3780;

wire  [0:23]  net3787;

wire  [0:7]  net4031;

wire  [0:7]  net3995;

wire  [0:23]  net4609;

wire  [0:23]  net3032;

wire  [0:7]  net3771;

wire  [0:23]  net4670;

wire  [0:47]  net2608;

wire  [0:23]  net2412;

wire  [0:7]  net3113;

wire  [0:47]  net3019;

wire  [0:7]  net3829;

wire  [0:7]  net2321;

wire  [0:47]  net4497;

wire  [0:23]  net3687;

wire  [0:23]  net3231;

wire  [0:47]  net3302;

wire  [0:7]  net4158;

wire  [0:23]  net4607;

wire  [0:47]  net2241;

wire  [0:7]  net3861;

wire  [0:47]  net4448;

wire  [0:7]  net4027;

wire  [0:47]  net3304;

wire  [0:47]  net4061;

wire  [0:47]  net2935;

wire  [0:47]  net2974;

wire  [0:23]  net3852;

wire  [0:23]  net3855;

wire  [0:47]  net4247;

wire  [0:23]  net3293;

wire  [0:7]  net4195;

wire  [0:23]  net4673;

wire  [0:47]  net2693;

wire  [0:47]  net4775;

wire  [0:47]  net3571;

wire  [0:7]  net3931;

wire  [0:7]  net4261;

wire  [0:47]  net4134;

wire  [0:47]  net2612;

wire  [0:47]  net4413;

wire  [0:47]  net4793;

wire  [0:7]  net4647;

wire  [0:47]  net3896;

wire  [0:7]  net2785;

wire  [0:7]  net4523;

wire  [0:47]  net3972;

wire  [0:47]  net2646;

wire  [0:23]  net3789;

wire  [0:23]  net2543;

wire  [0:47]  net4613;

wire  [0:23]  net2473;

wire  [0:47]  net2971;

wire  [0:47]  net3101;

wire  [0:47]  net2582;

wire  [0:47]  net4227;

wire  [0:47]  net4122;

wire  [0:7]  net3440;

wire  [0:47]  net4088;

wire  [0:47]  net2581;

wire  [0:23]  net3522;

wire  [0:7]  net2845;

wire  [0:47]  net3920;

wire  [0:23]  net2869;

wire  [0:47]  net4004;

wire  [0:23]  net3886;

wire  [0:47]  net3402;

wire  [0:23]  net3850;

wire  [0:23]  net4345;

wire  [0:23]  net3232;

wire  [0:7]  net4683;

wire  [0:7]  net3339;

wire  [0:23]  net4509;

wire  [0:23]  net2278;

wire  [0:7]  net2680;

wire  [0:47]  net4391;

wire  [0:47]  net2662;

wire  [0:47]  net3018;

wire  [0:23]  net4178;

wire  [0:23]  net2638;

wire  [0:47]  net3317;

wire  [0:7]  net4755;

wire  [0:7]  net3875;

wire  [0:23]  net3033;

wire  [0:47]  net4663;

wire  [0:47]  net3263;

wire  [0:23]  net4346;

wire  [0:23]  net4026;

wire  [0:23]  net4506;

wire  [0:47]  net3758;

wire  [0:47]  net3806;

wire  [0:23]  net3452;

wire  [0:23]  net2704;

wire  [0:7]  net3537;

wire  [0:47]  net3596;

wire  [0:7]  net4687;

wire  [0:47]  net3840;

wire  [0:23]  net3065;

wire  [0:47]  net4057;

wire  [0:47]  net2348;

wire  [0:7]  net2786;

wire  [0:47]  net2497;

wire  [0:7]  net3865;

wire  [0:23]  net4441;

wire  [0:7]  net2320;

wire  [0:47]  net4284;

wire  [0:47]  net4548;

wire  [0:47]  net2530;

wire  [0:7]  net3607;

wire  [0:7]  net3278;

wire  [0:47]  net4824;

wire  [0:47]  net3841;

wire  [0:7]  net2329;

wire  [0:47]  net4288;

wire  [0:23]  net2632;

wire  [0:7]  net4426;

wire  [0:47]  net4060;

wire  [0:7]  net3867;

wire  [0:23]  net3296;

wire  [0:47]  net4390;

wire  [0:47]  net4451;

wire  [0:23]  net3724;

wire  [0:47]  net2939;

wire  [0:23]  net3206;

wire  [0:47]  net4250;

wire  [0:47]  net3592;

wire  [0:47]  net2773;

wire  [0:7]  net3667;

wire  [0:47]  net4739;

wire  [0:23]  net4117;

wire  [0:47]  net3483;

wire  [0:23]  net2965;

wire  [0:47]  net4450;

wire  [0:47]  net3512;

wire  [0:23]  net3558;

wire  [0:47]  net2343;

wire  [0:47]  net3733;

wire  [0:23]  net3199;

wire  [0:23]  net3393;

wire  [0:47]  net2648;

wire  [0:7]  net4367;

wire  [0:47]  net3678;

wire  [0:23]  net3534;

wire  [0:7]  net3701;

wire  [0:23]  net4052;

wire  [0:47]  net4552;

wire  [0:7]  net2783;

wire  [0:47]  net4063;

wire  [0:23]  net2410;

wire  [0:47]  net4171;

wire  [0:47]  net4825;

wire  [0:7]  net3175;

wire  [0:47]  net4742;

wire  [0:47]  net2692;

wire  [0:7]  net2325;

wire  [0:47]  net2499;

wire  [0:7]  net3503;

wire  [0:47]  net3347;

wire  [0:23]  net2737;

wire  [0:7]  net4423;

wire  [0:47]  net2691;

wire  [0:47]  net3568;

wire  [0:23]  net2474;

wire  [0:47]  net3237;

wire  [0:7]  net2788;

wire  [0:47]  net2416;

wire  [0:7]  net4099;

wire  [0:47]  net3481;

wire  [0:47]  net3630;

wire  [0:47]  net4087;

wire  [0:23]  net2967;

wire  [0:7]  net2324;

wire  [0:7]  net4096;

wire  [0:47]  net3679;

wire  [0:23]  net2550;

wire  [0:7]  net2683;

wire  [0:47]  net3639;

wire  [0:47]  net2775;

wire  [0:23]  net2903;

wire  [0:47]  net3480;

wire  [0:23]  net2297;

wire  [0:47]  net3346;

wire  [0:23]  net4770;

wire  [0:47]  net4716;

wire  [0:23]  net3621;

wire  [0:23]  net2295;

wire  [0:23]  net4015;

wire  [0:7]  net3933;

wire  [0:47]  net2660;

wire  [0:47]  net3464;

wire  [0:47]  net3299;

wire  [0:23]  net2217;

wire  [0:7]  net2717;

wire  [0:47]  net2645;

wire  [0:7]  net3830;

wire  [0:47]  net2237;

wire  [0:47]  net2580;

wire  [0:47]  net3593;

wire  [0:47]  net2418;

wire  [0:47]  net3316;

wire  [0:47]  net4138;

wire  [0:7]  net2204;

wire  [0:47]  net3513;

wire  [0:23]  net4051;

wire  [0:47]  net3300;

wire  [0:47]  net2421;

wire  [0:7]  net2387;

wire  [0:7]  net3171;

wire  [0:47]  net2827;

wire  [0:47]  net4712;

wire  [0:47]  net2354;

wire  [0:7]  net2331;

wire  [0:23]  net4347;

wire  [0:7]  net4685;

wire  [0:23]  net4442;

wire  [0:47]  net3960;

wire  [0:23]  net3721;

wire  [0:47]  net4333;

wire  [0:47]  net3796;

wire  [0:23]  net4190;

wire  [0:47]  net2531;

wire  [0:7]  net4588;

wire  [0:47]  net3677;

wire  [0:47]  net2584;

wire  [0:23]  net3394;

wire  [0:7]  net2727;

wire  [0:47]  net2991;

wire  [0:7]  net2553;

wire  [0:23]  net3361;

wire  [0:7]  net4814;

wire  [0:47]  net3076;

wire  [0:47]  net4447;

wire  [0:7]  net3373;

wire  [0:47]  net4714;

wire  [0:47]  net3405;

wire  [0:47]  net4222;

wire  [0:47]  net2239;

wire  [0:7]  net3992;

wire  [0:23]  net2292;

wire  [0:47]  net3428;

wire  [0:7]  net4157;

wire  [0:47]  net3150;

wire  [0:47]  net2341;

wire  [0:7]  net2563;

wire  [0:47]  net3432;

wire  [0:23]  net3068;

wire  [0:47]  net2913;

wire  [0:7]  net2619;

wire  [0:47]  net4616;

wire  [0:47]  net3515;

wire  [0:47]  net2585;

wire  [0:23]  net3459;

wire  [0:7]  net3371;

wire  [0:7]  net3047;

wire  [0:47]  net3023;

wire  [0:47]  net3154;

wire  [0:47]  net3642;

wire  [0:47]  net3100;

wire  [0:7]  net4651;

wire  [0:23]  net4674;

wire  [0:47]  net3975;

wire  [0:47]  net3349;

wire  [0:23]  net4279;

wire  [0:47]  net2236;

wire  [0:47]  net2812;

wire  [0:7]  net3277;

wire  [0:23]  net3288;

wire  [0:47]  net4295;

wire  [0:47]  net2526;

wire  [0:7]  net4592;

wire  [0:47]  net3899;

wire  [0:23]  net3196;

wire  [0:47]  net2663;

wire  [0:47]  net4137;

wire  [0:23]  net2901;

wire  [0:47]  net4459;

wire  [0:47]  net3401;

wire  [0:7]  net4754;

wire  [0:47]  net3265;

wire  [0:47]  net2822;

wire  [0:7]  net4320;

wire  [0:7]  net2326;

wire  [0:23]  net3297;

wire  [0:7]  net3603;

wire  [0:47]  net3137;

wire  [0:7]  net3501;

wire  [0:47]  net4058;

wire  [0:7]  net4589;

wire  [0:23]  net4014;

wire  [0:7]  net3535;

wire  [0:23]  net4343;

wire  [0:47]  net2774;

wire  [0:47]  net4006;

wire  [0:23]  net2468;

wire  [0:47]  net2975;

wire  [0:47]  net3139;

wire  [0:23]  net4773;

wire  [0:7]  net3172;

wire  [0:47]  net3099;

wire  [0:23]  net4510;

wire  [0:47]  net3241;

wire  [0:23]  net3195;

wire  [0:47]  net4302;

wire  [0:23]  net3198;

wire  [0:23]  net2476;

wire  [0:23]  net2739;

wire  [0:23]  net4114;

wire  [0:23]  net2871;

wire  [0:23]  net2703;

wire  [0:47]  net4135;

wire  [0:23]  net4834;

wire  [0:7]  net2460;

wire  [0:47]  net4005;

wire  [0:47]  net3151;

wire  [0:47]  net3463;

wire  [0:7]  net2623;

wire  [0:7]  net3770;

wire  [0:47]  net3838;

wire  [0:47]  net3791;

wire  [0:47]  net4056;

wire  [0:7]  net4695;

wire  [0:23]  net2740;

wire  [0:23]  net3949;

wire  [0:47]  net4717;

wire  [0:47]  net3430;

wire  [0:7]  net4486;

wire  [0:47]  net2988;

wire  [0:47]  net3243;

wire  [0:47]  net3078;

wire  [0:47]  net4576;

wire  [0:23]  net3295;

wire  [0:47]  net3565;

wire  [0:7]  net2457;

wire  [0:47]  net3643;

wire  [0:23]  net3042;

wire  [0:7]  net4029;

wire  [0:7]  net2391;

wire  [0:47]  net3466;

wire  [0:7]  net4531;

wire  [0:23]  net4354;

wire  [0:47]  net3792;

wire  [0:23]  net2868;

wire  [0:47]  net4790;

wire  [0:47]  net3957;

wire  [0:23]  net4671;

wire  [0:47]  net2808;

wire  [0:23]  net3625;

wire  [0:47]  net2496;

wire  [0:7]  net4681;

wire  [0:7]  net4355;

wire  [0:23]  net4050;

wire  [0:7]  net3115;

wire  [0:47]  net2481;

wire  [0:23]  net3560;

wire  [0:47]  net2695;

wire  [0:47]  net3756;

wire  [0:7]  net2555;

wire  [0:7]  net3116;

wire  [0:47]  net3152;

wire  [0:7]  net4156;

wire  [0:23]  net3888;

wire  [0:47]  net4612;

wire  [0:23]  net4443;

wire  [0:47]  net4221;

wire  [0:23]  net4771;

wire  [0:47]  net4083;

wire  [0:47]  net3810;

wire  [0:47]  net4611;

wire  [0:47]  net4580;

wire  [0:7]  net3769;

wire  [0:47]  net2233;

wire  [0:7]  net3663;

wire  [0:23]  net3616;

wire  [0:47]  net4084;

wire  [0:47]  net4741;

wire  [0:7]  net3863;

wire  [0:47]  net4740;

wire  [0:7]  net3441;

wire  [0:7]  net3768;

wire  [0:23]  net2290;

wire  [0:47]  net3893;

wire  [0:23]  net3786;

wire  [0:47]  net4827;

wire  [0:47]  net2338;

wire  [0:7]  net2620;

wire  [0:47]  net4285;

wire  [0:47]  net4131;

wire  [0:47]  net2858;

wire  [0:47]  net3730;

wire  [0:7]  net2679;

wire  [0:47]  net3153;

wire  [0:23]  net3527;

wire  [0:7]  net2551;

wire  [0:23]  net4837;

wire  [0:23]  net2866;

wire  [0:7]  net4100;

wire  [0:23]  net4707;

wire  [0:47]  net4119;

wire  [0:23]  net2705;

wire  [0:23]  net3559;

wire  [0:47]  net4002;

wire  [0:23]  net2738;

wire  [0:23]  net2277;

wire  [0:47]  net4136;

wire  [0:23]  net3785;

wire  [0:7]  net3280;

wire  [0:23]  net3129;

wire  [0:23]  net4215;

wire  [0:47]  net2491;

wire  [0:47]  net2819;

wire  [0:47]  net4225;

wire  [0:23]  net3851;

wire  [0:7]  net2682;

wire  [0:47]  net2234;

wire  [0:47]  net4466;

wire  [0:23]  net3294;

wire  [0:47]  net3967;

wire  [0:23]  net3067;

wire  [0:47]  net3807;

wire  [0:47]  net4623;

wire  [0:47]  net3892;

wire  [0:47]  net2337;

wire  [0:23]  net4507;

wire  [0:47]  net4822;

wire  [0:47]  net3266;

wire  [0:7]  net2846;

wire  [0:47]  net4452;

wire  [0:47]  net4220;

wire  [0:23]  net3950;

wire  [0:23]  net2804;

wire  [0:47]  net4778;

wire  [0:7]  net2399;

wire  [0:47]  net3627;

wire  [0:7]  net3111;

wire  [0:47]  net2856;

wire  [0:47]  net2529;

wire  [0:47]  net3072;

wire  [0:47]  net2972;

wire  [0:7]  net4353;

wire  [0:47]  net3135;

wire  [0:7]  net3338;

wire  [0:23]  net2575;

wire  [0:47]  net2347;

wire  [0:23]  net4544;

wire  [0:47]  net4300;

wire  [0:47]  net4007;

wire  [0:47]  net2661;

wire  [0:23]  net2803;

wire  [0:23]  net4277;

wire  [0:23]  net2293;

wire  [0:47]  net3431;

wire  [0:47]  net3186;

wire  [0:47]  net4660;

wire  [0:7]  net4428;

wire  [0:7]  net3547;

wire  [0:23]  net2960;

wire  [0:23]  net4708;

wire  [0:47]  net2857;

wire  [0:23]  net3370;

wire  [0:47]  net4626;

wire  [0:47]  net4226;

wire  [0:7]  net3275;

wire  [0:7]  net4753;

wire  [0:23]  net4278;

wire  [0:47]  net2498;

wire  [0:47]  net2447;

wire  [0:47]  net4331;

wire  [0:23]  net4672;

wire  [0:7]  net3604;

wire  [0:47]  net3138;

wire  [0:7]  net4155;

wire  [0:23]  net2796;

wire  [0:47]  net4412;

wire  [0:47]  net3238;

wire  [0:47]  net4743;

wire  [0:7]  net3279;

wire  [0:47]  net4414;

wire  [0:23]  net4281;

wire  [0:47]  net3570;

wire  [0:47]  net4139;

wire  [0:47]  net4826;

wire  [0:23]  net4377;

wire  [0:47]  net4549;

wire  [0:7]  net2843;

wire  [0:7]  net3443;

wire  [0:47]  net2483;

wire  [0:47]  net3468;

wire  [0:47]  net2480;

wire  [0:23]  net4675;

wire  [0:47]  net2647;

wire  [0:47]  net4553;

wire  [0:7]  net2459;

wire  [0:47]  net4003;

wire  [0:47]  net2448;

wire  [0:23]  net4772;

wire  [0:47]  net3429;

wire  [0:47]  net4415;

wire  [0:47]  net4498;

wire  [0:47]  net2643;

wire  [0:47]  net4120;

wire  [0:47]  net2859;

wire  [0:7]  net4159;

wire  [0:23]  net2281;

wire  [0:47]  net2976;

wire  [0:23]  net4542;

wire  [0:47]  net3675;

wire  [0:7]  net3934;

wire  [0:23]  net2289;

wire  [0:7]  net2549;

wire  [0:23]  net2409;

wire  [0:47]  net3351;

wire  [0:23]  net2802;

wire  [0:47]  net2609;

wire  [0:47]  net3843;

wire  [0:47]  net3921;

wire  [0:47]  net4550;

wire  [0:47]  net2983;

wire  [0:23]  net3362;

wire  [0:47]  net4386;

wire  [0:23]  net3887;

wire  [0:47]  net3647;

wire  [0:7]  net2877;

wire  [0:47]  net2989;

wire  [0:7]  net3041;

wire  [0:7]  net3664;

wire  [0:47]  net2342;

wire  [0:7]  net3383;

wire  [0:23]  net2540;

wire  [0:47]  net3922;

wire  [0:47]  net3073;

wire  [0:47]  net2586;

wire  [0:47]  net4330;

wire  [0:47]  net4779;

wire  [0:47]  net3311;

wire  [0:23]  net2966;

wire  [0:47]  net2810;

wire  [0:23]  net4179;

wire  [0:47]  net3897;

wire  [0:23]  net2541;

wire  [0:23]  net4518;

wire  [0:23]  net4183;

wire  [0:47]  net2744;

wire  [0:7]  net4648;

wire  [0:7]  net4039;

wire  [0:47]  net4629;

wire  [0:7]  net4262;

wire  [0:23]  net4380;

wire  [0:23]  net3624;

wire  [0:7]  net3043;

wire  [0:23]  net3698;

wire  [0:47]  net3973;

wire  [0:47]  net2445;

wire  [0:47]  net3407;

wire  [0:47]  net3155;

wire  [0:23]  net4769;

wire  [0:47]  net2482;

wire  [0:23]  net3723;

wire  [0:23]  net4839;

wire  [0:7]  net2458;

wire  [0:47]  net3400;

wire  [0:47]  net4334;

wire  [0:7]  net3502;

wire  [0:47]  net4389;

wire  [0:47]  net4630;

wire  [0:47]  net4301;

wire  [0:7]  net4260;

wire  [0:23]  net3854;

wire  [0:47]  net3595;

wire  [0:47]  net3958;

wire  [0:47]  net2420;

wire  [0:47]  net2611;

wire  [0:47]  net4780;

wire  [0:47]  net3301;

wire  [0:23]  net4016;

wire  [0:7]  net4487;

wire  [0:23]  net4214;

wire  [0:47]  net4303;

wire  [0:23]  net2969;

wire  [0:23]  net3688;

wire  [0:47]  net3732;

wire  [0:47]  net2910;

wire  [0:7]  net4813;

wire  [0:47]  net4713;

wire  [0:47]  net4464;

wire  [0:7]  net4098;

wire  [0:7]  net4322;

wire  [0:47]  net4658;

wire  [0:7]  net2516;

wire  [0:47]  net2940;

wire  [0:23]  net4838;

wire  [0:47]  net2528;

wire  [0:47]  net2854;

wire  [0:47]  net2915;

wire  [0:7]  net4189;

wire  [0:47]  net4575;

wire  [0:7]  net3831;

wire  [0:7]  net3112;

wire  [0:47]  net4166;

wire  [0:23]  net2288;

wire  [0:47]  net3811;

wire  [0:23]  net4511;

wire  [0:47]  net3102;

wire  [0:47]  net4554;

wire  [0:23]  net2968;

wire  [0:47]  net2340;

wire  [0:47]  net4463;

wire  [0:47]  net4299;

wire  [0:7]  net3533;

wire  [0:23]  net3229;

wire  [0:47]  net3793;

wire  [0:23]  net2291;

wire  [0:47]  net4462;

wire  [0:47]  net3315;

wire  [0:47]  net4283;

wire  [0:23]  net2573;

wire  [0:47]  net2990;

wire  [0:47]  net3236;

wire  [0:7]  net3055;

wire  [0:7]  net2385;

wire  [0:7]  net3276;

wire  [0:7]  net3205;

wire  [0:47]  net3729;

wire  [0:47]  net2914;

wire  [0:7]  net4519;

wire  [0:47]  net2246;

wire  [0:47]  net2232;

wire  [0:7]  net4649;

wire  [0:7]  net2322;

wire  [0:47]  net3924;

wire  [0:23]  net3034;

wire  [0:47]  net4614;

wire  [0:7]  net2624;

wire  [0:23]  net2706;

wire  [0:23]  net3524;

wire  [0:47]  net4286;

wire  [0:47]  net4579;

wire  [0:23]  net4444;

wire  [0:23]  net2870;

wire  [0:47]  net3319;

wire  [0:23]  net3460;

wire  [0:23]  net4764;

wire  [0:23]  net3523;

wire  [0:7]  net3605;

wire  [0:23]  net4605;

wire  [0:47]  net3303;

wire  [0:47]  net2417;

wire  [0:23]  net2538;

wire  [0:23]  net2714;

wire  [0:23]  net4180;

wire  [0:23]  net2867;

wire  [0:47]  net3348;

wire  [0:7]  net3500;

wire  [0:47]  net2772;

wire  [0:47]  net3077;

wire  [0:7]  net3936;

wire  [0:47]  net3760;

wire  [0:47]  net4792;

wire  [0:7]  net4424;

wire  [0:7]  net3993;

wire  [0:23]  net4017;



lowla_modified I349 ( .clk(tclk_i), .min(net02082), .lao(net2191));
bram_bufferx4x6 I350 ( .in(sdi), .out(net02082));
tckbufx16 I242 ( .in(tclk_i), .out(net4849));
clk_colbuf8kx8 I_clktree_qdrv_tr ( .clko(clk_tree_drv[7:0]),
     .clki(glb_in[7:0]));
fabric_buf8k I343 ( .f_in(net2101), .f_out(fabric_out_33_18));
fabric_buf8k I344 ( .f_in(net2100), .f_out(fabric_out_33_17));
fabric_buf8k I345 ( .f_in(padin_r[28]), .f_out(padin_136));
array_RGT_IO_1x16top I_io_33top ( .sp4_v_b_00_17(sp4_v_b_33_17[15:0]),
     .sp4_v_t_00_32(net4847[0:15]), .ceb(net4846),
     .padin(padin_r[54:28]), .pado(pado_r[54:28]),
     .padeb(padeb_r[54:28]), .fabric_out_17(net2100),
     .fabric_out_18(net2101), .fabric_out_19(net5001),
     .fabric_out_21(net5002), .fabric_out_20(net2104),
     .fabric_out_25(net4996), .fabric_out_24(net5005),
     .fabric_out_22(net5003), .fabric_out_23(net5004),
     .fabric_out_27(net4999), .fabric_out_26(net4997),
     .fabric_out_28(net5000), .fabric_out_30(net4994),
     .fabric_out_29(net4995), .fabric_out_31(net4993),
     .fabric_out_32(net4992), .lft_op_00_17(slf_op_32_17[7:0]),
     .lft_op_00_18(net3539[0:7]), .lft_op_00_19(net3537[0:7]),
     .lft_op_00_20(net3547[0:7]), .lft_op_00_21(net3608[0:7]),
     .lft_op_00_22(net3607[0:7]), .lft_op_00_23(net3606[0:7]),
     .lft_op_00_24(net3605[0:7]), .lft_op_00_25(net3604[0:7]),
     .lft_op_00_26(net3603[0:7]), .lft_op_00_27(net3667[0:7]),
     .lft_op_00_28(net3665[0:7]), .lft_op_00_29(net3666[0:7]),
     .lft_op_00_30(net3663[0:7]), .lft_op_00_31(net3664[0:7]),
     .lft_op_00_32(net3535[0:7]),
     .cdone_in(end_of_startup_lft_b[16:1]),
     .tnl_op_00_17({slf_op_32_33[3], slf_op_32_33[2], slf_op_32_33[1],
     slf_op_32_33[0], slf_op_32_33[3], slf_op_32_33[2],
     slf_op_32_33[1], slf_op_32_33[0]}), .SP4_h_l_00_26(net2935[0:47]),
     .SP4_h_l_00_23(net2938[0:47]), .slf_op_00_29(slf_op_33_29[3:0]),
     .slf_op_00_28(slf_op_33_28[3:0]),
     .slf_op_00_27(slf_op_33_27[3:0]),
     .slf_op_00_26(slf_op_33_26[3:0]),
     .slf_op_00_25(slf_op_33_25[3:0]),
     .slf_op_00_24(slf_op_33_24[3:0]),
     .slf_op_00_23(slf_op_33_23[3:0]),
     .slf_op_00_22(slf_op_33_22[3:0]), .SP4_h_l_00_25(net2936[0:47]),
     .SP4_h_l_00_24(net2937[0:47]), .slf_op_00_17(slf_op_33_17[3:0]),
     .slf_op_00_18(slf_op_33_18[3:0]),
     .slf_op_00_19(slf_op_33_19[3:0]),
     .slf_op_00_20(slf_op_33_20[3:0]),
     .bnl_op_00_32(bnl_op_33_17[7:0]), .SP4_h_l_00_32(net2991[0:47]),
     .SP4_h_l_00_31(net2990[0:47]), .pgate(pgate_r[255:0]),
     .vdd_cntl(vdd_cntl_r[255:0]), .reset_b(reset_r[255:0]),
     .cf_l(cf_r[383:0]), .SP4_h_l_00_30(net2989[0:47]),
     .SP4_h_l_00_29(net2988[0:47]), .SP4_h_l_00_28(net2987[0:47]),
     .SP4_h_l_00_27(net2986[0:47]), .SP4_h_l_00_17(net2915[0:47]),
     .SP4_h_l_00_18(net2914[0:47]), .SP4_h_l_00_19(net2913[0:47]),
     .SP4_h_l_00_20(net2912[0:47]), .SP4_h_l_00_21(net2940[0:47]),
     .SP4_h_l_00_22(net2939[0:47]), .slf_op_00_31(slf_op_33_31[3:0]),
     .slf_op_00_32(slf_op_33_32[3:0]),
     .slf_op_00_21(slf_op_33_21[3:0]), .SP12_h_l_00_32(net3030[0:23]),
     .SP12_h_l_00_31(net3032[0:23]), .SP12_h_l_00_30(net3031[0:23]),
     .SP12_h_l_00_29(net3034[0:23]), .SP12_h_l_00_28(net3033[0:23]),
     .SP12_h_l_00_27(net3035[0:23]), .SP12_h_l_00_26(net2960[0:23]),
     .SP12_h_l_00_25(net2969[0:23]), .SP12_h_l_00_24(net2968[0:23]),
     .SP12_h_l_00_23(net2967[0:23]), .SP12_h_l_00_22(net2966[0:23]),
     .SP12_h_l_00_21(net2965[0:23]), .SP12_h_l_00_20(net2901[0:23]),
     .SP12_h_l_00_18(net2903[0:23]), .SP12_h_l_00_19(net2902[0:23]),
     .SP12_h_l_00_17(net2904[0:23]), .slf_op_00_30(slf_op_33_30[3:0]),
     .wl(wl_r[255:0]), .shift(net4851), .bs_en(net4854),
     .mode(net4850), .sdi(net2191), .hiz_b(net4853), .prog(prog),
     .hold(hold_r_t), .update(net4852),
     .glb_netwk_col(clk_tree_drv[7:0]), .r(net4855),
     .spi_ss_in_b(spi_ss_in_b_r[63:32]), .sdo(net4856),
     .bl(bl[1743:1726]), .tclk(net4849), .spioeb({tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}), .spiout({tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}));
array_BRAM_1x8top I_bram_25_top ( .glb_netwk(net2204[0:7]),
     .bm_sdo_i(bm_sdo_i), .bm_sclkrw_o(bm_sclkrw_o),
     .bm_sdi_o(bm_sdi_o), .bm_sweb_o(bm_sweb_o), .bm_sdo_o(bm_sdo_o),
     .bm_sweb_i(bm_sweb_i), .bm_sdi_i(bm_sdi_i),
     .bm_sclkrw_i(bm_sclkrw_i), .wl(wl_r[255:0]),
     .pgate(pgate_r[255:0]), .vdd_cntl(vdd_cntl_r[255:0]),
     .reset_b(reset_r[255:0]), .sp12_h_r_01(net2217[0:23]),
     .lft_op_10(net3931[0:7]), .sp4_h_l_04(net3404[0:47]),
     .sp4_h_l_06(net3431[0:47]), .lft_op_09(net3932[0:7]),
     .lft_op_08(net3933[0:7]), .lft_op_06(net3935[0:7]),
     .lft_op_07(net3934[0:7]), .lft_op_05(net3936[0:7]),
     .lft_op_03(net3865[0:7]), .lft_op_04(net3875[0:7]),
     .lft_op_02(net3867[0:7]), .sp4_h_r_09(net2229[0:47]),
     .bnr_op_01(bnr_op_25_17[7:0]), .sp4_r_v_b_01(sp4_v_b_26_17[47:0]),
     .sp4_r_v_b_02(net2232[0:47]), .sp4_r_v_b_03(net2233[0:47]),
     .sp4_r_v_b_04(net2234[0:47]), .sp4_r_v_b_05(net2235[0:47]),
     .sp4_r_v_b_06(net2236[0:47]), .sp4_r_v_b_07(net2237[0:47]),
     .sp4_r_v_b_08(net2238[0:47]), .sp4_r_v_b_09(net2239[0:47]),
     .sp4_r_v_b_10(net2240[0:47]), .sp4_r_v_b_11(net2241[0:47]),
     .sp4_r_v_b_12(net2242[0:47]), .sp4_r_v_b_13(net2243[0:47]),
     .sp4_r_v_b_14(net2244[0:47]), .sp4_r_v_b_16(net2245[0:47]),
     .sp4_r_v_b_15(net2246[0:47]), .bnl_op_01(bnl_op_25_17[7:0]),
     .lft_op_01(slf_op_24_17[7:0]), .bot_op_01(bot_op_25_17[7:0]),
     .sp12_v_b_01(sp12_v_b_25_17[23:0]), .sp4_v_b_16(net3510[0:47]),
     .sp4_v_b_15(net3511[0:47]), .sp4_v_b_14(net3513[0:47]),
     .sp4_v_b_13(net3512[0:47]), .sp4_v_b_12(net3514[0:47]),
     .sp4_v_b_11(net3515[0:47]), .sp4_v_b_10(net3468[0:47]),
     .sp4_v_b_09(net3467[0:47]), .sp4_v_b_08(net3466[0:47]),
     .sp4_v_b_07(net3465[0:47]), .sp4_v_b_06(net3464[0:47]),
     .sp4_v_b_05(net3463[0:47]), .sp4_v_b_04(net3400[0:47]),
     .sp4_v_b_03(net3401[0:47]), .sp4_v_b_02(net3402[0:47]),
     .sp4_v_b_01(sp4_v_b_25_17[47:0]), .sp12_h_l_10(net3452[0:23]),
     .sp12_h_l_09(net3461[0:23]), .sp12_h_l_08(net3460[0:23]),
     .sp12_h_l_07(net3459[0:23]), .sp12_h_l_06(net3458[0:23]),
     .sp12_h_l_05(net3457[0:23]), .sp12_h_l_04(net3393[0:23]),
     .sp12_h_l_03(net3394[0:23]), .sp12_h_l_02(net3395[0:23]),
     .sp12_h_l_01(net3396[0:23]), .sp12_h_r_10(net2277[0:23]),
     .sp12_h_r_15(net2278[0:23]), .sp12_h_l_15(net3524[0:23]),
     .sp12_h_l_14(net3523[0:23]), .sp12_h_r_14(net2281[0:23]),
     .sp12_h_r_16(net2282[0:23]), .sp12_h_l_16(net3522[0:23]),
     .sp12_h_l_13(net3526[0:23]), .sp12_h_l_12(net3525[0:23]),
     .sp12_h_l_11(net3527[0:23]), .sp12_h_r_13(net2287[0:23]),
     .sp12_h_r_12(net2288[0:23]), .sp12_h_r_11(net2289[0:23]),
     .sp12_h_r_09(net2290[0:23]), .sp12_h_r_08(net2291[0:23]),
     .sp12_h_r_07(net2292[0:23]), .sp12_h_r_06(net2293[0:23]),
     .sp12_h_r_05(net2294[0:23]), .sp12_h_r_04(net2295[0:23]),
     .sp12_h_r_03(net2296[0:23]), .sp12_h_r_02(net2297[0:23]),
     .lft_op_14(net3991[0:7]), .lft_op_13(net3994[0:7]),
     .lft_op_12(net3993[0:7]), .lft_op_11(net3995[0:7]),
     .lft_op_15(net3992[0:7]), .slf_op_15(net3500[0:7]),
     .slf_op_14(net3499[0:7]), .slf_op_13(net3502[0:7]),
     .slf_op_12(net3501[0:7]), .slf_op_11(net3503[0:7]),
     .slf_op_10(net3439[0:7]), .slf_op_09(net3440[0:7]),
     .slf_op_08(net3441[0:7]), .slf_op_07(net3442[0:7]),
     .slf_op_06(net3443[0:7]), .slf_op_05(net3444[0:7]),
     .slf_op_04(net3383[0:7]), .slf_op_03(net3373[0:7]),
     .slf_op_01(slf_op_25_17[7:0]), .slf_op_02(net3375[0:7]),
     .rgt_op_01(slf_op_26_17[7:0]), .rgt_op_02(net2319[0:7]),
     .rgt_op_03(net2320[0:7]), .rgt_op_04(net2321[0:7]),
     .rgt_op_05(net2322[0:7]), .rgt_op_06(net2323[0:7]),
     .rgt_op_07(net2324[0:7]), .rgt_op_08(net2325[0:7]),
     .rgt_op_09(net2326[0:7]), .rgt_op_10(net2327[0:7]),
     .rgt_op_11(net2328[0:7]), .rgt_op_12(net2329[0:7]),
     .rgt_op_13(net2330[0:7]), .rgt_op_14(net2331[0:7]),
     .rgt_op_15(net2332[0:7]), .sp4_h_l_05(net3432[0:47]),
     .sp4_h_l_02(net3406[0:47]), .sp4_h_l_03(net3405[0:47]),
     .sp4_h_l_01(net3407[0:47]), .sp4_h_r_01(net2337[0:47]),
     .sp4_h_r_02(net2338[0:47]), .sp4_h_r_03(net2339[0:47]),
     .sp4_h_r_04(net2340[0:47]), .sp4_h_r_05(net2341[0:47]),
     .sp4_h_r_06(net2342[0:47]), .sp4_h_r_07(net2343[0:47]),
     .sp4_h_r_08(net2344[0:47]), .sp4_h_r_10(net2345[0:47]),
     .sp4_h_r_11(net2346[0:47]), .sp4_h_r_12(net2347[0:47]),
     .sp4_h_r_13(net2348[0:47]), .sp4_h_r_14(net2349[0:47]),
     .sp4_h_r_15(net2350[0:47]), .sp4_h_r_16(net2351[0:47]),
     .lft_op_16(net3863[0:7]), .tnl_op_16({slf_op_24_33[3],
     slf_op_24_33[2], slf_op_24_33[1], slf_op_24_33[0],
     slf_op_24_33[3], slf_op_24_33[2], slf_op_24_33[1],
     slf_op_24_33[0]}), .sp4_v_t_16(net2354[0:47]),
     .top_op_16({slf_op_25_00[3], slf_op_25_00[2], slf_op_25_00[1],
     slf_op_25_00[0], slf_op_25_00[3], slf_op_25_00[2],
     slf_op_25_00[1], slf_op_25_00[0]}), .slf_op_16(net3371[0:7]),
     .tnr_op_16({slf_op_26_33[3], slf_op_26_33[2], slf_op_26_33[1],
     slf_op_26_33[0], slf_op_26_33[3], slf_op_26_33[2],
     slf_op_26_33[1], slf_op_26_33[0]}), .sp12_v_t_16(net2358[0:23]),
     .rgt_op_16(net2359[0:7]), .sp4_h_l_16(net3483[0:47]),
     .sp4_h_l_14(net3481[0:47]), .sp4_h_l_15(net3482[0:47]),
     .sp4_h_l_13(net3480[0:47]), .sp4_h_l_12(net3479[0:47]),
     .sp4_h_l_11(net3478[0:47]), .sp4_h_l_10(net3427[0:47]),
     .sp4_h_l_09(net3428[0:47]), .sp4_h_l_08(net3429[0:47]),
     .sp4_h_l_07(net3430[0:47]), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sreb_i(bm_sreb_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .bm_wdummymux_en_o(bm_wdummymux_en_o),
     .bm_sreb_o(bm_sreb_o), .bm_sclk_o(bm_sclk_o),
     .bm_sa_o(bm_sa_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_o),
     .bm_init_o(bm_init_o), .bl(bl[1347:1306]), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]));
array_LT1x16top I_it_21_top ( .glb_netwk(net2385[0:7]),
     .sp12_v_t_16(net2386[0:23]), .rgt_op_16(net2387[0:7]),
     .top_op_16({slf_op_21_33[3], slf_op_21_33[2], slf_op_21_33[1],
     slf_op_21_33[0], slf_op_21_33[3], slf_op_21_33[2],
     slf_op_21_33[1], slf_op_21_33[0]}), .rgt_op_03(net2389[0:7]),
     .slf_op_02(net4687[0:7]), .rgt_op_02(net2391[0:7]),
     .rgt_op_01(slf_op_22_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3219[0:7]), .lft_op_03(net3209[0:7]),
     .lft_op_02(net3211[0:7]), .lft_op_01(slf_op_20_17[7:0]),
     .rgt_op_04(net2399[0:7]), .carry_in(carry_in_21_17),
     .bnl_op_01(bnl_op_21_17[7:0]), .slf_op_04(net4695[0:7]),
     .slf_op_03(net4685[0:7]), .slf_op_01(slf_op_21_17[7:0]),
     .sp4_h_l_04(net4716[0:47]), .carry_out(net2406),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_21_17[23:0]),
     .sp12_h_r_04(net2409[0:23]), .sp12_h_r_03(net2410[0:23]),
     .sp12_h_r_02(net2411[0:23]), .sp12_h_r_01(net2412[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net4683[0:7]),
     .sp4_v_b_01(sp4_v_b_21_17[47:0]), .sp4_r_v_b_04(net2416[0:47]),
     .sp4_r_v_b_03(net2417[0:47]), .sp4_r_v_b_02(net2418[0:47]),
     .sp4_r_v_b_01(sp4_v_b_22_17[47:0]), .sp4_h_r_04(net2420[0:47]),
     .sp4_h_r_03(net2421[0:47]), .sp4_h_r_02(net2422[0:47]),
     .sp4_h_r_01(net2423[0:47]), .sp4_h_l_03(net4717[0:47]),
     .sp4_h_l_02(net4718[0:47]), .sp4_h_l_01(net4719[0:47]),
     .bl(bl[1143:1090]), .bot_op_01(bot_op_21_17[7:0]),
     .sp12_h_l_01(net4708[0:23]), .sp12_h_l_02(net4707[0:23]),
     .sp12_h_l_03(net4706[0:23]), .sp12_h_l_04(net4705[0:23]),
     .sp4_v_b_04(net4712[0:47]), .sp4_v_b_03(net4713[0:47]),
     .sp4_v_b_02(net4714[0:47]), .bnr_op_01(bnr_op_21_17[7:0]),
     .sp4_h_l_05(net4744[0:47]), .sp4_h_l_06(net4743[0:47]),
     .sp4_h_l_07(net4742[0:47]), .sp4_h_l_08(net4741[0:47]),
     .sp4_h_l_09(net4740[0:47]), .sp4_h_l_10(net4739[0:47]),
     .sp4_h_r_10(net2443[0:47]), .sp4_h_r_09(net2444[0:47]),
     .sp4_h_r_08(net2445[0:47]), .sp4_h_r_07(net2446[0:47]),
     .sp4_h_r_06(net2447[0:47]), .sp4_h_r_05(net2448[0:47]),
     .slf_op_05(net4756[0:7]), .slf_op_06(net4755[0:7]),
     .slf_op_07(net4754[0:7]), .slf_op_08(net4753[0:7]),
     .slf_op_09(net4752[0:7]), .slf_op_10(net4751[0:7]),
     .rgt_op_10(net2455[0:7]), .rgt_op_09(net2456[0:7]),
     .rgt_op_08(net2457[0:7]), .rgt_op_07(net2458[0:7]),
     .rgt_op_06(net2459[0:7]), .rgt_op_05(net2460[0:7]),
     .lft_op_10(net3275[0:7]), .lft_op_09(net3276[0:7]),
     .lft_op_08(net3277[0:7]), .lft_op_07(net3278[0:7]),
     .lft_op_06(net3279[0:7]), .lft_op_05(net3280[0:7]),
     .sp12_h_l_10(net4764[0:23]), .sp12_h_r_10(net2468[0:23]),
     .sp12_h_l_09(net4773[0:23]), .sp12_h_l_08(net4772[0:23]),
     .sp12_h_l_07(net4771[0:23]), .sp12_h_l_06(net4770[0:23]),
     .sp12_h_r_05(net2473[0:23]), .sp12_h_r_06(net2474[0:23]),
     .sp12_h_r_07(net2475[0:23]), .sp12_h_r_08(net2476[0:23]),
     .sp12_h_r_09(net2477[0:23]), .sp12_h_l_05(net4769[0:23]),
     .sp4_r_v_b_05(net2479[0:47]), .sp4_r_v_b_06(net2480[0:47]),
     .sp4_r_v_b_07(net2481[0:47]), .sp4_r_v_b_08(net2482[0:47]),
     .sp4_r_v_b_09(net2483[0:47]), .sp4_r_v_b_10(net2484[0:47]),
     .sp4_v_b_10(net4780[0:47]), .sp4_v_b_09(net4779[0:47]),
     .sp4_v_b_08(net4778[0:47]), .sp4_v_b_07(net4777[0:47]),
     .sp4_v_b_06(net4776[0:47]), .sp4_v_b_05(net4775[0:47]),
     .sp4_v_t_16(net2491[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net2494[0:47]),
     .sp4_h_r_12(net2495[0:47]), .sp4_h_r_13(net2496[0:47]),
     .sp4_h_r_14(net2497[0:47]), .sp4_h_r_15(net2498[0:47]),
     .sp4_h_r_16(net2499[0:47]), .sp4_h_l_16(net4795[0:47]),
     .sp4_h_l_15(net4794[0:47]), .sp4_h_l_14(net4793[0:47]),
     .sp4_h_l_13(net4792[0:47]), .sp4_h_l_12(net4791[0:47]),
     .sp4_h_l_11(net4790[0:47]), .tnr_op_16({slf_op_22_33[3],
     slf_op_22_33[2], slf_op_22_33[1], slf_op_22_33[0],
     slf_op_22_33[3], slf_op_22_33[2], slf_op_22_33[1],
     slf_op_22_33[0]}), .tnl_op_16({slf_op_20_33[3], slf_op_20_33[2],
     slf_op_20_33[1], slf_op_20_33[0], slf_op_20_33[3],
     slf_op_20_33[2], slf_op_20_33[1], slf_op_20_33[0]}),
     .lft_op_16(net3207[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net4812[0:7]), .slf_op_14(net4811[0:7]),
     .slf_op_13(net4814[0:7]), .slf_op_12(net4813[0:7]),
     .slf_op_11(net4815[0:7]), .rgt_op_14(net2515[0:7]),
     .rgt_op_15(net2516[0:7]), .rgt_op_12(net2517[0:7]),
     .rgt_op_13(net2518[0:7]), .rgt_op_11(net2519[0:7]),
     .sp4_v_b_16(net4822[0:47]), .sp4_v_b_14(net4825[0:47]),
     .sp4_v_b_15(net4823[0:47]), .sp4_v_b_13(net4824[0:47]),
     .sp4_v_b_11(net4827[0:47]), .sp4_v_b_12(net4826[0:47]),
     .sp4_r_v_b_16(net2526[0:47]), .sp4_r_v_b_15(net2527[0:47]),
     .sp4_r_v_b_13(net2528[0:47]), .sp4_r_v_b_14(net2529[0:47]),
     .sp4_r_v_b_12(net2530[0:47]), .sp4_r_v_b_11(net2531[0:47]),
     .sp12_h_l_16(net4834[0:23]), .sp12_h_l_15(net4836[0:23]),
     .sp12_h_l_14(net4835[0:23]), .sp12_h_l_13(net4838[0:23]),
     .sp12_h_l_12(net4837[0:23]), .sp12_h_l_11(net4839[0:23]),
     .sp12_h_r_16(net2538[0:23]), .sp12_h_r_14(net2539[0:23]),
     .sp12_h_r_15(net2540[0:23]), .sp12_h_r_12(net2541[0:23]),
     .sp12_h_r_13(net2542[0:23]), .sp12_h_r_11(net2543[0:23]),
     .lft_op_14(net3335[0:7]), .lft_op_15(net3336[0:7]),
     .lft_op_12(net3337[0:7]), .lft_op_11(net3339[0:7]),
     .lft_op_13(net3338[0:7]));
array_LT1x16top I_it_28_top ( .glb_netwk(net2549[0:7]),
     .sp12_v_t_16(net2550[0:23]), .rgt_op_16(net2551[0:7]),
     .top_op_16({slf_op_28_33[3], slf_op_28_33[2], slf_op_28_33[1],
     slf_op_28_33[0], slf_op_28_33[3], slf_op_28_33[2],
     slf_op_28_33[1], slf_op_28_33[0]}), .rgt_op_03(net2553[0:7]),
     .slf_op_02(net2719[0:7]), .rgt_op_02(net2555[0:7]),
     .rgt_op_01(slf_op_29_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4203[0:7]), .lft_op_03(net4193[0:7]),
     .lft_op_02(net4195[0:7]), .lft_op_01(slf_op_27_17[7:0]),
     .rgt_op_04(net2563[0:7]), .carry_in(carry_in_28_17),
     .bnl_op_01(bnl_op_28_17[7:0]), .slf_op_04(net2727[0:7]),
     .slf_op_03(net2717[0:7]), .slf_op_01(slf_op_28_17[7:0]),
     .sp4_h_l_04(net2748[0:47]), .carry_out(net2570),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_28_17[23:0]),
     .sp12_h_r_04(net2573[0:23]), .sp12_h_r_03(net2574[0:23]),
     .sp12_h_r_02(net2575[0:23]), .sp12_h_r_01(net2576[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2715[0:7]),
     .sp4_v_b_01(sp4_v_b_28_17[47:0]), .sp4_r_v_b_04(net2580[0:47]),
     .sp4_r_v_b_03(net2581[0:47]), .sp4_r_v_b_02(net2582[0:47]),
     .sp4_r_v_b_01(sp4_v_b_29_17[47:0]), .sp4_h_r_04(net2584[0:47]),
     .sp4_h_r_03(net2585[0:47]), .sp4_h_r_02(net2586[0:47]),
     .sp4_h_r_01(net2587[0:47]), .sp4_h_l_03(net2749[0:47]),
     .sp4_h_l_02(net2750[0:47]), .sp4_h_l_01(net2751[0:47]),
     .bl(bl[1509:1456]), .bot_op_01(bot_op_28_17[7:0]),
     .sp12_h_l_01(net2740[0:23]), .sp12_h_l_02(net2739[0:23]),
     .sp12_h_l_03(net2738[0:23]), .sp12_h_l_04(net2737[0:23]),
     .sp4_v_b_04(net2744[0:47]), .sp4_v_b_03(net2745[0:47]),
     .sp4_v_b_02(net2746[0:47]), .bnr_op_01(bnr_op_28_17[7:0]),
     .sp4_h_l_05(net2776[0:47]), .sp4_h_l_06(net2775[0:47]),
     .sp4_h_l_07(net2774[0:47]), .sp4_h_l_08(net2773[0:47]),
     .sp4_h_l_09(net2772[0:47]), .sp4_h_l_10(net2771[0:47]),
     .sp4_h_r_10(net2607[0:47]), .sp4_h_r_09(net2608[0:47]),
     .sp4_h_r_08(net2609[0:47]), .sp4_h_r_07(net2610[0:47]),
     .sp4_h_r_06(net2611[0:47]), .sp4_h_r_05(net2612[0:47]),
     .slf_op_05(net2788[0:7]), .slf_op_06(net2787[0:7]),
     .slf_op_07(net2786[0:7]), .slf_op_08(net2785[0:7]),
     .slf_op_09(net2784[0:7]), .slf_op_10(net2783[0:7]),
     .rgt_op_10(net2619[0:7]), .rgt_op_09(net2620[0:7]),
     .rgt_op_08(net2621[0:7]), .rgt_op_07(net2622[0:7]),
     .rgt_op_06(net2623[0:7]), .rgt_op_05(net2624[0:7]),
     .lft_op_10(net4259[0:7]), .lft_op_09(net4260[0:7]),
     .lft_op_08(net4261[0:7]), .lft_op_07(net4262[0:7]),
     .lft_op_06(net4263[0:7]), .lft_op_05(net4264[0:7]),
     .sp12_h_l_10(net2796[0:23]), .sp12_h_r_10(net2632[0:23]),
     .sp12_h_l_09(net2805[0:23]), .sp12_h_l_08(net2804[0:23]),
     .sp12_h_l_07(net2803[0:23]), .sp12_h_l_06(net2802[0:23]),
     .sp12_h_r_05(net2637[0:23]), .sp12_h_r_06(net2638[0:23]),
     .sp12_h_r_07(net2639[0:23]), .sp12_h_r_08(net2640[0:23]),
     .sp12_h_r_09(net2641[0:23]), .sp12_h_l_05(net2801[0:23]),
     .sp4_r_v_b_05(net2643[0:47]), .sp4_r_v_b_06(net2644[0:47]),
     .sp4_r_v_b_07(net2645[0:47]), .sp4_r_v_b_08(net2646[0:47]),
     .sp4_r_v_b_09(net2647[0:47]), .sp4_r_v_b_10(net2648[0:47]),
     .sp4_v_b_10(net2812[0:47]), .sp4_v_b_09(net2811[0:47]),
     .sp4_v_b_08(net2810[0:47]), .sp4_v_b_07(net2809[0:47]),
     .sp4_v_b_06(net2808[0:47]), .sp4_v_b_05(net2807[0:47]),
     .sp4_v_t_16(net2655[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net2658[0:47]),
     .sp4_h_r_12(net2659[0:47]), .sp4_h_r_13(net2660[0:47]),
     .sp4_h_r_14(net2661[0:47]), .sp4_h_r_15(net2662[0:47]),
     .sp4_h_r_16(net2663[0:47]), .sp4_h_l_16(net2827[0:47]),
     .sp4_h_l_15(net2826[0:47]), .sp4_h_l_14(net2825[0:47]),
     .sp4_h_l_13(net2824[0:47]), .sp4_h_l_12(net2823[0:47]),
     .sp4_h_l_11(net2822[0:47]), .tnr_op_16({slf_op_29_33[3],
     slf_op_29_33[2], slf_op_29_33[1], slf_op_29_33[0],
     slf_op_29_33[3], slf_op_29_33[2], slf_op_29_33[1],
     slf_op_29_33[0]}), .tnl_op_16({slf_op_27_33[3], slf_op_27_33[2],
     slf_op_27_33[1], slf_op_27_33[0], slf_op_27_33[3],
     slf_op_27_33[2], slf_op_27_33[1], slf_op_27_33[0]}),
     .lft_op_16(net4191[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net2844[0:7]), .slf_op_14(net2843[0:7]),
     .slf_op_13(net2846[0:7]), .slf_op_12(net2845[0:7]),
     .slf_op_11(net2847[0:7]), .rgt_op_14(net2679[0:7]),
     .rgt_op_15(net2680[0:7]), .rgt_op_12(net2681[0:7]),
     .rgt_op_13(net2682[0:7]), .rgt_op_11(net2683[0:7]),
     .sp4_v_b_16(net2854[0:47]), .sp4_v_b_14(net2857[0:47]),
     .sp4_v_b_15(net2855[0:47]), .sp4_v_b_13(net2856[0:47]),
     .sp4_v_b_11(net2859[0:47]), .sp4_v_b_12(net2858[0:47]),
     .sp4_r_v_b_16(net2690[0:47]), .sp4_r_v_b_15(net2691[0:47]),
     .sp4_r_v_b_13(net2692[0:47]), .sp4_r_v_b_14(net2693[0:47]),
     .sp4_r_v_b_12(net2694[0:47]), .sp4_r_v_b_11(net2695[0:47]),
     .sp12_h_l_16(net2866[0:23]), .sp12_h_l_15(net2868[0:23]),
     .sp12_h_l_14(net2867[0:23]), .sp12_h_l_13(net2870[0:23]),
     .sp12_h_l_12(net2869[0:23]), .sp12_h_l_11(net2871[0:23]),
     .sp12_h_r_16(net2702[0:23]), .sp12_h_r_14(net2703[0:23]),
     .sp12_h_r_15(net2704[0:23]), .sp12_h_r_12(net2705[0:23]),
     .sp12_h_r_13(net2706[0:23]), .sp12_h_r_11(net2707[0:23]),
     .lft_op_14(net4319[0:7]), .lft_op_15(net4320[0:7]),
     .lft_op_12(net4321[0:7]), .lft_op_11(net4323[0:7]),
     .lft_op_13(net4322[0:7]));
array_LT1x16top I_it_27_top ( .glb_netwk(net2713[0:7]),
     .sp12_v_t_16(net2714[0:23]), .rgt_op_16(net2715[0:7]),
     .top_op_16({slf_op_27_33[3], slf_op_27_33[2], slf_op_27_33[1],
     slf_op_27_33[0], slf_op_27_33[3], slf_op_27_33[2],
     slf_op_27_33[1], slf_op_27_33[0]}), .rgt_op_03(net2717[0:7]),
     .slf_op_02(net4195[0:7]), .rgt_op_02(net2719[0:7]),
     .rgt_op_01(slf_op_28_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2321[0:7]), .lft_op_03(net2320[0:7]),
     .lft_op_02(net2319[0:7]), .lft_op_01(slf_op_26_17[7:0]),
     .rgt_op_04(net2727[0:7]), .carry_in(carry_in_27_17),
     .bnl_op_01(bnl_op_27_17[7:0]), .slf_op_04(net4203[0:7]),
     .slf_op_03(net4193[0:7]), .slf_op_01(slf_op_27_17[7:0]),
     .sp4_h_l_04(net4224[0:47]), .carry_out(net2734),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_27_17[23:0]),
     .sp12_h_r_04(net2737[0:23]), .sp12_h_r_03(net2738[0:23]),
     .sp12_h_r_02(net2739[0:23]), .sp12_h_r_01(net2740[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net4191[0:7]),
     .sp4_v_b_01(sp4_v_b_27_17[47:0]), .sp4_r_v_b_04(net2744[0:47]),
     .sp4_r_v_b_03(net2745[0:47]), .sp4_r_v_b_02(net2746[0:47]),
     .sp4_r_v_b_01(sp4_v_b_28_17[47:0]), .sp4_h_r_04(net2748[0:47]),
     .sp4_h_r_03(net2749[0:47]), .sp4_h_r_02(net2750[0:47]),
     .sp4_h_r_01(net2751[0:47]), .sp4_h_l_03(net4225[0:47]),
     .sp4_h_l_02(net4226[0:47]), .sp4_h_l_01(net4227[0:47]),
     .bl(bl[1455:1402]), .bot_op_01(bot_op_27_17[7:0]),
     .sp12_h_l_01(net4216[0:23]), .sp12_h_l_02(net4215[0:23]),
     .sp12_h_l_03(net4214[0:23]), .sp12_h_l_04(net4213[0:23]),
     .sp4_v_b_04(net4220[0:47]), .sp4_v_b_03(net4221[0:47]),
     .sp4_v_b_02(net4222[0:47]), .bnr_op_01(bnr_op_27_17[7:0]),
     .sp4_h_l_05(net4252[0:47]), .sp4_h_l_06(net4251[0:47]),
     .sp4_h_l_07(net4250[0:47]), .sp4_h_l_08(net4249[0:47]),
     .sp4_h_l_09(net4248[0:47]), .sp4_h_l_10(net4247[0:47]),
     .sp4_h_r_10(net2771[0:47]), .sp4_h_r_09(net2772[0:47]),
     .sp4_h_r_08(net2773[0:47]), .sp4_h_r_07(net2774[0:47]),
     .sp4_h_r_06(net2775[0:47]), .sp4_h_r_05(net2776[0:47]),
     .slf_op_05(net4264[0:7]), .slf_op_06(net4263[0:7]),
     .slf_op_07(net4262[0:7]), .slf_op_08(net4261[0:7]),
     .slf_op_09(net4260[0:7]), .slf_op_10(net4259[0:7]),
     .rgt_op_10(net2783[0:7]), .rgt_op_09(net2784[0:7]),
     .rgt_op_08(net2785[0:7]), .rgt_op_07(net2786[0:7]),
     .rgt_op_06(net2787[0:7]), .rgt_op_05(net2788[0:7]),
     .lft_op_10(net2327[0:7]), .lft_op_09(net2326[0:7]),
     .lft_op_08(net2325[0:7]), .lft_op_07(net2324[0:7]),
     .lft_op_06(net2323[0:7]), .lft_op_05(net2322[0:7]),
     .sp12_h_l_10(net4272[0:23]), .sp12_h_r_10(net2796[0:23]),
     .sp12_h_l_09(net4281[0:23]), .sp12_h_l_08(net4280[0:23]),
     .sp12_h_l_07(net4279[0:23]), .sp12_h_l_06(net4278[0:23]),
     .sp12_h_r_05(net2801[0:23]), .sp12_h_r_06(net2802[0:23]),
     .sp12_h_r_07(net2803[0:23]), .sp12_h_r_08(net2804[0:23]),
     .sp12_h_r_09(net2805[0:23]), .sp12_h_l_05(net4277[0:23]),
     .sp4_r_v_b_05(net2807[0:47]), .sp4_r_v_b_06(net2808[0:47]),
     .sp4_r_v_b_07(net2809[0:47]), .sp4_r_v_b_08(net2810[0:47]),
     .sp4_r_v_b_09(net2811[0:47]), .sp4_r_v_b_10(net2812[0:47]),
     .sp4_v_b_10(net4288[0:47]), .sp4_v_b_09(net4287[0:47]),
     .sp4_v_b_08(net4286[0:47]), .sp4_v_b_07(net4285[0:47]),
     .sp4_v_b_06(net4284[0:47]), .sp4_v_b_05(net4283[0:47]),
     .sp4_v_t_16(net2819[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net2822[0:47]),
     .sp4_h_r_12(net2823[0:47]), .sp4_h_r_13(net2824[0:47]),
     .sp4_h_r_14(net2825[0:47]), .sp4_h_r_15(net2826[0:47]),
     .sp4_h_r_16(net2827[0:47]), .sp4_h_l_16(net4303[0:47]),
     .sp4_h_l_15(net4302[0:47]), .sp4_h_l_14(net4301[0:47]),
     .sp4_h_l_13(net4300[0:47]), .sp4_h_l_12(net4299[0:47]),
     .sp4_h_l_11(net4298[0:47]), .tnr_op_16({slf_op_28_33[3],
     slf_op_28_33[2], slf_op_28_33[1], slf_op_28_33[0],
     slf_op_28_33[3], slf_op_28_33[2], slf_op_28_33[1],
     slf_op_28_33[0]}), .tnl_op_16({slf_op_26_33[3], slf_op_26_33[2],
     slf_op_26_33[1], slf_op_26_33[0], slf_op_26_33[3],
     slf_op_26_33[2], slf_op_26_33[1], slf_op_26_33[0]}),
     .lft_op_16(net2359[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net4320[0:7]), .slf_op_14(net4319[0:7]),
     .slf_op_13(net4322[0:7]), .slf_op_12(net4321[0:7]),
     .slf_op_11(net4323[0:7]), .rgt_op_14(net2843[0:7]),
     .rgt_op_15(net2844[0:7]), .rgt_op_12(net2845[0:7]),
     .rgt_op_13(net2846[0:7]), .rgt_op_11(net2847[0:7]),
     .sp4_v_b_16(net4330[0:47]), .sp4_v_b_14(net4333[0:47]),
     .sp4_v_b_15(net4331[0:47]), .sp4_v_b_13(net4332[0:47]),
     .sp4_v_b_11(net4335[0:47]), .sp4_v_b_12(net4334[0:47]),
     .sp4_r_v_b_16(net2854[0:47]), .sp4_r_v_b_15(net2855[0:47]),
     .sp4_r_v_b_13(net2856[0:47]), .sp4_r_v_b_14(net2857[0:47]),
     .sp4_r_v_b_12(net2858[0:47]), .sp4_r_v_b_11(net2859[0:47]),
     .sp12_h_l_16(net4342[0:23]), .sp12_h_l_15(net4344[0:23]),
     .sp12_h_l_14(net4343[0:23]), .sp12_h_l_13(net4346[0:23]),
     .sp12_h_l_12(net4345[0:23]), .sp12_h_l_11(net4347[0:23]),
     .sp12_h_r_16(net2866[0:23]), .sp12_h_r_14(net2867[0:23]),
     .sp12_h_r_15(net2868[0:23]), .sp12_h_r_12(net2869[0:23]),
     .sp12_h_r_13(net2870[0:23]), .sp12_h_r_11(net2871[0:23]),
     .lft_op_14(net2331[0:7]), .lft_op_15(net2332[0:7]),
     .lft_op_12(net2329[0:7]), .lft_op_11(net2328[0:7]),
     .lft_op_13(net2330[0:7]));
array_LT1x16top I_it_32_top ( .glb_netwk(net2877[0:7]),
     .sp12_v_t_16(net2878[0:23]), .rgt_op_16({slf_op_33_32[3],
     slf_op_33_32[2], slf_op_33_32[1], slf_op_33_32[0],
     slf_op_33_32[3], slf_op_33_32[2], slf_op_33_32[1],
     slf_op_33_32[0]}), .top_op_16({slf_op_32_33[3], slf_op_32_33[2],
     slf_op_32_33[1], slf_op_32_33[0], slf_op_32_33[3],
     slf_op_32_33[2], slf_op_32_33[1], slf_op_32_33[0]}),
     .rgt_op_03({slf_op_33_19[3], slf_op_33_19[2], slf_op_33_19[1],
     slf_op_33_19[0], slf_op_33_19[3], slf_op_33_19[2],
     slf_op_33_19[1], slf_op_33_19[0]}), .slf_op_02(net3539[0:7]),
     .rgt_op_02({slf_op_33_18[3], slf_op_33_18[2], slf_op_33_18[1],
     slf_op_33_18[0], slf_op_33_18[3], slf_op_33_18[2],
     slf_op_33_18[1], slf_op_33_18[0]}), .rgt_op_01({slf_op_33_17[3],
     slf_op_33_17[2], slf_op_33_17[1], slf_op_33_17[0],
     slf_op_33_17[3], slf_op_33_17[2], slf_op_33_17[1],
     slf_op_33_17[0]}), .purst(purst), .prog(prog),
     .lft_op_04(net4039[0:7]), .lft_op_03(net4029[0:7]),
     .lft_op_02(net4031[0:7]), .lft_op_01(slf_op_31_17[7:0]),
     .rgt_op_04({slf_op_33_20[3], slf_op_33_20[2], slf_op_33_20[1],
     slf_op_33_20[0], slf_op_33_20[3], slf_op_33_20[2],
     slf_op_33_20[1], slf_op_33_20[0]}), .carry_in(carry_in_32_17),
     .bnl_op_01(bnl_op_32_17[7:0]), .slf_op_04(net3547[0:7]),
     .slf_op_03(net3537[0:7]), .slf_op_01(slf_op_32_17[7:0]),
     .sp4_h_l_04(net3568[0:47]), .carry_out(net2898),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_32_17[23:0]),
     .sp12_h_r_04(net2901[0:23]), .sp12_h_r_03(net2902[0:23]),
     .sp12_h_r_02(net2903[0:23]), .sp12_h_r_01(net2904[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net3535[0:7]),
     .sp4_v_b_01(sp4_v_b_32_17[47:0]), .sp4_r_v_b_04(net2908[0:47]),
     .sp4_r_v_b_03(net2909[0:47]), .sp4_r_v_b_02(net2910[0:47]),
     .sp4_r_v_b_01(net2911[0:47]), .sp4_h_r_04(net2912[0:47]),
     .sp4_h_r_03(net2913[0:47]), .sp4_h_r_02(net2914[0:47]),
     .sp4_h_r_01(net2915[0:47]), .sp4_h_l_03(net3569[0:47]),
     .sp4_h_l_02(net3570[0:47]), .sp4_h_l_01(net3571[0:47]),
     .bl(bl[1725:1672]), .bot_op_01(bot_op_32_17[7:0]),
     .sp12_h_l_01(net3560[0:23]), .sp12_h_l_02(net3559[0:23]),
     .sp12_h_l_03(net3558[0:23]), .sp12_h_l_04(net3557[0:23]),
     .sp4_v_b_04(net3564[0:47]), .sp4_v_b_03(net3565[0:47]),
     .sp4_v_b_02(net3566[0:47]), .bnr_op_01(bnr_op_32_17[7:0]),
     .sp4_h_l_05(net3596[0:47]), .sp4_h_l_06(net3595[0:47]),
     .sp4_h_l_07(net3594[0:47]), .sp4_h_l_08(net3593[0:47]),
     .sp4_h_l_09(net3592[0:47]), .sp4_h_l_10(net3591[0:47]),
     .sp4_h_r_10(net2935[0:47]), .sp4_h_r_09(net2936[0:47]),
     .sp4_h_r_08(net2937[0:47]), .sp4_h_r_07(net2938[0:47]),
     .sp4_h_r_06(net2939[0:47]), .sp4_h_r_05(net2940[0:47]),
     .slf_op_05(net3608[0:7]), .slf_op_06(net3607[0:7]),
     .slf_op_07(net3606[0:7]), .slf_op_08(net3605[0:7]),
     .slf_op_09(net3604[0:7]), .slf_op_10(net3603[0:7]),
     .rgt_op_10({slf_op_33_26[3], slf_op_33_26[2], slf_op_33_26[1],
     slf_op_33_26[0], slf_op_33_26[3], slf_op_33_26[2],
     slf_op_33_26[1], slf_op_33_26[0]}), .rgt_op_09({slf_op_33_25[3],
     slf_op_33_25[2], slf_op_33_25[1], slf_op_33_25[0],
     slf_op_33_25[3], slf_op_33_25[2], slf_op_33_25[1],
     slf_op_33_25[0]}), .rgt_op_08({slf_op_33_24[3], slf_op_33_24[2],
     slf_op_33_24[1], slf_op_33_24[0], slf_op_33_24[3],
     slf_op_33_24[2], slf_op_33_24[1], slf_op_33_24[0]}),
     .rgt_op_07({slf_op_33_23[3], slf_op_33_23[2], slf_op_33_23[1],
     slf_op_33_23[0], slf_op_33_23[3], slf_op_33_23[2],
     slf_op_33_23[1], slf_op_33_23[0]}), .rgt_op_06({slf_op_33_22[3],
     slf_op_33_22[2], slf_op_33_22[1], slf_op_33_22[0],
     slf_op_33_22[3], slf_op_33_22[2], slf_op_33_22[1],
     slf_op_33_22[0]}), .rgt_op_05({slf_op_33_21[3], slf_op_33_21[2],
     slf_op_33_21[1], slf_op_33_21[0], slf_op_33_21[3],
     slf_op_33_21[2], slf_op_33_21[1], slf_op_33_21[0]}),
     .lft_op_10(net4095[0:7]), .lft_op_09(net4096[0:7]),
     .lft_op_08(net4097[0:7]), .lft_op_07(net4098[0:7]),
     .lft_op_06(net4099[0:7]), .lft_op_05(net4100[0:7]),
     .sp12_h_l_10(net3616[0:23]), .sp12_h_r_10(net2960[0:23]),
     .sp12_h_l_09(net3625[0:23]), .sp12_h_l_08(net3624[0:23]),
     .sp12_h_l_07(net3623[0:23]), .sp12_h_l_06(net3622[0:23]),
     .sp12_h_r_05(net2965[0:23]), .sp12_h_r_06(net2966[0:23]),
     .sp12_h_r_07(net2967[0:23]), .sp12_h_r_08(net2968[0:23]),
     .sp12_h_r_09(net2969[0:23]), .sp12_h_l_05(net3621[0:23]),
     .sp4_r_v_b_05(net2971[0:47]), .sp4_r_v_b_06(net2972[0:47]),
     .sp4_r_v_b_07(net2973[0:47]), .sp4_r_v_b_08(net2974[0:47]),
     .sp4_r_v_b_09(net2975[0:47]), .sp4_r_v_b_10(net2976[0:47]),
     .sp4_v_b_10(net3632[0:47]), .sp4_v_b_09(net3631[0:47]),
     .sp4_v_b_08(net3630[0:47]), .sp4_v_b_07(net3629[0:47]),
     .sp4_v_b_06(net3628[0:47]), .sp4_v_b_05(net3627[0:47]),
     .sp4_v_t_16(net2983[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net2986[0:47]),
     .sp4_h_r_12(net2987[0:47]), .sp4_h_r_13(net2988[0:47]),
     .sp4_h_r_14(net2989[0:47]), .sp4_h_r_15(net2990[0:47]),
     .sp4_h_r_16(net2991[0:47]), .sp4_h_l_16(net3647[0:47]),
     .sp4_h_l_15(net3646[0:47]), .sp4_h_l_14(net3645[0:47]),
     .sp4_h_l_13(net3644[0:47]), .sp4_h_l_12(net3643[0:47]),
     .sp4_h_l_11(net3642[0:47]), .tnr_op_16({tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .tnl_op_16({slf_op_31_33[3], slf_op_31_33[2], slf_op_31_33[1],
     slf_op_31_33[0], slf_op_31_33[3], slf_op_31_33[2],
     slf_op_31_33[1], slf_op_31_33[0]}), .lft_op_16(net4027[0:7]),
     .wl(wl_r[255:0]), .slf_op_15(net3664[0:7]),
     .slf_op_14(net3663[0:7]), .slf_op_13(net3666[0:7]),
     .slf_op_12(net3665[0:7]), .slf_op_11(net3667[0:7]),
     .rgt_op_14({slf_op_33_30[3], slf_op_33_30[2], slf_op_33_30[1],
     slf_op_33_30[0], slf_op_33_30[3], slf_op_33_30[2],
     slf_op_33_30[1], slf_op_33_30[0]}), .rgt_op_15({slf_op_33_31[3],
     slf_op_33_31[2], slf_op_33_31[1], slf_op_33_31[0],
     slf_op_33_31[3], slf_op_33_31[2], slf_op_33_31[1],
     slf_op_33_31[0]}), .rgt_op_12({slf_op_33_28[3], slf_op_33_28[2],
     slf_op_33_28[1], slf_op_33_28[0], slf_op_33_28[3],
     slf_op_33_28[2], slf_op_33_28[1], slf_op_33_28[0]}),
     .rgt_op_13({slf_op_33_29[3], slf_op_33_29[2], slf_op_33_29[1],
     slf_op_33_29[0], slf_op_33_29[3], slf_op_33_29[2],
     slf_op_33_29[1], slf_op_33_29[0]}), .rgt_op_11({slf_op_33_27[3],
     slf_op_33_27[2], slf_op_33_27[1], slf_op_33_27[0],
     slf_op_33_27[3], slf_op_33_27[2], slf_op_33_27[1],
     slf_op_33_27[0]}), .sp4_v_b_16(net3674[0:47]),
     .sp4_v_b_14(net3677[0:47]), .sp4_v_b_15(net3675[0:47]),
     .sp4_v_b_13(net3676[0:47]), .sp4_v_b_11(net3679[0:47]),
     .sp4_v_b_12(net3678[0:47]), .sp4_r_v_b_16(net3018[0:47]),
     .sp4_r_v_b_15(net3019[0:47]), .sp4_r_v_b_13(net3020[0:47]),
     .sp4_r_v_b_14(net3021[0:47]), .sp4_r_v_b_12(net3022[0:47]),
     .sp4_r_v_b_11(net3023[0:47]), .sp12_h_l_16(net3686[0:23]),
     .sp12_h_l_15(net3688[0:23]), .sp12_h_l_14(net3687[0:23]),
     .sp12_h_l_13(net3690[0:23]), .sp12_h_l_12(net3689[0:23]),
     .sp12_h_l_11(net3691[0:23]), .sp12_h_r_16(net3030[0:23]),
     .sp12_h_r_14(net3031[0:23]), .sp12_h_r_15(net3032[0:23]),
     .sp12_h_r_12(net3033[0:23]), .sp12_h_r_13(net3034[0:23]),
     .sp12_h_r_11(net3035[0:23]), .lft_op_14(net4155[0:7]),
     .lft_op_15(net4156[0:7]), .lft_op_12(net4157[0:7]),
     .lft_op_11(net4159[0:7]), .lft_op_13(net4158[0:7]));
array_LT1x16top I_it_22_top ( .glb_netwk(net3041[0:7]),
     .sp12_v_t_16(net3042[0:23]), .rgt_op_16(net3043[0:7]),
     .top_op_16({slf_op_22_33[3], slf_op_22_33[2], slf_op_22_33[1],
     slf_op_22_33[0], slf_op_22_33[3], slf_op_22_33[2],
     slf_op_22_33[1], slf_op_22_33[0]}), .rgt_op_03(net3045[0:7]),
     .slf_op_02(net2391[0:7]), .rgt_op_02(net3047[0:7]),
     .rgt_op_01(slf_op_23_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4695[0:7]), .lft_op_03(net4685[0:7]),
     .lft_op_02(net4687[0:7]), .lft_op_01(slf_op_21_17[7:0]),
     .rgt_op_04(net3055[0:7]), .carry_in(carry_in_22_17),
     .bnl_op_01(bnl_op_22_17[7:0]), .slf_op_04(net2399[0:7]),
     .slf_op_03(net2389[0:7]), .slf_op_01(slf_op_22_17[7:0]),
     .sp4_h_l_04(net2420[0:47]), .carry_out(net3062),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_22_17[23:0]),
     .sp12_h_r_04(net3065[0:23]), .sp12_h_r_03(net3066[0:23]),
     .sp12_h_r_02(net3067[0:23]), .sp12_h_r_01(net3068[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2387[0:7]),
     .sp4_v_b_01(sp4_v_b_22_17[47:0]), .sp4_r_v_b_04(net3072[0:47]),
     .sp4_r_v_b_03(net3073[0:47]), .sp4_r_v_b_02(net3074[0:47]),
     .sp4_r_v_b_01(sp4_v_b_23_17[47:0]), .sp4_h_r_04(net3076[0:47]),
     .sp4_h_r_03(net3077[0:47]), .sp4_h_r_02(net3078[0:47]),
     .sp4_h_r_01(net3079[0:47]), .sp4_h_l_03(net2421[0:47]),
     .sp4_h_l_02(net2422[0:47]), .sp4_h_l_01(net2423[0:47]),
     .bl(bl[1197:1144]), .bot_op_01(bot_op_22_17[7:0]),
     .sp12_h_l_01(net2412[0:23]), .sp12_h_l_02(net2411[0:23]),
     .sp12_h_l_03(net2410[0:23]), .sp12_h_l_04(net2409[0:23]),
     .sp4_v_b_04(net2416[0:47]), .sp4_v_b_03(net2417[0:47]),
     .sp4_v_b_02(net2418[0:47]), .bnr_op_01(bnr_op_22_17[7:0]),
     .sp4_h_l_05(net2448[0:47]), .sp4_h_l_06(net2447[0:47]),
     .sp4_h_l_07(net2446[0:47]), .sp4_h_l_08(net2445[0:47]),
     .sp4_h_l_09(net2444[0:47]), .sp4_h_l_10(net2443[0:47]),
     .sp4_h_r_10(net3099[0:47]), .sp4_h_r_09(net3100[0:47]),
     .sp4_h_r_08(net3101[0:47]), .sp4_h_r_07(net3102[0:47]),
     .sp4_h_r_06(net3103[0:47]), .sp4_h_r_05(net3104[0:47]),
     .slf_op_05(net2460[0:7]), .slf_op_06(net2459[0:7]),
     .slf_op_07(net2458[0:7]), .slf_op_08(net2457[0:7]),
     .slf_op_09(net2456[0:7]), .slf_op_10(net2455[0:7]),
     .rgt_op_10(net3111[0:7]), .rgt_op_09(net3112[0:7]),
     .rgt_op_08(net3113[0:7]), .rgt_op_07(net3114[0:7]),
     .rgt_op_06(net3115[0:7]), .rgt_op_05(net3116[0:7]),
     .lft_op_10(net4751[0:7]), .lft_op_09(net4752[0:7]),
     .lft_op_08(net4753[0:7]), .lft_op_07(net4754[0:7]),
     .lft_op_06(net4755[0:7]), .lft_op_05(net4756[0:7]),
     .sp12_h_l_10(net2468[0:23]), .sp12_h_r_10(net3124[0:23]),
     .sp12_h_l_09(net2477[0:23]), .sp12_h_l_08(net2476[0:23]),
     .sp12_h_l_07(net2475[0:23]), .sp12_h_l_06(net2474[0:23]),
     .sp12_h_r_05(net3129[0:23]), .sp12_h_r_06(net3130[0:23]),
     .sp12_h_r_07(net3131[0:23]), .sp12_h_r_08(net3132[0:23]),
     .sp12_h_r_09(net3133[0:23]), .sp12_h_l_05(net2473[0:23]),
     .sp4_r_v_b_05(net3135[0:47]), .sp4_r_v_b_06(net3136[0:47]),
     .sp4_r_v_b_07(net3137[0:47]), .sp4_r_v_b_08(net3138[0:47]),
     .sp4_r_v_b_09(net3139[0:47]), .sp4_r_v_b_10(net3140[0:47]),
     .sp4_v_b_10(net2484[0:47]), .sp4_v_b_09(net2483[0:47]),
     .sp4_v_b_08(net2482[0:47]), .sp4_v_b_07(net2481[0:47]),
     .sp4_v_b_06(net2480[0:47]), .sp4_v_b_05(net2479[0:47]),
     .sp4_v_t_16(net3147[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net3150[0:47]),
     .sp4_h_r_12(net3151[0:47]), .sp4_h_r_13(net3152[0:47]),
     .sp4_h_r_14(net3153[0:47]), .sp4_h_r_15(net3154[0:47]),
     .sp4_h_r_16(net3155[0:47]), .sp4_h_l_16(net2499[0:47]),
     .sp4_h_l_15(net2498[0:47]), .sp4_h_l_14(net2497[0:47]),
     .sp4_h_l_13(net2496[0:47]), .sp4_h_l_12(net2495[0:47]),
     .sp4_h_l_11(net2494[0:47]), .tnr_op_16({slf_op_23_33[3],
     slf_op_23_33[2], slf_op_23_33[1], slf_op_23_33[0],
     slf_op_23_33[3], slf_op_23_33[2], slf_op_23_33[1],
     slf_op_23_33[0]}), .tnl_op_16({slf_op_21_33[3], slf_op_21_33[2],
     slf_op_21_33[1], slf_op_21_33[0], slf_op_21_33[3],
     slf_op_21_33[2], slf_op_21_33[1], slf_op_21_33[0]}),
     .lft_op_16(net4683[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net2516[0:7]), .slf_op_14(net2515[0:7]),
     .slf_op_13(net2518[0:7]), .slf_op_12(net2517[0:7]),
     .slf_op_11(net2519[0:7]), .rgt_op_14(net3171[0:7]),
     .rgt_op_15(net3172[0:7]), .rgt_op_12(net3173[0:7]),
     .rgt_op_13(net3174[0:7]), .rgt_op_11(net3175[0:7]),
     .sp4_v_b_16(net2526[0:47]), .sp4_v_b_14(net2529[0:47]),
     .sp4_v_b_15(net2527[0:47]), .sp4_v_b_13(net2528[0:47]),
     .sp4_v_b_11(net2531[0:47]), .sp4_v_b_12(net2530[0:47]),
     .sp4_r_v_b_16(net3182[0:47]), .sp4_r_v_b_15(net3183[0:47]),
     .sp4_r_v_b_13(net3184[0:47]), .sp4_r_v_b_14(net3185[0:47]),
     .sp4_r_v_b_12(net3186[0:47]), .sp4_r_v_b_11(net3187[0:47]),
     .sp12_h_l_16(net2538[0:23]), .sp12_h_l_15(net2540[0:23]),
     .sp12_h_l_14(net2539[0:23]), .sp12_h_l_13(net2542[0:23]),
     .sp12_h_l_12(net2541[0:23]), .sp12_h_l_11(net2543[0:23]),
     .sp12_h_r_16(net3194[0:23]), .sp12_h_r_14(net3195[0:23]),
     .sp12_h_r_15(net3196[0:23]), .sp12_h_r_12(net3197[0:23]),
     .sp12_h_r_13(net3198[0:23]), .sp12_h_r_11(net3199[0:23]),
     .lft_op_14(net4811[0:7]), .lft_op_15(net4812[0:7]),
     .lft_op_12(net4813[0:7]), .lft_op_11(net4815[0:7]),
     .lft_op_13(net4814[0:7]));
array_LT1x16top I_it_19_top ( .glb_netwk(net3205[0:7]),
     .sp12_v_t_16(net3206[0:23]), .rgt_op_16(net3207[0:7]),
     .top_op_16({slf_op_19_33[3], slf_op_19_33[2], slf_op_19_33[1],
     slf_op_19_33[0], slf_op_19_33[3], slf_op_19_33[2],
     slf_op_19_33[1], slf_op_19_33[0]}), .rgt_op_03(net3209[0:7]),
     .slf_op_02(net4359[0:7]), .rgt_op_02(net3211[0:7]),
     .rgt_op_01(slf_op_20_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4531[0:7]), .lft_op_03(net4521[0:7]),
     .lft_op_02(net4523[0:7]), .lft_op_01(slf_op_18_17[7:0]),
     .rgt_op_04(net3219[0:7]), .carry_in(carry_in_19_17),
     .bnl_op_01(bnl_op_19_17[7:0]), .slf_op_04(net4367[0:7]),
     .slf_op_03(net4357[0:7]), .slf_op_01(slf_op_19_17[7:0]),
     .sp4_h_l_04(net4388[0:47]), .carry_out(net3226),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_19_17[23:0]),
     .sp12_h_r_04(net3229[0:23]), .sp12_h_r_03(net3230[0:23]),
     .sp12_h_r_02(net3231[0:23]), .sp12_h_r_01(net3232[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net4355[0:7]),
     .sp4_v_b_01(sp4_v_b_19_17[47:0]), .sp4_r_v_b_04(net3236[0:47]),
     .sp4_r_v_b_03(net3237[0:47]), .sp4_r_v_b_02(net3238[0:47]),
     .sp4_r_v_b_01(sp4_v_b_20_17[47:0]), .sp4_h_r_04(net3240[0:47]),
     .sp4_h_r_03(net3241[0:47]), .sp4_h_r_02(net3242[0:47]),
     .sp4_h_r_01(net3243[0:47]), .sp4_h_l_03(net4389[0:47]),
     .sp4_h_l_02(net4390[0:47]), .sp4_h_l_01(net4391[0:47]),
     .bl(bl[1035:982]), .bot_op_01(bot_op_19_17[7:0]),
     .sp12_h_l_01(net4380[0:23]), .sp12_h_l_02(net4379[0:23]),
     .sp12_h_l_03(net4378[0:23]), .sp12_h_l_04(net4377[0:23]),
     .sp4_v_b_04(net4384[0:47]), .sp4_v_b_03(net4385[0:47]),
     .sp4_v_b_02(net4386[0:47]), .bnr_op_01(bnr_op_19_17[7:0]),
     .sp4_h_l_05(net4416[0:47]), .sp4_h_l_06(net4415[0:47]),
     .sp4_h_l_07(net4414[0:47]), .sp4_h_l_08(net4413[0:47]),
     .sp4_h_l_09(net4412[0:47]), .sp4_h_l_10(net4411[0:47]),
     .sp4_h_r_10(net3263[0:47]), .sp4_h_r_09(net3264[0:47]),
     .sp4_h_r_08(net3265[0:47]), .sp4_h_r_07(net3266[0:47]),
     .sp4_h_r_06(net3267[0:47]), .sp4_h_r_05(net3268[0:47]),
     .slf_op_05(net4428[0:7]), .slf_op_06(net4427[0:7]),
     .slf_op_07(net4426[0:7]), .slf_op_08(net4425[0:7]),
     .slf_op_09(net4424[0:7]), .slf_op_10(net4423[0:7]),
     .rgt_op_10(net3275[0:7]), .rgt_op_09(net3276[0:7]),
     .rgt_op_08(net3277[0:7]), .rgt_op_07(net3278[0:7]),
     .rgt_op_06(net3279[0:7]), .rgt_op_05(net3280[0:7]),
     .lft_op_10(net4587[0:7]), .lft_op_09(net4588[0:7]),
     .lft_op_08(net4589[0:7]), .lft_op_07(net4590[0:7]),
     .lft_op_06(net4591[0:7]), .lft_op_05(net4592[0:7]),
     .sp12_h_l_10(net4436[0:23]), .sp12_h_r_10(net3288[0:23]),
     .sp12_h_l_09(net4445[0:23]), .sp12_h_l_08(net4444[0:23]),
     .sp12_h_l_07(net4443[0:23]), .sp12_h_l_06(net4442[0:23]),
     .sp12_h_r_05(net3293[0:23]), .sp12_h_r_06(net3294[0:23]),
     .sp12_h_r_07(net3295[0:23]), .sp12_h_r_08(net3296[0:23]),
     .sp12_h_r_09(net3297[0:23]), .sp12_h_l_05(net4441[0:23]),
     .sp4_r_v_b_05(net3299[0:47]), .sp4_r_v_b_06(net3300[0:47]),
     .sp4_r_v_b_07(net3301[0:47]), .sp4_r_v_b_08(net3302[0:47]),
     .sp4_r_v_b_09(net3303[0:47]), .sp4_r_v_b_10(net3304[0:47]),
     .sp4_v_b_10(net4452[0:47]), .sp4_v_b_09(net4451[0:47]),
     .sp4_v_b_08(net4450[0:47]), .sp4_v_b_07(net4449[0:47]),
     .sp4_v_b_06(net4448[0:47]), .sp4_v_b_05(net4447[0:47]),
     .sp4_v_t_16(net3311[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net3314[0:47]),
     .sp4_h_r_12(net3315[0:47]), .sp4_h_r_13(net3316[0:47]),
     .sp4_h_r_14(net3317[0:47]), .sp4_h_r_15(net3318[0:47]),
     .sp4_h_r_16(net3319[0:47]), .sp4_h_l_16(net4467[0:47]),
     .sp4_h_l_15(net4466[0:47]), .sp4_h_l_14(net4465[0:47]),
     .sp4_h_l_13(net4464[0:47]), .sp4_h_l_12(net4463[0:47]),
     .sp4_h_l_11(net4462[0:47]), .tnr_op_16({slf_op_20_33[3],
     slf_op_20_33[2], slf_op_20_33[1], slf_op_20_33[0],
     slf_op_20_33[3], slf_op_20_33[2], slf_op_20_33[1],
     slf_op_20_33[0]}), .tnl_op_16({slf_op_18_33[3], slf_op_18_33[2],
     slf_op_18_33[1], slf_op_18_33[0], slf_op_18_33[3],
     slf_op_18_33[2], slf_op_18_33[1], slf_op_18_33[0]}),
     .lft_op_16(net4519[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net4484[0:7]), .slf_op_14(net4483[0:7]),
     .slf_op_13(net4486[0:7]), .slf_op_12(net4485[0:7]),
     .slf_op_11(net4487[0:7]), .rgt_op_14(net3335[0:7]),
     .rgt_op_15(net3336[0:7]), .rgt_op_12(net3337[0:7]),
     .rgt_op_13(net3338[0:7]), .rgt_op_11(net3339[0:7]),
     .sp4_v_b_16(net4494[0:47]), .sp4_v_b_14(net4497[0:47]),
     .sp4_v_b_15(net4495[0:47]), .sp4_v_b_13(net4496[0:47]),
     .sp4_v_b_11(net4499[0:47]), .sp4_v_b_12(net4498[0:47]),
     .sp4_r_v_b_16(net3346[0:47]), .sp4_r_v_b_15(net3347[0:47]),
     .sp4_r_v_b_13(net3348[0:47]), .sp4_r_v_b_14(net3349[0:47]),
     .sp4_r_v_b_12(net3350[0:47]), .sp4_r_v_b_11(net3351[0:47]),
     .sp12_h_l_16(net4506[0:23]), .sp12_h_l_15(net4508[0:23]),
     .sp12_h_l_14(net4507[0:23]), .sp12_h_l_13(net4510[0:23]),
     .sp12_h_l_12(net4509[0:23]), .sp12_h_l_11(net4511[0:23]),
     .sp12_h_r_16(net3358[0:23]), .sp12_h_r_14(net3359[0:23]),
     .sp12_h_r_15(net3360[0:23]), .sp12_h_r_12(net3361[0:23]),
     .sp12_h_r_13(net3362[0:23]), .sp12_h_r_11(net3363[0:23]),
     .lft_op_14(net4647[0:7]), .lft_op_15(net4648[0:7]),
     .lft_op_12(net4649[0:7]), .lft_op_11(net4651[0:7]),
     .lft_op_13(net4650[0:7]));
array_LT1x16top I_it_24_top ( .glb_netwk(net3369[0:7]),
     .sp12_v_t_16(net3370[0:23]), .rgt_op_16(net3371[0:7]),
     .top_op_16({slf_op_24_33[3], slf_op_24_33[2], slf_op_24_33[1],
     slf_op_24_33[0], slf_op_24_33[3], slf_op_24_33[2],
     slf_op_24_33[1], slf_op_24_33[0]}), .rgt_op_03(net3373[0:7]),
     .slf_op_02(net3867[0:7]), .rgt_op_02(net3375[0:7]),
     .rgt_op_01(slf_op_25_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3055[0:7]), .lft_op_03(net3045[0:7]),
     .lft_op_02(net3047[0:7]), .lft_op_01(slf_op_23_17[7:0]),
     .rgt_op_04(net3383[0:7]), .carry_in(carry_in_24_17),
     .bnl_op_01(bnl_op_24_17[7:0]), .slf_op_04(net3875[0:7]),
     .slf_op_03(net3865[0:7]), .slf_op_01(slf_op_24_17[7:0]),
     .sp4_h_l_04(net3896[0:47]), .carry_out(net3390),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_24_17[23:0]),
     .sp12_h_r_04(net3393[0:23]), .sp12_h_r_03(net3394[0:23]),
     .sp12_h_r_02(net3395[0:23]), .sp12_h_r_01(net3396[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net3863[0:7]),
     .sp4_v_b_01(sp4_v_b_24_17[47:0]), .sp4_r_v_b_04(net3400[0:47]),
     .sp4_r_v_b_03(net3401[0:47]), .sp4_r_v_b_02(net3402[0:47]),
     .sp4_r_v_b_01(sp4_v_b_25_17[47:0]), .sp4_h_r_04(net3404[0:47]),
     .sp4_h_r_03(net3405[0:47]), .sp4_h_r_02(net3406[0:47]),
     .sp4_h_r_01(net3407[0:47]), .sp4_h_l_03(net3897[0:47]),
     .sp4_h_l_02(net3898[0:47]), .sp4_h_l_01(net3899[0:47]),
     .bl(bl[1305:1252]), .bot_op_01(bot_op_24_17[7:0]),
     .sp12_h_l_01(net3888[0:23]), .sp12_h_l_02(net3887[0:23]),
     .sp12_h_l_03(net3886[0:23]), .sp12_h_l_04(net3885[0:23]),
     .sp4_v_b_04(net3892[0:47]), .sp4_v_b_03(net3893[0:47]),
     .sp4_v_b_02(net3894[0:47]), .bnr_op_01(bnr_op_24_17[7:0]),
     .sp4_h_l_05(net3924[0:47]), .sp4_h_l_06(net3923[0:47]),
     .sp4_h_l_07(net3922[0:47]), .sp4_h_l_08(net3921[0:47]),
     .sp4_h_l_09(net3920[0:47]), .sp4_h_l_10(net3919[0:47]),
     .sp4_h_r_10(net3427[0:47]), .sp4_h_r_09(net3428[0:47]),
     .sp4_h_r_08(net3429[0:47]), .sp4_h_r_07(net3430[0:47]),
     .sp4_h_r_06(net3431[0:47]), .sp4_h_r_05(net3432[0:47]),
     .slf_op_05(net3936[0:7]), .slf_op_06(net3935[0:7]),
     .slf_op_07(net3934[0:7]), .slf_op_08(net3933[0:7]),
     .slf_op_09(net3932[0:7]), .slf_op_10(net3931[0:7]),
     .rgt_op_10(net3439[0:7]), .rgt_op_09(net3440[0:7]),
     .rgt_op_08(net3441[0:7]), .rgt_op_07(net3442[0:7]),
     .rgt_op_06(net3443[0:7]), .rgt_op_05(net3444[0:7]),
     .lft_op_10(net3111[0:7]), .lft_op_09(net3112[0:7]),
     .lft_op_08(net3113[0:7]), .lft_op_07(net3114[0:7]),
     .lft_op_06(net3115[0:7]), .lft_op_05(net3116[0:7]),
     .sp12_h_l_10(net3944[0:23]), .sp12_h_r_10(net3452[0:23]),
     .sp12_h_l_09(net3953[0:23]), .sp12_h_l_08(net3952[0:23]),
     .sp12_h_l_07(net3951[0:23]), .sp12_h_l_06(net3950[0:23]),
     .sp12_h_r_05(net3457[0:23]), .sp12_h_r_06(net3458[0:23]),
     .sp12_h_r_07(net3459[0:23]), .sp12_h_r_08(net3460[0:23]),
     .sp12_h_r_09(net3461[0:23]), .sp12_h_l_05(net3949[0:23]),
     .sp4_r_v_b_05(net3463[0:47]), .sp4_r_v_b_06(net3464[0:47]),
     .sp4_r_v_b_07(net3465[0:47]), .sp4_r_v_b_08(net3466[0:47]),
     .sp4_r_v_b_09(net3467[0:47]), .sp4_r_v_b_10(net3468[0:47]),
     .sp4_v_b_10(net3960[0:47]), .sp4_v_b_09(net3959[0:47]),
     .sp4_v_b_08(net3958[0:47]), .sp4_v_b_07(net3957[0:47]),
     .sp4_v_b_06(net3956[0:47]), .sp4_v_b_05(net3955[0:47]),
     .sp4_v_t_16(net3475[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net3478[0:47]),
     .sp4_h_r_12(net3479[0:47]), .sp4_h_r_13(net3480[0:47]),
     .sp4_h_r_14(net3481[0:47]), .sp4_h_r_15(net3482[0:47]),
     .sp4_h_r_16(net3483[0:47]), .sp4_h_l_16(net3975[0:47]),
     .sp4_h_l_15(net3974[0:47]), .sp4_h_l_14(net3973[0:47]),
     .sp4_h_l_13(net3972[0:47]), .sp4_h_l_12(net3971[0:47]),
     .sp4_h_l_11(net3970[0:47]), .tnr_op_16({slf_op_25_00[3],
     slf_op_25_00[2], slf_op_25_00[1], slf_op_25_00[0],
     slf_op_25_00[3], slf_op_25_00[2], slf_op_25_00[1],
     slf_op_25_00[0]}), .tnl_op_16({slf_op_23_33[3], slf_op_23_33[2],
     slf_op_23_33[1], slf_op_23_33[0], slf_op_23_33[3],
     slf_op_23_33[2], slf_op_23_33[1], slf_op_23_33[0]}),
     .lft_op_16(net3043[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net3992[0:7]), .slf_op_14(net3991[0:7]),
     .slf_op_13(net3994[0:7]), .slf_op_12(net3993[0:7]),
     .slf_op_11(net3995[0:7]), .rgt_op_14(net3499[0:7]),
     .rgt_op_15(net3500[0:7]), .rgt_op_12(net3501[0:7]),
     .rgt_op_13(net3502[0:7]), .rgt_op_11(net3503[0:7]),
     .sp4_v_b_16(net4002[0:47]), .sp4_v_b_14(net4005[0:47]),
     .sp4_v_b_15(net4003[0:47]), .sp4_v_b_13(net4004[0:47]),
     .sp4_v_b_11(net4007[0:47]), .sp4_v_b_12(net4006[0:47]),
     .sp4_r_v_b_16(net3510[0:47]), .sp4_r_v_b_15(net3511[0:47]),
     .sp4_r_v_b_13(net3512[0:47]), .sp4_r_v_b_14(net3513[0:47]),
     .sp4_r_v_b_12(net3514[0:47]), .sp4_r_v_b_11(net3515[0:47]),
     .sp12_h_l_16(net4014[0:23]), .sp12_h_l_15(net4016[0:23]),
     .sp12_h_l_14(net4015[0:23]), .sp12_h_l_13(net4018[0:23]),
     .sp12_h_l_12(net4017[0:23]), .sp12_h_l_11(net4019[0:23]),
     .sp12_h_r_16(net3522[0:23]), .sp12_h_r_14(net3523[0:23]),
     .sp12_h_r_15(net3524[0:23]), .sp12_h_r_12(net3525[0:23]),
     .sp12_h_r_13(net3526[0:23]), .sp12_h_r_11(net3527[0:23]),
     .lft_op_14(net3171[0:7]), .lft_op_15(net3172[0:7]),
     .lft_op_12(net3173[0:7]), .lft_op_11(net3175[0:7]),
     .lft_op_13(net3174[0:7]));
array_LT1x16top I_it_31_top ( .glb_netwk(net3533[0:7]),
     .sp12_v_t_16(net3534[0:23]), .rgt_op_16(net3535[0:7]),
     .top_op_16({slf_op_31_33[3], slf_op_31_33[2], slf_op_31_33[1],
     slf_op_31_33[0], slf_op_31_33[3], slf_op_31_33[2],
     slf_op_31_33[1], slf_op_31_33[0]}), .rgt_op_03(net3537[0:7]),
     .slf_op_02(net4031[0:7]), .rgt_op_02(net3539[0:7]),
     .rgt_op_01(slf_op_32_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3711[0:7]), .lft_op_03(net3701[0:7]),
     .lft_op_02(net3703[0:7]), .lft_op_01(slf_op_30_17[7:0]),
     .rgt_op_04(net3547[0:7]), .carry_in(carry_in_31_17),
     .bnl_op_01(bnl_op_31_17[7:0]), .slf_op_04(net4039[0:7]),
     .slf_op_03(net4029[0:7]), .slf_op_01(slf_op_31_17[7:0]),
     .sp4_h_l_04(net4060[0:47]), .carry_out(net3554),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_31_17[23:0]),
     .sp12_h_r_04(net3557[0:23]), .sp12_h_r_03(net3558[0:23]),
     .sp12_h_r_02(net3559[0:23]), .sp12_h_r_01(net3560[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net4027[0:7]),
     .sp4_v_b_01(sp4_v_b_31_17[47:0]), .sp4_r_v_b_04(net3564[0:47]),
     .sp4_r_v_b_03(net3565[0:47]), .sp4_r_v_b_02(net3566[0:47]),
     .sp4_r_v_b_01(sp4_v_b_32_17[47:0]), .sp4_h_r_04(net3568[0:47]),
     .sp4_h_r_03(net3569[0:47]), .sp4_h_r_02(net3570[0:47]),
     .sp4_h_r_01(net3571[0:47]), .sp4_h_l_03(net4061[0:47]),
     .sp4_h_l_02(net4062[0:47]), .sp4_h_l_01(net4063[0:47]),
     .bl(bl[1671:1618]), .bot_op_01(bot_op_31_17[7:0]),
     .sp12_h_l_01(net4052[0:23]), .sp12_h_l_02(net4051[0:23]),
     .sp12_h_l_03(net4050[0:23]), .sp12_h_l_04(net4049[0:23]),
     .sp4_v_b_04(net4056[0:47]), .sp4_v_b_03(net4057[0:47]),
     .sp4_v_b_02(net4058[0:47]), .bnr_op_01(bnr_op_31_17[7:0]),
     .sp4_h_l_05(net4088[0:47]), .sp4_h_l_06(net4087[0:47]),
     .sp4_h_l_07(net4086[0:47]), .sp4_h_l_08(net4085[0:47]),
     .sp4_h_l_09(net4084[0:47]), .sp4_h_l_10(net4083[0:47]),
     .sp4_h_r_10(net3591[0:47]), .sp4_h_r_09(net3592[0:47]),
     .sp4_h_r_08(net3593[0:47]), .sp4_h_r_07(net3594[0:47]),
     .sp4_h_r_06(net3595[0:47]), .sp4_h_r_05(net3596[0:47]),
     .slf_op_05(net4100[0:7]), .slf_op_06(net4099[0:7]),
     .slf_op_07(net4098[0:7]), .slf_op_08(net4097[0:7]),
     .slf_op_09(net4096[0:7]), .slf_op_10(net4095[0:7]),
     .rgt_op_10(net3603[0:7]), .rgt_op_09(net3604[0:7]),
     .rgt_op_08(net3605[0:7]), .rgt_op_07(net3606[0:7]),
     .rgt_op_06(net3607[0:7]), .rgt_op_05(net3608[0:7]),
     .lft_op_10(net3767[0:7]), .lft_op_09(net3768[0:7]),
     .lft_op_08(net3769[0:7]), .lft_op_07(net3770[0:7]),
     .lft_op_06(net3771[0:7]), .lft_op_05(net3772[0:7]),
     .sp12_h_l_10(net4108[0:23]), .sp12_h_r_10(net3616[0:23]),
     .sp12_h_l_09(net4117[0:23]), .sp12_h_l_08(net4116[0:23]),
     .sp12_h_l_07(net4115[0:23]), .sp12_h_l_06(net4114[0:23]),
     .sp12_h_r_05(net3621[0:23]), .sp12_h_r_06(net3622[0:23]),
     .sp12_h_r_07(net3623[0:23]), .sp12_h_r_08(net3624[0:23]),
     .sp12_h_r_09(net3625[0:23]), .sp12_h_l_05(net4113[0:23]),
     .sp4_r_v_b_05(net3627[0:47]), .sp4_r_v_b_06(net3628[0:47]),
     .sp4_r_v_b_07(net3629[0:47]), .sp4_r_v_b_08(net3630[0:47]),
     .sp4_r_v_b_09(net3631[0:47]), .sp4_r_v_b_10(net3632[0:47]),
     .sp4_v_b_10(net4124[0:47]), .sp4_v_b_09(net4123[0:47]),
     .sp4_v_b_08(net4122[0:47]), .sp4_v_b_07(net4121[0:47]),
     .sp4_v_b_06(net4120[0:47]), .sp4_v_b_05(net4119[0:47]),
     .sp4_v_t_16(net3639[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net3642[0:47]),
     .sp4_h_r_12(net3643[0:47]), .sp4_h_r_13(net3644[0:47]),
     .sp4_h_r_14(net3645[0:47]), .sp4_h_r_15(net3646[0:47]),
     .sp4_h_r_16(net3647[0:47]), .sp4_h_l_16(net4139[0:47]),
     .sp4_h_l_15(net4138[0:47]), .sp4_h_l_14(net4137[0:47]),
     .sp4_h_l_13(net4136[0:47]), .sp4_h_l_12(net4135[0:47]),
     .sp4_h_l_11(net4134[0:47]), .tnr_op_16({slf_op_32_33[3],
     slf_op_32_33[2], slf_op_32_33[1], slf_op_32_33[0],
     slf_op_32_33[3], slf_op_32_33[2], slf_op_32_33[1],
     slf_op_32_33[0]}), .tnl_op_16({slf_op_30_33[3], slf_op_30_33[2],
     slf_op_30_33[1], slf_op_30_33[0], slf_op_30_33[3],
     slf_op_30_33[2], slf_op_30_33[1], slf_op_30_33[0]}),
     .lft_op_16(net3699[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net4156[0:7]), .slf_op_14(net4155[0:7]),
     .slf_op_13(net4158[0:7]), .slf_op_12(net4157[0:7]),
     .slf_op_11(net4159[0:7]), .rgt_op_14(net3663[0:7]),
     .rgt_op_15(net3664[0:7]), .rgt_op_12(net3665[0:7]),
     .rgt_op_13(net3666[0:7]), .rgt_op_11(net3667[0:7]),
     .sp4_v_b_16(net4166[0:47]), .sp4_v_b_14(net4169[0:47]),
     .sp4_v_b_15(net4167[0:47]), .sp4_v_b_13(net4168[0:47]),
     .sp4_v_b_11(net4171[0:47]), .sp4_v_b_12(net4170[0:47]),
     .sp4_r_v_b_16(net3674[0:47]), .sp4_r_v_b_15(net3675[0:47]),
     .sp4_r_v_b_13(net3676[0:47]), .sp4_r_v_b_14(net3677[0:47]),
     .sp4_r_v_b_12(net3678[0:47]), .sp4_r_v_b_11(net3679[0:47]),
     .sp12_h_l_16(net4178[0:23]), .sp12_h_l_15(net4180[0:23]),
     .sp12_h_l_14(net4179[0:23]), .sp12_h_l_13(net4182[0:23]),
     .sp12_h_l_12(net4181[0:23]), .sp12_h_l_11(net4183[0:23]),
     .sp12_h_r_16(net3686[0:23]), .sp12_h_r_14(net3687[0:23]),
     .sp12_h_r_15(net3688[0:23]), .sp12_h_r_12(net3689[0:23]),
     .sp12_h_r_13(net3690[0:23]), .sp12_h_r_11(net3691[0:23]),
     .lft_op_14(net3827[0:7]), .lft_op_15(net3828[0:7]),
     .lft_op_12(net3829[0:7]), .lft_op_11(net3831[0:7]),
     .lft_op_13(net3830[0:7]));
array_LT1x16top I_it_29_top ( .glb_netwk(net3697[0:7]),
     .sp12_v_t_16(net3698[0:23]), .rgt_op_16(net3699[0:7]),
     .top_op_16({slf_op_29_33[3], slf_op_29_33[2], slf_op_29_33[1],
     slf_op_29_33[0], slf_op_29_33[3], slf_op_29_33[2],
     slf_op_29_33[1], slf_op_29_33[0]}), .rgt_op_03(net3701[0:7]),
     .slf_op_02(net2555[0:7]), .rgt_op_02(net3703[0:7]),
     .rgt_op_01(slf_op_30_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2727[0:7]), .lft_op_03(net2717[0:7]),
     .lft_op_02(net2719[0:7]), .lft_op_01(slf_op_28_17[7:0]),
     .rgt_op_04(net3711[0:7]), .carry_in(carry_in_29_17),
     .bnl_op_01(bnl_op_29_17[7:0]), .slf_op_04(net2563[0:7]),
     .slf_op_03(net2553[0:7]), .slf_op_01(slf_op_29_17[7:0]),
     .sp4_h_l_04(net2584[0:47]), .carry_out(net3718),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_29_17[23:0]),
     .sp12_h_r_04(net3721[0:23]), .sp12_h_r_03(net3722[0:23]),
     .sp12_h_r_02(net3723[0:23]), .sp12_h_r_01(net3724[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2551[0:7]),
     .sp4_v_b_01(sp4_v_b_29_17[47:0]), .sp4_r_v_b_04(net3728[0:47]),
     .sp4_r_v_b_03(net3729[0:47]), .sp4_r_v_b_02(net3730[0:47]),
     .sp4_r_v_b_01(sp4_v_b_30_17[47:0]), .sp4_h_r_04(net3732[0:47]),
     .sp4_h_r_03(net3733[0:47]), .sp4_h_r_02(net3734[0:47]),
     .sp4_h_r_01(net3735[0:47]), .sp4_h_l_03(net2585[0:47]),
     .sp4_h_l_02(net2586[0:47]), .sp4_h_l_01(net2587[0:47]),
     .bl(bl[1563:1510]), .bot_op_01(bot_op_29_17[7:0]),
     .sp12_h_l_01(net2576[0:23]), .sp12_h_l_02(net2575[0:23]),
     .sp12_h_l_03(net2574[0:23]), .sp12_h_l_04(net2573[0:23]),
     .sp4_v_b_04(net2580[0:47]), .sp4_v_b_03(net2581[0:47]),
     .sp4_v_b_02(net2582[0:47]), .bnr_op_01(bnr_op_29_17[7:0]),
     .sp4_h_l_05(net2612[0:47]), .sp4_h_l_06(net2611[0:47]),
     .sp4_h_l_07(net2610[0:47]), .sp4_h_l_08(net2609[0:47]),
     .sp4_h_l_09(net2608[0:47]), .sp4_h_l_10(net2607[0:47]),
     .sp4_h_r_10(net3755[0:47]), .sp4_h_r_09(net3756[0:47]),
     .sp4_h_r_08(net3757[0:47]), .sp4_h_r_07(net3758[0:47]),
     .sp4_h_r_06(net3759[0:47]), .sp4_h_r_05(net3760[0:47]),
     .slf_op_05(net2624[0:7]), .slf_op_06(net2623[0:7]),
     .slf_op_07(net2622[0:7]), .slf_op_08(net2621[0:7]),
     .slf_op_09(net2620[0:7]), .slf_op_10(net2619[0:7]),
     .rgt_op_10(net3767[0:7]), .rgt_op_09(net3768[0:7]),
     .rgt_op_08(net3769[0:7]), .rgt_op_07(net3770[0:7]),
     .rgt_op_06(net3771[0:7]), .rgt_op_05(net3772[0:7]),
     .lft_op_10(net2783[0:7]), .lft_op_09(net2784[0:7]),
     .lft_op_08(net2785[0:7]), .lft_op_07(net2786[0:7]),
     .lft_op_06(net2787[0:7]), .lft_op_05(net2788[0:7]),
     .sp12_h_l_10(net2632[0:23]), .sp12_h_r_10(net3780[0:23]),
     .sp12_h_l_09(net2641[0:23]), .sp12_h_l_08(net2640[0:23]),
     .sp12_h_l_07(net2639[0:23]), .sp12_h_l_06(net2638[0:23]),
     .sp12_h_r_05(net3785[0:23]), .sp12_h_r_06(net3786[0:23]),
     .sp12_h_r_07(net3787[0:23]), .sp12_h_r_08(net3788[0:23]),
     .sp12_h_r_09(net3789[0:23]), .sp12_h_l_05(net2637[0:23]),
     .sp4_r_v_b_05(net3791[0:47]), .sp4_r_v_b_06(net3792[0:47]),
     .sp4_r_v_b_07(net3793[0:47]), .sp4_r_v_b_08(net3794[0:47]),
     .sp4_r_v_b_09(net3795[0:47]), .sp4_r_v_b_10(net3796[0:47]),
     .sp4_v_b_10(net2648[0:47]), .sp4_v_b_09(net2647[0:47]),
     .sp4_v_b_08(net2646[0:47]), .sp4_v_b_07(net2645[0:47]),
     .sp4_v_b_06(net2644[0:47]), .sp4_v_b_05(net2643[0:47]),
     .sp4_v_t_16(net3803[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net3806[0:47]),
     .sp4_h_r_12(net3807[0:47]), .sp4_h_r_13(net3808[0:47]),
     .sp4_h_r_14(net3809[0:47]), .sp4_h_r_15(net3810[0:47]),
     .sp4_h_r_16(net3811[0:47]), .sp4_h_l_16(net2663[0:47]),
     .sp4_h_l_15(net2662[0:47]), .sp4_h_l_14(net2661[0:47]),
     .sp4_h_l_13(net2660[0:47]), .sp4_h_l_12(net2659[0:47]),
     .sp4_h_l_11(net2658[0:47]), .tnr_op_16({slf_op_30_33[3],
     slf_op_30_33[2], slf_op_30_33[1], slf_op_30_33[0],
     slf_op_30_33[3], slf_op_30_33[2], slf_op_30_33[1],
     slf_op_30_33[0]}), .tnl_op_16({slf_op_28_33[3], slf_op_28_33[2],
     slf_op_28_33[1], slf_op_28_33[0], slf_op_28_33[3],
     slf_op_28_33[2], slf_op_28_33[1], slf_op_28_33[0]}),
     .lft_op_16(net2715[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net2680[0:7]), .slf_op_14(net2679[0:7]),
     .slf_op_13(net2682[0:7]), .slf_op_12(net2681[0:7]),
     .slf_op_11(net2683[0:7]), .rgt_op_14(net3827[0:7]),
     .rgt_op_15(net3828[0:7]), .rgt_op_12(net3829[0:7]),
     .rgt_op_13(net3830[0:7]), .rgt_op_11(net3831[0:7]),
     .sp4_v_b_16(net2690[0:47]), .sp4_v_b_14(net2693[0:47]),
     .sp4_v_b_15(net2691[0:47]), .sp4_v_b_13(net2692[0:47]),
     .sp4_v_b_11(net2695[0:47]), .sp4_v_b_12(net2694[0:47]),
     .sp4_r_v_b_16(net3838[0:47]), .sp4_r_v_b_15(net3839[0:47]),
     .sp4_r_v_b_13(net3840[0:47]), .sp4_r_v_b_14(net3841[0:47]),
     .sp4_r_v_b_12(net3842[0:47]), .sp4_r_v_b_11(net3843[0:47]),
     .sp12_h_l_16(net2702[0:23]), .sp12_h_l_15(net2704[0:23]),
     .sp12_h_l_14(net2703[0:23]), .sp12_h_l_13(net2706[0:23]),
     .sp12_h_l_12(net2705[0:23]), .sp12_h_l_11(net2707[0:23]),
     .sp12_h_r_16(net3850[0:23]), .sp12_h_r_14(net3851[0:23]),
     .sp12_h_r_15(net3852[0:23]), .sp12_h_r_12(net3853[0:23]),
     .sp12_h_r_13(net3854[0:23]), .sp12_h_r_11(net3855[0:23]),
     .lft_op_14(net2843[0:7]), .lft_op_15(net2844[0:7]),
     .lft_op_12(net2845[0:7]), .lft_op_11(net2847[0:7]),
     .lft_op_13(net2846[0:7]));
array_LT1x16top I_it_23_top ( .glb_netwk(net3861[0:7]),
     .sp12_v_t_16(net3862[0:23]), .rgt_op_16(net3863[0:7]),
     .top_op_16({slf_op_23_33[3], slf_op_23_33[2], slf_op_23_33[1],
     slf_op_23_33[0], slf_op_23_33[3], slf_op_23_33[2],
     slf_op_23_33[1], slf_op_23_33[0]}), .rgt_op_03(net3865[0:7]),
     .slf_op_02(net3047[0:7]), .rgt_op_02(net3867[0:7]),
     .rgt_op_01(slf_op_24_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2399[0:7]), .lft_op_03(net2389[0:7]),
     .lft_op_02(net2391[0:7]), .lft_op_01(slf_op_22_17[7:0]),
     .rgt_op_04(net3875[0:7]), .carry_in(carry_in_23_17),
     .bnl_op_01(bnl_op_23_17[7:0]), .slf_op_04(net3055[0:7]),
     .slf_op_03(net3045[0:7]), .slf_op_01(slf_op_23_17[7:0]),
     .sp4_h_l_04(net3076[0:47]), .carry_out(net3882),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_23_17[23:0]),
     .sp12_h_r_04(net3885[0:23]), .sp12_h_r_03(net3886[0:23]),
     .sp12_h_r_02(net3887[0:23]), .sp12_h_r_01(net3888[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net3043[0:7]),
     .sp4_v_b_01(sp4_v_b_23_17[47:0]), .sp4_r_v_b_04(net3892[0:47]),
     .sp4_r_v_b_03(net3893[0:47]), .sp4_r_v_b_02(net3894[0:47]),
     .sp4_r_v_b_01(sp4_v_b_24_17[47:0]), .sp4_h_r_04(net3896[0:47]),
     .sp4_h_r_03(net3897[0:47]), .sp4_h_r_02(net3898[0:47]),
     .sp4_h_r_01(net3899[0:47]), .sp4_h_l_03(net3077[0:47]),
     .sp4_h_l_02(net3078[0:47]), .sp4_h_l_01(net3079[0:47]),
     .bl(bl[1251:1198]), .bot_op_01(bot_op_23_17[7:0]),
     .sp12_h_l_01(net3068[0:23]), .sp12_h_l_02(net3067[0:23]),
     .sp12_h_l_03(net3066[0:23]), .sp12_h_l_04(net3065[0:23]),
     .sp4_v_b_04(net3072[0:47]), .sp4_v_b_03(net3073[0:47]),
     .sp4_v_b_02(net3074[0:47]), .bnr_op_01(bnr_op_23_17[7:0]),
     .sp4_h_l_05(net3104[0:47]), .sp4_h_l_06(net3103[0:47]),
     .sp4_h_l_07(net3102[0:47]), .sp4_h_l_08(net3101[0:47]),
     .sp4_h_l_09(net3100[0:47]), .sp4_h_l_10(net3099[0:47]),
     .sp4_h_r_10(net3919[0:47]), .sp4_h_r_09(net3920[0:47]),
     .sp4_h_r_08(net3921[0:47]), .sp4_h_r_07(net3922[0:47]),
     .sp4_h_r_06(net3923[0:47]), .sp4_h_r_05(net3924[0:47]),
     .slf_op_05(net3116[0:7]), .slf_op_06(net3115[0:7]),
     .slf_op_07(net3114[0:7]), .slf_op_08(net3113[0:7]),
     .slf_op_09(net3112[0:7]), .slf_op_10(net3111[0:7]),
     .rgt_op_10(net3931[0:7]), .rgt_op_09(net3932[0:7]),
     .rgt_op_08(net3933[0:7]), .rgt_op_07(net3934[0:7]),
     .rgt_op_06(net3935[0:7]), .rgt_op_05(net3936[0:7]),
     .lft_op_10(net2455[0:7]), .lft_op_09(net2456[0:7]),
     .lft_op_08(net2457[0:7]), .lft_op_07(net2458[0:7]),
     .lft_op_06(net2459[0:7]), .lft_op_05(net2460[0:7]),
     .sp12_h_l_10(net3124[0:23]), .sp12_h_r_10(net3944[0:23]),
     .sp12_h_l_09(net3133[0:23]), .sp12_h_l_08(net3132[0:23]),
     .sp12_h_l_07(net3131[0:23]), .sp12_h_l_06(net3130[0:23]),
     .sp12_h_r_05(net3949[0:23]), .sp12_h_r_06(net3950[0:23]),
     .sp12_h_r_07(net3951[0:23]), .sp12_h_r_08(net3952[0:23]),
     .sp12_h_r_09(net3953[0:23]), .sp12_h_l_05(net3129[0:23]),
     .sp4_r_v_b_05(net3955[0:47]), .sp4_r_v_b_06(net3956[0:47]),
     .sp4_r_v_b_07(net3957[0:47]), .sp4_r_v_b_08(net3958[0:47]),
     .sp4_r_v_b_09(net3959[0:47]), .sp4_r_v_b_10(net3960[0:47]),
     .sp4_v_b_10(net3140[0:47]), .sp4_v_b_09(net3139[0:47]),
     .sp4_v_b_08(net3138[0:47]), .sp4_v_b_07(net3137[0:47]),
     .sp4_v_b_06(net3136[0:47]), .sp4_v_b_05(net3135[0:47]),
     .sp4_v_t_16(net3967[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net3970[0:47]),
     .sp4_h_r_12(net3971[0:47]), .sp4_h_r_13(net3972[0:47]),
     .sp4_h_r_14(net3973[0:47]), .sp4_h_r_15(net3974[0:47]),
     .sp4_h_r_16(net3975[0:47]), .sp4_h_l_16(net3155[0:47]),
     .sp4_h_l_15(net3154[0:47]), .sp4_h_l_14(net3153[0:47]),
     .sp4_h_l_13(net3152[0:47]), .sp4_h_l_12(net3151[0:47]),
     .sp4_h_l_11(net3150[0:47]), .tnr_op_16({slf_op_24_33[3],
     slf_op_24_33[2], slf_op_24_33[1], slf_op_24_33[0],
     slf_op_24_33[3], slf_op_24_33[2], slf_op_24_33[1],
     slf_op_24_33[0]}), .tnl_op_16({slf_op_22_33[3], slf_op_22_33[2],
     slf_op_22_33[1], slf_op_22_33[0], slf_op_22_33[3],
     slf_op_22_33[2], slf_op_22_33[1], slf_op_22_33[0]}),
     .lft_op_16(net2387[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net3172[0:7]), .slf_op_14(net3171[0:7]),
     .slf_op_13(net3174[0:7]), .slf_op_12(net3173[0:7]),
     .slf_op_11(net3175[0:7]), .rgt_op_14(net3991[0:7]),
     .rgt_op_15(net3992[0:7]), .rgt_op_12(net3993[0:7]),
     .rgt_op_13(net3994[0:7]), .rgt_op_11(net3995[0:7]),
     .sp4_v_b_16(net3182[0:47]), .sp4_v_b_14(net3185[0:47]),
     .sp4_v_b_15(net3183[0:47]), .sp4_v_b_13(net3184[0:47]),
     .sp4_v_b_11(net3187[0:47]), .sp4_v_b_12(net3186[0:47]),
     .sp4_r_v_b_16(net4002[0:47]), .sp4_r_v_b_15(net4003[0:47]),
     .sp4_r_v_b_13(net4004[0:47]), .sp4_r_v_b_14(net4005[0:47]),
     .sp4_r_v_b_12(net4006[0:47]), .sp4_r_v_b_11(net4007[0:47]),
     .sp12_h_l_16(net3194[0:23]), .sp12_h_l_15(net3196[0:23]),
     .sp12_h_l_14(net3195[0:23]), .sp12_h_l_13(net3198[0:23]),
     .sp12_h_l_12(net3197[0:23]), .sp12_h_l_11(net3199[0:23]),
     .sp12_h_r_16(net4014[0:23]), .sp12_h_r_14(net4015[0:23]),
     .sp12_h_r_15(net4016[0:23]), .sp12_h_r_12(net4017[0:23]),
     .sp12_h_r_13(net4018[0:23]), .sp12_h_r_11(net4019[0:23]),
     .lft_op_14(net2515[0:7]), .lft_op_15(net2516[0:7]),
     .lft_op_12(net2517[0:7]), .lft_op_11(net2519[0:7]),
     .lft_op_13(net2518[0:7]));
array_LT1x16top I_it_30_top ( .glb_netwk(net4025[0:7]),
     .sp12_v_t_16(net4026[0:23]), .rgt_op_16(net4027[0:7]),
     .top_op_16({slf_op_30_33[3], slf_op_30_33[2], slf_op_30_33[1],
     slf_op_30_33[0], slf_op_30_33[3], slf_op_30_33[2],
     slf_op_30_33[1], slf_op_30_33[0]}), .rgt_op_03(net4029[0:7]),
     .slf_op_02(net3703[0:7]), .rgt_op_02(net4031[0:7]),
     .rgt_op_01(slf_op_31_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2563[0:7]), .lft_op_03(net2553[0:7]),
     .lft_op_02(net2555[0:7]), .lft_op_01(slf_op_29_17[7:0]),
     .rgt_op_04(net4039[0:7]), .carry_in(carry_in_30_17),
     .bnl_op_01(bnl_op_30_17[7:0]), .slf_op_04(net3711[0:7]),
     .slf_op_03(net3701[0:7]), .slf_op_01(slf_op_30_17[7:0]),
     .sp4_h_l_04(net3732[0:47]), .carry_out(net4046),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_30_17[23:0]),
     .sp12_h_r_04(net4049[0:23]), .sp12_h_r_03(net4050[0:23]),
     .sp12_h_r_02(net4051[0:23]), .sp12_h_r_01(net4052[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net3699[0:7]),
     .sp4_v_b_01(sp4_v_b_30_17[47:0]), .sp4_r_v_b_04(net4056[0:47]),
     .sp4_r_v_b_03(net4057[0:47]), .sp4_r_v_b_02(net4058[0:47]),
     .sp4_r_v_b_01(sp4_v_b_31_17[47:0]), .sp4_h_r_04(net4060[0:47]),
     .sp4_h_r_03(net4061[0:47]), .sp4_h_r_02(net4062[0:47]),
     .sp4_h_r_01(net4063[0:47]), .sp4_h_l_03(net3733[0:47]),
     .sp4_h_l_02(net3734[0:47]), .sp4_h_l_01(net3735[0:47]),
     .bl(bl[1617:1564]), .bot_op_01(bot_op_30_17[7:0]),
     .sp12_h_l_01(net3724[0:23]), .sp12_h_l_02(net3723[0:23]),
     .sp12_h_l_03(net3722[0:23]), .sp12_h_l_04(net3721[0:23]),
     .sp4_v_b_04(net3728[0:47]), .sp4_v_b_03(net3729[0:47]),
     .sp4_v_b_02(net3730[0:47]), .bnr_op_01(bnr_op_30_17[7:0]),
     .sp4_h_l_05(net3760[0:47]), .sp4_h_l_06(net3759[0:47]),
     .sp4_h_l_07(net3758[0:47]), .sp4_h_l_08(net3757[0:47]),
     .sp4_h_l_09(net3756[0:47]), .sp4_h_l_10(net3755[0:47]),
     .sp4_h_r_10(net4083[0:47]), .sp4_h_r_09(net4084[0:47]),
     .sp4_h_r_08(net4085[0:47]), .sp4_h_r_07(net4086[0:47]),
     .sp4_h_r_06(net4087[0:47]), .sp4_h_r_05(net4088[0:47]),
     .slf_op_05(net3772[0:7]), .slf_op_06(net3771[0:7]),
     .slf_op_07(net3770[0:7]), .slf_op_08(net3769[0:7]),
     .slf_op_09(net3768[0:7]), .slf_op_10(net3767[0:7]),
     .rgt_op_10(net4095[0:7]), .rgt_op_09(net4096[0:7]),
     .rgt_op_08(net4097[0:7]), .rgt_op_07(net4098[0:7]),
     .rgt_op_06(net4099[0:7]), .rgt_op_05(net4100[0:7]),
     .lft_op_10(net2619[0:7]), .lft_op_09(net2620[0:7]),
     .lft_op_08(net2621[0:7]), .lft_op_07(net2622[0:7]),
     .lft_op_06(net2623[0:7]), .lft_op_05(net2624[0:7]),
     .sp12_h_l_10(net3780[0:23]), .sp12_h_r_10(net4108[0:23]),
     .sp12_h_l_09(net3789[0:23]), .sp12_h_l_08(net3788[0:23]),
     .sp12_h_l_07(net3787[0:23]), .sp12_h_l_06(net3786[0:23]),
     .sp12_h_r_05(net4113[0:23]), .sp12_h_r_06(net4114[0:23]),
     .sp12_h_r_07(net4115[0:23]), .sp12_h_r_08(net4116[0:23]),
     .sp12_h_r_09(net4117[0:23]), .sp12_h_l_05(net3785[0:23]),
     .sp4_r_v_b_05(net4119[0:47]), .sp4_r_v_b_06(net4120[0:47]),
     .sp4_r_v_b_07(net4121[0:47]), .sp4_r_v_b_08(net4122[0:47]),
     .sp4_r_v_b_09(net4123[0:47]), .sp4_r_v_b_10(net4124[0:47]),
     .sp4_v_b_10(net3796[0:47]), .sp4_v_b_09(net3795[0:47]),
     .sp4_v_b_08(net3794[0:47]), .sp4_v_b_07(net3793[0:47]),
     .sp4_v_b_06(net3792[0:47]), .sp4_v_b_05(net3791[0:47]),
     .sp4_v_t_16(net4131[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net4134[0:47]),
     .sp4_h_r_12(net4135[0:47]), .sp4_h_r_13(net4136[0:47]),
     .sp4_h_r_14(net4137[0:47]), .sp4_h_r_15(net4138[0:47]),
     .sp4_h_r_16(net4139[0:47]), .sp4_h_l_16(net3811[0:47]),
     .sp4_h_l_15(net3810[0:47]), .sp4_h_l_14(net3809[0:47]),
     .sp4_h_l_13(net3808[0:47]), .sp4_h_l_12(net3807[0:47]),
     .sp4_h_l_11(net3806[0:47]), .tnr_op_16({slf_op_31_33[3],
     slf_op_31_33[2], slf_op_31_33[1], slf_op_31_33[0],
     slf_op_31_33[3], slf_op_31_33[2], slf_op_31_33[1],
     slf_op_31_33[0]}), .tnl_op_16({slf_op_29_33[3], slf_op_29_33[2],
     slf_op_29_33[1], slf_op_29_33[0], slf_op_29_33[3],
     slf_op_29_33[2], slf_op_29_33[1], slf_op_29_33[0]}),
     .lft_op_16(net2551[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net3828[0:7]), .slf_op_14(net3827[0:7]),
     .slf_op_13(net3830[0:7]), .slf_op_12(net3829[0:7]),
     .slf_op_11(net3831[0:7]), .rgt_op_14(net4155[0:7]),
     .rgt_op_15(net4156[0:7]), .rgt_op_12(net4157[0:7]),
     .rgt_op_13(net4158[0:7]), .rgt_op_11(net4159[0:7]),
     .sp4_v_b_16(net3838[0:47]), .sp4_v_b_14(net3841[0:47]),
     .sp4_v_b_15(net3839[0:47]), .sp4_v_b_13(net3840[0:47]),
     .sp4_v_b_11(net3843[0:47]), .sp4_v_b_12(net3842[0:47]),
     .sp4_r_v_b_16(net4166[0:47]), .sp4_r_v_b_15(net4167[0:47]),
     .sp4_r_v_b_13(net4168[0:47]), .sp4_r_v_b_14(net4169[0:47]),
     .sp4_r_v_b_12(net4170[0:47]), .sp4_r_v_b_11(net4171[0:47]),
     .sp12_h_l_16(net3850[0:23]), .sp12_h_l_15(net3852[0:23]),
     .sp12_h_l_14(net3851[0:23]), .sp12_h_l_13(net3854[0:23]),
     .sp12_h_l_12(net3853[0:23]), .sp12_h_l_11(net3855[0:23]),
     .sp12_h_r_16(net4178[0:23]), .sp12_h_r_14(net4179[0:23]),
     .sp12_h_r_15(net4180[0:23]), .sp12_h_r_12(net4181[0:23]),
     .sp12_h_r_13(net4182[0:23]), .sp12_h_r_11(net4183[0:23]),
     .lft_op_14(net2679[0:7]), .lft_op_15(net2680[0:7]),
     .lft_op_12(net2681[0:7]), .lft_op_11(net2683[0:7]),
     .lft_op_13(net2682[0:7]));
array_LT1x16top I_it_26_top ( .glb_netwk(net4189[0:7]),
     .sp12_v_t_16(net4190[0:23]), .rgt_op_16(net4191[0:7]),
     .top_op_16({slf_op_26_33[3], slf_op_26_33[2], slf_op_26_33[1],
     slf_op_26_33[0], slf_op_26_33[3], slf_op_26_33[2],
     slf_op_26_33[1], slf_op_26_33[0]}), .rgt_op_03(net4193[0:7]),
     .slf_op_02(net2319[0:7]), .rgt_op_02(net4195[0:7]),
     .rgt_op_01(slf_op_27_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3383[0:7]), .lft_op_03(net3373[0:7]),
     .lft_op_02(net3375[0:7]), .lft_op_01(slf_op_25_17[7:0]),
     .rgt_op_04(net4203[0:7]), .carry_in(carry_in_26_17),
     .bnl_op_01(bnl_op_26_17[7:0]), .slf_op_04(net2321[0:7]),
     .slf_op_03(net2320[0:7]), .slf_op_01(slf_op_26_17[7:0]),
     .sp4_h_l_04(net2340[0:47]), .carry_out(net4210),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_26_17[23:0]),
     .sp12_h_r_04(net4213[0:23]), .sp12_h_r_03(net4214[0:23]),
     .sp12_h_r_02(net4215[0:23]), .sp12_h_r_01(net4216[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2359[0:7]),
     .sp4_v_b_01(sp4_v_b_26_17[47:0]), .sp4_r_v_b_04(net4220[0:47]),
     .sp4_r_v_b_03(net4221[0:47]), .sp4_r_v_b_02(net4222[0:47]),
     .sp4_r_v_b_01(sp4_v_b_27_17[47:0]), .sp4_h_r_04(net4224[0:47]),
     .sp4_h_r_03(net4225[0:47]), .sp4_h_r_02(net4226[0:47]),
     .sp4_h_r_01(net4227[0:47]), .sp4_h_l_03(net2339[0:47]),
     .sp4_h_l_02(net2338[0:47]), .sp4_h_l_01(net2337[0:47]),
     .bl(bl[1401:1348]), .bot_op_01(bot_op_26_17[7:0]),
     .sp12_h_l_01(net2217[0:23]), .sp12_h_l_02(net2297[0:23]),
     .sp12_h_l_03(net2296[0:23]), .sp12_h_l_04(net2295[0:23]),
     .sp4_v_b_04(net2234[0:47]), .sp4_v_b_03(net2233[0:47]),
     .sp4_v_b_02(net2232[0:47]), .bnr_op_01(bnr_op_26_17[7:0]),
     .sp4_h_l_05(net2341[0:47]), .sp4_h_l_06(net2342[0:47]),
     .sp4_h_l_07(net2343[0:47]), .sp4_h_l_08(net2344[0:47]),
     .sp4_h_l_09(net2229[0:47]), .sp4_h_l_10(net2345[0:47]),
     .sp4_h_r_10(net4247[0:47]), .sp4_h_r_09(net4248[0:47]),
     .sp4_h_r_08(net4249[0:47]), .sp4_h_r_07(net4250[0:47]),
     .sp4_h_r_06(net4251[0:47]), .sp4_h_r_05(net4252[0:47]),
     .slf_op_05(net2322[0:7]), .slf_op_06(net2323[0:7]),
     .slf_op_07(net2324[0:7]), .slf_op_08(net2325[0:7]),
     .slf_op_09(net2326[0:7]), .slf_op_10(net2327[0:7]),
     .rgt_op_10(net4259[0:7]), .rgt_op_09(net4260[0:7]),
     .rgt_op_08(net4261[0:7]), .rgt_op_07(net4262[0:7]),
     .rgt_op_06(net4263[0:7]), .rgt_op_05(net4264[0:7]),
     .lft_op_10(net3439[0:7]), .lft_op_09(net3440[0:7]),
     .lft_op_08(net3441[0:7]), .lft_op_07(net3442[0:7]),
     .lft_op_06(net3443[0:7]), .lft_op_05(net3444[0:7]),
     .sp12_h_l_10(net2277[0:23]), .sp12_h_r_10(net4272[0:23]),
     .sp12_h_l_09(net2290[0:23]), .sp12_h_l_08(net2291[0:23]),
     .sp12_h_l_07(net2292[0:23]), .sp12_h_l_06(net2293[0:23]),
     .sp12_h_r_05(net4277[0:23]), .sp12_h_r_06(net4278[0:23]),
     .sp12_h_r_07(net4279[0:23]), .sp12_h_r_08(net4280[0:23]),
     .sp12_h_r_09(net4281[0:23]), .sp12_h_l_05(net2294[0:23]),
     .sp4_r_v_b_05(net4283[0:47]), .sp4_r_v_b_06(net4284[0:47]),
     .sp4_r_v_b_07(net4285[0:47]), .sp4_r_v_b_08(net4286[0:47]),
     .sp4_r_v_b_09(net4287[0:47]), .sp4_r_v_b_10(net4288[0:47]),
     .sp4_v_b_10(net2240[0:47]), .sp4_v_b_09(net2239[0:47]),
     .sp4_v_b_08(net2238[0:47]), .sp4_v_b_07(net2237[0:47]),
     .sp4_v_b_06(net2236[0:47]), .sp4_v_b_05(net2235[0:47]),
     .sp4_v_t_16(net4295[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net4298[0:47]),
     .sp4_h_r_12(net4299[0:47]), .sp4_h_r_13(net4300[0:47]),
     .sp4_h_r_14(net4301[0:47]), .sp4_h_r_15(net4302[0:47]),
     .sp4_h_r_16(net4303[0:47]), .sp4_h_l_16(net2351[0:47]),
     .sp4_h_l_15(net2350[0:47]), .sp4_h_l_14(net2349[0:47]),
     .sp4_h_l_13(net2348[0:47]), .sp4_h_l_12(net2347[0:47]),
     .sp4_h_l_11(net2346[0:47]), .tnr_op_16({slf_op_27_33[3],
     slf_op_27_33[2], slf_op_27_33[1], slf_op_27_33[0],
     slf_op_27_33[3], slf_op_27_33[2], slf_op_27_33[1],
     slf_op_27_33[0]}), .tnl_op_16({slf_op_25_00[3], slf_op_25_00[2],
     slf_op_25_00[1], slf_op_25_00[0], slf_op_25_00[3],
     slf_op_25_00[2], slf_op_25_00[1], slf_op_25_00[0]}),
     .lft_op_16(net3371[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net2332[0:7]), .slf_op_14(net2331[0:7]),
     .slf_op_13(net2330[0:7]), .slf_op_12(net2329[0:7]),
     .slf_op_11(net2328[0:7]), .rgt_op_14(net4319[0:7]),
     .rgt_op_15(net4320[0:7]), .rgt_op_12(net4321[0:7]),
     .rgt_op_13(net4322[0:7]), .rgt_op_11(net4323[0:7]),
     .sp4_v_b_16(net2245[0:47]), .sp4_v_b_14(net2244[0:47]),
     .sp4_v_b_15(net2246[0:47]), .sp4_v_b_13(net2243[0:47]),
     .sp4_v_b_11(net2241[0:47]), .sp4_v_b_12(net2242[0:47]),
     .sp4_r_v_b_16(net4330[0:47]), .sp4_r_v_b_15(net4331[0:47]),
     .sp4_r_v_b_13(net4332[0:47]), .sp4_r_v_b_14(net4333[0:47]),
     .sp4_r_v_b_12(net4334[0:47]), .sp4_r_v_b_11(net4335[0:47]),
     .sp12_h_l_16(net2282[0:23]), .sp12_h_l_15(net2278[0:23]),
     .sp12_h_l_14(net2281[0:23]), .sp12_h_l_13(net2287[0:23]),
     .sp12_h_l_12(net2288[0:23]), .sp12_h_l_11(net2289[0:23]),
     .sp12_h_r_16(net4342[0:23]), .sp12_h_r_14(net4343[0:23]),
     .sp12_h_r_15(net4344[0:23]), .sp12_h_r_12(net4345[0:23]),
     .sp12_h_r_13(net4346[0:23]), .sp12_h_r_11(net4347[0:23]),
     .lft_op_14(net3499[0:7]), .lft_op_15(net3500[0:7]),
     .lft_op_12(net3501[0:7]), .lft_op_11(net3503[0:7]),
     .lft_op_13(net3502[0:7]));
array_LT1x16top I_lt_18_top ( .glb_netwk(net4353[0:7]),
     .sp12_v_t_16(net4354[0:23]), .rgt_op_16(net4355[0:7]),
     .top_op_16({slf_op_18_33[3], slf_op_18_33[2], slf_op_18_33[1],
     slf_op_18_33[0], slf_op_18_33[3], slf_op_18_33[2],
     slf_op_18_33[1], slf_op_18_33[0]}), .rgt_op_03(net4357[0:7]),
     .slf_op_02(net4523[0:7]), .rgt_op_02(net4359[0:7]),
     .rgt_op_01(slf_op_19_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(slf_op_17_20[7:0]), .lft_op_03(slf_op_17_19[7:0]),
     .lft_op_02(slf_op_17_18[7:0]), .lft_op_01(slf_op_17_17[7:0]),
     .rgt_op_04(net4367[0:7]), .carry_in(carry_in_18_17),
     .bnl_op_01(bnl_op_18_17[7:0]), .slf_op_04(net4531[0:7]),
     .slf_op_03(net4521[0:7]), .slf_op_01(slf_op_18_17[7:0]),
     .sp4_h_l_04(net4552[0:47]), .carry_out(net4374),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_18_17[23:0]),
     .sp12_h_r_04(net4377[0:23]), .sp12_h_r_03(net4378[0:23]),
     .sp12_h_r_02(net4379[0:23]), .sp12_h_r_01(net4380[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net4519[0:7]),
     .sp4_v_b_01(sp4_v_b_18_17[47:0]), .sp4_r_v_b_04(net4384[0:47]),
     .sp4_r_v_b_03(net4385[0:47]), .sp4_r_v_b_02(net4386[0:47]),
     .sp4_r_v_b_01(sp4_v_b_19_17[47:0]), .sp4_h_r_04(net4388[0:47]),
     .sp4_h_r_03(net4389[0:47]), .sp4_h_r_02(net4390[0:47]),
     .sp4_h_r_01(net4391[0:47]), .sp4_h_l_03(net4553[0:47]),
     .sp4_h_l_02(net4554[0:47]), .sp4_h_l_01(net4555[0:47]),
     .bl(bl[981:928]), .bot_op_01(bot_op_18_17[7:0]),
     .sp12_h_l_01(net4544[0:23]), .sp12_h_l_02(net4543[0:23]),
     .sp12_h_l_03(net4542[0:23]), .sp12_h_l_04(net4541[0:23]),
     .sp4_v_b_04(net4548[0:47]), .sp4_v_b_03(net4549[0:47]),
     .sp4_v_b_02(net4550[0:47]), .bnr_op_01(bnr_op_18_17[7:0]),
     .sp4_h_l_05(net4580[0:47]), .sp4_h_l_06(net4579[0:47]),
     .sp4_h_l_07(net4578[0:47]), .sp4_h_l_08(net4577[0:47]),
     .sp4_h_l_09(net4576[0:47]), .sp4_h_l_10(net4575[0:47]),
     .sp4_h_r_10(net4411[0:47]), .sp4_h_r_09(net4412[0:47]),
     .sp4_h_r_08(net4413[0:47]), .sp4_h_r_07(net4414[0:47]),
     .sp4_h_r_06(net4415[0:47]), .sp4_h_r_05(net4416[0:47]),
     .slf_op_05(net4592[0:7]), .slf_op_06(net4591[0:7]),
     .slf_op_07(net4590[0:7]), .slf_op_08(net4589[0:7]),
     .slf_op_09(net4588[0:7]), .slf_op_10(net4587[0:7]),
     .rgt_op_10(net4423[0:7]), .rgt_op_09(net4424[0:7]),
     .rgt_op_08(net4425[0:7]), .rgt_op_07(net4426[0:7]),
     .rgt_op_06(net4427[0:7]), .rgt_op_05(net4428[0:7]),
     .lft_op_10(slf_op_17_26[7:0]), .lft_op_09(slf_op_17_25[7:0]),
     .lft_op_08(slf_op_17_24[7:0]), .lft_op_07(slf_op_17_23[7:0]),
     .lft_op_06(slf_op_17_22[7:0]), .lft_op_05(slf_op_17_21[7:0]),
     .sp12_h_l_10(net4600[0:23]), .sp12_h_r_10(net4436[0:23]),
     .sp12_h_l_09(net4609[0:23]), .sp12_h_l_08(net4608[0:23]),
     .sp12_h_l_07(net4607[0:23]), .sp12_h_l_06(net4606[0:23]),
     .sp12_h_r_05(net4441[0:23]), .sp12_h_r_06(net4442[0:23]),
     .sp12_h_r_07(net4443[0:23]), .sp12_h_r_08(net4444[0:23]),
     .sp12_h_r_09(net4445[0:23]), .sp12_h_l_05(net4605[0:23]),
     .sp4_r_v_b_05(net4447[0:47]), .sp4_r_v_b_06(net4448[0:47]),
     .sp4_r_v_b_07(net4449[0:47]), .sp4_r_v_b_08(net4450[0:47]),
     .sp4_r_v_b_09(net4451[0:47]), .sp4_r_v_b_10(net4452[0:47]),
     .sp4_v_b_10(net4616[0:47]), .sp4_v_b_09(net4615[0:47]),
     .sp4_v_b_08(net4614[0:47]), .sp4_v_b_07(net4613[0:47]),
     .sp4_v_b_06(net4612[0:47]), .sp4_v_b_05(net4611[0:47]),
     .sp4_v_t_16(net4459[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net4462[0:47]),
     .sp4_h_r_12(net4463[0:47]), .sp4_h_r_13(net4464[0:47]),
     .sp4_h_r_14(net4465[0:47]), .sp4_h_r_15(net4466[0:47]),
     .sp4_h_r_16(net4467[0:47]), .sp4_h_l_16(net4631[0:47]),
     .sp4_h_l_15(net4630[0:47]), .sp4_h_l_14(net4629[0:47]),
     .sp4_h_l_13(net4628[0:47]), .sp4_h_l_12(net4627[0:47]),
     .sp4_h_l_11(net4626[0:47]), .tnr_op_16({slf_op_19_33[3],
     slf_op_19_33[2], slf_op_19_33[1], slf_op_19_33[0],
     slf_op_19_33[3], slf_op_19_33[2], slf_op_19_33[1],
     slf_op_19_33[0]}), .tnl_op_16({slf_op_17_33[3], slf_op_17_33[2],
     slf_op_17_33[1], slf_op_17_33[0], slf_op_17_33[3],
     slf_op_17_33[2], slf_op_17_33[1], slf_op_17_33[0]}),
     .lft_op_16(slf_op_17_32[7:0]), .wl(wl_r[255:0]),
     .slf_op_15(net4648[0:7]), .slf_op_14(net4647[0:7]),
     .slf_op_13(net4650[0:7]), .slf_op_12(net4649[0:7]),
     .slf_op_11(net4651[0:7]), .rgt_op_14(net4483[0:7]),
     .rgt_op_15(net4484[0:7]), .rgt_op_12(net4485[0:7]),
     .rgt_op_13(net4486[0:7]), .rgt_op_11(net4487[0:7]),
     .sp4_v_b_16(net4658[0:47]), .sp4_v_b_14(net4661[0:47]),
     .sp4_v_b_15(net4659[0:47]), .sp4_v_b_13(net4660[0:47]),
     .sp4_v_b_11(net4663[0:47]), .sp4_v_b_12(net4662[0:47]),
     .sp4_r_v_b_16(net4494[0:47]), .sp4_r_v_b_15(net4495[0:47]),
     .sp4_r_v_b_13(net4496[0:47]), .sp4_r_v_b_14(net4497[0:47]),
     .sp4_r_v_b_12(net4498[0:47]), .sp4_r_v_b_11(net4499[0:47]),
     .sp12_h_l_16(net4670[0:23]), .sp12_h_l_15(net4672[0:23]),
     .sp12_h_l_14(net4671[0:23]), .sp12_h_l_13(net4674[0:23]),
     .sp12_h_l_12(net4673[0:23]), .sp12_h_l_11(net4675[0:23]),
     .sp12_h_r_16(net4506[0:23]), .sp12_h_r_14(net4507[0:23]),
     .sp12_h_r_15(net4508[0:23]), .sp12_h_r_12(net4509[0:23]),
     .sp12_h_r_13(net4510[0:23]), .sp12_h_r_11(net4511[0:23]),
     .lft_op_14(slf_op_17_30[7:0]), .lft_op_15(slf_op_17_31[7:0]),
     .lft_op_12(slf_op_17_28[7:0]), .lft_op_11(slf_op_17_27[7:0]),
     .lft_op_13(slf_op_17_29[7:0]));
array_LT1x16top I_lt_17_top ( .glb_netwk(net4517[0:7]),
     .sp12_v_t_16(net4518[0:23]), .rgt_op_16(net4519[0:7]),
     .top_op_16({slf_op_17_33[3], slf_op_17_33[2], slf_op_17_33[1],
     slf_op_17_33[0], slf_op_17_33[3], slf_op_17_33[2],
     slf_op_17_33[1], slf_op_17_33[0]}), .rgt_op_03(net4521[0:7]),
     .slf_op_02(slf_op_17_18[7:0]), .rgt_op_02(net4523[0:7]),
     .rgt_op_01(slf_op_18_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(lft_op_17_20[7:0]), .lft_op_03(lft_op_17_19[7:0]),
     .lft_op_02(lft_op_17_18[7:0]), .lft_op_01(lft_op_17_17[7:0]),
     .rgt_op_04(net4531[0:7]), .carry_in(carry_in_17_17),
     .bnl_op_01(bnl_op_17_17[7:0]), .slf_op_04(slf_op_17_20[7:0]),
     .slf_op_03(slf_op_17_19[7:0]), .slf_op_01(slf_op_17_17[7:0]),
     .sp4_h_l_04(sp4_h_l_17_20[47:0]), .carry_out(net4538),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_17_17[23:0]),
     .sp12_h_r_04(net4541[0:23]), .sp12_h_r_03(net4542[0:23]),
     .sp12_h_r_02(net4543[0:23]), .sp12_h_r_01(net4544[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(slf_op_17_32[7:0]),
     .sp4_v_b_01(sp4_v_b_17_17[47:0]), .sp4_r_v_b_04(net4548[0:47]),
     .sp4_r_v_b_03(net4549[0:47]), .sp4_r_v_b_02(net4550[0:47]),
     .sp4_r_v_b_01(sp4_v_b_18_17[47:0]), .sp4_h_r_04(net4552[0:47]),
     .sp4_h_r_03(net4553[0:47]), .sp4_h_r_02(net4554[0:47]),
     .sp4_h_r_01(net4555[0:47]), .sp4_h_l_03(sp4_h_l_17_19[47:0]),
     .sp4_h_l_02(sp4_h_l_17_18[47:0]),
     .sp4_h_l_01(sp4_h_l_17_17[47:0]), .bl(bl[927:874]),
     .bot_op_01(bot_op_17_17[7:0]), .sp12_h_l_01(sp12_h_l_17_17[23:0]),
     .sp12_h_l_02(sp12_h_l_17_18[23:0]),
     .sp12_h_l_03(sp12_h_l_17_19[23:0]),
     .sp12_h_l_04(sp12_h_l_17_20[23:0]),
     .sp4_v_b_04(sp4_v_b_17_20[47:0]),
     .sp4_v_b_03(sp4_v_b_17_19[47:0]),
     .sp4_v_b_02(sp4_v_b_17_18[47:0]), .bnr_op_01(bnr_op_17_17[7:0]),
     .sp4_h_l_05(sp4_h_l_17_21[47:0]),
     .sp4_h_l_06(sp4_h_l_17_22[47:0]),
     .sp4_h_l_07(sp4_h_l_17_23[47:0]),
     .sp4_h_l_08(sp4_h_l_17_24[47:0]),
     .sp4_h_l_09(sp4_h_l_17_25[47:0]),
     .sp4_h_l_10(sp4_h_l_17_26[47:0]), .sp4_h_r_10(net4575[0:47]),
     .sp4_h_r_09(net4576[0:47]), .sp4_h_r_08(net4577[0:47]),
     .sp4_h_r_07(net4578[0:47]), .sp4_h_r_06(net4579[0:47]),
     .sp4_h_r_05(net4580[0:47]), .slf_op_05(slf_op_17_21[7:0]),
     .slf_op_06(slf_op_17_22[7:0]), .slf_op_07(slf_op_17_23[7:0]),
     .slf_op_08(slf_op_17_24[7:0]), .slf_op_09(slf_op_17_25[7:0]),
     .slf_op_10(slf_op_17_26[7:0]), .rgt_op_10(net4587[0:7]),
     .rgt_op_09(net4588[0:7]), .rgt_op_08(net4589[0:7]),
     .rgt_op_07(net4590[0:7]), .rgt_op_06(net4591[0:7]),
     .rgt_op_05(net4592[0:7]), .lft_op_10(lft_op_17_26[7:0]),
     .lft_op_09(lft_op_17_25[7:0]), .lft_op_08(lft_op_17_24[7:0]),
     .lft_op_07(lft_op_17_23[7:0]), .lft_op_06(lft_op_17_22[7:0]),
     .lft_op_05(lft_op_17_21[7:0]), .sp12_h_l_10(sp12_h_l_17_26[23:0]),
     .sp12_h_r_10(net4600[0:23]), .sp12_h_l_09(sp12_h_l_17_25[23:0]),
     .sp12_h_l_08(sp12_h_l_17_24[23:0]),
     .sp12_h_l_07(sp12_h_l_17_23[23:0]),
     .sp12_h_l_06(sp12_h_l_17_22[23:0]), .sp12_h_r_05(net4605[0:23]),
     .sp12_h_r_06(net4606[0:23]), .sp12_h_r_07(net4607[0:23]),
     .sp12_h_r_08(net4608[0:23]), .sp12_h_r_09(net4609[0:23]),
     .sp12_h_l_05(sp12_h_l_17_21[23:0]), .sp4_r_v_b_05(net4611[0:47]),
     .sp4_r_v_b_06(net4612[0:47]), .sp4_r_v_b_07(net4613[0:47]),
     .sp4_r_v_b_08(net4614[0:47]), .sp4_r_v_b_09(net4615[0:47]),
     .sp4_r_v_b_10(net4616[0:47]), .sp4_v_b_10(sp4_v_b_17_26[47:0]),
     .sp4_v_b_09(sp4_v_b_17_25[47:0]),
     .sp4_v_b_08(sp4_v_b_17_24[47:0]),
     .sp4_v_b_07(sp4_v_b_17_23[47:0]),
     .sp4_v_b_06(sp4_v_b_17_22[47:0]),
     .sp4_v_b_05(sp4_v_b_17_21[47:0]), .sp4_v_t_16(net4623[0:47]),
     .pgate(pgate_r[255:0]), .reset_b(reset_r[255:0]),
     .sp4_h_r_11(net4626[0:47]), .sp4_h_r_12(net4627[0:47]),
     .sp4_h_r_13(net4628[0:47]), .sp4_h_r_14(net4629[0:47]),
     .sp4_h_r_15(net4630[0:47]), .sp4_h_r_16(net4631[0:47]),
     .sp4_h_l_16(sp4_h_l_17_32[47:0]),
     .sp4_h_l_15(sp4_h_l_17_31[47:0]),
     .sp4_h_l_14(sp4_h_l_17_30[47:0]),
     .sp4_h_l_13(sp4_h_l_17_29[47:0]),
     .sp4_h_l_12(sp4_h_l_17_28[47:0]),
     .sp4_h_l_11(sp4_h_l_17_27[47:0]), .tnr_op_16({slf_op_18_33[3],
     slf_op_18_33[2], slf_op_18_33[1], slf_op_18_33[0],
     slf_op_18_33[3], slf_op_18_33[2], slf_op_18_33[1],
     slf_op_18_33[0]}), .tnl_op_16({tnl_op_17_32[3], tnl_op_17_32[2],
     tnl_op_17_32[1], tnl_op_17_32[0], tnl_op_17_32[3],
     tnl_op_17_32[2], tnl_op_17_32[1], tnl_op_17_32[0]}),
     .lft_op_16(lft_op_17_32[7:0]), .wl(wl_r[255:0]),
     .slf_op_15(slf_op_17_31[7:0]), .slf_op_14(slf_op_17_30[7:0]),
     .slf_op_13(slf_op_17_29[7:0]), .slf_op_12(slf_op_17_28[7:0]),
     .slf_op_11(slf_op_17_27[7:0]), .rgt_op_14(net4647[0:7]),
     .rgt_op_15(net4648[0:7]), .rgt_op_12(net4649[0:7]),
     .rgt_op_13(net4650[0:7]), .rgt_op_11(net4651[0:7]),
     .sp4_v_b_16(sp4_v_b_17_32[47:0]),
     .sp4_v_b_14(sp4_v_b_17_30[47:0]),
     .sp4_v_b_15(sp4_v_b_17_31[47:0]),
     .sp4_v_b_13(sp4_v_b_17_29[47:0]),
     .sp4_v_b_11(sp4_v_b_17_27[47:0]),
     .sp4_v_b_12(sp4_v_b_17_28[47:0]), .sp4_r_v_b_16(net4658[0:47]),
     .sp4_r_v_b_15(net4659[0:47]), .sp4_r_v_b_13(net4660[0:47]),
     .sp4_r_v_b_14(net4661[0:47]), .sp4_r_v_b_12(net4662[0:47]),
     .sp4_r_v_b_11(net4663[0:47]), .sp12_h_l_16(sp12_h_l_17_32[23:0]),
     .sp12_h_l_15(sp12_h_l_17_31[23:0]),
     .sp12_h_l_14(sp12_h_l_17_30[23:0]),
     .sp12_h_l_13(sp12_h_l_17_29[23:0]),
     .sp12_h_l_12(sp12_h_l_17_28[23:0]),
     .sp12_h_l_11(sp12_h_l_17_27[23:0]), .sp12_h_r_16(net4670[0:23]),
     .sp12_h_r_14(net4671[0:23]), .sp12_h_r_15(net4672[0:23]),
     .sp12_h_r_12(net4673[0:23]), .sp12_h_r_13(net4674[0:23]),
     .sp12_h_r_11(net4675[0:23]), .lft_op_14(lft_op_17_30[7:0]),
     .lft_op_15(lft_op_17_31[7:0]), .lft_op_12(lft_op_17_28[7:0]),
     .lft_op_11(lft_op_17_27[7:0]), .lft_op_13(lft_op_17_29[7:0]));
array_LT1x16top I_it_20_top ( .glb_netwk(net4681[0:7]),
     .sp12_v_t_16(net4682[0:23]), .rgt_op_16(net4683[0:7]),
     .top_op_16({slf_op_20_33[3], slf_op_20_33[2], slf_op_20_33[1],
     slf_op_20_33[0], slf_op_20_33[3], slf_op_20_33[2],
     slf_op_20_33[1], slf_op_20_33[0]}), .rgt_op_03(net4685[0:7]),
     .slf_op_02(net3211[0:7]), .rgt_op_02(net4687[0:7]),
     .rgt_op_01(slf_op_21_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4367[0:7]), .lft_op_03(net4357[0:7]),
     .lft_op_02(net4359[0:7]), .lft_op_01(slf_op_19_17[7:0]),
     .rgt_op_04(net4695[0:7]), .carry_in(carry_in_20_17),
     .bnl_op_01(bnl_op_20_17[7:0]), .slf_op_04(net3219[0:7]),
     .slf_op_03(net3209[0:7]), .slf_op_01(slf_op_20_17[7:0]),
     .sp4_h_l_04(net3240[0:47]), .carry_out(net4702),
     .vdd_cntl(vdd_cntl_r[255:0]), .sp12_v_b__01(sp12_v_b_20_17[23:0]),
     .sp12_h_r_04(net4705[0:23]), .sp12_h_r_03(net4706[0:23]),
     .sp12_h_r_02(net4707[0:23]), .sp12_h_r_01(net4708[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net3207[0:7]),
     .sp4_v_b_01(sp4_v_b_20_17[47:0]), .sp4_r_v_b_04(net4712[0:47]),
     .sp4_r_v_b_03(net4713[0:47]), .sp4_r_v_b_02(net4714[0:47]),
     .sp4_r_v_b_01(sp4_v_b_21_17[47:0]), .sp4_h_r_04(net4716[0:47]),
     .sp4_h_r_03(net4717[0:47]), .sp4_h_r_02(net4718[0:47]),
     .sp4_h_r_01(net4719[0:47]), .sp4_h_l_03(net3241[0:47]),
     .sp4_h_l_02(net3242[0:47]), .sp4_h_l_01(net3243[0:47]),
     .bl(bl[1089:1036]), .bot_op_01(bot_op_20_17[7:0]),
     .sp12_h_l_01(net3232[0:23]), .sp12_h_l_02(net3231[0:23]),
     .sp12_h_l_03(net3230[0:23]), .sp12_h_l_04(net3229[0:23]),
     .sp4_v_b_04(net3236[0:47]), .sp4_v_b_03(net3237[0:47]),
     .sp4_v_b_02(net3238[0:47]), .bnr_op_01(bnr_op_20_17[7:0]),
     .sp4_h_l_05(net3268[0:47]), .sp4_h_l_06(net3267[0:47]),
     .sp4_h_l_07(net3266[0:47]), .sp4_h_l_08(net3265[0:47]),
     .sp4_h_l_09(net3264[0:47]), .sp4_h_l_10(net3263[0:47]),
     .sp4_h_r_10(net4739[0:47]), .sp4_h_r_09(net4740[0:47]),
     .sp4_h_r_08(net4741[0:47]), .sp4_h_r_07(net4742[0:47]),
     .sp4_h_r_06(net4743[0:47]), .sp4_h_r_05(net4744[0:47]),
     .slf_op_05(net3280[0:7]), .slf_op_06(net3279[0:7]),
     .slf_op_07(net3278[0:7]), .slf_op_08(net3277[0:7]),
     .slf_op_09(net3276[0:7]), .slf_op_10(net3275[0:7]),
     .rgt_op_10(net4751[0:7]), .rgt_op_09(net4752[0:7]),
     .rgt_op_08(net4753[0:7]), .rgt_op_07(net4754[0:7]),
     .rgt_op_06(net4755[0:7]), .rgt_op_05(net4756[0:7]),
     .lft_op_10(net4423[0:7]), .lft_op_09(net4424[0:7]),
     .lft_op_08(net4425[0:7]), .lft_op_07(net4426[0:7]),
     .lft_op_06(net4427[0:7]), .lft_op_05(net4428[0:7]),
     .sp12_h_l_10(net3288[0:23]), .sp12_h_r_10(net4764[0:23]),
     .sp12_h_l_09(net3297[0:23]), .sp12_h_l_08(net3296[0:23]),
     .sp12_h_l_07(net3295[0:23]), .sp12_h_l_06(net3294[0:23]),
     .sp12_h_r_05(net4769[0:23]), .sp12_h_r_06(net4770[0:23]),
     .sp12_h_r_07(net4771[0:23]), .sp12_h_r_08(net4772[0:23]),
     .sp12_h_r_09(net4773[0:23]), .sp12_h_l_05(net3293[0:23]),
     .sp4_r_v_b_05(net4775[0:47]), .sp4_r_v_b_06(net4776[0:47]),
     .sp4_r_v_b_07(net4777[0:47]), .sp4_r_v_b_08(net4778[0:47]),
     .sp4_r_v_b_09(net4779[0:47]), .sp4_r_v_b_10(net4780[0:47]),
     .sp4_v_b_10(net3304[0:47]), .sp4_v_b_09(net3303[0:47]),
     .sp4_v_b_08(net3302[0:47]), .sp4_v_b_07(net3301[0:47]),
     .sp4_v_b_06(net3300[0:47]), .sp4_v_b_05(net3299[0:47]),
     .sp4_v_t_16(net4787[0:47]), .pgate(pgate_r[255:0]),
     .reset_b(reset_r[255:0]), .sp4_h_r_11(net4790[0:47]),
     .sp4_h_r_12(net4791[0:47]), .sp4_h_r_13(net4792[0:47]),
     .sp4_h_r_14(net4793[0:47]), .sp4_h_r_15(net4794[0:47]),
     .sp4_h_r_16(net4795[0:47]), .sp4_h_l_16(net3319[0:47]),
     .sp4_h_l_15(net3318[0:47]), .sp4_h_l_14(net3317[0:47]),
     .sp4_h_l_13(net3316[0:47]), .sp4_h_l_12(net3315[0:47]),
     .sp4_h_l_11(net3314[0:47]), .tnr_op_16({slf_op_21_33[3],
     slf_op_21_33[2], slf_op_21_33[1], slf_op_21_33[0],
     slf_op_21_33[3], slf_op_21_33[2], slf_op_21_33[1],
     slf_op_21_33[0]}), .tnl_op_16({slf_op_19_33[3], slf_op_19_33[2],
     slf_op_19_33[1], slf_op_19_33[0], slf_op_19_33[3],
     slf_op_19_33[2], slf_op_19_33[1], slf_op_19_33[0]}),
     .lft_op_16(net4355[0:7]), .wl(wl_r[255:0]),
     .slf_op_15(net3336[0:7]), .slf_op_14(net3335[0:7]),
     .slf_op_13(net3338[0:7]), .slf_op_12(net3337[0:7]),
     .slf_op_11(net3339[0:7]), .rgt_op_14(net4811[0:7]),
     .rgt_op_15(net4812[0:7]), .rgt_op_12(net4813[0:7]),
     .rgt_op_13(net4814[0:7]), .rgt_op_11(net4815[0:7]),
     .sp4_v_b_16(net3346[0:47]), .sp4_v_b_14(net3349[0:47]),
     .sp4_v_b_15(net3347[0:47]), .sp4_v_b_13(net3348[0:47]),
     .sp4_v_b_11(net3351[0:47]), .sp4_v_b_12(net3350[0:47]),
     .sp4_r_v_b_16(net4822[0:47]), .sp4_r_v_b_15(net4823[0:47]),
     .sp4_r_v_b_13(net4824[0:47]), .sp4_r_v_b_14(net4825[0:47]),
     .sp4_r_v_b_12(net4826[0:47]), .sp4_r_v_b_11(net4827[0:47]),
     .sp12_h_l_16(net3358[0:23]), .sp12_h_l_15(net3360[0:23]),
     .sp12_h_l_14(net3359[0:23]), .sp12_h_l_13(net3362[0:23]),
     .sp12_h_l_12(net3361[0:23]), .sp12_h_l_11(net3363[0:23]),
     .sp12_h_r_16(net4834[0:23]), .sp12_h_r_14(net4835[0:23]),
     .sp12_h_r_15(net4836[0:23]), .sp12_h_r_12(net4837[0:23]),
     .sp12_h_r_13(net4838[0:23]), .sp12_h_r_11(net4839[0:23]),
     .lft_op_14(net4483[0:7]), .lft_op_15(net4484[0:7]),
     .lft_op_12(net4485[0:7]), .lft_op_11(net4487[0:7]),
     .lft_op_13(net4486[0:7]));
preio_top_r I_preio_top_r ( .ceb_o(ceb_o), .ceb_i(net4846),
     .sp4_h_r_32_33(net4847[0:15]), .bl_25(bl[1347:1306]),
     .tclk_i(net4849), .mode_i(net4850), .shift_i(net4851),
     .update_i(net4852), .hiz_b_i(net4853), .bs_en_i(net4854),
     .r_i(net4855), .sdi(net4856), .sp4_h_l_17_33(sp4_h_l_17_33[15:0]),
     .wl_r({wl_r[270], wl_r[271], wl_r[269], wl_r[268], wl_r[266],
     wl_r[267], wl_r[265], wl_r[264], wl_r[262], wl_r[263], wl_r[261],
     wl_r[260], wl_r[258], wl_r[259], wl_r[257], wl_r[256]}),
     .vdd_cntl_r({vdd_cntl_r[270], vdd_cntl_r[271], vdd_cntl_r[269],
     vdd_cntl_r[268], vdd_cntl_r[266], vdd_cntl_r[267],
     vdd_cntl_r[265], vdd_cntl_r[264], vdd_cntl_r[262],
     vdd_cntl_r[263], vdd_cntl_r[261], vdd_cntl_r[260],
     vdd_cntl_r[258], vdd_cntl_r[259], vdd_cntl_r[257],
     vdd_cntl_r[256]}), .tievdd(tievdd), .tiegnd(tiegnd),
     .reset_r({reset_r[270], reset_r[271], reset_r[269], reset_r[268],
     reset_r[266], reset_r[267], reset_r[265], reset_r[264],
     reset_r[262], reset_r[263], reset_r[261], reset_r[260],
     reset_r[258], reset_r[259], reset_r[257], reset_r[256]}),
     .prog(prog), .pgate_r({pgate_r[270], pgate_r[271], pgate_r[269],
     pgate_r[268], pgate_r[266], pgate_r[267], pgate_r[265],
     pgate_r[264], pgate_r[262], pgate_r[263], pgate_r[261],
     pgate_r[260], pgate_r[258], pgate_r[259], pgate_r[257],
     pgate_r[256]}), .padin_t(padin_t[59:30]), .hold_t_r(hold_t_r),
     .end_of_startup_top_r(end_of_startup_top_r[32:17]),
     .update_o(update_o), .tclk_o(tclk_o), .shift_o(shift_o),
     .sdo(sdo), .r_o(r_o), .pado_t(pado_t[59:30]),
     .padin_192(padin_192), .padeb_t(padeb_t[59:30]), .mode_o(mode_o),
     .hiz_b_o(hiz_b_o), .fabric_out_17_33(fabric_out_17_33),
     .cf_t(cf_t[383:0]), .bs_en_o(bs_en_o),
     .bnl_op_17_33(lft_op_17_32[7:0]),
     .slf_op_17_33(slf_op_17_33[3:0]), .glb_net_17(net4517[0:7]),
     .bl_17(bl[927:874]), .lft_op_17_33(slf_op_17_32[7:0]),
     .sp12_v_b_17_33(net4518[0:23]), .sp4_v_b_17_33(net4623[0:47]),
     .slf_op_18_33(slf_op_18_33[3:0]), .glb_net_18(net4353[0:7]),
     .bl_18(bl[981:928]), .lft_op_18_33(net4519[0:7]),
     .sp12_v_b_18_33(net4354[0:23]), .sp4_v_b_18_33(net4459[0:47]),
     .slf_op_19_33(slf_op_19_33[3:0]), .glb_net_19(net3205[0:7]),
     .bl_19(bl[1035:982]), .lft_op_19_33(net4355[0:7]),
     .sp12_v_b_19_33(net3206[0:23]), .sp4_v_b_19_33(net3311[0:47]),
     .slf_op_20_33(slf_op_20_33[3:0]), .glb_net_20(net4681[0:7]),
     .bl_20(bl[1089:1036]), .lft_op_20_33(net3207[0:7]),
     .sp12_v_b_20_33(net4682[0:23]), .sp4_v_b_20_33(net4787[0:47]),
     .slf_op_21_33(slf_op_21_33[3:0]), .glb_net_21(net2385[0:7]),
     .bl_21(bl[1143:1090]), .lft_op_21_33(net4683[0:7]),
     .sp12_v_b_21_33(net2386[0:23]), .sp4_v_b_21_33(net2491[0:47]),
     .slf_op_22_33(slf_op_22_33[3:0]), .glb_net_22(net3041[0:7]),
     .bl_22(bl[1197:1144]), .lft_op_22_33(net2387[0:7]),
     .sp12_v_b_22_33(net3042[0:23]), .sp4_v_b_22_33(net3147[0:47]),
     .slf_op_23_33(slf_op_23_33[3:0]), .glb_net_23(net3861[0:7]),
     .bl_23(bl[1251:1198]), .lft_op_23_33(net3043[0:7]),
     .sp12_v_b_23_33(net3862[0:23]), .sp4_v_b_23_33(net3967[0:47]),
     .slf_op_24_33(slf_op_24_33[3:0]), .glb_net_24(net3369[0:7]),
     .bl_24(bl[1305:1252]), .lft_op_24_33(net3863[0:7]),
     .sp4_v_b_24_33(net3475[0:47]), .slf_op_25_33(slf_op_25_00[3:0]),
     .glb_net_25(net2204[0:7]), .lft_op_25_33(net3371[0:7]),
     .sp4_v_b_25_33(net2354[0:47]), .slf_op_26_33(slf_op_26_33[3:0]),
     .glb_net_26(net4189[0:7]), .bl_26(bl[1401:1348]),
     .lft_op_26_33(net2359[0:7]), .sp4_v_b_26_33(net4295[0:47]),
     .sp12_v_b_26_33(net4190[0:23]), .sp12_v_b_25_33(net2358[0:23]),
     .sp12_v_b_24_33(net3370[0:23]), .slf_op_27_33(slf_op_27_33[3:0]),
     .glb_net_27(net2713[0:7]), .bl_27(bl[1455:1402]),
     .lft_op_27_33(net4191[0:7]), .sp12_v_b_27_33(net2714[0:23]),
     .sp4_v_b_27_33(net2819[0:47]), .slf_op_28_33(slf_op_28_33[3:0]),
     .glb_net_28(net2549[0:7]), .bl_28(bl[1509:1456]),
     .lft_op_28_33(net2715[0:7]), .sp12_v_b_28_33(net2550[0:23]),
     .sp4_v_b_28_33(net2655[0:47]), .slf_op_29_33(slf_op_29_33[3:0]),
     .glb_net_29(net3697[0:7]), .bl_29(bl[1563:1510]),
     .lft_op_29_33(net2551[0:7]), .sp12_v_b_29_33(net3698[0:23]),
     .sp4_v_b_29_33(net3803[0:47]), .slf_op_30_33(slf_op_30_33[3:0]),
     .glb_net_30(net4025[0:7]), .bl_30(bl[1617:1564]),
     .lft_op_30_33(net3699[0:7]), .sp12_v_b_30_33(net4026[0:23]),
     .sp4_v_b_30_33(net4131[0:47]), .slf_op_31_33(slf_op_31_33[3:0]),
     .glb_net_31(net3533[0:7]), .bl_31(bl[1671:1618]),
     .lft_op_31_33(net4027[0:7]), .sp12_v_b_31_33(net3534[0:23]),
     .sp4_v_b_31_33(net3639[0:47]), .bnr_op_32_33({slf_op_33_32[3],
     slf_op_33_32[2], slf_op_33_32[1], slf_op_33_32[0],
     slf_op_33_32[3], slf_op_33_32[2], slf_op_33_32[1],
     slf_op_33_32[0]}), .slf_op_32_33(slf_op_32_33[3:0]),
     .glb_net_32(net2877[0:7]), .bl_32(bl[1725:1672]),
     .lft_op_32_33(net3535[0:7]), .sp12_v_b_32_33(net2878[0:23]),
     .sp4_v_b_32_33(net2983[0:47]));
bram_bufferx4 I348 ( .in(ceb_i), .out(net4846));
bram_bufferx4 I250 ( .in(hiz_b_i), .out(net4853));
bram_bufferx4 I244 ( .in(mode_i), .out(net4850));
bram_bufferx4 I245 ( .in(update_i), .out(net4852));
bram_bufferx4 I246 ( .in(shift_i), .out(net4851));
bram_bufferx4 I247 ( .in(bs_en_i), .out(net4854));
bram_bufferx4 I249 ( .in(r_i), .out(net4855));

endmodule
// Library - leafcell, Cell - preio_top_l, View - schematic
// LAST TIME SAVED: Oct 16 14:27:51 2008
// NETLIST TIME: Nov 14 16:17:19 2008
`timescale 1ns / 1ns 

module preio_top_l ( bs_en_o, ceb_o, cf_top_l, fabric_out_15_33,
     fabric_out_16_33, hiz_b_o, mode_o, padeb_t_l, padin_193, pado_t_l,
     r_o, sdo, shift_o, slf_op_01_33, slf_op_02_33, slf_op_03_33,
     slf_op_04_33, slf_op_05_33, slf_op_06_33, slf_op_07_33,
     slf_op_08_33, slf_op_09_33, slf_op_10_33, slf_op_11_33,
     slf_op_12_33, slf_op_13_33, slf_op_14_33, slf_op_15_33,
     slf_op_16_33, tclk_o, update_o, bl_01, bl_02, bl_03, bl_04, bl_05,
     bl_06, bl_07, bl_08, bl_09, bl_10, bl_11, bl_12, bl_13, bl_14,
     bl_15, bl_16, sp4_h_l_01_33, sp4_h_r_16_33, sp4_v_b_01_33,
     sp4_v_b_02_33, sp4_v_b_03_33, sp4_v_b_04_33, sp4_v_b_05_33,
     sp4_v_b_06_33, sp4_v_b_07_33, sp4_v_b_08_33, sp4_v_b_09_33,
     sp4_v_b_10_33, sp4_v_b_11_33, sp4_v_b_12_33, sp4_v_b_13_33,
     sp4_v_b_14_33, sp4_v_b_15_33, sp4_v_b_16_33, sp12_v_b_01_33,
     sp12_v_b_02_33, sp12_v_b_03_33, sp12_v_b_04_33, sp12_v_b_05_33,
     sp12_v_b_06_33, sp12_v_b_07_33, sp12_v_b_08_33, sp12_v_b_09_33,
     sp12_v_b_10_33, sp12_v_b_11_33, sp12_v_b_12_33, sp12_v_b_13_33,
     sp12_v_b_14_33, sp12_v_b_15_33, sp12_v_b_16_33, bnl_op_01_33,
     bnr_op_16_33, bs_en_i, ceb_i, end_of_startup_top_l, glb_net_01,
     glb_net_02, glb_net_03, glb_net_04, glb_net_05, glb_net_06,
     glb_net_07, glb_net_08, glb_net_09, glb_net_10, glb_net_11,
     glb_net_12, glb_net_13, glb_net_14, glb_net_15, glb_net_16,
     hiz_b_i, hold_t_l, lft_op_01_33, lft_op_02_33, lft_op_03_33,
     lft_op_04_33, lft_op_05_33, lft_op_06_33, lft_op_07_33,
     lft_op_08_33, lft_op_09_33, lft_op_10_33, lft_op_11_33,
     lft_op_12_33, lft_op_13_33, lft_op_14_33, lft_op_15_33,
     lft_op_16_33, mode_i, padin_t_l, pgate_l, prog, r_i, reset_l, sdi,
     shift_i, tclk_i, tiegnd, tievdd, update_i, vdd_cntl_l, wl_l );
output  bs_en_o, ceb_o, fabric_out_15_33, fabric_out_16_33, hiz_b_o,
     mode_o, padin_193, r_o, sdo, shift_o, tclk_o, update_o;


input  bs_en_i, ceb_i, hiz_b_i, hold_t_l, mode_i, prog, r_i, sdi,
     shift_i, tclk_i, tiegnd, tievdd, update_i;

output [3:0]  slf_op_02_33;
output [3:0]  slf_op_05_33;
output [3:0]  slf_op_06_33;
output [3:0]  slf_op_16_33;
output [3:0]  slf_op_13_33;
output [3:0]  slf_op_07_33;
output [3:0]  slf_op_03_33;
output [3:0]  slf_op_15_33;
output [3:0]  slf_op_01_33;
output [3:0]  slf_op_10_33;
output [3:0]  slf_op_12_33;
output [3:0]  slf_op_04_33;
output [3:0]  slf_op_11_33;
output [29:0]  padeb_t_l;
output [29:0]  pado_t_l;
output [383:0]  cf_top_l;
output [3:0]  slf_op_09_33;
output [3:0]  slf_op_14_33;
output [3:0]  slf_op_08_33;

inout [47:0]  sp4_v_b_02_33;
inout [47:0]  sp4_v_b_11_33;
inout [23:0]  sp12_v_b_12_33;
inout [47:0]  sp4_v_b_16_33;
inout [23:0]  sp12_v_b_16_33;
inout [23:0]  sp12_v_b_15_33;
inout [23:0]  sp12_v_b_01_33;
inout [23:0]  sp12_v_b_04_33;
inout [23:0]  sp12_v_b_14_33;
inout [47:0]  sp4_v_b_14_33;
inout [23:0]  sp12_v_b_03_33;
inout [23:0]  sp12_v_b_07_33;
inout [53:0]  bl_10;
inout [23:0]  sp12_v_b_06_33;
inout [47:0]  sp4_v_b_12_33;
inout [15:0]  sp4_h_r_16_33;
inout [47:0]  sp4_v_b_10_33;
inout [53:0]  bl_13;
inout [53:0]  bl_11;
inout [23:0]  sp12_v_b_10_33;
inout [23:0]  sp12_v_b_05_33;
inout [47:0]  sp4_v_b_15_33;
inout [53:0]  bl_06;
inout [53:0]  bl_04;
inout [53:0]  bl_02;
inout [47:0]  sp4_v_b_07_33;
inout [47:0]  sp4_v_b_05_33;
inout [47:0]  sp4_v_b_13_33;
inout [23:0]  sp12_v_b_09_33;
inout [23:0]  sp12_v_b_08_33;
inout [53:0]  bl_07;
inout [47:0]  sp4_v_b_01_33;
inout [53:0]  bl_12;
inout [23:0]  sp12_v_b_11_33;
inout [47:0]  sp4_v_b_09_33;
inout [47:0]  sp4_v_b_03_33;
inout [53:0]  bl_15;
inout [53:0]  bl_03;
inout [47:0]  sp4_v_b_06_33;
inout [15:0]  sp4_h_l_01_33;
inout [23:0]  sp12_v_b_13_33;
inout [53:0]  bl_16;
inout [23:0]  sp12_v_b_02_33;
inout [53:0]  bl_05;
inout [47:0]  sp4_v_b_04_33;
inout [53:0]  bl_09;
inout [53:0]  bl_14;
inout [53:0]  bl_01;
inout [41:0]  bl_08;
inout [47:0]  sp4_v_b_08_33;

input [15:0]  vdd_cntl_l;
input [7:0]  glb_net_10;
input [7:0]  lft_op_06_33;
input [7:0]  glb_net_07;
input [7:0]  lft_op_14_33;
input [15:0]  reset_l;
input [7:0]  glb_net_13;
input [7:0]  lft_op_02_33;
input [7:0]  lft_op_10_33;
input [7:0]  lft_op_08_33;
input [7:0]  glb_net_16;
input [7:0]  lft_op_05_33;
input [7:0]  lft_op_16_33;
input [15:0]  pgate_l;
input [7:0]  lft_op_03_33;
input [7:0]  lft_op_01_33;
input [7:0]  glb_net_01;
input [7:0]  glb_net_08;
input [7:0]  bnr_op_16_33;
input [7:0]  lft_op_13_33;
input [7:0]  glb_net_12;
input [7:0]  glb_net_11;
input [7:0]  lft_op_15_33;
input [7:0]  lft_op_12_33;
input [7:0]  glb_net_14;
input [7:0]  glb_net_04;
input [7:0]  glb_net_05;
input [7:0]  lft_op_04_33;
input [7:0]  glb_net_02;
input [7:0]  lft_op_09_33;
input [15:0]  wl_l;
input [16:1]  end_of_startup_top_l;
input [29:0]  padin_t_l;
input [7:0]  lft_op_07_33;
input [7:0]  lft_op_11_33;
input [7:0]  glb_net_09;
input [7:0]  glb_net_15;
input [7:0]  glb_net_06;
input [7:0]  bnl_op_01_33;
input [7:0]  glb_net_03;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:15]  net1134;

wire  [0:15]  net854;

wire  [0:1]  net1188;

wire  [0:15]  net924;

wire  [0:15]  net714;

wire  [0:15]  net644;

wire  [0:1]  net1193;

wire  [0:1]  net1190;

wire  [0:15]  net994;

wire  [0:15]  net1064;

wire  [0:1]  net735;

wire  [0:15]  net679;

wire  [0:1]  net1203;

wire  [0:1]  net1205;

wire  [0:1]  net910;

wire  [0:1]  net801;

wire  [0:15]  net784;

wire  [0:15]  net959;

wire  [0:15]  net819;

wire  [0:1]  net1155;

wire  [0:1]  net1207;

wire  [0:1]  net1195;

wire  [0:1]  net1201;

wire  [0:1]  net1204;

wire  [0:1]  net1206;

wire  [0:1]  net1212;

wire  [0:1]  net805;

wire  [0:15]  net889;

wire  [0:1]  net1185;

wire  [0:15]  net1029;

wire  [0:15]  net1099;

wire  [0:1]  net799;

wire  [0:15]  net749;



lowla_modified I330 ( .clk(tclk_i), .min(net0599), .lao(net1138));
bram_bufferx4x6 I333 ( .in(sdi), .out(net0599));
tckbufx16 I257 ( .in(tclk_i), .out(tclk_o));
fabric_buf8k I332 ( .f_in(net817), .f_out(fabric_out_15_33));
fabric_buf8k I331 ( .f_in(net1167), .f_out(fabric_out_16_33));
fabric_buf8k I328 ( .f_in(padin_t_l[29]), .f_out(padin_193));
io_col4_BRAM_TOP I_IO_08_33bram ( .ceb(ceb_o), .bl({bl_08[5], bl_08[4],
     bl_08[37], bl_08[36], bl_08[35], bl_08[34], bl_08[33], bl_08[32],
     bl_08[14], bl_08[20], bl_08[19], bl_08[18], bl_08[17], bl_08[16],
     bl_08[27], bl_08[26], bl_08[25], bl_08[23]}), .sdo(net858),
     .sdi(net613), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[8]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[15:14]), .pado(pado_t_l[15:14]),
     .padeb(padeb_t_l[15:14]), .sp4_h_l(sp4_v_b_08_33[47:0]),
     .sp12_h_l(sp12_v_b_08_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1204[0:1]), .tnl_op(lft_op_07_33[7:0]),
     .lft_op(lft_op_08_33[7:0]), .bnl_op(lft_op_09_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[191:168]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_08_33[3:0]), .glb_netwk(glb_net_08[7:0]),
     .hold(hold_t_l), .fabric_out(net1196), .sp4_v_t(net889[0:15]),
     .sp4_v_b(net644[0:15]));
io_col4_TOP I_IO_02_33 ( .ceb(ceb_o), .bl({bl_02[5], bl_02[4],
     bl_02[37], bl_02[36], bl_02[35], bl_02[34], bl_02[33], bl_02[32],
     bl_02[14], bl_02[20], bl_02[19], bl_02[18], bl_02[17], bl_02[16],
     bl_02[27], bl_02[26], bl_02[25], bl_02[23]}), .sdo(net718),
     .sdi(net648), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[2]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[3:2]), .pado(pado_t_l[3:2]),
     .padeb(padeb_t_l[3:2]), .sp4_h_l(sp4_v_b_02_33[47:0]),
     .sp12_h_l(sp12_v_b_02_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1195[0:1]), .tnl_op(lft_op_01_33[7:0]),
     .lft_op(lft_op_02_33[7:0]), .bnl_op(lft_op_03_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[47:24]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_02_33[3:0]), .glb_netwk(glb_net_02[7:0]),
     .hold(hold_t_l), .fabric_out(net1208), .sp4_v_t(net749[0:15]),
     .sp4_v_b(net679[0:15]));
io_col4_TOP I_IO_11_33 ( .ceb(ceb_o), .bl({bl_11[5], bl_11[4],
     bl_11[37], bl_11[36], bl_11[35], bl_11[34], bl_11[33], bl_11[32],
     bl_11[14], bl_11[20], bl_11[19], bl_11[18], bl_11[17], bl_11[16],
     bl_11[27], bl_11[26], bl_11[25], bl_11[23]}), .sdo(net753),
     .sdi(net683), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[11]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[21:20]), .pado(pado_t_l[21:20]),
     .padeb(padeb_t_l[21:20]), .sp4_h_l(sp4_v_b_11_33[47:0]),
     .sp12_h_l(sp12_v_b_11_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1205[0:1]), .tnl_op(lft_op_10_33[7:0]),
     .lft_op(lft_op_11_33[7:0]), .bnl_op(lft_op_12_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[263:240]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_11_33[3:0]), .glb_netwk(glb_net_11[7:0]),
     .hold(hold_t_l), .fabric_out(net1209), .sp4_v_t(net784[0:15]),
     .sp4_v_b(net714[0:15]));
io_col4_TOP I_IO_01_33 ( .ceb(ceb_o), .bl({bl_01[5], bl_01[4],
     bl_01[37], bl_01[36], bl_01[35], bl_01[34], bl_01[33], bl_01[32],
     bl_01[14], bl_01[20], bl_01[19], bl_01[18], bl_01[17], bl_01[16],
     bl_01[27], bl_01[26], bl_01[25], bl_01[23]}), .sdo(sdo),
     .sdi(net718), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[1]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[1:0]), .pado(pado_t_l[1:0]),
     .padeb(padeb_t_l[1:0]), .sp4_h_l(sp4_v_b_01_33[47:0]),
     .sp12_h_l(sp12_v_b_01_33[23:0]), .prog(prog),
     .spi_ss_in_b(net735[0:1]), .tnl_op(bnl_op_01_33[7:0]),
     .lft_op(lft_op_01_33[7:0]), .bnl_op(lft_op_02_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[23:0]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_01_33[3:0]), .glb_netwk(glb_net_01[7:0]),
     .hold(hold_t_l), .fabric_out(net747),
     .sp4_v_t(sp4_h_l_01_33[15:0]), .sp4_v_b(net749[0:15]));
io_col4_TOP I_IO_10_33 ( .ceb(ceb_o), .bl({bl_10[5], bl_10[4],
     bl_10[37], bl_10[36], bl_10[35], bl_10[34], bl_10[33], bl_10[32],
     bl_10[14], bl_10[20], bl_10[19], bl_10[18], bl_10[17], bl_10[16],
     bl_10[27], bl_10[26], bl_10[25], bl_10[23]}), .sdo(net1103),
     .sdi(net753), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[10]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[19:18]), .pado(pado_t_l[19:18]),
     .padeb(padeb_t_l[19:18]), .sp4_h_l(sp4_v_b_10_33[47:0]),
     .sp12_h_l(sp12_v_b_10_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1201[0:1]), .tnl_op(lft_op_09_33[7:0]),
     .lft_op(lft_op_10_33[7:0]), .bnl_op(lft_op_11_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[239:216]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_10_33[3:0]), .glb_netwk(glb_net_10[7:0]),
     .hold(hold_t_l), .fabric_out(net1191), .sp4_v_t(net1134[0:15]),
     .sp4_v_b(net784[0:15]));
io_col4_TOP I_IO_15_33 ( .ceb(ceb_o), .bl({bl_15[5], bl_15[4],
     bl_15[37], bl_15[36], bl_15[35], bl_15[34], bl_15[33], bl_15[32],
     bl_15[14], bl_15[20], bl_15[19], bl_15[18], bl_15[17], bl_15[16],
     bl_15[27], bl_15[26], bl_15[25], bl_15[23]}), .sdo(net1033),
     .sdi(net788), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[15]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(net799[0:1]), .pado(net799[0:1]), .padeb(net801[0:1]),
     .sp4_h_l(sp4_v_b_15_33[47:0]), .sp12_h_l(sp12_v_b_15_33[23:0]),
     .prog(prog), .spi_ss_in_b(net805[0:1]),
     .tnl_op(lft_op_14_33[7:0]), .lft_op(lft_op_15_33[7:0]),
     .bnl_op(lft_op_16_33[7:0]), .pgate(pgate_l[15:0]),
     .reset(reset_l[15:0]), .wl(wl_l[15:0]), .cf(cf_top_l[359:336]),
     .vdd_cntl(vdd_cntl_l[15:0]), .slf_op(slf_op_15_33[3:0]),
     .glb_netwk(glb_net_15[7:0]), .hold(hold_t_l), .fabric_out(net817),
     .sp4_v_t(net1064[0:15]), .sp4_v_b(net819[0:15]));
io_col4_TOP I_IO_05_33 ( .ceb(ceb_o), .bl({bl_05[5], bl_05[4],
     bl_05[37], bl_05[36], bl_05[35], bl_05[34], bl_05[33], bl_05[32],
     bl_05[14], bl_05[20], bl_05[19], bl_05[18], bl_05[17], bl_05[16],
     bl_05[27], bl_05[26], bl_05[25], bl_05[23]}), .sdo(net1068),
     .sdi(net823), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[5]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[9:8]), .pado(pado_t_l[9:8]),
     .padeb(padeb_t_l[9:8]), .sp4_h_l(sp4_v_b_05_33[47:0]),
     .sp12_h_l(sp12_v_b_05_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1207[0:1]), .tnl_op(lft_op_04_33[7:0]),
     .lft_op(lft_op_05_33[7:0]), .bnl_op(lft_op_06_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[119:96]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_05_33[3:0]), .glb_netwk(glb_net_05[7:0]),
     .hold(hold_t_l), .fabric_out(net852), .sp4_v_t(net1099[0:15]),
     .sp4_v_b(net854[0:15]));
io_col4_TOP I_IO_07_33 ( .ceb(ceb_o), .bl({bl_07[5], bl_07[4],
     bl_07[37], bl_07[36], bl_07[35], bl_07[34], bl_07[33], bl_07[32],
     bl_07[14], bl_07[20], bl_07[19], bl_07[18], bl_07[17], bl_07[16],
     bl_07[27], bl_07[26], bl_07[25], bl_07[23]}), .sdo(net893),
     .sdi(net858), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[7]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[13:12]), .pado(pado_t_l[13:12]),
     .padeb(padeb_t_l[13:12]), .sp4_h_l(sp4_v_b_07_33[47:0]),
     .sp12_h_l(sp12_v_b_07_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1190[0:1]), .tnl_op(lft_op_06_33[7:0]),
     .lft_op(lft_op_07_33[7:0]), .bnl_op(lft_op_08_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[167:144]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_07_33[3:0]), .glb_netwk(glb_net_07[7:0]),
     .hold(hold_t_l), .fabric_out(net887), .sp4_v_t(net924[0:15]),
     .sp4_v_b(net889[0:15]));
io_col4_TOP I_IO_06_33 ( .ceb(ceb_o), .bl({bl_06[5], bl_06[4],
     bl_06[37], bl_06[36], bl_06[35], bl_06[34], bl_06[33], bl_06[32],
     bl_06[14], bl_06[20], bl_06[19], bl_06[18], bl_06[17], bl_06[16],
     bl_06[27], bl_06[26], bl_06[25], bl_06[23]}), .sdo(net823),
     .sdi(net893), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[6]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[11:10]), .pado(pado_t_l[11:10]),
     .padeb(padeb_t_l[11:10]), .sp4_h_l(sp4_v_b_06_33[47:0]),
     .sp12_h_l(sp12_v_b_06_33[23:0]), .prog(prog),
     .spi_ss_in_b(net910[0:1]), .tnl_op(lft_op_05_33[7:0]),
     .lft_op(lft_op_06_33[7:0]), .bnl_op(lft_op_07_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[143:120]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_06_33[3:0]), .glb_netwk(glb_net_06[7:0]),
     .hold(hold_t_l), .fabric_out(net922), .sp4_v_t(net854[0:15]),
     .sp4_v_b(net924[0:15]));
io_col4_TOP I_IO_03_33 ( .ceb(ceb_o), .bl({bl_03[5], bl_03[4],
     bl_03[37], bl_03[36], bl_03[35], bl_03[34], bl_03[33], bl_03[32],
     bl_03[14], bl_03[20], bl_03[19], bl_03[18], bl_03[17], bl_03[16],
     bl_03[27], bl_03[26], bl_03[25], bl_03[23]}), .sdo(net648),
     .sdi(net928), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[3]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[5:4]), .pado(pado_t_l[5:4]),
     .padeb(padeb_t_l[5:4]), .sp4_h_l(sp4_v_b_03_33[47:0]),
     .sp12_h_l(sp12_v_b_03_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1203[0:1]), .tnl_op(lft_op_02_33[7:0]),
     .lft_op(lft_op_03_33[7:0]), .bnl_op(lft_op_04_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[71:48]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_03_33[3:0]), .glb_netwk(glb_net_03[7:0]),
     .hold(hold_t_l), .fabric_out(net1199), .sp4_v_t(net679[0:15]),
     .sp4_v_b(net959[0:15]));
io_col4_TOP I_IO_13_33 ( .ceb(ceb_o), .bl({bl_13[5], bl_13[4],
     bl_13[37], bl_13[36], bl_13[35], bl_13[34], bl_13[33], bl_13[32],
     bl_13[14], bl_13[20], bl_13[19], bl_13[18], bl_13[17], bl_13[16],
     bl_13[27], bl_13[26], bl_13[25], bl_13[23]}), .sdo(net998),
     .sdi(net963), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[13]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[25:24]), .pado(pado_t_l[25:24]),
     .padeb(padeb_t_l[25:24]), .sp4_h_l(sp4_v_b_13_33[47:0]),
     .sp12_h_l(sp12_v_b_13_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1212[0:1]), .tnl_op(lft_op_12_33[7:0]),
     .lft_op(lft_op_13_33[7:0]), .bnl_op(lft_op_14_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[311:288]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_13_33[3:0]), .glb_netwk(glb_net_13[7:0]),
     .hold(hold_t_l), .fabric_out(net1211), .sp4_v_t(net1029[0:15]),
     .sp4_v_b(net994[0:15]));
io_col4_TOP I_IO_12_33 ( .ceb(ceb_o), .bl({bl_12[5], bl_12[4],
     bl_12[37], bl_12[36], bl_12[35], bl_12[34], bl_12[33], bl_12[32],
     bl_12[14], bl_12[20], bl_12[19], bl_12[18], bl_12[17], bl_12[16],
     bl_12[27], bl_12[26], bl_12[25], bl_12[23]}), .sdo(net683),
     .sdi(net998), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[12]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[23:22]), .pado(pado_t_l[23:22]),
     .padeb(padeb_t_l[23:22]), .sp4_h_l(sp4_v_b_12_33[47:0]),
     .sp12_h_l(sp12_v_b_12_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1206[0:1]), .tnl_op(lft_op_11_33[7:0]),
     .lft_op(lft_op_12_33[7:0]), .bnl_op(lft_op_13_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[287:264]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_12_33[3:0]), .glb_netwk(glb_net_12[7:0]),
     .hold(hold_t_l), .fabric_out(net1214), .sp4_v_t(net714[0:15]),
     .sp4_v_b(net1029[0:15]));
io_col4_TOP I_IO_14_33 ( .ceb(ceb_o), .bl({bl_14[5], bl_14[4],
     bl_14[37], bl_14[36], bl_14[35], bl_14[34], bl_14[33], bl_14[32],
     bl_14[14], bl_14[20], bl_14[19], bl_14[18], bl_14[17], bl_14[16],
     bl_14[27], bl_14[26], bl_14[25], bl_14[23]}), .sdo(net963),
     .sdi(net1033), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[14]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[27:26]), .pado(pado_t_l[27:26]),
     .padeb(padeb_t_l[27:26]), .sp4_h_l(sp4_v_b_14_33[47:0]),
     .sp12_h_l(sp12_v_b_14_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1185[0:1]), .tnl_op(lft_op_13_33[7:0]),
     .lft_op(lft_op_14_33[7:0]), .bnl_op(lft_op_15_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[335:312]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_14_33[3:0]), .glb_netwk(glb_net_14[7:0]),
     .hold(hold_t_l), .fabric_out(net1213), .sp4_v_t(net994[0:15]),
     .sp4_v_b(net1064[0:15]));
io_col4_TOP I_IO_04_33 ( .ceb(ceb_o), .bl({bl_04[5], bl_04[4],
     bl_04[37], bl_04[36], bl_04[35], bl_04[34], bl_04[33], bl_04[32],
     bl_04[14], bl_04[20], bl_04[19], bl_04[18], bl_04[17], bl_04[16],
     bl_04[27], bl_04[26], bl_04[25], bl_04[23]}), .sdo(net928),
     .sdi(net1068), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[4]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[7:6]), .pado(pado_t_l[7:6]),
     .padeb(padeb_t_l[7:6]), .sp4_h_l(sp4_v_b_04_33[47:0]),
     .sp12_h_l(sp12_v_b_04_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1193[0:1]), .tnl_op(lft_op_03_33[7:0]),
     .lft_op(lft_op_04_33[7:0]), .bnl_op(lft_op_05_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[95:72]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_04_33[3:0]), .glb_netwk(glb_net_04[7:0]),
     .hold(hold_t_l), .fabric_out(net1194), .sp4_v_t(net959[0:15]),
     .sp4_v_b(net1099[0:15]));
io_col4_TOP I_IO_09_33 ( .ceb(ceb_o), .bl({bl_09[5], bl_09[4],
     bl_09[37], bl_09[36], bl_09[35], bl_09[34], bl_09[33], bl_09[32],
     bl_09[14], bl_09[20], bl_09[19], bl_09[18], bl_09[17], bl_09[16],
     bl_09[27], bl_09[26], bl_09[25], bl_09[23]}), .sdo(net613),
     .sdi(net1103), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[9]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[17:16]), .pado(pado_t_l[17:16]),
     .padeb(padeb_t_l[17:16]), .sp4_h_l(sp4_v_b_09_33[47:0]),
     .sp12_h_l(sp12_v_b_09_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1188[0:1]), .tnl_op(lft_op_08_33[7:0]),
     .lft_op(lft_op_09_33[7:0]), .bnl_op(lft_op_10_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[215:192]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_09_33[3:0]), .glb_netwk(glb_net_09[7:0]),
     .hold(hold_t_l), .fabric_out(net1202), .sp4_v_t(net644[0:15]),
     .sp4_v_b(net1134[0:15]));
io_col4_TOP I_IO_16_33 ( .ceb(ceb_o), .bl({bl_16[5], bl_16[4],
     bl_16[37], bl_16[36], bl_16[35], bl_16[34], bl_16[33], bl_16[32],
     bl_16[14], bl_16[20], bl_16[19], bl_16[18], bl_16[17], bl_16[16],
     bl_16[27], bl_16[26], bl_16[25], bl_16[23]}), .sdo(net788),
     .sdi(net1138), .spiout({tiegnd, tiegnd}),
     .cdone_in(end_of_startup_top_l[16]), .spioeb({tievdd, tievdd}),
     .mode(mode_o), .shift(shift_o), .hiz_b(hiz_b_o), .r(r_o),
     .bs_en(bs_en_o), .tclk(tclk_o), .update(update_o),
     .padin(padin_t_l[29:28]), .pado(pado_t_l[29:28]),
     .padeb(padeb_t_l[29:28]), .sp4_h_l(sp4_v_b_16_33[47:0]),
     .sp12_h_l(sp12_v_b_16_33[23:0]), .prog(prog),
     .spi_ss_in_b(net1155[0:1]), .tnl_op(lft_op_15_33[7:0]),
     .lft_op(lft_op_16_33[7:0]), .bnl_op(bnr_op_16_33[7:0]),
     .pgate(pgate_l[15:0]), .reset(reset_l[15:0]), .wl(wl_l[15:0]),
     .cf(cf_top_l[383:360]), .vdd_cntl(vdd_cntl_l[15:0]),
     .slf_op(slf_op_16_33[3:0]), .glb_netwk(glb_net_16[7:0]),
     .hold(hold_t_l), .fabric_out(net1167), .sp4_v_t(net819[0:15]),
     .sp4_v_b(sp4_h_r_16_33[15:0]));
bram_bufferx4 I329 ( .in(ceb_i), .out(ceb_o));
bram_bufferx4 I251 ( .in(r_i), .out(r_o));
bram_bufferx4 I253 ( .in(hiz_b_i), .out(hiz_b_o));
bram_bufferx4 I256 ( .in(shift_i), .out(shift_o));
bram_bufferx4 I255 ( .in(update_i), .out(update_o));
bram_bufferx4 I252 ( .in(bs_en_i), .out(bs_en_o));
bram_bufferx4 I254 ( .in(mode_i), .out(mode_o));

endmodule
// Library - leafcell, Cell - array_LFT_IO_1x16top, View - schematic
// LAST TIME SAVED: Feb  4 15:29:08 2008
// NETLIST TIME: Nov 14 16:17:19 2008
`timescale 1ns / 1ns 

module array_LFT_IO_1x16top ( cf_l, fabric_out_17, fabric_out_18,
     fabric_out_19, fabric_out_20, fabric_out_21, fabric_out_22,
     fabric_out_23, fabric_out_24, fabric_out_25, fabric_out_26,
     fabric_out_27, fabric_out_28, fabric_out_29, fabric_out_30,
     fabric_out_31, fabric_out_32, padeb, pado, sdo, slf_op_00_17,
     slf_op_00_18, slf_op_00_19, slf_op_00_20, slf_op_00_21,
     slf_op_00_22, slf_op_00_23, slf_op_00_24, slf_op_00_25,
     slf_op_00_26, slf_op_00_27, slf_op_00_28, slf_op_00_29,
     slf_op_00_30, slf_op_00_31, slf_op_00_32, spi_ss_in_b,
     SP4_h_l_00_17, SP4_h_l_00_18, SP4_h_l_00_19, SP4_h_l_00_20,
     SP4_h_l_00_21, SP4_h_l_00_22, SP4_h_l_00_23, SP4_h_l_00_24,
     SP4_h_l_00_25, SP4_h_l_00_26, SP4_h_l_00_27, SP4_h_l_00_28,
     SP4_h_l_00_29, SP4_h_l_00_30, SP4_h_l_00_31, SP4_h_l_00_32,
     SP12_h_l_00_17, SP12_h_l_00_18, SP12_h_l_00_19, SP12_h_l_00_20,
     SP12_h_l_00_21, SP12_h_l_00_22, SP12_h_l_00_23, SP12_h_l_00_24,
     SP12_h_l_00_25, SP12_h_l_00_26, SP12_h_l_00_27, SP12_h_l_00_28,
     SP12_h_l_00_29, SP12_h_l_00_30, SP12_h_l_00_31, SP12_h_l_00_32,
     bl, pgate, reset_b, sp4_v_b_00_17, sp4_v_t_00_32, vdd_cntl, wl,
     bnl_op_00_17, bs_en, cdone_in, ceb, glb_netwk_col, hiz_b, hold,
     mode, padin, prog, r, rgt_op_00_17, rgt_op_00_18, rgt_op_00_19,
     rgt_op_00_20, rgt_op_00_21, rgt_op_00_22, rgt_op_00_23,
     rgt_op_00_24, rgt_op_00_25, rgt_op_00_26, rgt_op_00_27,
     rgt_op_00_28, rgt_op_00_29, rgt_op_00_30, rgt_op_00_31,
     rgt_op_00_32, sdi, shift, spioeb, spiout, tclk, tnl_op_00_32,
     update );
output  fabric_out_17, fabric_out_18, fabric_out_19, fabric_out_20,
     fabric_out_21, fabric_out_22, fabric_out_23, fabric_out_24,
     fabric_out_25, fabric_out_26, fabric_out_27, fabric_out_28,
     fabric_out_29, fabric_out_30, fabric_out_31, fabric_out_32, sdo;


input  bs_en, ceb, hiz_b, hold, mode, prog, r, sdi, shift, tclk,
     update;

output [3:0]  slf_op_00_26;
output [3:0]  slf_op_00_18;
output [3:0]  slf_op_00_25;
output [3:0]  slf_op_00_21;
output [3:0]  slf_op_00_27;
output [3:0]  slf_op_00_28;
output [3:0]  slf_op_00_23;
output [3:0]  slf_op_00_30;
output [49:24]  padeb;
output [31:0]  spi_ss_in_b;
output [3:0]  slf_op_00_17;
output [3:0]  slf_op_00_22;
output [3:0]  slf_op_00_31;
output [3:0]  slf_op_00_29;
output [3:0]  slf_op_00_24;
output [3:0]  slf_op_00_20;
output [383:0]  cf_l;
output [3:0]  slf_op_00_32;
output [3:0]  slf_op_00_19;
output [49:24]  pado;

inout [23:0]  SP12_h_l_00_30;
inout [47:0]  SP4_h_l_00_19;
inout [23:0]  SP12_h_l_00_31;
inout [23:0]  SP12_h_l_00_27;
inout [23:0]  SP12_h_l_00_28;
inout [47:0]  SP4_h_l_00_17;
inout [47:0]  SP4_h_l_00_20;
inout [23:0]  SP12_h_l_00_26;
inout [23:0]  SP12_h_l_00_32;
inout [47:0]  SP4_h_l_00_24;
inout [47:0]  SP4_h_l_00_25;
inout [47:0]  SP4_h_l_00_21;
inout [23:0]  SP12_h_l_00_29;
inout [23:0]  SP12_h_l_00_24;
inout [47:0]  SP4_h_l_00_22;
inout [47:0]  SP4_h_l_00_18;
inout [23:0]  SP12_h_l_00_21;
inout [47:0]  SP4_h_l_00_27;
inout [15:0]  sp4_v_b_00_17;
inout [23:0]  SP12_h_l_00_18;
inout [47:0]  SP4_h_l_00_23;
inout [47:0]  SP4_h_l_00_32;
inout [23:0]  SP12_h_l_00_20;
inout [17:0]  bl;
inout [23:0]  SP12_h_l_00_22;
inout [47:0]  SP4_h_l_00_28;
inout [23:0]  SP12_h_l_00_25;
inout [47:0]  SP4_h_l_00_26;
inout [47:0]  SP4_h_l_00_30;
inout [23:0]  SP12_h_l_00_19;
inout [47:0]  SP4_h_l_00_31;
inout [15:0]  sp4_v_t_00_32;
inout [271:16]  pgate;
inout [271:16]  vdd_cntl;
inout [271:16]  reset_b;
inout [23:0]  SP12_h_l_00_23;
inout [23:0]  SP12_h_l_00_17;
inout [271:16]  wl;
inout [47:0]  SP4_h_l_00_29;

input [7:0]  rgt_op_00_21;
input [7:0]  rgt_op_00_25;
input [7:0]  rgt_op_00_18;
input [7:0]  rgt_op_00_19;
input [7:0]  rgt_op_00_24;
input [7:0]  rgt_op_00_32;
input [7:0]  tnl_op_00_32;
input [7:0]  rgt_op_00_31;
input [7:0]  rgt_op_00_17;
input [32:17]  cdone_in;
input [31:0]  spiout;
input [7:0]  rgt_op_00_26;
input [7:0]  bnl_op_00_17;
input [49:24]  padin;
input [31:0]  spioeb;
input [7:0]  rgt_op_00_29;
input [7:0]  rgt_op_00_28;
input [7:0]  rgt_op_00_30;
input [7:0]  rgt_op_00_27;
input [7:0]  rgt_op_00_22;
input [7:0]  rgt_op_00_20;
input [7:0]  glb_netwk_col;
input [7:0]  rgt_op_00_23;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net892;

wire  [0:15]  net690;

wire  [0:1]  net1131;

wire  [0:15]  net860;

wire  [0:15]  net1098;

wire  [0:15]  net1132;

wire  [0:15]  net656;

wire  [0:1]  net1130;

wire  [0:15]  net758;

wire  [0:15]  net928;

wire  [0:1]  net1187;

wire  [0:15]  net1030;

wire  [0:15]  net1166;

wire  [0:15]  net792;

wire  [0:15]  net724;

wire  [0:1]  net824;

wire  [0:15]  net826;

wire  [0:1]  net825;

wire  [0:15]  net996;

wire  [7:0]  glb_netwk;

wire  [0:15]  net1064;

wire  [0:15]  net962;



clk_colbuf8kx8 I106 ( .clko(glb_netwk[7:0]),
     .clki(glb_netwk_col[7:0]));
io_col4_LFT I_io_00_25 ( .ceb(ceb), .sdo(net676), .sdi(net642),
     .spiout(spiout[17:16]), .cdone_in(cdone_in[25]),
     .spioeb(spioeb[17:16]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[41:40]), .pado(pado[41:40]), .padeb(padeb[41:40]),
     .sp4_v_t(net656[0:15]), .spi_ss_in_b(spi_ss_in_b[17:16]),
     .reset(reset_b[159:144]), .sp4_v_b(net690[0:15]),
     .cf(cf_l[215:192]), .bl(bl[17:0]), .slf_op(slf_op_00_25[3:0]),
     .hold(hold), .fabric_out(fabric_out_25), .prog(prog),
     .lft_op(rgt_op_00_25[7:0]), .sp12_h_l(SP12_h_l_00_25[23:0]),
     .sp4_h_l(SP4_h_l_00_25[47:0]), .wl(wl[159:144]),
     .vdd_cntl(vdd_cntl[159:144]), .glb_netwk(glb_netwk[7:0]),
     .pgate(pgate[159:144]), .bnl_op(rgt_op_00_24[7:0]),
     .tnl_op(rgt_op_00_26[7:0]));
io_col4_LFT I_io_00_24 ( .ceb(ceb), .sdo(net710), .sdi(net676),
     .spiout(spiout[15:14]), .cdone_in(cdone_in[24]),
     .spioeb(spioeb[15:14]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[39:38]), .pado(pado[39:38]), .padeb(padeb[39:38]),
     .sp4_v_t(net690[0:15]), .sp4_h_l(SP4_h_l_00_24[47:0]),
     .sp12_h_l(SP12_h_l_00_24[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[15:14]), .tnl_op(rgt_op_00_25[7:0]),
     .lft_op(rgt_op_00_24[7:0]), .bnl_op(rgt_op_00_23[7:0]),
     .pgate(pgate[143:128]), .reset(reset_b[143:128]),
     .sp4_v_b(net724[0:15]), .wl(wl[143:128]), .cf(cf_l[191:168]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[143:128]),
     .slf_op(slf_op_00_24[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_24));
io_col4_LFT I_io_00_23 ( .ceb(ceb), .sdo(net948), .sdi(net710),
     .spiout(spiout[13:12]), .cdone_in(cdone_in[23]),
     .spioeb(spioeb[13:12]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[37:36]), .pado(pado[37:36]), .padeb(padeb[37:36]),
     .sp4_v_t(net724[0:15]), .sp4_h_l(SP4_h_l_00_23[47:0]),
     .sp12_h_l(SP12_h_l_00_23[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[13:12]), .tnl_op(rgt_op_00_24[7:0]),
     .lft_op(rgt_op_00_23[7:0]), .bnl_op(rgt_op_00_22[7:0]),
     .pgate(pgate[127:112]), .reset(reset_b[127:112]),
     .sp4_v_b(net962[0:15]), .wl(wl[127:112]), .cf(cf_l[167:144]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[127:112]),
     .slf_op(slf_op_00_23[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_23));
io_col4_LFT I_io_00_31 ( .ceb(ceb), .sdo(net778), .sdi(net744),
     .spiout(spiout[29:28]), .cdone_in(cdone_in[31]),
     .spioeb(spioeb[29:28]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[49:48]), .pado(pado[49:48]), .padeb(padeb[49:48]),
     .sp4_v_t(net758[0:15]), .sp4_h_l(SP4_h_l_00_31[47:0]),
     .sp12_h_l(SP12_h_l_00_31[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[29:28]), .tnl_op(rgt_op_00_32[7:0]),
     .lft_op(rgt_op_00_31[7:0]), .bnl_op(rgt_op_00_30[7:0]),
     .pgate(pgate[255:240]), .reset(reset_b[255:240]),
     .sp4_v_b(net792[0:15]), .wl(wl[255:240]), .cf(cf_l[359:336]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[255:240]),
     .slf_op(slf_op_00_31[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_31));
io_col4_LFT I_io_00_30 ( .ceb(ceb), .sdo(net812), .sdi(net778),
     .spiout(spiout[27:26]), .cdone_in(cdone_in[30]),
     .spioeb(spioeb[27:26]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[47:46]), .pado(pado[47:46]), .padeb(padeb[47:46]),
     .sp4_v_t(net792[0:15]), .sp4_h_l(SP4_h_l_00_30[47:0]),
     .sp12_h_l(SP12_h_l_00_30[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[27:26]), .tnl_op(rgt_op_00_31[7:0]),
     .lft_op(rgt_op_00_30[7:0]), .bnl_op(rgt_op_00_29[7:0]),
     .pgate(pgate[239:224]), .reset(reset_b[239:224]),
     .sp4_v_b(net826[0:15]), .wl(wl[239:224]), .cf(cf_l[335:312]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[239:224]),
     .slf_op(slf_op_00_30[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_30));
io_col4_LFT I_io_00_29 ( .ceb(ceb), .sdo(net846), .sdi(net812),
     .spiout(spiout[25:24]), .cdone_in(cdone_in[29]),
     .spioeb(spioeb[25:24]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net824[0:1]), .pado(net824[0:1]), .padeb(net825[0:1]),
     .sp4_v_t(net826[0:15]), .sp4_h_l(SP4_h_l_00_29[47:0]),
     .sp12_h_l(SP12_h_l_00_29[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[25:24]), .tnl_op(rgt_op_00_30[7:0]),
     .lft_op(rgt_op_00_29[7:0]), .bnl_op(rgt_op_00_28[7:0]),
     .pgate(pgate[223:208]), .reset(reset_b[223:208]),
     .sp4_v_b(net860[0:15]), .wl(wl[223:208]), .cf(cf_l[311:288]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[223:208]),
     .slf_op(slf_op_00_29[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_29));
io_col4_LFT I_io_00_28 ( .ceb(ceb), .sdo(net1152), .sdi(net846),
     .spiout(spiout[23:22]), .cdone_in(cdone_in[28]),
     .spioeb(spioeb[23:22]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[45:44]), .pado(pado[45:44]), .padeb(padeb[45:44]),
     .sp4_v_t(net860[0:15]), .sp4_h_l(SP4_h_l_00_28[47:0]),
     .sp12_h_l(SP12_h_l_00_28[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[23:22]), .tnl_op(rgt_op_00_29[7:0]),
     .lft_op(rgt_op_00_28[7:0]), .bnl_op(rgt_op_00_27[7:0]),
     .pgate(pgate[207:192]), .reset(reset_b[207:192]),
     .sp4_v_b(net1166[0:15]), .wl(wl[207:192]), .cf(cf_l[287:264]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[207:192]),
     .slf_op(slf_op_00_28[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_28));
io_col4_LFT I_io_00_32 ( .ceb(ceb), .sdo(net744), .sdi(sdi),
     .spiout(spiout[31:30]), .cdone_in(cdone_in[32]),
     .spioeb(spioeb[31:30]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net892[0:1]), .pado(net892[0:1]), .padeb(net1187[0:1]),
     .sp4_v_t(sp4_v_t_00_32[15:0]), .sp4_h_l(SP4_h_l_00_32[47:0]),
     .sp12_h_l(SP12_h_l_00_32[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[31:30]), .tnl_op(tnl_op_00_32[7:0]),
     .lft_op(rgt_op_00_32[7:0]), .bnl_op(rgt_op_00_31[7:0]),
     .pgate(pgate[271:256]), .reset(reset_b[271:256]),
     .sp4_v_b(net758[0:15]), .wl(wl[271:256]), .cf(cf_l[383:360]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[271:256]),
     .slf_op(slf_op_00_32[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_32));
io_col4_LFT I_io_00_21 ( .ceb(ceb), .sdo(net1084), .sdi(net914),
     .spiout(spiout[9:8]), .cdone_in(cdone_in[21]),
     .spioeb(spioeb[9:8]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[33:32]), .pado(pado[33:32]), .padeb(padeb[33:32]),
     .sp4_v_t(net928[0:15]), .sp4_h_l(SP4_h_l_00_21[47:0]),
     .sp12_h_l(SP12_h_l_00_21[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[9:8]), .tnl_op(rgt_op_00_22[7:0]),
     .lft_op(rgt_op_00_21[7:0]), .bnl_op(rgt_op_00_20[7:0]),
     .pgate(pgate[95:80]), .reset(reset_b[95:80]),
     .sp4_v_b(net1098[0:15]), .wl(wl[95:80]), .cf(cf_l[119:96]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[95:80]),
     .slf_op(slf_op_00_21[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_21));
io_col4_LFT I_io_00_22 ( .ceb(ceb), .sdo(net914), .sdi(net948),
     .spiout(spiout[11:10]), .cdone_in(cdone_in[22]),
     .spioeb(spioeb[11:10]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[35:34]), .pado(pado[35:34]), .padeb(padeb[35:34]),
     .sp4_v_t(net962[0:15]), .sp4_h_l(SP4_h_l_00_22[47:0]),
     .sp12_h_l(SP12_h_l_00_22[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[11:10]), .tnl_op(rgt_op_00_23[7:0]),
     .lft_op(rgt_op_00_22[7:0]), .bnl_op(rgt_op_00_21[7:0]),
     .pgate(pgate[111:96]), .reset(reset_b[111:96]),
     .sp4_v_b(net928[0:15]), .wl(wl[111:96]), .cf(cf_l[143:120]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[111:96]),
     .slf_op(slf_op_00_22[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_22));
io_col4_LFT I_io_00_18 ( .ceb(ceb), .sdo(net1016), .sdi(net982),
     .spiout(spiout[3:2]), .cdone_in(cdone_in[18]),
     .spioeb(spioeb[3:2]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[27:26]), .pado(pado[27:26]), .padeb(padeb[27:26]),
     .sp4_v_t(net996[0:15]), .sp4_h_l(SP4_h_l_00_18[47:0]),
     .sp12_h_l(SP12_h_l_00_18[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[3:2]), .tnl_op(rgt_op_00_19[7:0]),
     .lft_op(rgt_op_00_18[7:0]), .bnl_op(rgt_op_00_17[7:0]),
     .pgate(pgate[47:32]), .reset(reset_b[47:32]),
     .sp4_v_b(net1030[0:15]), .wl(wl[47:32]), .cf(cf_l[47:24]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[47:32]),
     .slf_op(slf_op_00_18[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_18));
io_col4_LFT I_io_00_17 ( .ceb(ceb), .sdo(sdo), .sdi(net1016),
     .spiout(spiout[1:0]), .cdone_in(cdone_in[17]),
     .spioeb(spioeb[1:0]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[25:24]), .pado(pado[25:24]), .padeb(padeb[25:24]),
     .sp4_v_t(net1030[0:15]), .sp4_h_l(SP4_h_l_00_17[47:0]),
     .sp12_h_l(SP12_h_l_00_17[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[1:0]), .tnl_op(rgt_op_00_18[7:0]),
     .lft_op(rgt_op_00_17[7:0]), .bnl_op(bnl_op_00_17[7:0]),
     .pgate(pgate[31:16]), .reset(reset_b[31:16]),
     .sp4_v_b(sp4_v_b_00_17[15:0]), .wl(wl[31:16]), .cf(cf_l[23:0]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[31:16]),
     .slf_op(slf_op_00_17[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_17));
io_col4_LFT I_io_00_19 ( .ceb(ceb), .sdo(net982), .sdi(net1050),
     .spiout(spiout[5:4]), .cdone_in(cdone_in[19]),
     .spioeb(spioeb[5:4]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[29:28]), .pado(pado[29:28]), .padeb(padeb[29:28]),
     .sp4_v_t(net1064[0:15]), .sp4_h_l(SP4_h_l_00_19[47:0]),
     .sp12_h_l(SP12_h_l_00_19[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[5:4]), .tnl_op(rgt_op_00_20[7:0]),
     .lft_op(rgt_op_00_19[7:0]), .bnl_op(rgt_op_00_18[7:0]),
     .pgate(pgate[63:48]), .reset(reset_b[63:48]),
     .sp4_v_b(net996[0:15]), .wl(wl[63:48]), .cf(cf_l[71:48]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[63:48]),
     .slf_op(slf_op_00_19[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_19));
io_col4_LFT I_io_00_20 ( .ceb(ceb), .sdo(net1050), .sdi(net1084),
     .spiout(spiout[7:6]), .cdone_in(cdone_in[20]),
     .spioeb(spioeb[7:6]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[31:30]), .pado(pado[31:30]), .padeb(padeb[31:30]),
     .sp4_v_t(net1098[0:15]), .sp4_h_l(SP4_h_l_00_20[47:0]),
     .sp12_h_l(SP12_h_l_00_20[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[7:6]), .tnl_op(rgt_op_00_21[7:0]),
     .lft_op(rgt_op_00_20[7:0]), .bnl_op(rgt_op_00_19[7:0]),
     .pgate(pgate[79:64]), .reset(reset_b[79:64]),
     .sp4_v_b(net1064[0:15]), .wl(wl[79:64]), .cf(cf_l[95:72]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[79:64]),
     .slf_op(slf_op_00_20[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_20));
io_col4_LFT I_io_00_26 ( .ceb(ceb), .sdo(net642), .sdi(net1118),
     .spiout(spiout[19:18]), .cdone_in(cdone_in[26]),
     .spioeb(spioeb[19:18]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(net1130[0:1]), .pado(net1130[0:1]), .padeb(net1131[0:1]),
     .sp4_v_t(net1132[0:15]), .sp4_h_l(SP4_h_l_00_26[47:0]),
     .sp12_h_l(SP12_h_l_00_26[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[19:18]), .tnl_op(rgt_op_00_27[7:0]),
     .lft_op(rgt_op_00_26[7:0]), .bnl_op(rgt_op_00_25[7:0]),
     .pgate(pgate[175:160]), .reset(reset_b[175:160]),
     .sp4_v_b(net656[0:15]), .wl(wl[175:160]), .cf(cf_l[239:216]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[175:160]),
     .slf_op(slf_op_00_26[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_26));
io_col4_LFT I_io_00_27 ( .ceb(ceb), .sdo(net1118), .sdi(net1152),
     .spiout(spiout[21:20]), .cdone_in(cdone_in[27]),
     .spioeb(spioeb[21:20]), .mode(mode), .shift(shift), .hiz_b(hiz_b),
     .r(r), .bs_en(bs_en), .tclk(tclk), .update(update),
     .padin(padin[43:42]), .pado(pado[43:42]), .padeb(padeb[43:42]),
     .sp4_v_t(net1166[0:15]), .sp4_h_l(SP4_h_l_00_27[47:0]),
     .sp12_h_l(SP12_h_l_00_27[23:0]), .prog(prog),
     .spi_ss_in_b(spi_ss_in_b[21:20]), .tnl_op(rgt_op_00_28[7:0]),
     .lft_op(rgt_op_00_27[7:0]), .bnl_op(rgt_op_00_26[7:0]),
     .pgate(pgate[191:176]), .reset(reset_b[191:176]),
     .sp4_v_b(net1132[0:15]), .wl(wl[191:176]), .cf(cf_l[263:240]),
     .bl(bl[17:0]), .vdd_cntl(vdd_cntl[191:176]),
     .slf_op(slf_op_00_27[3:0]), .glb_netwk(glb_netwk[7:0]),
     .hold(hold), .fabric_out(fabric_out_27));

endmodule
// Library - leafcell, Cell - quad_tl_ice8, View - schematic
// LAST TIME SAVED: Oct 16 13:40:13 2008
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module quad_tl_ice8 ( bm_init_o, bm_rcapmux_en_o, bm_sa_o, bm_sclk_o,
     bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o, bs_en_o, ceb_o, cf_l, cf_t, fabric_out_00_17,
     fabric_out_15_33, fabric_out_16_33, hiz_b_o, mode_o, padeb_l_t,
     padeb_t_l, padin_26, padin_193, pado_l_t, pado_t_l, r_o, sdo,
     shift_o, slf_op_00_17, slf_op_01_17, slf_op_02_17, slf_op_03_17,
     slf_op_04_17, slf_op_05_17, slf_op_06_17, slf_op_07_17,
     slf_op_08_17, slf_op_09_17, slf_op_10_17, slf_op_11_17,
     slf_op_12_17, slf_op_13_17, slf_op_14_17, slf_op_15_17,
     slf_op_16_17, slf_op_16_18, slf_op_16_19, slf_op_16_20,
     slf_op_16_21, slf_op_16_22, slf_op_16_23, slf_op_16_24,
     slf_op_16_25, slf_op_16_26, slf_op_16_27, slf_op_16_28,
     slf_op_16_29, slf_op_16_30, slf_op_16_31, slf_op_16_32,
     slf_op_16_33, tclk_o, update_o, bl, pgate_l, reset_l,
     sp4_h_r_16_17, sp4_h_r_16_18, sp4_h_r_16_19, sp4_h_r_16_20,
     sp4_h_r_16_21, sp4_h_r_16_22, sp4_h_r_16_23, sp4_h_r_16_24,
     sp4_h_r_16_25, sp4_h_r_16_26, sp4_h_r_16_27, sp4_h_r_16_28,
     sp4_h_r_16_29, sp4_h_r_16_30, sp4_h_r_16_31, sp4_h_r_16_32,
     sp4_h_r_16_33, sp4_r_v_b_16_17, sp4_r_v_b_16_18, sp4_r_v_b_16_19,
     sp4_r_v_b_16_20, sp4_r_v_b_16_21, sp4_r_v_b_16_22,
     sp4_r_v_b_16_23, sp4_r_v_b_16_24, sp4_r_v_b_16_25,
     sp4_r_v_b_16_26, sp4_r_v_b_16_27, sp4_r_v_b_16_28,
     sp4_r_v_b_16_29, sp4_r_v_b_16_30, sp4_r_v_b_16_31,
     sp4_r_v_b_16_32, sp4_v_b_00_17, sp4_v_b_01_17, sp4_v_b_02_17,
     sp4_v_b_03_17, sp4_v_b_04_17, sp4_v_b_05_17, sp4_v_b_06_17,
     sp4_v_b_07_17, sp4_v_b_08_17, sp4_v_b_09_17, sp4_v_b_10_17,
     sp4_v_b_11_17, sp4_v_b_12_17, sp4_v_b_13_17, sp4_v_b_14_17,
     sp4_v_b_15_17, sp4_v_b_16_17, sp12_h_r_16_17, sp12_h_r_16_18,
     sp12_h_r_16_19, sp12_h_r_16_20, sp12_h_r_16_21, sp12_h_r_16_22,
     sp12_h_r_16_23, sp12_h_r_16_24, sp12_h_r_16_25, sp12_h_r_16_26,
     sp12_h_r_16_27, sp12_h_r_16_28, sp12_h_r_16_29, sp12_h_r_16_30,
     sp12_h_r_16_31, sp12_h_r_16_32, sp12_v_b_01_17, sp12_v_b_02_17,
     sp12_v_b_03_17, sp12_v_b_04_17, sp12_v_b_05_17, sp12_v_b_06_17,
     sp12_v_b_07_17, sp12_v_b_08_17, sp12_v_b_09_17, sp12_v_b_10_17,
     sp12_v_b_11_17, sp12_v_b_12_17, sp12_v_b_13_17, sp12_v_b_14_17,
     sp12_v_b_15_17, sp12_v_b_16_17, vdd_cntl_l, wl_l, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bnl_op_01_17,
     bnl_op_02_17, bnl_op_03_17, bnl_op_04_17, bnl_op_05_17,
     bnl_op_06_17, bnl_op_07_17, bnl_op_08_17, bnl_op_09_17,
     bnl_op_10_17, bnl_op_11_17, bnl_op_12_17, bnl_op_13_17,
     bnl_op_14_17, bnl_op_15_17, bnl_op_16_17, bnr_op_00_17,
     bnr_op_01_17, bnr_op_02_17, bnr_op_03_17, bnr_op_04_17,
     bnr_op_05_17, bnr_op_06_17, bnr_op_07_17, bnr_op_08_17,
     bnr_op_09_17, bnr_op_10_17, bnr_op_11_17, bnr_op_12_17,
     bnr_op_13_17, bnr_op_14_17, bnr_op_15_17, bnr_op_16_17,
     bot_op_01_17, bot_op_02_17, bot_op_03_17, bot_op_04_17,
     bot_op_05_17, bot_op_06_17, bot_op_07_17, bot_op_08_17,
     bot_op_09_17, bot_op_10_17, bot_op_11_17, bot_op_12_17,
     bot_op_13_17, bot_op_14_17, bot_op_15_17, bot_op_16_17, bs_en_i,
     carry_in_01_17, carry_in_02_17, carry_in_03_17, carry_in_04_17,
     carry_in_05_17, carry_in_06_17, carry_in_07_17, carry_in_09_17,
     carry_in_10_17, carry_in_11_17, carry_in_12_17, carry_in_13_17,
     carry_in_14_17, carry_in_15_17, carry_in_16_17, ceb_i,
     end_of_startup_lft_t, end_of_startup_top_l, glb_in, hiz_b_i,
     hold_l_t, hold_t_l, mode_i, padin_l_t, padin_t_l, prog, purst,
     r_i, rgt_op_16_17, rgt_op_16_18, rgt_op_16_19, rgt_op_16_20,
     rgt_op_16_21, rgt_op_16_22, rgt_op_16_23, rgt_op_16_24,
     rgt_op_16_25, rgt_op_16_26, rgt_op_16_27, rgt_op_16_28,
     rgt_op_16_29, rgt_op_16_30, rgt_op_16_31, rgt_op_16_32, sdi,
     shift_i, tclk_i, tiegnd, tievdd, tnr_op_16_32, update_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bs_en_o, ceb_o,
     fabric_out_00_17, fabric_out_15_33, fabric_out_16_33, hiz_b_o,
     mode_o, padin_26, padin_193, r_o, sdo, shift_o, tclk_o, update_o;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en_i,
     carry_in_01_17, carry_in_02_17, carry_in_03_17, carry_in_04_17,
     carry_in_05_17, carry_in_06_17, carry_in_07_17, carry_in_09_17,
     carry_in_10_17, carry_in_11_17, carry_in_12_17, carry_in_13_17,
     carry_in_14_17, carry_in_15_17, carry_in_16_17, ceb_i, hiz_b_i,
     hold_l_t, hold_t_l, mode_i, prog, purst, r_i, sdi, shift_i,
     tclk_i, tiegnd, tievdd, update_i;

output [7:0]  slf_op_16_31;
output [383:0]  cf_l;
output [7:0]  slf_op_16_27;
output [7:0]  bm_sa_o;
output [7:0]  slf_op_09_17;
output [7:0]  slf_op_16_29;
output [7:0]  slf_op_16_28;
output [383:0]  cf_t;
output [7:0]  slf_op_12_17;
output [7:0]  slf_op_16_32;
output [49:24]  padeb_l_t;
output [7:0]  slf_op_16_25;
output [7:0]  slf_op_13_17;
output [7:0]  slf_op_08_17;
output [7:0]  slf_op_07_17;
output [7:0]  slf_op_16_22;
output [7:0]  slf_op_10_17;
output [7:0]  slf_op_16_30;
output [7:0]  slf_op_16_19;
output [7:0]  slf_op_02_17;
output [49:24]  pado_l_t;
output [7:0]  slf_op_11_17;
output [7:0]  slf_op_05_17;
output [7:0]  slf_op_16_26;
output [7:0]  slf_op_16_23;
output [7:0]  slf_op_04_17;
output [7:0]  slf_op_16_17;
output [7:0]  slf_op_03_17;
output [7:0]  slf_op_16_21;
output [3:0]  slf_op_16_33;
output [7:0]  slf_op_06_17;
output [7:0]  slf_op_16_20;
output [7:0]  slf_op_15_17;
output [3:0]  slf_op_00_17;
output [7:0]  slf_op_16_18;
output [29:0]  pado_t_l;
output [7:0]  slf_op_16_24;
output [7:0]  slf_op_01_17;
output [7:0]  slf_op_14_17;
output [29:0]  padeb_t_l;

inout [23:0]  sp12_h_r_16_23;
inout [23:0]  sp12_h_r_16_22;
inout [47:0]  sp4_h_r_16_18;
inout [23:0]  sp12_h_r_16_17;
inout [47:0]  sp4_v_b_12_17;
inout [23:0]  sp12_h_r_16_21;
inout [47:0]  sp4_v_b_06_17;
inout [23:0]  sp12_v_b_11_17;
inout [47:0]  sp4_v_b_09_17;
inout [47:0]  sp4_r_v_b_16_27;
inout [47:0]  sp4_v_b_13_17;
inout [47:0]  sp4_v_b_11_17;
inout [47:0]  sp4_h_r_16_31;
inout [47:0]  sp4_h_r_16_30;
inout [47:0]  sp4_r_v_b_16_18;
inout [47:0]  sp4_v_b_10_17;
inout [47:0]  sp4_h_r_16_22;
inout [23:0]  sp12_h_r_16_20;
inout [47:0]  sp4_r_v_b_16_20;
inout [47:0]  sp4_r_v_b_16_28;
inout [47:0]  sp4_r_v_b_16_25;
inout [23:0]  sp12_h_r_16_28;
inout [47:0]  sp4_r_v_b_16_21;
inout [23:0]  sp12_h_r_16_31;
inout [23:0]  sp12_h_r_16_19;
inout [47:0]  sp4_r_v_b_16_26;
inout [47:0]  sp4_h_r_16_20;
inout [47:0]  sp4_h_r_16_32;
inout [23:0]  sp12_h_r_16_18;
inout [47:0]  sp4_h_r_16_24;
inout [23:0]  sp12_v_b_01_17;
inout [47:0]  sp4_v_b_02_17;
inout [23:0]  sp12_v_b_02_17;
inout [47:0]  sp4_h_r_16_23;
inout [47:0]  sp4_r_v_b_16_17;
inout [47:0]  sp4_r_v_b_16_30;
inout [23:0]  sp12_v_b_15_17;
inout [23:0]  sp12_h_r_16_25;
inout [23:0]  sp12_h_r_16_32;
inout [47:0]  sp4_h_r_16_27;
inout [47:0]  sp4_v_b_03_17;
inout [23:0]  sp12_v_b_09_17;
inout [23:0]  sp12_v_b_16_17;
inout [47:0]  sp4_h_r_16_26;
inout [15:0]  sp4_h_r_16_33;
inout [23:0]  sp12_v_b_13_17;
inout [23:0]  sp12_v_b_07_17;
inout [23:0]  sp12_h_r_16_26;
inout [47:0]  sp4_h_r_16_29;
inout [47:0]  sp4_h_r_16_25;
inout [47:0]  sp4_h_r_16_28;
inout [47:0]  sp4_v_b_05_17;
inout [47:0]  sp4_v_b_04_17;
inout [47:0]  sp4_r_v_b_16_31;
inout [47:0]  sp4_v_b_16_17;
inout [47:0]  sp4_r_v_b_16_24;
inout [23:0]  sp12_v_b_10_17;
inout [23:0]  sp12_v_b_03_17;
inout [47:0]  sp4_r_v_b_16_32;
inout [23:0]  sp12_h_r_16_27;
inout [47:0]  sp4_h_r_16_17;
inout [23:0]  sp12_v_b_06_17;
inout [23:0]  sp12_v_b_05_17;
inout [47:0]  sp4_v_b_07_17;
inout [47:0]  sp4_h_r_16_21;
inout [23:0]  sp12_v_b_08_17;
inout [271:0]  vdd_cntl_l;
inout [23:0]  sp12_v_b_12_17;
inout [47:0]  sp4_h_r_16_19;
inout [271:0]  wl_l;
inout [47:0]  sp4_v_b_14_17;
inout [271:0]  reset_l;
inout [15:0]  sp4_v_b_00_17;
inout [47:0]  sp4_r_v_b_16_22;
inout [47:0]  sp4_v_b_15_17;
inout [47:0]  sp4_r_v_b_16_23;
inout [869:0]  bl;
inout [23:0]  sp12_h_r_16_29;
inout [23:0]  sp12_v_b_04_17;
inout [23:0]  sp12_h_r_16_30;
inout [271:0]  pgate_l;
inout [47:0]  sp4_v_b_01_17;
inout [47:0]  sp4_r_v_b_16_19;
inout [23:0]  sp12_h_r_16_24;
inout [47:0]  sp4_r_v_b_16_29;
inout [47:0]  sp4_v_b_08_17;
inout [23:0]  sp12_v_b_14_17;

input [7:0]  bot_op_05_17;
input [7:0]  rgt_op_16_26;
input [7:0]  bnr_op_16_17;
input [7:0]  bnl_op_08_17;
input [7:0]  rgt_op_16_17;
input [7:0]  rgt_op_16_20;
input [16:1]  end_of_startup_top_l;
input [7:0]  bnl_op_05_17;
input [7:0]  bnr_op_14_17;
input [7:0]  rgt_op_16_31;
input [7:0]  rgt_op_16_19;
input [7:0]  bot_op_02_17;
input [7:0]  bnr_op_05_17;
input [7:0]  bnr_op_08_17;
input [7:0]  bnr_op_00_17;
input [7:0]  rgt_op_16_22;
input [7:0]  rgt_op_16_25;
input [7:0]  bnr_op_13_17;
input [7:0]  rgt_op_16_32;
input [7:0]  bnl_op_10_17;
input [7:0]  bnr_op_04_17;
input [7:0]  bnl_op_13_17;
input [7:0]  glb_in;
input [7:0]  bnl_op_16_17;
input [7:0]  bnr_op_06_17;
input [7:0]  bnl_op_06_17;
input [7:0]  bot_op_04_17;
input [7:0]  bot_op_16_17;
input [7:0]  bnl_op_02_17;
input [7:0]  rgt_op_16_30;
input [7:0]  bot_op_14_17;
input [7:0]  bnr_op_12_17;
input [7:0]  bnr_op_09_17;
input [7:0]  bot_op_03_17;
input [7:0]  bnl_op_09_17;
input [7:0]  rgt_op_16_23;
input [7:0]  bnl_op_01_17;
input [7:0]  bnl_op_15_17;
input [7:0]  rgt_op_16_21;
input [7:0]  bnr_op_10_17;
input [7:0]  bot_op_11_17;
input [7:0]  bnl_op_14_17;
input [7:0]  bot_op_06_17;
input [7:0]  rgt_op_16_29;
input [7:0]  bnl_op_04_17;
input [7:0]  bot_op_13_17;
input [7:0]  bnr_op_11_17;
input [7:0]  rgt_op_16_27;
input [7:0]  bnr_op_02_17;
input [7:0]  bot_op_01_17;
input [7:0]  bot_op_07_17;
input [7:0]  bnl_op_03_17;
input [7:0]  rgt_op_16_24;
input [7:0]  bnr_op_07_17;
input [7:0]  bnr_op_15_17;
input [7:0]  bm_sa_i;
input [7:0]  bot_op_12_17;
input [16:1]  end_of_startup_lft_t;
input [7:0]  bot_op_08_17;
input [7:0]  bot_op_15_17;
input [7:0]  bnl_op_11_17;
input [7:0]  bnl_op_12_17;
input [49:24]  padin_l_t;
input [7:0]  bnr_op_01_17;
input [7:0]  rgt_op_16_28;
input [29:0]  padin_t_l;
input [7:0]  rgt_op_16_18;
input [7:0]  bot_op_09_17;
input [3:0]  tnr_op_16_32;
input [7:0]  bnl_op_07_17;
input [7:0]  bnr_op_03_17;
input [7:0]  bot_op_10_17;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:47]  net2619;

wire  [0:47]  net3554;

wire  [0:23]  net3939;

wire  [0:7]  net2874;

wire  [0:47]  net4051;

wire  [0:47]  net3112;

wire  [0:47]  net3389;

wire  [0:47]  net3820;

wire  [0:23]  net3383;

wire  [0:47]  net3168;

wire  [0:47]  net4367;

wire  [0:47]  net2402;

wire  [0:47]  net4571;

wire  [0:47]  net2343;

wire  [0:47]  net3076;

wire  [0:47]  net3073;

wire  [0:47]  net2335;

wire  [0:7]  net4892;

wire  [0:7]  net4343;

wire  [0:47]  net4901;

wire  [0:47]  net3562;

wire  [0:23]  net4525;

wire  [0:47]  net4090;

wire  [0:47]  net2622;

wire  [0:23]  net3480;

wire  [0:23]  net2280;

wire  [0:47]  net3570;

wire  [0:7]  net3527;

wire  [0:47]  net4385;

wire  [0:47]  net3729;

wire  [0:7]  net2259;

wire  [0:7]  net3788;

wire  [0:7]  net4112;

wire  [0:23]  net2959;

wire  [0:47]  net3978;

wire  [0:47]  net3819;

wire  [0:47]  net3841;

wire  [0:23]  net4517;

wire  [0:47]  net3166;

wire  [0:7]  net2398;

wire  [0:23]  net3710;

wire  [0:7]  net2164;

wire  [0:23]  net2633;

wire  [0:47]  net2864;

wire  [0:47]  net4331;

wire  [0:47]  net4250;

wire  [0:23]  net3809;

wire  [0:23]  net3222;

wire  [0:47]  net2587;

wire  [0:47]  net2678;

wire  [0:7]  net4835;

wire  [0:47]  net4465;

wire  [0:47]  net2787;

wire  [0:7]  net3854;

wire  [0:47]  net4495;

wire  [0:7]  net2160;

wire  [0:47]  net3193;

wire  [0:23]  net4297;

wire  [0:47]  net4202;

wire  [0:7]  net2611;

wire  [0:23]  net3645;

wire  [0:7]  net4832;

wire  [0:47]  net4220;

wire  [0:23]  net2634;

wire  [0:47]  net3896;

wire  [0:7]  net3750;

wire  [0:47]  net2289;

wire  [0:47]  net2320;

wire  [0:23]  net3457;

wire  [0:47]  net4795;

wire  [0:23]  net4361;

wire  [0:23]  net4848;

wire  [0:7]  net3647;

wire  [0:47]  net3555;

wire  [0:23]  net3219;

wire  [0:23]  net4429;

wire  [0:23]  net2730;

wire  [0:47]  net2592;

wire  [0:7]  net2316;

wire  [0:23]  net2342;

wire  [0:7]  net2713;

wire  [0:47]  net2429;

wire  [0:23]  net4592;

wire  [0:47]  net2699;

wire  [0:7]  net4077;

wire  [0:23]  net2448;

wire  [0:7]  net2434;

wire  [0:47]  net2902;

wire  [0:47]  net3679;

wire  [0:23]  net3050;

wire  [0:23]  net3449;

wire  [0:47]  net4334;

wire  [0:7]  net4566;

wire  [0:47]  net3877;

wire  [0:47]  net3928;

wire  [0:23]  net2567;

wire  [0:7]  net4438;

wire  [0:47]  net3715;

wire  [0:47]  net3568;

wire  [0:47]  net3109;

wire  [0:23]  net4589;

wire  [0:47]  net4166;

wire  [0:47]  net3390;

wire  [0:47]  net2238;

wire  [0:7]  net3205;

wire  [0:47]  net4413;

wire  [0:47]  net4042;

wire  [0:47]  net2324;

wire  [0:23]  net2505;

wire  [0:47]  net3391;

wire  [0:23]  net3612;

wire  [0:7]  net3973;

wire  [0:7]  net3753;

wire  [0:47]  net4171;

wire  [0:7]  net3264;

wire  [0:7]  net3364;

wire  [0:7]  net4891;

wire  [0:47]  net3434;

wire  [0:23]  net2235;

wire  [0:47]  net4249;

wire  [0:7]  net2818;

wire  [0:47]  net3552;

wire  [0:23]  net3613;

wire  [0:47]  net3515;

wire  [0:7]  net2492;

wire  [0:7]  net2775;

wire  [0:47]  net3388;

wire  [0:7]  net4016;

wire  [0:7]  net4890;

wire  [0:47]  net3227;

wire  [0:23]  net3446;

wire  [0:47]  net3329;

wire  [0:23]  net4191;

wire  [0:23]  net2351;

wire  [0:7]  net2876;

wire  [0:47]  net3655;

wire  [0:47]  net4384;

wire  [0:7]  net3526;

wire  [0:47]  net2515;

wire  [0:7]  net4625;

wire  [0:23]  net2668;

wire  [0:23]  net4098;

wire  [0:47]  net2223;

wire  [0:23]  net3451;

wire  [0:47]  net2901;

wire  [0:47]  net4547;

wire  [0:47]  net4543;

wire  [0:47]  net3844;

wire  [0:7]  net4405;

wire  [0:47]  net2315;

wire  [0:23]  net2454;

wire  [0:23]  net4035;

wire  [0:7]  net2712;

wire  [0:7]  net2549;

wire  [0:47]  net3763;

wire  [0:47]  net3244;

wire  [0:47]  net2865;

wire  [0:23]  net4034;

wire  [0:7]  net2875;

wire  [0:23]  net4852;

wire  [0:23]  net4354;

wire  [0:23]  net2570;

wire  [0:47]  net2673;

wire  [0:23]  net3874;

wire  [0:23]  net3772;

wire  [0:23]  net4918;

wire  [0:47]  net4056;

wire  [0:47]  net3725;

wire  [0:7]  net3853;

wire  [0:23]  net3610;

wire  [0:47]  net4791;

wire  [0:23]  net2449;

wire  [0:23]  net4849;

wire  [0:7]  net2655;

wire  [0:7]  net2397;

wire  [0:23]  net2724;

wire  [0:23]  net2796;

wire  [0:47]  net2623;

wire  [0:47]  net2899;

wire  [0:23]  net4132;

wire  [0:47]  net3728;

wire  [0:47]  net4537;

wire  [0:7]  net3530;

wire  [0:7]  net2399;

wire  [0:47]  net2916;

wire  [0:31]  net4979;

wire  [0:47]  net3002;

wire  [0:23]  net4028;

wire  [0:23]  net2446;

wire  [0:47]  net2703;

wire  [0:47]  net2786;

wire  [0:47]  net3402;

wire  [0:23]  net3122;

wire  [0:23]  net4135;

wire  [0:23]  net4914;

wire  [0:47]  net2624;

wire  [0:47]  net4168;

wire  [0:47]  net4007;

wire  [0:23]  net3644;

wire  [0:47]  net3519;

wire  [0:47]  net2739;

wire  [0:7]  net4788;

wire  [0:47]  net3657;

wire  [0:23]  net4425;

wire  [0:23]  net2277;

wire  [0:47]  net3926;

wire  [0:7]  net2610;

wire  [0:23]  net2962;

wire  [0:23]  net4266;

wire  [0:23]  net2457;

wire  [0:23]  net2828;

wire  [0:23]  net2896;

wire  [0:47]  net4467;

wire  [0:47]  net3682;

wire  [0:23]  net2993;

wire  [0:23]  net2479;

wire  [0:47]  net4041;

wire  [0:47]  net3399;

wire  [0:47]  net3351;

wire  [0:23]  net4913;

wire  [0:23]  net3972;

wire  [0:7]  net2936;

wire  [0:47]  net2419;

wire  [0:23]  net4523;

wire  [0:47]  net3879;

wire  [0:47]  net4903;

wire  [0:23]  net3057;

wire  [0:47]  net2704;

wire  [0:47]  net3161;

wire  [0:23]  net3711;

wire  [0:47]  net2413;

wire  [0:23]  net4786;

wire  [0:7]  net2257;

wire  [0:7]  net3752;

wire  [0:23]  net3609;

wire  [0:47]  net4332;

wire  [0:47]  net4902;

wire  [0:47]  net3678;

wire  [0:23]  net4200;

wire  [0:47]  net3923;

wire  [0:23]  net4101;

wire  [0:23]  net4587;

wire  [0:23]  net3056;

wire  [0:7]  net3531;

wire  [0:47]  net4055;

wire  [0:7]  net2612;

wire  [0:23]  net4459;

wire  [0:23]  net4526;

wire  [0:23]  net2968;

wire  [0:7]  net4182;

wire  [0:7]  net2199;

wire  [0:7]  net3623;

wire  [0:47]  net3842;

wire  [0:7]  net3691;

wire  [0:47]  net3271;

wire  [0:7]  net2552;

wire  [0:47]  net3681;

wire  [0:7]  net4240;

wire  [0:23]  net3709;

wire  [0:47]  net3518;

wire  [0:7]  net2482;

wire  [0:23]  net4591;

wire  [0:47]  net2513;

wire  [0:47]  net3925;

wire  [0:7]  net2771;

wire  [0:23]  net3319;

wire  [0:23]  net3774;

wire  [0:47]  net2286;

wire  [0:23]  net3448;

wire  [0:23]  net3544;

wire  [0:47]  net3602;

wire  [0:7]  net3914;

wire  [0:47]  net4482;

wire  [0:47]  net4469;

wire  [0:7]  net3810;

wire  [0:7]  net3912;

wire  [0:47]  net3435;

wire  [0:23]  net4426;

wire  [0:7]  net3134;

wire  [0:47]  net4470;

wire  [0:47]  net2841;

wire  [0:47]  net2573;

wire  [0:47]  net4870;

wire  [0:23]  net2451;

wire  [0:47]  net3113;

wire  [0:47]  net3065;

wire  [0:47]  net2577;

wire  [0:47]  net4905;

wire  [0:7]  net3625;

wire  [0:7]  net2251;

wire  [0:7]  net2548;

wire  [0:7]  net3690;

wire  [0:23]  net3120;

wire  [0:47]  net2401;

wire  [0:47]  net3654;

wire  [0:47]  net2900;

wire  [0:23]  net4850;

wire  [0:47]  net2412;

wire  [0:47]  net4492;

wire  [0:47]  net3407;

wire  [0:7]  net3915;

wire  [0:23]  net3447;

wire  [0:7]  net4402;

wire  [0:47]  net4329;

wire  [0:47]  net4416;

wire  [0:23]  net4458;

wire  [0:23]  net3971;

wire  [0:7]  net4181;

wire  [0:47]  net3062;

wire  [0:23]  net2447;

wire  [0:47]  net4580;

wire  [0:47]  net3652;

wire  [0:7]  net2669;

wire  [0:23]  net2450;

wire  [0:23]  net2569;

wire  [0:23]  net3614;

wire  [0:23]  net3318;

wire  [0:23]  net3620;

wire  [0:7]  net3856;

wire  [0:47]  net2425;

wire  [0:7]  net3424;

wire  [0:23]  net4363;

wire  [0:7]  net2506;

wire  [0:7]  net3144;

wire  [0:47]  net3878;

wire  [0:47]  net3732;

wire  [0:23]  net3287;

wire  [0:47]  net2218;

wire  [0:47]  net3567;

wire  [0:47]  net4866;

wire  [0:23]  net2958;

wire  [0:7]  net4122;

wire  [0:23]  net3483;

wire  [0:23]  net4435;

wire  [0:7]  net4504;

wire  [0:47]  net3030;

wire  [0:23]  net4265;

wire  [0:47]  net2591;

wire  [0:47]  net4139;

wire  [0:47]  net3225;

wire  [0:7]  net3913;

wire  [0:47]  net2288;

wire  [0:47]  net3027;

wire  [0:47]  net4304;

wire  [0:47]  net3353;

wire  [0:47]  net3228;

wire  [0:47]  net2753;

wire  [0:7]  net3796;

wire  [0:47]  net2418;

wire  [0:47]  net2700;

wire  [0:7]  net4509;

wire  [0:47]  net4088;

wire  [0:47]  net4484;

wire  [0:7]  net4242;

wire  [0:47]  net4904;

wire  [0:47]  net2840;

wire  [0:23]  net2568;

wire  [0:7]  net3484;

wire  [0:47]  net3760;

wire  [0:47]  net3111;

wire  [0:23]  net2460;

wire  [0:47]  net4855;

wire  [0:23]  net4461;

wire  [0:47]  net4792;

wire  [0:47]  net3491;

wire  [0:47]  net4572;

wire  [0:7]  net4183;

wire  [0:47]  net3714;

wire  [0:47]  net3891;

wire  [0:23]  net3873;

wire  [0:47]  net3274;

wire  [0:7]  net3749;

wire  [0:7]  net3427;

wire  [0:7]  net3321;

wire  [0:7]  net3916;

wire  [0:47]  net2621;

wire  [0:47]  net2738;

wire  [0:7]  net3423;

wire  [0:47]  net3239;

wire  [0:47]  net3078;

wire  [0:23]  net2635;

wire  [0:47]  net3356;

wire  [0:47]  net4005;

wire  [0:47]  net4253;

wire  [0:23]  net4103;

wire  [0:47]  net4308;

wire  [0:47]  net3192;

wire  [0:23]  net3946;

wire  [0:47]  net2430;

wire  [0:47]  net3162;

wire  [0:47]  net3080;

wire  [0:23]  net2636;

wire  [0:23]  net3643;

wire  [0:47]  net3881;

wire  [0:47]  net2246;

wire  [0:23]  net4522;

wire  [0:7]  net4508;

wire  [0:47]  net4797;

wire  [0:47]  net4466;

wire  [0:47]  net2428;

wire  [0:47]  net4170;

wire  [0:7]  net4436;

wire  [0:47]  net3876;

wire  [0:23]  net2458;

wire  [0:23]  net2794;

wire  [0:47]  net2538;

wire  [0:7]  net3460;

wire  [0:23]  net4264;

wire  [0:47]  net3081;

wire  [0:47]  net4415;

wire  [0:7]  net2162;

wire  [0:23]  net4197;

wire  [0:47]  net3079;

wire  [0:47]  net4528;

wire  [0:47]  net2516;

wire  [0:47]  net4703;

wire  [0:23]  net3221;

wire  [0:23]  net3376;

wire  [0:47]  net2539;

wire  [0:23]  net3381;

wire  [0:47]  net3813;

wire  [0:23]  net2281;

wire  [0:23]  net2733;

wire  [0:47]  net3189;

wire  [0:7]  net3307;

wire  [0:7]  net2553;

wire  [0:7]  net2832;

wire  [0:7]  net4018;

wire  [0:7]  net3693;

wire  [0:47]  net4533;

wire  [0:7]  net2393;

wire  [0:7]  net3367;

wire  [0:47]  net2747;

wire  [0:23]  net3546;

wire  [0:47]  net3565;

wire  [0:47]  net4569;

wire  [0:23]  net3806;

wire  [0:47]  net4545;

wire  [0:23]  net2665;

wire  [0:23]  net3940;

wire  [0:7]  net4299;

wire  [0:47]  net4003;

wire  [0:7]  net4404;

wire  [0:47]  net2839;

wire  [0:47]  net3387;

wire  [0:23]  net3482;

wire  [0:7]  net2266;

wire  [0:47]  net4793;

wire  [0:23]  net4588;

wire  [0:23]  net2503;

wire  [0:47]  net4869;

wire  [0:7]  net4342;

wire  [0:47]  net3005;

wire  [0:47]  net4309;

wire  [0:47]  net4548;

wire  [0:7]  net3586;

wire  [0:47]  net4412;

wire  [0:23]  net3320;

wire  [0:47]  net2679;

wire  [0:47]  net4169;

wire  [0:47]  net2590;

wire  [0:47]  net3063;

wire  [0:23]  net4843;

wire  [0:47]  net3355;

wire  [0:47]  net4536;

wire  [0:47]  net3680;

wire  [0:47]  net2537;

wire  [0:23]  net2795;

wire  [0:47]  net3980;

wire  [0:47]  net3817;

wire  [0:47]  net2755;

wire  [0:47]  net2917;

wire  [0:7]  net4136;

wire  [0:47]  net3025;

wire  [0:7]  net3949;

wire  [0:7]  net2436;

wire  [0:23]  net3808;

wire  [0:47]  net3492;

wire  [0:47]  net4141;

wire  [0:7]  net4075;

wire  [0:47]  net2576;

wire  [0:7]  net2714;

wire  [0:47]  net3437;

wire  [0:23]  net3286;

wire  [0:7]  net3852;

wire  [0:47]  net2903;

wire  [0:47]  net4579;

wire  [0:7]  net4505;

wire  [0:7]  net2773;

wire  [0:47]  net4820;

wire  [0:47]  net2245;

wire  [0:7]  net2879;

wire  [0:23]  net2732;

wire  [0:23]  net3055;

wire  [0:47]  net4859;

wire  [0:7]  net2609;

wire  [0:23]  net3870;

wire  [0:47]  net4496;

wire  [0:7]  net3365;

wire  [0:47]  net2285;

wire  [0:7]  net3633;

wire  [0:23]  net2561;

wire  [3:0]  slf_op_09_33;

wire  [0:7]  net2435;

wire  [0:23]  net3157;

wire  [0:47]  net3731;

wire  [3:0]  slf_op_07_33;

wire  [0:23]  net4272;

wire  [0:23]  net4102;

wire  [0:7]  net2177;

wire  [0:23]  net3123;

wire  [0:7]  net2608;

wire  [0:23]  net3969;

wire  [0:47]  net2784;

wire  [0:47]  net3716;

wire  [0:23]  net4460;

wire  [0:47]  net4008;

wire  [0:47]  net4497;

wire  [0:47]  net4143;

wire  [0:23]  net2631;

wire  [0:47]  net2426;

wire  [0:47]  net2322;

wire  [0:47]  net3326;

wire  [0:23]  net3218;

wire  [0:7]  net2711;

wire  [0:7]  net4834;

wire  [0:7]  net3368;

wire  [0:7]  net4015;

wire  [0:7]  net4241;

wire  [0:23]  net2893;

wire  [0:7]  net3204;

wire  [3:0]  slf_op_00_18;

wire  [3:0]  slf_op_00_25;

wire  [3:0]  slf_op_13_33;

wire  [0:23]  net4037;

wire  [0:47]  net4382;

wire  [0:47]  net2862;

wire  [0:23]  net3288;

wire  [0:47]  net2536;

wire  [0:47]  net4383;

wire  [0:47]  net4471;

wire  [3:0]  slf_op_10_33;

wire  [0:47]  net4307;

wire  [0:47]  net2740;

wire  [0:47]  net3713;

wire  [0:7]  net2395;

wire  [0:47]  net2291;

wire  [0:7]  net2810;

wire  [0:47]  net3489;

wire  [0:47]  net2948;

wire  [0:47]  net4823;

wire  [0:47]  net3977;

wire  [0:47]  net3229;

wire  [0:7]  net3528;

wire  [0:47]  net2783;

wire  [0:47]  net3517;

wire  [0:47]  net3880;

wire  [0:7]  net2937;

wire  [0:23]  net3783;

wire  [0:47]  net4534;

wire  [0:47]  net3814;

wire  [0:47]  net3892;

wire  [0:47]  net2837;

wire  [0:7]  net3694;

wire  [0:23]  net3708;

wire  [0:47]  net2945;

wire  [0:7]  net4506;

wire  [0:47]  net2998;

wire  [0:47]  net2290;

wire  [0:47]  net2337;

wire  [0:47]  net4380;

wire  [0:23]  net2991;

wire  [0:47]  net4798;

wire  [0:7]  net3692;

wire  [0:47]  net2947;

wire  [0:23]  net4263;

wire  [0:7]  net4764;

wire  [0:7]  net2772;

wire  [0:47]  net3976;

wire  [3:0]  slf_op_06_33;

wire  [0:47]  net2782;

wire  [0:7]  net4440;

wire  [0:23]  net2798;

wire  [0:7]  net3363;

wire  [0:7]  net4238;

wire  [0:23]  net3871;

wire  [0:23]  net3872;

wire  [0:47]  net4203;

wire  [0:7]  net2643;

wire  [0:23]  net3317;

wire  [0:47]  net3191;

wire  [0:7]  net3751;

wire  [0:7]  net4285;

wire  [0:47]  net3439;

wire  [0:47]  net3328;

wire  [0:47]  net2867;

wire  [0:7]  net4076;

wire  [0:23]  net3775;

wire  [0:7]  net4277;

wire  [0:23]  net2805;

wire  [0:47]  net4059;

wire  [0:47]  net3598;

wire  [0:47]  net3188;

wire  [3:0]  slf_op_00_19;

wire  [0:47]  net4578;

wire  [0:7]  net4568;

wire  [3:0]  slf_op_00_31;

wire  [0:47]  net3165;

wire  [0:47]  net4206;

wire  [0:23]  net3285;

wire  [0:47]  net3240;

wire  [0:7]  net2433;

wire  [0:23]  net3707;

wire  [0:47]  net3599;

wire  [0:23]  net3156;

wire  [0:23]  net4598;

wire  [0:23]  net2354;

wire  [0:47]  net4857;

wire  [0:23]  net3938;

wire  [0:47]  net4217;

wire  [0:7]  net2163;

wire  [0:23]  net2445;

wire  [0:7]  net4766;

wire  [0:23]  net3776;

wire  [0:47]  net4540;

wire  [0:47]  net2918;

wire  [0:47]  net3924;

wire  [0:47]  net3241;

wire  [0:47]  net4574;

wire  [0:47]  net2735;

wire  [0:47]  net4532;

wire  [0:47]  net3843;

wire  [0:23]  net2452;

wire  [0:7]  net3587;

wire  [0:7]  net4180;

wire  [0:7]  net2551;

wire  [0:23]  net2459;

wire  [0:47]  net4365;

wire  [0:47]  net3352;

wire  [0:47]  net4222;

wire  [0:47]  net4251;

wire  [0:47]  net2511;

wire  [0:47]  net3004;

wire  [0:7]  net3200;

wire  [0:47]  net3840;

wire  [0:47]  net3064;

wire  [0:47]  net4821;

wire  [0:47]  net3600;

wire  [0:47]  net4575;

wire  [3:0]  slf_op_14_33;

wire  [0:47]  net4089;

wire  [0:47]  net4854;

wire  [0:47]  net4573;

wire  [0:23]  net4262;

wire  [0:23]  net3702;

wire  [0:47]  net2431;

wire  [0:7]  net3786;

wire  [0:47]  net2540;

wire  [0:47]  net4146;

wire  [0:47]  net4306;

wire  [0:47]  net3108;

wire  [0:7]  net3590;

wire  [0:47]  net3981;

wire  [0:7]  net2396;

wire  [0:23]  net4787;

wire  [0:47]  net3895;

wire  [3:0]  slf_op_00_28;

wire  [0:7]  net2438;

wire  [0:7]  net2250;

wire  [0:47]  net3487;

wire  [0:47]  net3275;

wire  [0:7]  net2934;

wire  [0:23]  net4261;

wire  [0:23]  net4295;

wire  [0:23]  net3450;

wire  [3:0]  slf_op_04_33;

wire  [0:7]  net4894;

wire  [0:23]  net2231;

wire  [0:23]  net2887;

wire  [0:47]  net3601;

wire  [0:47]  net3066;

wire  [0:7]  net2394;

wire  [0:7]  net4403;

wire  [0:47]  net3392;

wire  [0:47]  net4366;

wire  [0:47]  net3488;

wire  [0:47]  net4546;

wire  [0:47]  net2541;

wire  [0:47]  net3226;

wire  [0:7]  net4567;

wire  [0:47]  net4377;

wire  [3:0]  slf_op_00_29;

wire  [0:47]  net3730;

wire  [0:23]  net4916;

wire  [0:23]  net4133;

wire  [0:47]  net4539;

wire  [0:7]  net4178;

wire  [0:7]  net2260;

wire  [0:47]  net4535;

wire  [0:23]  net2279;

wire  [0:47]  net2949;

wire  [0:7]  net4341;

wire  [0:47]  net4370;

wire  [0:47]  net4207;

wire  [0:23]  net3547;

wire  [0:47]  net3325;

wire  [0:23]  net2642;

wire  [0:47]  net3677;

wire  [3:0]  slf_op_00_21;

wire  [0:7]  net4462;

wire  [0:7]  net2484;

wire  [0:7]  net2332;

wire  [0:7]  net3260;

wire  [0:7]  net2184;

wire  [0:23]  net2356;

wire  [0:47]  net2750;

wire  [0:23]  net4198;

wire  [0:23]  net3481;

wire  [0:47]  net4167;

wire  [0:47]  net2672;

wire  [0:7]  net4564;

wire  [0:23]  net3213;

wire  [0:47]  net3982;

wire  [0:7]  net3458;

wire  [0:23]  net2892;

wire  [0:47]  net3764;

wire  [0:23]  net2349;

wire  [0:47]  net3331;

wire  [0:7]  net4774;

wire  [0:7]  net3529;

wire  [0:23]  net3154;

wire  [3:0]  slf_op_12_33;

wire  [0:47]  net4472;

wire  [0:47]  net3403;

wire  [0:23]  net2229;

wire  [3:0]  slf_op_08_33;

wire  [0:23]  net3807;

wire  [3:0]  slf_op_00_22;

wire  [0:23]  net2632;

wire  [0:47]  net2215;

wire  [0:47]  net4039;

wire  [0:47]  net2240;

wire  [0:47]  net2292;

wire  [0:47]  net4330;

wire  [0:23]  net3865;

wire  [0:7]  net3203;

wire  [0:47]  net2441;

wire  [0:47]  net4858;

wire  [0:47]  net4004;

wire  [0:7]  net4565;

wire  [0:47]  net4254;

wire  [0:23]  net2829;

wire  [0:47]  net4087;

wire  [0:23]  net2992;

wire  [0:47]  net2751;

wire  [0:7]  net4833;

wire  [0:47]  net3762;

wire  [0:23]  net2353;

wire  [0:47]  net3224;

wire  [0:7]  net2331;

wire  [0:23]  net3294;

wire  [0:47]  net3003;

wire  [0:47]  net4874;

wire  [0:47]  net2913;

wire  [0:47]  net4140;

wire  [0:23]  net4427;

wire  [0:23]  net2894;

wire  [0:7]  net2774;

wire  [3:0]  slf_op_00_20;

wire  [0:47]  net4043;

wire  [0:7]  net4893;

wire  [0:47]  net4057;

wire  [0:7]  net3959;

wire  [0:23]  net3058;

wire  [0:47]  net4044;

wire  [0:47]  net2224;

wire  [0:47]  net2842;

wire  [3:0]  slf_op_02_33;

wire  [0:47]  net2283;

wire  [0:7]  net4345;

wire  [0:7]  net4020;

wire  [0:47]  net4529;

wire  [0:7]  net3462;

wire  [0:7]  net3366;

wire  [0:47]  net3845;

wire  [0:7]  net3202;

wire  [0:47]  net2584;

wire  [3:0]  slf_op_03_33;

wire  [0:47]  net3110;

wire  [0:23]  net4785;

wire  [3:0]  slf_op_01_33;

wire  [0:7]  net4017;

wire  [0:23]  net2731;

wire  [0:7]  net2647;

wire  [0:47]  net4214;

wire  [3:0]  slf_op_05_33;

wire  [0:7]  net2188;

wire  [0:47]  net2319;

wire  [0:47]  net3354;

wire  [0:23]  net3125;

wire  [0:23]  net3545;

wire  [0:7]  net4401;

wire  [0:7]  net4830;

wire  [0:47]  net3167;

wire  [0:23]  net2504;

wire  [0:47]  net4218;

wire  [0:7]  net4114;

wire  [0:47]  net4906;

wire  [0:7]  net3589;

wire  [0:23]  net2957;

wire  [0:23]  net2960;

wire  [0:23]  net2994;

wire  [0:23]  net2895;

wire  [3:0]  slf_op_00_27;

wire  [0:47]  net4221;

wire  [0:47]  net4303;

wire  [0:7]  net3425;

wire  [0:47]  net4494;

wire  [0:47]  net3815;

wire  [0:23]  net3539;

wire  [0:7]  net3261;

wire  [0:47]  net3765;

wire  [0:47]  net2588;

wire  [0:47]  net4333;

wire  [0:7]  net4079;

wire  [0:47]  net4414;

wire  [0:47]  net3718;

wire  [0:7]  net3588;

wire  [0:47]  net4058;

wire  [0:47]  net3276;

wire  [0:23]  net3937;

wire  [0:23]  net4298;

wire  [0:47]  net2340;

wire  [0:47]  net3243;

wire  [0:47]  net3550;

wire  [0:23]  net4424;

wire  [0:23]  net2831;

wire  [0:23]  net2729;

wire  [0:7]  net2175;

wire  [0:23]  net4761;

wire  [0:47]  net4531;

wire  [0:7]  net4019;

wire  [0:47]  net2835;

wire  [0:23]  net3155;

wire  [0:47]  net3438;

wire  [0:23]  net3548;

wire  [0:7]  net2995;

wire  [0:47]  net3404;

wire  [0:47]  net2440;

wire  [0:47]  net2287;

wire  [0:23]  net4109;

wire  [0:47]  net4145;

wire  [0:7]  net2333;

wire  [0:7]  net4239;

wire  [0:47]  net2222;

wire  [0:7]  net2317;

wire  [0:23]  net2666;

wire  [0:23]  net4851;

wire  [0:7]  net3855;

wire  [0:47]  net3272;

wire  [0:7]  net3262;

wire  [0:23]  net3121;

wire  [0:47]  net4204;

wire  [0:47]  net3514;

wire  [0:47]  net3190;

wire  [0:7]  net3470;

wire  [0:47]  net4302;

wire  [0:47]  net4483;

wire  [0:47]  net4577;

wire  [0:23]  net2453;

wire  [0:47]  net4873;

wire  [0:47]  net3597;

wire  [0:47]  net2914;

wire  [0:47]  net3566;

wire  [0:47]  net2427;

wire  [0:47]  net3893;

wire  [0:23]  net4100;

wire  [0:47]  net4219;

wire  [0:47]  net4381;

wire  [0:47]  net2785;

wire  [0:47]  net3436;

wire  [0:7]  net2437;

wire  [0:23]  net4915;

wire  [0:23]  net4784;

wire  [0:23]  net4428;

wire  [0:47]  net3553;

wire  [0:7]  net2550;

wire  [0:7]  net3426;

wire  [0:23]  net4360;

wire  [0:47]  net3405;

wire  [0:7]  net2400;

wire  [0:23]  net2797;

wire  [0:47]  net2946;

wire  [0:23]  net4359;

wire  [0:47]  net4856;

wire  [0:7]  net4275;

wire  [0:47]  net2836;

wire  [0:47]  net3163;

wire  [0:23]  net2667;

wire  [0:7]  net2808;

wire  [0:7]  net4831;

wire  [0:47]  net3927;

wire  [0:23]  net2455;

wire  [0:23]  net3284;

wire  [0:47]  net3656;

wire  [0:47]  net4252;

wire  [0:15]  net2411;

wire  [0:47]  net2910;

wire  [3:0]  slf_op_00_32;

wire  [0:23]  net2502;

wire  [0:47]  net4544;

wire  [0:47]  net2674;

wire  [0:47]  net3651;

wire  [0:23]  net4036;

wire  [0:47]  net3077;

wire  [0:47]  net2999;

wire  [0:47]  net2737;

wire  [0:23]  net4917;

wire  [0:47]  net2572;

wire  [0:47]  net3330;

wire  [3:0]  slf_op_00_26;

wire  [0:23]  net2226;

wire  [0:47]  net3029;

wire  [0:47]  net2346;

wire  [0:23]  net4199;

wire  [0:23]  net3611;

wire  [0:7]  net3857;

wire  [0:47]  net4538;

wire  [0:7]  net4507;

wire  [0:47]  net2736;

wire  [0:7]  net4078;

wire  [0:7]  net2878;

wire  [0:47]  net4871;

wire  [0:47]  net2754;

wire  [0:7]  net2715;

wire  [0:47]  net4091;

wire  [0:23]  net2228;

wire  [0:47]  net4368;

wire  [0:47]  net2898;

wire  [0:47]  net2950;

wire  [0:47]  net4822;

wire  [0:47]  net4570;

wire  [0:7]  net4344;

wire  [0:47]  net3717;

wire  [0:47]  net2574;

wire  [0:47]  net3000;

wire  [0:23]  net3646;

wire  [0:47]  net2247;

wire  [0:7]  net3263;

wire  [0:47]  net3894;

wire  [0:23]  net2799;

wire  [0:7]  net2330;

wire  [0:7]  net3689;

wire  [3:0]  slf_op_00_24;

wire  [0:23]  net4134;

wire  [0:7]  net4346;

wire  [0:23]  net2830;

wire  [0:23]  net4362;

wire  [0:47]  net4369;

wire  [0:23]  net4033;

wire  [0:47]  net4144;

wire  [0:47]  net3061;

wire  [0:47]  net2702;

wire  [0:7]  net3201;

wire  [0:7]  net3299;

wire  [0:47]  net3324;

wire  [0:47]  net2213;

wire  [0:47]  net3761;

wire  [0:47]  net3569;

wire  [0:7]  net2716;

wire  [0:47]  net2677;

wire  [0:23]  net3384;

wire  [0:7]  net3136;

wire  [0:47]  net2915;

wire  [0:47]  net4818;

wire  [0:7]  net2167;

wire  [0:23]  net3124;

wire  [0:23]  net3773;

wire  [0:7]  net4179;

wire  [0:47]  net2676;

wire  [0:23]  net4196;

wire  [0:7]  net2265;

wire  [0:47]  net2424;

wire  [0:47]  net3650;

wire  [0:47]  net2863;

wire  [0:47]  net3242;

wire  [0:7]  net2179;

wire  [0:23]  net2961;

wire  [0:23]  net3220;

wire  [0:23]  net4099;

wire  [3:0]  slf_op_00_30;

wire  [7:0]  clk_tree_drv;

wire  [0:47]  net3818;

wire  [0:47]  net3888;

wire  [0:7]  net3158;

wire  [0:7]  net2268;

wire  [0:47]  net2575;

wire  [0:47]  net2248;

wire  [0:47]  net3026;

wire  [0:47]  net3273;

wire  [0:47]  net4872;

wire  [0:47]  net2509;

wire  [0:7]  net2935;

wire  [0:47]  net3983;

wire  [0:47]  net4417;

wire  [0:47]  net3406;

wire  [0:47]  net3733;

wire  [3:0]  slf_op_00_23;

wire  [0:23]  net3283;

wire  [0:47]  net4054;

wire  [0:23]  net3385;

wire  [0:47]  net2701;

wire  [0:47]  net3028;

wire  [0:23]  net4296;

wire  [0:7]  net2169;

wire  [0:7]  net4448;

wire  [0:47]  net4530;

wire  [0:7]  net3951;

wire  [0:47]  net2510;

wire  [0:47]  net4040;

wire  [0:47]  net2514;

wire  [0:47]  net4086;

wire  [0:7]  net2938;

wire  [0:47]  net3516;

wire  [0:23]  net2282;

wire  [0:47]  net2338;

wire  [0:23]  net2566;

wire  [0:47]  net2752;

wire  [0:7]  net2267;

wire  [0:23]  net3970;

wire  [0:7]  net3297;

wire  [0:47]  net4576;

wire  [0:23]  net4590;

wire  [0:47]  net4006;

wire  [0:47]  net4819;

wire  [3:0]  slf_op_11_33;

wire  [0:23]  net4524;

wire  [0:47]  net3236;

wire  [0:23]  net3059;

wire  [0:23]  net2456;

wire  [0:23]  net3935;

wire  [0:23]  net3936;

wire  [0:47]  net2866;

wire  [0:23]  net2236;

wire  [0:47]  net2620;

wire  [0:47]  net3494;

wire  [3:0]  slf_op_15_33;

wire  [0:47]  net3493;

wire  [0:47]  net4205;

wire  [0:7]  net2877;

wire  [0:23]  net3777;

wire  [0:47]  net4493;

wire  [0:47]  net2589;

wire  [0:23]  net3131;

wire  [0:47]  net4796;

wire  [0:23]  net3382;

wire  [0:47]  net3551;

wire  [0:7]  net2645;



lowla_modified I333 ( .clk(net2044), .min(net02084), .lao(net2389));
bram_bufferx4x6 I334 ( .in(net4932), .out(net02084));
tckbufx16 I285 ( .in(net2044), .out(tclk_o));
clk_colbuf8kx8 I_clktree_qdrv_tl ( .clko(clk_tree_drv[7:0]),
     .clki(glb_in[7:0]));
fabric_buf8k I328 ( .f_in(padin_l_t[24]), .f_out(padin_26));
fabric_buf8k I327 ( .f_in(net4926), .f_out(fabric_out_00_17));
preio_top_l I_preio_top_l ( .ceb_i(ceb_i), .ceb_o(net02116),
     .wl_l({wl_l[270], wl_l[271], wl_l[269], wl_l[268], wl_l[266],
     wl_l[267], wl_l[265], wl_l[264], wl_l[262], wl_l[263], wl_l[261],
     wl_l[260], wl_l[258], wl_l[259], wl_l[257], wl_l[256]}),
     .sp4_h_r_16_33(sp4_h_r_16_33[15:0]), .vdd_cntl_l({vdd_cntl_l[270],
     vdd_cntl_l[271], vdd_cntl_l[269], vdd_cntl_l[268],
     vdd_cntl_l[266], vdd_cntl_l[267], vdd_cntl_l[265],
     vdd_cntl_l[264], vdd_cntl_l[262], vdd_cntl_l[263],
     vdd_cntl_l[261], vdd_cntl_l[260], vdd_cntl_l[258],
     vdd_cntl_l[259], vdd_cntl_l[257], vdd_cntl_l[256]}),
     .update_i(update_i), .tievdd(tievdd), .tiegnd(tiegnd),
     .tclk_i(tclk_i), .shift_i(shift_i), .sdi(sdi),
     .reset_l({reset_l[270], reset_l[271], reset_l[269], reset_l[268],
     reset_l[266], reset_l[267], reset_l[265], reset_l[264],
     reset_l[262], reset_l[263], reset_l[261], reset_l[260],
     reset_l[258], reset_l[259], reset_l[257], reset_l[256]}),
     .r_i(r_i), .prog(prog), .pgate_l({pgate_l[270], pgate_l[271],
     pgate_l[269], pgate_l[268], pgate_l[266], pgate_l[267],
     pgate_l[265], pgate_l[264], pgate_l[262], pgate_l[263],
     pgate_l[261], pgate_l[260], pgate_l[258], pgate_l[259],
     pgate_l[257], pgate_l[256]}), .mode_i(mode_i), .hiz_b_i(hiz_b_i),
     .bs_en_i(bs_en_i), .update_o(net2043), .tclk_o(net2044),
     .shift_o(net4938), .sdo(net4932), .r_o(net2047), .mode_o(net4940),
     .hiz_b_o(net2049), .glb_net_16(net4625[0:7]),
     .glb_net_15(net2995[0:7]), .glb_net_14(net3484[0:7]),
     .glb_net_13(net3973[0:7]), .glb_net_12(net3647[0:7]),
     .glb_net_11(net2669[0:7]), .glb_net_10(net2832[0:7]),
     .glb_net_09(net4136[0:7]), .glb_net_08(net2199[0:7]),
     .glb_net_07(net3810[0:7]), .glb_net_06(net3158[0:7]),
     .glb_net_05(net2506[0:7]), .glb_net_04(net4788[0:7]),
     .glb_net_03(net3321[0:7]), .glb_net_02(net4299[0:7]),
     .glb_net_01(net4462[0:7]), .bs_en_o(net2066), .bl_16(bl[869:816]),
     .bl_15(bl[815:762]), .bl_14(bl[761:708]), .bl_13(bl[707:654]),
     .bl_12(bl[653:600]), .bl_11(bl[599:546]), .bl_10(bl[545:492]),
     .bl_09(bl[491:438]), .bl_08(bl[437:396]), .bl_07(bl[395:342]),
     .bl_06(bl[341:288]), .bl_05(bl[287:234]), .bl_04(bl[233:180]),
     .bl_03(bl[179:126]), .bl_02(bl[125:72]), .bl_01(bl[71:18]),
     .sp12_v_b_10_33(net2805[0:23]), .slf_op_09_33(slf_op_09_33[3:0]),
     .sp4_v_b_10_33(net2910[0:47]), .lft_op_09_33(net2316[0:7]),
     .sp12_v_b_11_33(net2642[0:23]), .slf_op_10_33(slf_op_10_33[3:0]),
     .sp4_v_b_11_33(net2747[0:47]), .lft_op_10_33(net2184[0:7]),
     .sp12_v_b_12_33(net3620[0:23]), .slf_op_11_33(slf_op_11_33[3:0]),
     .sp4_v_b_12_33(net3725[0:47]), .lft_op_11_33(net2167[0:7]),
     .sp12_v_b_13_33(net3946[0:23]), .slf_op_12_33(slf_op_12_33[3:0]),
     .sp4_v_b_13_33(net4051[0:47]), .lft_op_12_33(net2643[0:7]),
     .sp12_v_b_14_33(net3457[0:23]), .slf_op_13_33(slf_op_13_33[3:0]),
     .sp4_v_b_14_33(net3562[0:47]), .lft_op_13_33(net2169[0:7]),
     .sp12_v_b_15_33(net2968[0:23]), .slf_op_14_33(slf_op_14_33[3:0]),
     .sp4_v_b_15_33(net3073[0:47]), .lft_op_14_33(net2188[0:7]),
     .sp12_v_b_16_33(net4598[0:23]), .slf_op_15_33(slf_op_15_33[3:0]),
     .sp4_v_b_16_33(net4703[0:47]), .lft_op_15_33(net3458[0:7]),
     .slf_op_16_33(slf_op_16_33[3:0]), .sp4_v_b_01_33(net4540[0:47]),
     .sp12_v_b_01_33(net4435[0:23]), .lft_op_16_33(slf_op_16_32[7:0]),
     .sp4_v_b_03_33(net3399[0:47]), .sp12_v_b_03_33(net3294[0:23]),
     .slf_op_02_33(slf_op_02_33[3:0]),
     .slf_op_04_33(slf_op_04_33[3:0]), .sp12_v_b_05_33(net2479[0:23]),
     .sp4_v_b_05_33(net2584[0:47]), .lft_op_04_33(net2160[0:7]),
     .lft_op_02_33(net4436[0:7]), .lft_op_05_33(net2179[0:7]),
     .sp4_v_b_06_33(net3236[0:47]), .sp12_v_b_07_33(net3783[0:23]),
     .sp4_v_b_04_33(net4866[0:47]), .sp12_v_b_04_33(net4761[0:23]),
     .slf_op_03_33(slf_op_03_33[3:0]), .lft_op_01_33(net2175[0:7]),
     .slf_op_01_33(slf_op_01_33[3:0]), .sp12_v_b_02_33(net4272[0:23]),
     .lft_op_03_33(net2177[0:7]), .sp4_v_b_02_33(net4377[0:47]),
     .slf_op_05_33(slf_op_05_33[3:0]), .sp12_v_b_06_33(net3131[0:23]),
     .lft_op_06_33(net2162[0:7]), .sp4_v_b_07_33(net3888[0:47]),
     .slf_op_06_33(slf_op_06_33[3:0]), .lft_op_08_33(net2164[0:7]),
     .sp4_v_b_09_33(net4214[0:47]), .slf_op_08_33(slf_op_08_33[3:0]),
     .sp12_v_b_09_33(net4109[0:23]), .lft_op_07_33(net2163[0:7]),
     .sp4_v_b_08_33(net2283[0:47]), .slf_op_07_33(slf_op_07_33[3:0]),
     .sp12_v_b_08_33(net2277[0:23]), .sp4_h_l_01_33(net2411[0:15]),
     .cf_top_l(cf_t[383:0]), .hold_t_l(hold_t_l),
     .padin_t_l(padin_t_l[29:0]), .padeb_t_l(padeb_t_l[29:0]),
     .pado_t_l(pado_t_l[29:0]),
     .end_of_startup_top_l(end_of_startup_top_l[16:1]),
     .padin_193(padin_193), .fabric_out_16_33(fabric_out_16_33),
     .fabric_out_15_33(fabric_out_15_33),
     .bnr_op_16_33(rgt_op_16_32[7:0]), .bnl_op_01_33({slf_op_00_32[3],
     slf_op_00_32[2], slf_op_00_32[1], slf_op_00_32[0],
     slf_op_00_32[3], slf_op_00_32[2], slf_op_00_32[1],
     slf_op_00_32[0]}));
array_LFT_IO_1x16top I_io_00top ( .sp4_v_b_00_17(sp4_v_b_00_17[15:0]),
     .sp4_v_t_00_32(net2411[0:15]), .ceb(ceb_o),
     .padin(padin_l_t[49:24]), .padeb(padeb_l_t[49:24]),
     .pado(pado_l_t[49:24]), .fabric_out_17(net4926),
     .fabric_out_18(net4957), .fabric_out_19(net4956),
     .fabric_out_20(net4970), .fabric_out_21(net4962),
     .fabric_out_22(net4972), .fabric_out_23(net4968),
     .fabric_out_24(net4963), .fabric_out_25(net4964),
     .fabric_out_26(net4965), .fabric_out_27(net4969),
     .fabric_out_28(net4966), .fabric_out_29(net4948),
     .fabric_out_30(net4967), .fabric_out_31(net5011),
     .fabric_out_32(net4971), .sdi(net2389),
     .tnl_op_00_32({slf_op_01_33[3], slf_op_01_33[2], slf_op_01_33[1],
     slf_op_01_33[0], slf_op_01_33[3], slf_op_01_33[2],
     slf_op_01_33[1], slf_op_01_33[0]}),
     .bnl_op_00_17(bnr_op_00_17[7:0]),
     .cdone_in(end_of_startup_lft_t[16:1]),
     .rgt_op_00_30(net2393[0:7]), .rgt_op_00_29(net2394[0:7]),
     .rgt_op_00_28(net2395[0:7]), .rgt_op_00_27(net2396[0:7]),
     .rgt_op_00_26(net2397[0:7]), .rgt_op_00_25(net2398[0:7]),
     .rgt_op_00_24(net2399[0:7]), .rgt_op_00_23(net2400[0:7]),
     .SP4_h_l_00_26(net2401[0:47]), .SP4_h_l_00_23(net2402[0:47]),
     .slf_op_00_29(slf_op_00_29[3:0]),
     .slf_op_00_28(slf_op_00_28[3:0]),
     .slf_op_00_27(slf_op_00_27[3:0]),
     .slf_op_00_26(slf_op_00_26[3:0]),
     .slf_op_00_25(slf_op_00_25[3:0]),
     .slf_op_00_24(slf_op_00_24[3:0]),
     .slf_op_00_23(slf_op_00_23[3:0]),
     .slf_op_00_22(slf_op_00_22[3:0]), .SP4_h_l_00_25(net2412[0:47]),
     .SP4_h_l_00_24(net2413[0:47]), .slf_op_00_17(slf_op_00_17[3:0]),
     .slf_op_00_18(slf_op_00_18[3:0]),
     .slf_op_00_19(slf_op_00_19[3:0]),
     .slf_op_00_20(slf_op_00_20[3:0]), .SP4_h_l_00_32(net2418[0:47]),
     .SP4_h_l_00_31(net2419[0:47]), .pgate(pgate_l[255:0]),
     .vdd_cntl(vdd_cntl_l[255:0]), .reset_b(reset_l[255:0]),
     .SP4_h_l_00_30(net2424[0:47]), .SP4_h_l_00_29(net2425[0:47]),
     .SP4_h_l_00_28(net2426[0:47]), .SP4_h_l_00_27(net2427[0:47]),
     .SP4_h_l_00_17(net2428[0:47]), .SP4_h_l_00_18(net2429[0:47]),
     .SP4_h_l_00_19(net2430[0:47]), .SP4_h_l_00_20(net2431[0:47]),
     .rgt_op_00_32(net2175[0:7]), .rgt_op_00_31(net2433[0:7]),
     .rgt_op_00_22(net2434[0:7]), .rgt_op_00_21(net2435[0:7]),
     .rgt_op_00_20(net2436[0:7]), .rgt_op_00_19(net2437[0:7]),
     .rgt_op_00_18(net2438[0:7]), .rgt_op_00_17(slf_op_01_17[7:0]),
     .SP4_h_l_00_21(net2440[0:47]), .SP4_h_l_00_22(net2441[0:47]),
     .slf_op_00_31(slf_op_00_31[3:0]),
     .slf_op_00_32(slf_op_00_32[3:0]),
     .slf_op_00_21(slf_op_00_21[3:0]), .SP12_h_l_00_32(net2445[0:23]),
     .SP12_h_l_00_31(net2446[0:23]), .SP12_h_l_00_30(net2447[0:23]),
     .SP12_h_l_00_29(net2448[0:23]), .SP12_h_l_00_28(net2449[0:23]),
     .SP12_h_l_00_27(net2450[0:23]), .SP12_h_l_00_26(net2451[0:23]),
     .SP12_h_l_00_25(net2452[0:23]), .SP12_h_l_00_24(net2453[0:23]),
     .SP12_h_l_00_23(net2454[0:23]), .SP12_h_l_00_22(net2455[0:23]),
     .SP12_h_l_00_21(net2456[0:23]), .SP12_h_l_00_20(net2457[0:23]),
     .SP12_h_l_00_18(net2458[0:23]), .SP12_h_l_00_19(net2459[0:23]),
     .SP12_h_l_00_17(net2460[0:23]), .slf_op_00_30(slf_op_00_30[3:0]),
     .wl(wl_l[255:0]), .shift(shift_o), .bs_en(bs_en_o), .mode(mode_o),
     .hiz_b(hiz_b_o), .prog(prog), .hold(hold_l_t), .update(update_o),
     .glb_netwk_col(clk_tree_drv[7:0]), .r(r_o),
     .spi_ss_in_b(net4979[0:31]), .sdo(sdo), .bl({bl[0], bl[1], bl[2],
     bl[3], bl[4], bl[5], bl[6], bl[7], bl[8], bl[9], bl[10], bl[11],
     bl[12], bl[13], bl[14], bl[15], bl[16], bl[17]}), .tclk(tclk_o),
     .cf_l(cf_l[383:0]), .spioeb({tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd}), .spiout({tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}));
array_BRAM_1x8top I_bram_08_top ( .glb_netwk(net2199[0:7]),
     .bm_sdo_o(bm_sdo_o), .bm_sweb_i(bm_sweb_i), .bm_sdi_i(bm_sdi_i),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sweb_o(bm_sweb_o),
     .bm_sclkrw_o(bm_sclkrw_o), .bm_sdi_o(bm_sdi_o),
     .bm_sdo_i(bm_sdo_i), .prog(prog),
     .glb_netwk_col(clk_tree_drv[7:0]),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bm_wdummymux_en_o(bm_wdummymux_en_o), .bm_sreb_o(bm_sreb_o),
     .bm_sclk_o(bm_sclk_o), .bm_sa_o(bm_sa_o[7:0]),
     .bm_rcapmux_en_o(bm_rcapmux_en_o), .bm_init_o(bm_init_o),
     .bl(bl[437:396]), .sp4_r_v_b_12(net2213[0:47]),
     .sp4_v_b_12(net3927[0:47]), .sp4_r_v_b_11(net2215[0:47]),
     .sp4_v_b_11(net3928[0:47]), .sp4_v_b_13(net3925[0:47]),
     .sp4_r_v_b_13(net2218[0:47]), .sp4_v_b_14(net3926[0:47]),
     .sp4_v_b_16(net3923[0:47]), .sp4_v_b_15(net3924[0:47]),
     .sp4_r_v_b_14(net2222[0:47]), .sp4_r_v_b_15(net2223[0:47]),
     .sp4_r_v_b_16(net2224[0:47]), .sp12_h_l_13(net3939[0:23]),
     .sp12_h_r_13(net2226[0:23]), .sp12_h_l_12(net3938[0:23]),
     .sp12_h_r_12(net2228[0:23]), .sp12_h_r_15(net2229[0:23]),
     .sp12_h_l_15(net3937[0:23]), .sp12_h_r_16(net2231[0:23]),
     .sp12_h_l_16(net3935[0:23]), .sp12_h_l_14(net3936[0:23]),
     .sp12_h_l_11(net3940[0:23]), .sp12_h_r_14(net2235[0:23]),
     .sp12_h_r_11(net2236[0:23]), .sp4_h_l_05(net3845[0:47]),
     .sp4_h_r_05(net2238[0:47]), .sp4_h_l_06(net3844[0:47]),
     .sp4_h_r_06(net2240[0:47]), .sp4_h_l_01(net3820[0:47]),
     .sp4_h_l_02(net3819[0:47]), .sp4_h_l_03(net3818[0:47]),
     .sp4_h_l_04(net3817[0:47]), .sp4_h_r_01(net2245[0:47]),
     .sp4_h_r_02(net2246[0:47]), .sp4_h_r_03(net2247[0:47]),
     .sp4_h_r_04(net2248[0:47]), .slf_op_05(net3857[0:7]),
     .rgt_op_06(net2250[0:7]), .rgt_op_05(net2251[0:7]),
     .slf_op_06(net3856[0:7]), .slf_op_01(slf_op_08_17[7:0]),
     .slf_op_02(net3788[0:7]), .slf_op_03(net3786[0:7]),
     .slf_op_04(net3796[0:7]), .rgt_op_04(net2257[0:7]),
     .rgt_op_01(slf_op_09_17[7:0]), .rgt_op_02(net2259[0:7]),
     .rgt_op_03(net2260[0:7]), .top_op_16({slf_op_08_33[3],
     slf_op_08_33[2], slf_op_08_33[1], slf_op_08_33[0],
     slf_op_08_33[3], slf_op_08_33[2], slf_op_08_33[1],
     slf_op_08_33[0]}), .bot_op_01(bot_op_08_17[7:0]),
     .tnr_op_16({slf_op_09_33[3], slf_op_09_33[2], slf_op_09_33[1],
     slf_op_09_33[0], slf_op_09_33[3], slf_op_09_33[2],
     slf_op_09_33[1], slf_op_09_33[0]}), .tnl_op_16({slf_op_07_33[3],
     slf_op_07_33[2], slf_op_07_33[1], slf_op_07_33[0],
     slf_op_07_33[3], slf_op_07_33[2], slf_op_07_33[1],
     slf_op_07_33[0]}), .rgt_op_09(net2265[0:7]),
     .rgt_op_08(net2266[0:7]), .rgt_op_07(net2267[0:7]),
     .rgt_op_10(net2268[0:7]), .lft_op_04(net3144[0:7]),
     .lft_op_03(net3134[0:7]), .lft_op_02(net3136[0:7]),
     .lft_op_01(slf_op_07_17[7:0]), .bnl_op_01(bnl_op_08_17[7:0]),
     .pgate(pgate_l[255:0]), .wl(wl_l[255:0]),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_t_16(net2277[0:23]),
     .sp12_v_b_01(sp12_v_b_08_17[23:0]), .sp12_h_r_04(net2279[0:23]),
     .sp12_h_r_02(net2280[0:23]), .sp12_h_r_10(net2281[0:23]),
     .sp12_h_r_01(net2282[0:23]), .sp4_v_t_16(net2283[0:47]),
     .sp4_v_b_01(sp4_v_b_08_17[47:0]), .sp4_r_v_b_10(net2285[0:47]),
     .sp4_r_v_b_09(net2286[0:47]), .sp4_r_v_b_08(net2287[0:47]),
     .sp4_r_v_b_07(net2288[0:47]), .sp4_h_r_10(net2289[0:47]),
     .sp4_h_r_09(net2290[0:47]), .sp4_h_r_08(net2291[0:47]),
     .sp4_h_r_07(net2292[0:47]), .sp4_h_l_10(net3840[0:47]),
     .sp4_h_l_09(net3841[0:47]), .sp4_h_l_08(net3842[0:47]),
     .sp4_h_l_07(net3843[0:47]), .reset_b(reset_l[255:0]),
     .slf_op_10(net3852[0:7]), .slf_op_09(net3853[0:7]),
     .slf_op_08(net3854[0:7]), .slf_op_07(net3855[0:7]),
     .slf_op_16(net2164[0:7]), .sp12_h_l_01(net3809[0:23]),
     .sp12_h_l_02(net3808[0:23]), .sp12_h_l_04(net3806[0:23]),
     .sp12_h_l_03(net3807[0:23]), .sp4_v_b_07(net3878[0:47]),
     .lft_op_10(net3200[0:7]), .lft_op_09(net3201[0:7]),
     .lft_op_05(net3205[0:7]), .lft_op_06(net3204[0:7]),
     .lft_op_07(net3203[0:7]), .lft_op_08(net3202[0:7]),
     .sp4_v_b_05(net3876[0:47]), .sp4_r_v_b_05(net2315[0:47]),
     .rgt_op_16(net2316[0:7]), .rgt_op_15(net2317[0:7]),
     .sp4_v_b_06(net3877[0:47]), .sp4_r_v_b_06(net2319[0:47]),
     .sp4_r_v_b_04(net2320[0:47]), .sp4_v_b_04(net3813[0:47]),
     .sp4_r_v_b_03(net2322[0:47]), .sp4_v_b_03(net3814[0:47]),
     .sp4_r_v_b_02(net2324[0:47]), .sp4_v_b_02(net3815[0:47]),
     .sp4_r_v_b_01(sp4_v_b_09_17[47:0]), .slf_op_15(net3913[0:7]),
     .slf_op_12(net3914[0:7]), .slf_op_13(net3915[0:7]),
     .rgt_op_11(net2330[0:7]), .rgt_op_12(net2331[0:7]),
     .rgt_op_13(net2332[0:7]), .rgt_op_14(net2333[0:7]),
     .sp4_h_l_15(net3895[0:47]), .sp4_h_r_15(net2335[0:47]),
     .sp4_h_l_16(net3896[0:47]), .sp4_h_r_16(net2337[0:47]),
     .sp4_h_r_14(net2338[0:47]), .sp4_h_l_14(net3894[0:47]),
     .sp4_h_r_13(net2340[0:47]), .sp4_h_l_13(net3893[0:47]),
     .sp12_h_r_07(net2342[0:23]), .sp4_h_r_12(net2343[0:47]),
     .sp4_h_l_12(net3892[0:47]), .sp12_h_l_05(net3870[0:23]),
     .sp4_h_r_11(net2346[0:47]), .sp12_h_l_08(net3873[0:23]),
     .sp4_h_l_11(net3891[0:47]), .sp12_h_r_03(net2349[0:23]),
     .sp12_h_l_10(net3865[0:23]), .sp12_h_r_09(net2351[0:23]),
     .sp12_h_l_09(net3874[0:23]), .sp12_h_r_08(net2353[0:23]),
     .sp12_h_r_05(net2354[0:23]), .sp12_h_l_06(net3871[0:23]),
     .sp12_h_r_06(net2356[0:23]), .bnr_op_01(bnr_op_08_17[7:0]),
     .lft_op_16(net2163[0:7]), .slf_op_14(net3912[0:7]),
     .slf_op_11(net3916[0:7]), .sp4_v_b_09(net3880[0:47]),
     .sp4_v_b_10(net3881[0:47]), .sp4_v_b_08(net3879[0:47]),
     .sp12_h_l_07(net3872[0:23]), .lft_op_14(net3260[0:7]),
     .lft_op_13(net3263[0:7]), .lft_op_12(net3262[0:7]),
     .lft_op_11(net3264[0:7]), .lft_op_15(net3261[0:7]));
array_LT1x16top I_it_05_top ( .glb_netwk(net2506[0:7]),
     .sp12_v_t_16(net2479[0:23]), .rgt_op_16(net2162[0:7]),
     .top_op_16({slf_op_05_33[3], slf_op_05_33[2], slf_op_05_33[1],
     slf_op_05_33[0], slf_op_05_33[3], slf_op_05_33[2],
     slf_op_05_33[1], slf_op_05_33[0]}), .rgt_op_03(net2482[0:7]),
     .slf_op_02(net4766[0:7]), .rgt_op_02(net2484[0:7]),
     .rgt_op_01(slf_op_06_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3307[0:7]), .lft_op_03(net3297[0:7]),
     .lft_op_02(net3299[0:7]), .lft_op_01(slf_op_04_17[7:0]),
     .rgt_op_04(net2492[0:7]), .carry_in(carry_in_05_17),
     .bnl_op_01(bnl_op_05_17[7:0]), .slf_op_04(net4774[0:7]),
     .slf_op_03(net4764[0:7]), .slf_op_01(slf_op_05_17[7:0]),
     .sp4_h_l_04(net4795[0:47]), .carry_out(net2499),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_05_17[23:0]),
     .sp12_h_r_04(net2502[0:23]), .sp12_h_r_03(net2503[0:23]),
     .sp12_h_r_02(net2504[0:23]), .sp12_h_r_01(net2505[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2179[0:7]),
     .sp4_v_b_01(sp4_v_b_05_17[47:0]), .sp4_r_v_b_04(net2509[0:47]),
     .sp4_r_v_b_03(net2510[0:47]), .sp4_r_v_b_02(net2511[0:47]),
     .sp4_r_v_b_01(sp4_v_b_06_17[47:0]), .sp4_h_r_04(net2513[0:47]),
     .sp4_h_r_03(net2514[0:47]), .sp4_h_r_02(net2515[0:47]),
     .sp4_h_r_01(net2516[0:47]), .sp4_h_l_03(net4796[0:47]),
     .sp4_h_l_02(net4797[0:47]), .sp4_h_l_01(net4798[0:47]),
     .bl(bl[287:234]), .bot_op_01(bot_op_05_17[7:0]),
     .sp12_h_l_01(net4787[0:23]), .sp12_h_l_02(net4786[0:23]),
     .sp12_h_l_03(net4785[0:23]), .sp12_h_l_04(net4784[0:23]),
     .sp4_v_b_04(net4791[0:47]), .sp4_v_b_03(net4792[0:47]),
     .sp4_v_b_02(net4793[0:47]), .bnr_op_01(bnr_op_05_17[7:0]),
     .sp4_h_l_05(net4823[0:47]), .sp4_h_l_06(net4822[0:47]),
     .sp4_h_l_07(net4821[0:47]), .sp4_h_l_08(net4820[0:47]),
     .sp4_h_l_09(net4819[0:47]), .sp4_h_l_10(net4818[0:47]),
     .sp4_h_r_10(net2536[0:47]), .sp4_h_r_09(net2537[0:47]),
     .sp4_h_r_08(net2538[0:47]), .sp4_h_r_07(net2539[0:47]),
     .sp4_h_r_06(net2540[0:47]), .sp4_h_r_05(net2541[0:47]),
     .slf_op_05(net4835[0:7]), .slf_op_06(net4834[0:7]),
     .slf_op_07(net4833[0:7]), .slf_op_08(net4832[0:7]),
     .slf_op_09(net4831[0:7]), .slf_op_10(net4830[0:7]),
     .rgt_op_10(net2548[0:7]), .rgt_op_09(net2549[0:7]),
     .rgt_op_08(net2550[0:7]), .rgt_op_07(net2551[0:7]),
     .rgt_op_06(net2552[0:7]), .rgt_op_05(net2553[0:7]),
     .lft_op_10(net3363[0:7]), .lft_op_09(net3364[0:7]),
     .lft_op_08(net3365[0:7]), .lft_op_07(net3366[0:7]),
     .lft_op_06(net3367[0:7]), .lft_op_05(net3368[0:7]),
     .sp12_h_l_10(net4843[0:23]), .sp12_h_r_10(net2561[0:23]),
     .sp12_h_l_09(net4852[0:23]), .sp12_h_l_08(net4851[0:23]),
     .sp12_h_l_07(net4850[0:23]), .sp12_h_l_06(net4849[0:23]),
     .sp12_h_r_05(net2566[0:23]), .sp12_h_r_06(net2567[0:23]),
     .sp12_h_r_07(net2568[0:23]), .sp12_h_r_08(net2569[0:23]),
     .sp12_h_r_09(net2570[0:23]), .sp12_h_l_05(net4848[0:23]),
     .sp4_r_v_b_05(net2572[0:47]), .sp4_r_v_b_06(net2573[0:47]),
     .sp4_r_v_b_07(net2574[0:47]), .sp4_r_v_b_08(net2575[0:47]),
     .sp4_r_v_b_09(net2576[0:47]), .sp4_r_v_b_10(net2577[0:47]),
     .sp4_v_b_10(net4859[0:47]), .sp4_v_b_09(net4858[0:47]),
     .sp4_v_b_08(net4857[0:47]), .sp4_v_b_07(net4856[0:47]),
     .sp4_v_b_06(net4855[0:47]), .sp4_v_b_05(net4854[0:47]),
     .sp4_v_t_16(net2584[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net2587[0:47]),
     .sp4_h_r_12(net2588[0:47]), .sp4_h_r_13(net2589[0:47]),
     .sp4_h_r_14(net2590[0:47]), .sp4_h_r_15(net2591[0:47]),
     .sp4_h_r_16(net2592[0:47]), .sp4_h_l_16(net4874[0:47]),
     .sp4_h_l_15(net4873[0:47]), .sp4_h_l_14(net4872[0:47]),
     .sp4_h_l_13(net4871[0:47]), .sp4_h_l_12(net4870[0:47]),
     .sp4_h_l_11(net4869[0:47]), .tnr_op_16({slf_op_06_33[3],
     slf_op_06_33[2], slf_op_06_33[1], slf_op_06_33[0],
     slf_op_06_33[3], slf_op_06_33[2], slf_op_06_33[1],
     slf_op_06_33[0]}), .tnl_op_16({slf_op_04_33[3], slf_op_04_33[2],
     slf_op_04_33[1], slf_op_04_33[0], slf_op_04_33[3],
     slf_op_04_33[2], slf_op_04_33[1], slf_op_04_33[0]}),
     .lft_op_16(net2160[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net4891[0:7]), .slf_op_14(net4890[0:7]),
     .slf_op_13(net4893[0:7]), .slf_op_12(net4892[0:7]),
     .slf_op_11(net4894[0:7]), .rgt_op_14(net2608[0:7]),
     .rgt_op_15(net2609[0:7]), .rgt_op_12(net2610[0:7]),
     .rgt_op_13(net2611[0:7]), .rgt_op_11(net2612[0:7]),
     .sp4_v_b_16(net4901[0:47]), .sp4_v_b_14(net4904[0:47]),
     .sp4_v_b_15(net4902[0:47]), .sp4_v_b_13(net4903[0:47]),
     .sp4_v_b_11(net4906[0:47]), .sp4_v_b_12(net4905[0:47]),
     .sp4_r_v_b_16(net2619[0:47]), .sp4_r_v_b_15(net2620[0:47]),
     .sp4_r_v_b_13(net2621[0:47]), .sp4_r_v_b_14(net2622[0:47]),
     .sp4_r_v_b_12(net2623[0:47]), .sp4_r_v_b_11(net2624[0:47]),
     .sp12_h_l_16(net4913[0:23]), .sp12_h_l_15(net4915[0:23]),
     .sp12_h_l_14(net4914[0:23]), .sp12_h_l_13(net4917[0:23]),
     .sp12_h_l_12(net4916[0:23]), .sp12_h_l_11(net4918[0:23]),
     .sp12_h_r_16(net2631[0:23]), .sp12_h_r_14(net2632[0:23]),
     .sp12_h_r_15(net2633[0:23]), .sp12_h_r_12(net2634[0:23]),
     .sp12_h_r_13(net2635[0:23]), .sp12_h_r_11(net2636[0:23]),
     .lft_op_14(net3423[0:7]), .lft_op_15(net3424[0:7]),
     .lft_op_12(net3425[0:7]), .lft_op_11(net3427[0:7]),
     .lft_op_13(net3426[0:7]));
array_LT1x16top I_it_11_top ( .glb_netwk(net2669[0:7]),
     .sp12_v_t_16(net2642[0:23]), .rgt_op_16(net2643[0:7]),
     .top_op_16({slf_op_11_33[3], slf_op_11_33[2], slf_op_11_33[1],
     slf_op_11_33[0], slf_op_11_33[3], slf_op_11_33[2],
     slf_op_11_33[1], slf_op_11_33[0]}), .rgt_op_03(net2645[0:7]),
     .slf_op_02(net2810[0:7]), .rgt_op_02(net2647[0:7]),
     .rgt_op_01(slf_op_12_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4122[0:7]), .lft_op_03(net4112[0:7]),
     .lft_op_02(net4114[0:7]), .lft_op_01(slf_op_10_17[7:0]),
     .rgt_op_04(net2655[0:7]), .carry_in(carry_in_11_17),
     .bnl_op_01(bnl_op_11_17[7:0]), .slf_op_04(net2818[0:7]),
     .slf_op_03(net2808[0:7]), .slf_op_01(slf_op_11_17[7:0]),
     .sp4_h_l_04(net2839[0:47]), .carry_out(net2662),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_11_17[23:0]),
     .sp12_h_r_04(net2665[0:23]), .sp12_h_r_03(net2666[0:23]),
     .sp12_h_r_02(net2667[0:23]), .sp12_h_r_01(net2668[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2167[0:7]),
     .sp4_v_b_01(sp4_v_b_11_17[47:0]), .sp4_r_v_b_04(net2672[0:47]),
     .sp4_r_v_b_03(net2673[0:47]), .sp4_r_v_b_02(net2674[0:47]),
     .sp4_r_v_b_01(sp4_v_b_12_17[47:0]), .sp4_h_r_04(net2676[0:47]),
     .sp4_h_r_03(net2677[0:47]), .sp4_h_r_02(net2678[0:47]),
     .sp4_h_r_01(net2679[0:47]), .sp4_h_l_03(net2840[0:47]),
     .sp4_h_l_02(net2841[0:47]), .sp4_h_l_01(net2842[0:47]),
     .bl(bl[599:546]), .bot_op_01(bot_op_11_17[7:0]),
     .sp12_h_l_01(net2831[0:23]), .sp12_h_l_02(net2830[0:23]),
     .sp12_h_l_03(net2829[0:23]), .sp12_h_l_04(net2828[0:23]),
     .sp4_v_b_04(net2835[0:47]), .sp4_v_b_03(net2836[0:47]),
     .sp4_v_b_02(net2837[0:47]), .bnr_op_01(bnr_op_11_17[7:0]),
     .sp4_h_l_05(net2867[0:47]), .sp4_h_l_06(net2866[0:47]),
     .sp4_h_l_07(net2865[0:47]), .sp4_h_l_08(net2864[0:47]),
     .sp4_h_l_09(net2863[0:47]), .sp4_h_l_10(net2862[0:47]),
     .sp4_h_r_10(net2699[0:47]), .sp4_h_r_09(net2700[0:47]),
     .sp4_h_r_08(net2701[0:47]), .sp4_h_r_07(net2702[0:47]),
     .sp4_h_r_06(net2703[0:47]), .sp4_h_r_05(net2704[0:47]),
     .slf_op_05(net2879[0:7]), .slf_op_06(net2878[0:7]),
     .slf_op_07(net2877[0:7]), .slf_op_08(net2876[0:7]),
     .slf_op_09(net2875[0:7]), .slf_op_10(net2874[0:7]),
     .rgt_op_10(net2711[0:7]), .rgt_op_09(net2712[0:7]),
     .rgt_op_08(net2713[0:7]), .rgt_op_07(net2714[0:7]),
     .rgt_op_06(net2715[0:7]), .rgt_op_05(net2716[0:7]),
     .lft_op_10(net4178[0:7]), .lft_op_09(net4179[0:7]),
     .lft_op_08(net4180[0:7]), .lft_op_07(net4181[0:7]),
     .lft_op_06(net4182[0:7]), .lft_op_05(net4183[0:7]),
     .sp12_h_l_10(net2887[0:23]), .sp12_h_r_10(net2724[0:23]),
     .sp12_h_l_09(net2896[0:23]), .sp12_h_l_08(net2895[0:23]),
     .sp12_h_l_07(net2894[0:23]), .sp12_h_l_06(net2893[0:23]),
     .sp12_h_r_05(net2729[0:23]), .sp12_h_r_06(net2730[0:23]),
     .sp12_h_r_07(net2731[0:23]), .sp12_h_r_08(net2732[0:23]),
     .sp12_h_r_09(net2733[0:23]), .sp12_h_l_05(net2892[0:23]),
     .sp4_r_v_b_05(net2735[0:47]), .sp4_r_v_b_06(net2736[0:47]),
     .sp4_r_v_b_07(net2737[0:47]), .sp4_r_v_b_08(net2738[0:47]),
     .sp4_r_v_b_09(net2739[0:47]), .sp4_r_v_b_10(net2740[0:47]),
     .sp4_v_b_10(net2903[0:47]), .sp4_v_b_09(net2902[0:47]),
     .sp4_v_b_08(net2901[0:47]), .sp4_v_b_07(net2900[0:47]),
     .sp4_v_b_06(net2899[0:47]), .sp4_v_b_05(net2898[0:47]),
     .sp4_v_t_16(net2747[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net2750[0:47]),
     .sp4_h_r_12(net2751[0:47]), .sp4_h_r_13(net2752[0:47]),
     .sp4_h_r_14(net2753[0:47]), .sp4_h_r_15(net2754[0:47]),
     .sp4_h_r_16(net2755[0:47]), .sp4_h_l_16(net2918[0:47]),
     .sp4_h_l_15(net2917[0:47]), .sp4_h_l_14(net2916[0:47]),
     .sp4_h_l_13(net2915[0:47]), .sp4_h_l_12(net2914[0:47]),
     .sp4_h_l_11(net2913[0:47]), .tnr_op_16({slf_op_12_33[3],
     slf_op_12_33[2], slf_op_12_33[1], slf_op_12_33[0],
     slf_op_12_33[3], slf_op_12_33[2], slf_op_12_33[1],
     slf_op_12_33[0]}), .tnl_op_16({slf_op_10_33[3], slf_op_10_33[2],
     slf_op_10_33[1], slf_op_10_33[0], slf_op_10_33[3],
     slf_op_10_33[2], slf_op_10_33[1], slf_op_10_33[0]}),
     .lft_op_16(net2184[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net2935[0:7]), .slf_op_14(net2934[0:7]),
     .slf_op_13(net2937[0:7]), .slf_op_12(net2936[0:7]),
     .slf_op_11(net2938[0:7]), .rgt_op_14(net2771[0:7]),
     .rgt_op_15(net2772[0:7]), .rgt_op_12(net2773[0:7]),
     .rgt_op_13(net2774[0:7]), .rgt_op_11(net2775[0:7]),
     .sp4_v_b_16(net2945[0:47]), .sp4_v_b_14(net2948[0:47]),
     .sp4_v_b_15(net2946[0:47]), .sp4_v_b_13(net2947[0:47]),
     .sp4_v_b_11(net2950[0:47]), .sp4_v_b_12(net2949[0:47]),
     .sp4_r_v_b_16(net2782[0:47]), .sp4_r_v_b_15(net2783[0:47]),
     .sp4_r_v_b_13(net2784[0:47]), .sp4_r_v_b_14(net2785[0:47]),
     .sp4_r_v_b_12(net2786[0:47]), .sp4_r_v_b_11(net2787[0:47]),
     .sp12_h_l_16(net2957[0:23]), .sp12_h_l_15(net2959[0:23]),
     .sp12_h_l_14(net2958[0:23]), .sp12_h_l_13(net2961[0:23]),
     .sp12_h_l_12(net2960[0:23]), .sp12_h_l_11(net2962[0:23]),
     .sp12_h_r_16(net2794[0:23]), .sp12_h_r_14(net2795[0:23]),
     .sp12_h_r_15(net2796[0:23]), .sp12_h_r_12(net2797[0:23]),
     .sp12_h_r_13(net2798[0:23]), .sp12_h_r_11(net2799[0:23]),
     .lft_op_14(net4238[0:7]), .lft_op_15(net4239[0:7]),
     .lft_op_12(net4240[0:7]), .lft_op_11(net4242[0:7]),
     .lft_op_13(net4241[0:7]));
array_LT1x16top I_it_10_top ( .glb_netwk(net2832[0:7]),
     .sp12_v_t_16(net2805[0:23]), .rgt_op_16(net2167[0:7]),
     .top_op_16({slf_op_10_33[3], slf_op_10_33[2], slf_op_10_33[1],
     slf_op_10_33[0], slf_op_10_33[3], slf_op_10_33[2],
     slf_op_10_33[1], slf_op_10_33[0]}), .rgt_op_03(net2808[0:7]),
     .slf_op_02(net4114[0:7]), .rgt_op_02(net2810[0:7]),
     .rgt_op_01(slf_op_11_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2257[0:7]), .lft_op_03(net2260[0:7]),
     .lft_op_02(net2259[0:7]), .lft_op_01(slf_op_09_17[7:0]),
     .rgt_op_04(net2818[0:7]), .carry_in(carry_in_10_17),
     .bnl_op_01(bnl_op_10_17[7:0]), .slf_op_04(net4122[0:7]),
     .slf_op_03(net4112[0:7]), .slf_op_01(slf_op_10_17[7:0]),
     .sp4_h_l_04(net4143[0:47]), .carry_out(net2825),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_10_17[23:0]),
     .sp12_h_r_04(net2828[0:23]), .sp12_h_r_03(net2829[0:23]),
     .sp12_h_r_02(net2830[0:23]), .sp12_h_r_01(net2831[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2184[0:7]),
     .sp4_v_b_01(sp4_v_b_10_17[47:0]), .sp4_r_v_b_04(net2835[0:47]),
     .sp4_r_v_b_03(net2836[0:47]), .sp4_r_v_b_02(net2837[0:47]),
     .sp4_r_v_b_01(sp4_v_b_11_17[47:0]), .sp4_h_r_04(net2839[0:47]),
     .sp4_h_r_03(net2840[0:47]), .sp4_h_r_02(net2841[0:47]),
     .sp4_h_r_01(net2842[0:47]), .sp4_h_l_03(net4144[0:47]),
     .sp4_h_l_02(net4145[0:47]), .sp4_h_l_01(net4146[0:47]),
     .bl(bl[545:492]), .bot_op_01(bot_op_10_17[7:0]),
     .sp12_h_l_01(net4135[0:23]), .sp12_h_l_02(net4134[0:23]),
     .sp12_h_l_03(net4133[0:23]), .sp12_h_l_04(net4132[0:23]),
     .sp4_v_b_04(net4139[0:47]), .sp4_v_b_03(net4140[0:47]),
     .sp4_v_b_02(net4141[0:47]), .bnr_op_01(bnr_op_10_17[7:0]),
     .sp4_h_l_05(net4171[0:47]), .sp4_h_l_06(net4170[0:47]),
     .sp4_h_l_07(net4169[0:47]), .sp4_h_l_08(net4168[0:47]),
     .sp4_h_l_09(net4167[0:47]), .sp4_h_l_10(net4166[0:47]),
     .sp4_h_r_10(net2862[0:47]), .sp4_h_r_09(net2863[0:47]),
     .sp4_h_r_08(net2864[0:47]), .sp4_h_r_07(net2865[0:47]),
     .sp4_h_r_06(net2866[0:47]), .sp4_h_r_05(net2867[0:47]),
     .slf_op_05(net4183[0:7]), .slf_op_06(net4182[0:7]),
     .slf_op_07(net4181[0:7]), .slf_op_08(net4180[0:7]),
     .slf_op_09(net4179[0:7]), .slf_op_10(net4178[0:7]),
     .rgt_op_10(net2874[0:7]), .rgt_op_09(net2875[0:7]),
     .rgt_op_08(net2876[0:7]), .rgt_op_07(net2877[0:7]),
     .rgt_op_06(net2878[0:7]), .rgt_op_05(net2879[0:7]),
     .lft_op_10(net2268[0:7]), .lft_op_09(net2265[0:7]),
     .lft_op_08(net2266[0:7]), .lft_op_07(net2267[0:7]),
     .lft_op_06(net2250[0:7]), .lft_op_05(net2251[0:7]),
     .sp12_h_l_10(net4191[0:23]), .sp12_h_r_10(net2887[0:23]),
     .sp12_h_l_09(net4200[0:23]), .sp12_h_l_08(net4199[0:23]),
     .sp12_h_l_07(net4198[0:23]), .sp12_h_l_06(net4197[0:23]),
     .sp12_h_r_05(net2892[0:23]), .sp12_h_r_06(net2893[0:23]),
     .sp12_h_r_07(net2894[0:23]), .sp12_h_r_08(net2895[0:23]),
     .sp12_h_r_09(net2896[0:23]), .sp12_h_l_05(net4196[0:23]),
     .sp4_r_v_b_05(net2898[0:47]), .sp4_r_v_b_06(net2899[0:47]),
     .sp4_r_v_b_07(net2900[0:47]), .sp4_r_v_b_08(net2901[0:47]),
     .sp4_r_v_b_09(net2902[0:47]), .sp4_r_v_b_10(net2903[0:47]),
     .sp4_v_b_10(net4207[0:47]), .sp4_v_b_09(net4206[0:47]),
     .sp4_v_b_08(net4205[0:47]), .sp4_v_b_07(net4204[0:47]),
     .sp4_v_b_06(net4203[0:47]), .sp4_v_b_05(net4202[0:47]),
     .sp4_v_t_16(net2910[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net2913[0:47]),
     .sp4_h_r_12(net2914[0:47]), .sp4_h_r_13(net2915[0:47]),
     .sp4_h_r_14(net2916[0:47]), .sp4_h_r_15(net2917[0:47]),
     .sp4_h_r_16(net2918[0:47]), .sp4_h_l_16(net4222[0:47]),
     .sp4_h_l_15(net4221[0:47]), .sp4_h_l_14(net4220[0:47]),
     .sp4_h_l_13(net4219[0:47]), .sp4_h_l_12(net4218[0:47]),
     .sp4_h_l_11(net4217[0:47]), .tnr_op_16({slf_op_11_33[3],
     slf_op_11_33[2], slf_op_11_33[1], slf_op_11_33[0],
     slf_op_11_33[3], slf_op_11_33[2], slf_op_11_33[1],
     slf_op_11_33[0]}), .tnl_op_16({slf_op_09_33[3], slf_op_09_33[2],
     slf_op_09_33[1], slf_op_09_33[0], slf_op_09_33[3],
     slf_op_09_33[2], slf_op_09_33[1], slf_op_09_33[0]}),
     .lft_op_16(net2316[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net4239[0:7]), .slf_op_14(net4238[0:7]),
     .slf_op_13(net4241[0:7]), .slf_op_12(net4240[0:7]),
     .slf_op_11(net4242[0:7]), .rgt_op_14(net2934[0:7]),
     .rgt_op_15(net2935[0:7]), .rgt_op_12(net2936[0:7]),
     .rgt_op_13(net2937[0:7]), .rgt_op_11(net2938[0:7]),
     .sp4_v_b_16(net4249[0:47]), .sp4_v_b_14(net4252[0:47]),
     .sp4_v_b_15(net4250[0:47]), .sp4_v_b_13(net4251[0:47]),
     .sp4_v_b_11(net4254[0:47]), .sp4_v_b_12(net4253[0:47]),
     .sp4_r_v_b_16(net2945[0:47]), .sp4_r_v_b_15(net2946[0:47]),
     .sp4_r_v_b_13(net2947[0:47]), .sp4_r_v_b_14(net2948[0:47]),
     .sp4_r_v_b_12(net2949[0:47]), .sp4_r_v_b_11(net2950[0:47]),
     .sp12_h_l_16(net4261[0:23]), .sp12_h_l_15(net4263[0:23]),
     .sp12_h_l_14(net4262[0:23]), .sp12_h_l_13(net4265[0:23]),
     .sp12_h_l_12(net4264[0:23]), .sp12_h_l_11(net4266[0:23]),
     .sp12_h_r_16(net2957[0:23]), .sp12_h_r_14(net2958[0:23]),
     .sp12_h_r_15(net2959[0:23]), .sp12_h_r_12(net2960[0:23]),
     .sp12_h_r_13(net2961[0:23]), .sp12_h_r_11(net2962[0:23]),
     .lft_op_14(net2333[0:7]), .lft_op_15(net2317[0:7]),
     .lft_op_12(net2331[0:7]), .lft_op_11(net2330[0:7]),
     .lft_op_13(net2332[0:7]));
array_LT1x16top I_it_15_top ( .glb_netwk(net2995[0:7]),
     .sp12_v_t_16(net2968[0:23]), .rgt_op_16(slf_op_16_32[7:0]),
     .top_op_16({slf_op_15_33[3], slf_op_15_33[2], slf_op_15_33[1],
     slf_op_15_33[0], slf_op_15_33[3], slf_op_15_33[2],
     slf_op_15_33[1], slf_op_15_33[0]}), .rgt_op_03(slf_op_16_19[7:0]),
     .slf_op_02(net3462[0:7]), .rgt_op_02(slf_op_16_18[7:0]),
     .rgt_op_01(slf_op_16_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3959[0:7]), .lft_op_03(net3949[0:7]),
     .lft_op_02(net3951[0:7]), .lft_op_01(slf_op_14_17[7:0]),
     .rgt_op_04(slf_op_16_20[7:0]), .carry_in(carry_in_15_17),
     .bnl_op_01(bnl_op_15_17[7:0]), .slf_op_04(net3470[0:7]),
     .slf_op_03(net3460[0:7]), .slf_op_01(slf_op_15_17[7:0]),
     .sp4_h_l_04(net3491[0:47]), .carry_out(net2988),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_15_17[23:0]),
     .sp12_h_r_04(net2991[0:23]), .sp12_h_r_03(net2992[0:23]),
     .sp12_h_r_02(net2993[0:23]), .sp12_h_r_01(net2994[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net3458[0:7]),
     .sp4_v_b_01(sp4_v_b_15_17[47:0]), .sp4_r_v_b_04(net2998[0:47]),
     .sp4_r_v_b_03(net2999[0:47]), .sp4_r_v_b_02(net3000[0:47]),
     .sp4_r_v_b_01(sp4_v_b_16_17[47:0]), .sp4_h_r_04(net3002[0:47]),
     .sp4_h_r_03(net3003[0:47]), .sp4_h_r_02(net3004[0:47]),
     .sp4_h_r_01(net3005[0:47]), .sp4_h_l_03(net3492[0:47]),
     .sp4_h_l_02(net3493[0:47]), .sp4_h_l_01(net3494[0:47]),
     .bl(bl[815:762]), .bot_op_01(bot_op_15_17[7:0]),
     .sp12_h_l_01(net3483[0:23]), .sp12_h_l_02(net3482[0:23]),
     .sp12_h_l_03(net3481[0:23]), .sp12_h_l_04(net3480[0:23]),
     .sp4_v_b_04(net3487[0:47]), .sp4_v_b_03(net3488[0:47]),
     .sp4_v_b_02(net3489[0:47]), .bnr_op_01(bnr_op_15_17[7:0]),
     .sp4_h_l_05(net3519[0:47]), .sp4_h_l_06(net3518[0:47]),
     .sp4_h_l_07(net3517[0:47]), .sp4_h_l_08(net3516[0:47]),
     .sp4_h_l_09(net3515[0:47]), .sp4_h_l_10(net3514[0:47]),
     .sp4_h_r_10(net3025[0:47]), .sp4_h_r_09(net3026[0:47]),
     .sp4_h_r_08(net3027[0:47]), .sp4_h_r_07(net3028[0:47]),
     .sp4_h_r_06(net3029[0:47]), .sp4_h_r_05(net3030[0:47]),
     .slf_op_05(net3531[0:7]), .slf_op_06(net3530[0:7]),
     .slf_op_07(net3529[0:7]), .slf_op_08(net3528[0:7]),
     .slf_op_09(net3527[0:7]), .slf_op_10(net3526[0:7]),
     .rgt_op_10(slf_op_16_26[7:0]), .rgt_op_09(slf_op_16_25[7:0]),
     .rgt_op_08(slf_op_16_24[7:0]), .rgt_op_07(slf_op_16_23[7:0]),
     .rgt_op_06(slf_op_16_22[7:0]), .rgt_op_05(slf_op_16_21[7:0]),
     .lft_op_10(net4015[0:7]), .lft_op_09(net4016[0:7]),
     .lft_op_08(net4017[0:7]), .lft_op_07(net4018[0:7]),
     .lft_op_06(net4019[0:7]), .lft_op_05(net4020[0:7]),
     .sp12_h_l_10(net3539[0:23]), .sp12_h_r_10(net3050[0:23]),
     .sp12_h_l_09(net3548[0:23]), .sp12_h_l_08(net3547[0:23]),
     .sp12_h_l_07(net3546[0:23]), .sp12_h_l_06(net3545[0:23]),
     .sp12_h_r_05(net3055[0:23]), .sp12_h_r_06(net3056[0:23]),
     .sp12_h_r_07(net3057[0:23]), .sp12_h_r_08(net3058[0:23]),
     .sp12_h_r_09(net3059[0:23]), .sp12_h_l_05(net3544[0:23]),
     .sp4_r_v_b_05(net3061[0:47]), .sp4_r_v_b_06(net3062[0:47]),
     .sp4_r_v_b_07(net3063[0:47]), .sp4_r_v_b_08(net3064[0:47]),
     .sp4_r_v_b_09(net3065[0:47]), .sp4_r_v_b_10(net3066[0:47]),
     .sp4_v_b_10(net3555[0:47]), .sp4_v_b_09(net3554[0:47]),
     .sp4_v_b_08(net3553[0:47]), .sp4_v_b_07(net3552[0:47]),
     .sp4_v_b_06(net3551[0:47]), .sp4_v_b_05(net3550[0:47]),
     .sp4_v_t_16(net3073[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net3076[0:47]),
     .sp4_h_r_12(net3077[0:47]), .sp4_h_r_13(net3078[0:47]),
     .sp4_h_r_14(net3079[0:47]), .sp4_h_r_15(net3080[0:47]),
     .sp4_h_r_16(net3081[0:47]), .sp4_h_l_16(net3570[0:47]),
     .sp4_h_l_15(net3569[0:47]), .sp4_h_l_14(net3568[0:47]),
     .sp4_h_l_13(net3567[0:47]), .sp4_h_l_12(net3566[0:47]),
     .sp4_h_l_11(net3565[0:47]), .tnr_op_16({slf_op_16_33[3],
     slf_op_16_33[2], slf_op_16_33[1], slf_op_16_33[0],
     slf_op_16_33[3], slf_op_16_33[2], slf_op_16_33[1],
     slf_op_16_33[0]}), .tnl_op_16({slf_op_14_33[3], slf_op_14_33[2],
     slf_op_14_33[1], slf_op_14_33[0], slf_op_14_33[3],
     slf_op_14_33[2], slf_op_14_33[1], slf_op_14_33[0]}),
     .lft_op_16(net2188[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net3587[0:7]), .slf_op_14(net3586[0:7]),
     .slf_op_13(net3589[0:7]), .slf_op_12(net3588[0:7]),
     .slf_op_11(net3590[0:7]), .rgt_op_14(slf_op_16_30[7:0]),
     .rgt_op_15(slf_op_16_31[7:0]), .rgt_op_12(slf_op_16_28[7:0]),
     .rgt_op_13(slf_op_16_29[7:0]), .rgt_op_11(slf_op_16_27[7:0]),
     .sp4_v_b_16(net3597[0:47]), .sp4_v_b_14(net3600[0:47]),
     .sp4_v_b_15(net3598[0:47]), .sp4_v_b_13(net3599[0:47]),
     .sp4_v_b_11(net3602[0:47]), .sp4_v_b_12(net3601[0:47]),
     .sp4_r_v_b_16(net3108[0:47]), .sp4_r_v_b_15(net3109[0:47]),
     .sp4_r_v_b_13(net3110[0:47]), .sp4_r_v_b_14(net3111[0:47]),
     .sp4_r_v_b_12(net3112[0:47]), .sp4_r_v_b_11(net3113[0:47]),
     .sp12_h_l_16(net3609[0:23]), .sp12_h_l_15(net3611[0:23]),
     .sp12_h_l_14(net3610[0:23]), .sp12_h_l_13(net3613[0:23]),
     .sp12_h_l_12(net3612[0:23]), .sp12_h_l_11(net3614[0:23]),
     .sp12_h_r_16(net3120[0:23]), .sp12_h_r_14(net3121[0:23]),
     .sp12_h_r_15(net3122[0:23]), .sp12_h_r_12(net3123[0:23]),
     .sp12_h_r_13(net3124[0:23]), .sp12_h_r_11(net3125[0:23]),
     .lft_op_14(net4075[0:7]), .lft_op_15(net4076[0:7]),
     .lft_op_12(net4077[0:7]), .lft_op_11(net4079[0:7]),
     .lft_op_13(net4078[0:7]));
array_LT1x16top I_it_06_top ( .glb_netwk(net3158[0:7]),
     .sp12_v_t_16(net3131[0:23]), .rgt_op_16(net2163[0:7]),
     .top_op_16({slf_op_06_33[3], slf_op_06_33[2], slf_op_06_33[1],
     slf_op_06_33[0], slf_op_06_33[3], slf_op_06_33[2],
     slf_op_06_33[1], slf_op_06_33[0]}), .rgt_op_03(net3134[0:7]),
     .slf_op_02(net2484[0:7]), .rgt_op_02(net3136[0:7]),
     .rgt_op_01(slf_op_07_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4774[0:7]), .lft_op_03(net4764[0:7]),
     .lft_op_02(net4766[0:7]), .lft_op_01(slf_op_05_17[7:0]),
     .rgt_op_04(net3144[0:7]), .carry_in(carry_in_06_17),
     .bnl_op_01(bnl_op_06_17[7:0]), .slf_op_04(net2492[0:7]),
     .slf_op_03(net2482[0:7]), .slf_op_01(slf_op_06_17[7:0]),
     .sp4_h_l_04(net2513[0:47]), .carry_out(net3151),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_06_17[23:0]),
     .sp12_h_r_04(net3154[0:23]), .sp12_h_r_03(net3155[0:23]),
     .sp12_h_r_02(net3156[0:23]), .sp12_h_r_01(net3157[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2162[0:7]),
     .sp4_v_b_01(sp4_v_b_06_17[47:0]), .sp4_r_v_b_04(net3161[0:47]),
     .sp4_r_v_b_03(net3162[0:47]), .sp4_r_v_b_02(net3163[0:47]),
     .sp4_r_v_b_01(sp4_v_b_07_17[47:0]), .sp4_h_r_04(net3165[0:47]),
     .sp4_h_r_03(net3166[0:47]), .sp4_h_r_02(net3167[0:47]),
     .sp4_h_r_01(net3168[0:47]), .sp4_h_l_03(net2514[0:47]),
     .sp4_h_l_02(net2515[0:47]), .sp4_h_l_01(net2516[0:47]),
     .bl(bl[341:288]), .bot_op_01(bot_op_06_17[7:0]),
     .sp12_h_l_01(net2505[0:23]), .sp12_h_l_02(net2504[0:23]),
     .sp12_h_l_03(net2503[0:23]), .sp12_h_l_04(net2502[0:23]),
     .sp4_v_b_04(net2509[0:47]), .sp4_v_b_03(net2510[0:47]),
     .sp4_v_b_02(net2511[0:47]), .bnr_op_01(bnr_op_06_17[7:0]),
     .sp4_h_l_05(net2541[0:47]), .sp4_h_l_06(net2540[0:47]),
     .sp4_h_l_07(net2539[0:47]), .sp4_h_l_08(net2538[0:47]),
     .sp4_h_l_09(net2537[0:47]), .sp4_h_l_10(net2536[0:47]),
     .sp4_h_r_10(net3188[0:47]), .sp4_h_r_09(net3189[0:47]),
     .sp4_h_r_08(net3190[0:47]), .sp4_h_r_07(net3191[0:47]),
     .sp4_h_r_06(net3192[0:47]), .sp4_h_r_05(net3193[0:47]),
     .slf_op_05(net2553[0:7]), .slf_op_06(net2552[0:7]),
     .slf_op_07(net2551[0:7]), .slf_op_08(net2550[0:7]),
     .slf_op_09(net2549[0:7]), .slf_op_10(net2548[0:7]),
     .rgt_op_10(net3200[0:7]), .rgt_op_09(net3201[0:7]),
     .rgt_op_08(net3202[0:7]), .rgt_op_07(net3203[0:7]),
     .rgt_op_06(net3204[0:7]), .rgt_op_05(net3205[0:7]),
     .lft_op_10(net4830[0:7]), .lft_op_09(net4831[0:7]),
     .lft_op_08(net4832[0:7]), .lft_op_07(net4833[0:7]),
     .lft_op_06(net4834[0:7]), .lft_op_05(net4835[0:7]),
     .sp12_h_l_10(net2561[0:23]), .sp12_h_r_10(net3213[0:23]),
     .sp12_h_l_09(net2570[0:23]), .sp12_h_l_08(net2569[0:23]),
     .sp12_h_l_07(net2568[0:23]), .sp12_h_l_06(net2567[0:23]),
     .sp12_h_r_05(net3218[0:23]), .sp12_h_r_06(net3219[0:23]),
     .sp12_h_r_07(net3220[0:23]), .sp12_h_r_08(net3221[0:23]),
     .sp12_h_r_09(net3222[0:23]), .sp12_h_l_05(net2566[0:23]),
     .sp4_r_v_b_05(net3224[0:47]), .sp4_r_v_b_06(net3225[0:47]),
     .sp4_r_v_b_07(net3226[0:47]), .sp4_r_v_b_08(net3227[0:47]),
     .sp4_r_v_b_09(net3228[0:47]), .sp4_r_v_b_10(net3229[0:47]),
     .sp4_v_b_10(net2577[0:47]), .sp4_v_b_09(net2576[0:47]),
     .sp4_v_b_08(net2575[0:47]), .sp4_v_b_07(net2574[0:47]),
     .sp4_v_b_06(net2573[0:47]), .sp4_v_b_05(net2572[0:47]),
     .sp4_v_t_16(net3236[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net3239[0:47]),
     .sp4_h_r_12(net3240[0:47]), .sp4_h_r_13(net3241[0:47]),
     .sp4_h_r_14(net3242[0:47]), .sp4_h_r_15(net3243[0:47]),
     .sp4_h_r_16(net3244[0:47]), .sp4_h_l_16(net2592[0:47]),
     .sp4_h_l_15(net2591[0:47]), .sp4_h_l_14(net2590[0:47]),
     .sp4_h_l_13(net2589[0:47]), .sp4_h_l_12(net2588[0:47]),
     .sp4_h_l_11(net2587[0:47]), .tnr_op_16({slf_op_07_33[3],
     slf_op_07_33[2], slf_op_07_33[1], slf_op_07_33[0],
     slf_op_07_33[3], slf_op_07_33[2], slf_op_07_33[1],
     slf_op_07_33[0]}), .tnl_op_16({slf_op_05_33[3], slf_op_05_33[2],
     slf_op_05_33[1], slf_op_05_33[0], slf_op_05_33[3],
     slf_op_05_33[2], slf_op_05_33[1], slf_op_05_33[0]}),
     .lft_op_16(net2179[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net2609[0:7]), .slf_op_14(net2608[0:7]),
     .slf_op_13(net2611[0:7]), .slf_op_12(net2610[0:7]),
     .slf_op_11(net2612[0:7]), .rgt_op_14(net3260[0:7]),
     .rgt_op_15(net3261[0:7]), .rgt_op_12(net3262[0:7]),
     .rgt_op_13(net3263[0:7]), .rgt_op_11(net3264[0:7]),
     .sp4_v_b_16(net2619[0:47]), .sp4_v_b_14(net2622[0:47]),
     .sp4_v_b_15(net2620[0:47]), .sp4_v_b_13(net2621[0:47]),
     .sp4_v_b_11(net2624[0:47]), .sp4_v_b_12(net2623[0:47]),
     .sp4_r_v_b_16(net3271[0:47]), .sp4_r_v_b_15(net3272[0:47]),
     .sp4_r_v_b_13(net3273[0:47]), .sp4_r_v_b_14(net3274[0:47]),
     .sp4_r_v_b_12(net3275[0:47]), .sp4_r_v_b_11(net3276[0:47]),
     .sp12_h_l_16(net2631[0:23]), .sp12_h_l_15(net2633[0:23]),
     .sp12_h_l_14(net2632[0:23]), .sp12_h_l_13(net2635[0:23]),
     .sp12_h_l_12(net2634[0:23]), .sp12_h_l_11(net2636[0:23]),
     .sp12_h_r_16(net3283[0:23]), .sp12_h_r_14(net3284[0:23]),
     .sp12_h_r_15(net3285[0:23]), .sp12_h_r_12(net3286[0:23]),
     .sp12_h_r_13(net3287[0:23]), .sp12_h_r_11(net3288[0:23]),
     .lft_op_14(net4890[0:7]), .lft_op_15(net4891[0:7]),
     .lft_op_12(net4892[0:7]), .lft_op_11(net4894[0:7]),
     .lft_op_13(net4893[0:7]));
array_LT1x16top I_it_03_top ( .glb_netwk(net3321[0:7]),
     .sp12_v_t_16(net3294[0:23]), .rgt_op_16(net2160[0:7]),
     .top_op_16({slf_op_03_33[3], slf_op_03_33[2], slf_op_03_33[1],
     slf_op_03_33[0], slf_op_03_33[3], slf_op_03_33[2],
     slf_op_03_33[1], slf_op_03_33[0]}), .rgt_op_03(net3297[0:7]),
     .slf_op_02(net4277[0:7]), .rgt_op_02(net3299[0:7]),
     .rgt_op_01(slf_op_04_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4448[0:7]), .lft_op_03(net4438[0:7]),
     .lft_op_02(net4440[0:7]), .lft_op_01(slf_op_02_17[7:0]),
     .rgt_op_04(net3307[0:7]), .carry_in(carry_in_03_17),
     .bnl_op_01(bnl_op_03_17[7:0]), .slf_op_04(net4285[0:7]),
     .slf_op_03(net4275[0:7]), .slf_op_01(slf_op_03_17[7:0]),
     .sp4_h_l_04(net4306[0:47]), .carry_out(net3314),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_03_17[23:0]),
     .sp12_h_r_04(net3317[0:23]), .sp12_h_r_03(net3318[0:23]),
     .sp12_h_r_02(net3319[0:23]), .sp12_h_r_01(net3320[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2177[0:7]),
     .sp4_v_b_01(sp4_v_b_03_17[47:0]), .sp4_r_v_b_04(net3324[0:47]),
     .sp4_r_v_b_03(net3325[0:47]), .sp4_r_v_b_02(net3326[0:47]),
     .sp4_r_v_b_01(sp4_v_b_04_17[47:0]), .sp4_h_r_04(net3328[0:47]),
     .sp4_h_r_03(net3329[0:47]), .sp4_h_r_02(net3330[0:47]),
     .sp4_h_r_01(net3331[0:47]), .sp4_h_l_03(net4307[0:47]),
     .sp4_h_l_02(net4308[0:47]), .sp4_h_l_01(net4309[0:47]),
     .bl(bl[179:126]), .bot_op_01(bot_op_03_17[7:0]),
     .sp12_h_l_01(net4298[0:23]), .sp12_h_l_02(net4297[0:23]),
     .sp12_h_l_03(net4296[0:23]), .sp12_h_l_04(net4295[0:23]),
     .sp4_v_b_04(net4302[0:47]), .sp4_v_b_03(net4303[0:47]),
     .sp4_v_b_02(net4304[0:47]), .bnr_op_01(bnr_op_03_17[7:0]),
     .sp4_h_l_05(net4334[0:47]), .sp4_h_l_06(net4333[0:47]),
     .sp4_h_l_07(net4332[0:47]), .sp4_h_l_08(net4331[0:47]),
     .sp4_h_l_09(net4330[0:47]), .sp4_h_l_10(net4329[0:47]),
     .sp4_h_r_10(net3351[0:47]), .sp4_h_r_09(net3352[0:47]),
     .sp4_h_r_08(net3353[0:47]), .sp4_h_r_07(net3354[0:47]),
     .sp4_h_r_06(net3355[0:47]), .sp4_h_r_05(net3356[0:47]),
     .slf_op_05(net4346[0:7]), .slf_op_06(net4345[0:7]),
     .slf_op_07(net4344[0:7]), .slf_op_08(net4343[0:7]),
     .slf_op_09(net4342[0:7]), .slf_op_10(net4341[0:7]),
     .rgt_op_10(net3363[0:7]), .rgt_op_09(net3364[0:7]),
     .rgt_op_08(net3365[0:7]), .rgt_op_07(net3366[0:7]),
     .rgt_op_06(net3367[0:7]), .rgt_op_05(net3368[0:7]),
     .lft_op_10(net4504[0:7]), .lft_op_09(net4505[0:7]),
     .lft_op_08(net4506[0:7]), .lft_op_07(net4507[0:7]),
     .lft_op_06(net4508[0:7]), .lft_op_05(net4509[0:7]),
     .sp12_h_l_10(net4354[0:23]), .sp12_h_r_10(net3376[0:23]),
     .sp12_h_l_09(net4363[0:23]), .sp12_h_l_08(net4362[0:23]),
     .sp12_h_l_07(net4361[0:23]), .sp12_h_l_06(net4360[0:23]),
     .sp12_h_r_05(net3381[0:23]), .sp12_h_r_06(net3382[0:23]),
     .sp12_h_r_07(net3383[0:23]), .sp12_h_r_08(net3384[0:23]),
     .sp12_h_r_09(net3385[0:23]), .sp12_h_l_05(net4359[0:23]),
     .sp4_r_v_b_05(net3387[0:47]), .sp4_r_v_b_06(net3388[0:47]),
     .sp4_r_v_b_07(net3389[0:47]), .sp4_r_v_b_08(net3390[0:47]),
     .sp4_r_v_b_09(net3391[0:47]), .sp4_r_v_b_10(net3392[0:47]),
     .sp4_v_b_10(net4370[0:47]), .sp4_v_b_09(net4369[0:47]),
     .sp4_v_b_08(net4368[0:47]), .sp4_v_b_07(net4367[0:47]),
     .sp4_v_b_06(net4366[0:47]), .sp4_v_b_05(net4365[0:47]),
     .sp4_v_t_16(net3399[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net3402[0:47]),
     .sp4_h_r_12(net3403[0:47]), .sp4_h_r_13(net3404[0:47]),
     .sp4_h_r_14(net3405[0:47]), .sp4_h_r_15(net3406[0:47]),
     .sp4_h_r_16(net3407[0:47]), .sp4_h_l_16(net4385[0:47]),
     .sp4_h_l_15(net4384[0:47]), .sp4_h_l_14(net4383[0:47]),
     .sp4_h_l_13(net4382[0:47]), .sp4_h_l_12(net4381[0:47]),
     .sp4_h_l_11(net4380[0:47]), .tnr_op_16({slf_op_04_33[3],
     slf_op_04_33[2], slf_op_04_33[1], slf_op_04_33[0],
     slf_op_04_33[3], slf_op_04_33[2], slf_op_04_33[1],
     slf_op_04_33[0]}), .tnl_op_16({slf_op_02_33[3], slf_op_02_33[2],
     slf_op_02_33[1], slf_op_02_33[0], slf_op_02_33[3],
     slf_op_02_33[2], slf_op_02_33[1], slf_op_02_33[0]}),
     .lft_op_16(net4436[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net4402[0:7]), .slf_op_14(net4401[0:7]),
     .slf_op_13(net4404[0:7]), .slf_op_12(net4403[0:7]),
     .slf_op_11(net4405[0:7]), .rgt_op_14(net3423[0:7]),
     .rgt_op_15(net3424[0:7]), .rgt_op_12(net3425[0:7]),
     .rgt_op_13(net3426[0:7]), .rgt_op_11(net3427[0:7]),
     .sp4_v_b_16(net4412[0:47]), .sp4_v_b_14(net4415[0:47]),
     .sp4_v_b_15(net4413[0:47]), .sp4_v_b_13(net4414[0:47]),
     .sp4_v_b_11(net4417[0:47]), .sp4_v_b_12(net4416[0:47]),
     .sp4_r_v_b_16(net3434[0:47]), .sp4_r_v_b_15(net3435[0:47]),
     .sp4_r_v_b_13(net3436[0:47]), .sp4_r_v_b_14(net3437[0:47]),
     .sp4_r_v_b_12(net3438[0:47]), .sp4_r_v_b_11(net3439[0:47]),
     .sp12_h_l_16(net4424[0:23]), .sp12_h_l_15(net4426[0:23]),
     .sp12_h_l_14(net4425[0:23]), .sp12_h_l_13(net4428[0:23]),
     .sp12_h_l_12(net4427[0:23]), .sp12_h_l_11(net4429[0:23]),
     .sp12_h_r_16(net3446[0:23]), .sp12_h_r_14(net3447[0:23]),
     .sp12_h_r_15(net3448[0:23]), .sp12_h_r_12(net3449[0:23]),
     .sp12_h_r_13(net3450[0:23]), .sp12_h_r_11(net3451[0:23]),
     .lft_op_14(net4564[0:7]), .lft_op_15(net4565[0:7]),
     .lft_op_12(net4566[0:7]), .lft_op_11(net4568[0:7]),
     .lft_op_13(net4567[0:7]));
array_LT1x16top I_it_14_top ( .glb_netwk(net3484[0:7]),
     .sp12_v_t_16(net3457[0:23]), .rgt_op_16(net3458[0:7]),
     .top_op_16({slf_op_14_33[3], slf_op_14_33[2], slf_op_14_33[1],
     slf_op_14_33[0], slf_op_14_33[3], slf_op_14_33[2],
     slf_op_14_33[1], slf_op_14_33[0]}), .rgt_op_03(net3460[0:7]),
     .slf_op_02(net3951[0:7]), .rgt_op_02(net3462[0:7]),
     .rgt_op_01(slf_op_15_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3633[0:7]), .lft_op_03(net3623[0:7]),
     .lft_op_02(net3625[0:7]), .lft_op_01(slf_op_13_17[7:0]),
     .rgt_op_04(net3470[0:7]), .carry_in(carry_in_14_17),
     .bnl_op_01(bnl_op_14_17[7:0]), .slf_op_04(net3959[0:7]),
     .slf_op_03(net3949[0:7]), .slf_op_01(slf_op_14_17[7:0]),
     .sp4_h_l_04(net3980[0:47]), .carry_out(net3477),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_14_17[23:0]),
     .sp12_h_r_04(net3480[0:23]), .sp12_h_r_03(net3481[0:23]),
     .sp12_h_r_02(net3482[0:23]), .sp12_h_r_01(net3483[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2188[0:7]),
     .sp4_v_b_01(sp4_v_b_14_17[47:0]), .sp4_r_v_b_04(net3487[0:47]),
     .sp4_r_v_b_03(net3488[0:47]), .sp4_r_v_b_02(net3489[0:47]),
     .sp4_r_v_b_01(sp4_v_b_15_17[47:0]), .sp4_h_r_04(net3491[0:47]),
     .sp4_h_r_03(net3492[0:47]), .sp4_h_r_02(net3493[0:47]),
     .sp4_h_r_01(net3494[0:47]), .sp4_h_l_03(net3981[0:47]),
     .sp4_h_l_02(net3982[0:47]), .sp4_h_l_01(net3983[0:47]),
     .bl(bl[761:708]), .bot_op_01(bot_op_14_17[7:0]),
     .sp12_h_l_01(net3972[0:23]), .sp12_h_l_02(net3971[0:23]),
     .sp12_h_l_03(net3970[0:23]), .sp12_h_l_04(net3969[0:23]),
     .sp4_v_b_04(net3976[0:47]), .sp4_v_b_03(net3977[0:47]),
     .sp4_v_b_02(net3978[0:47]), .bnr_op_01(bnr_op_14_17[7:0]),
     .sp4_h_l_05(net4008[0:47]), .sp4_h_l_06(net4007[0:47]),
     .sp4_h_l_07(net4006[0:47]), .sp4_h_l_08(net4005[0:47]),
     .sp4_h_l_09(net4004[0:47]), .sp4_h_l_10(net4003[0:47]),
     .sp4_h_r_10(net3514[0:47]), .sp4_h_r_09(net3515[0:47]),
     .sp4_h_r_08(net3516[0:47]), .sp4_h_r_07(net3517[0:47]),
     .sp4_h_r_06(net3518[0:47]), .sp4_h_r_05(net3519[0:47]),
     .slf_op_05(net4020[0:7]), .slf_op_06(net4019[0:7]),
     .slf_op_07(net4018[0:7]), .slf_op_08(net4017[0:7]),
     .slf_op_09(net4016[0:7]), .slf_op_10(net4015[0:7]),
     .rgt_op_10(net3526[0:7]), .rgt_op_09(net3527[0:7]),
     .rgt_op_08(net3528[0:7]), .rgt_op_07(net3529[0:7]),
     .rgt_op_06(net3530[0:7]), .rgt_op_05(net3531[0:7]),
     .lft_op_10(net3689[0:7]), .lft_op_09(net3690[0:7]),
     .lft_op_08(net3691[0:7]), .lft_op_07(net3692[0:7]),
     .lft_op_06(net3693[0:7]), .lft_op_05(net3694[0:7]),
     .sp12_h_l_10(net4028[0:23]), .sp12_h_r_10(net3539[0:23]),
     .sp12_h_l_09(net4037[0:23]), .sp12_h_l_08(net4036[0:23]),
     .sp12_h_l_07(net4035[0:23]), .sp12_h_l_06(net4034[0:23]),
     .sp12_h_r_05(net3544[0:23]), .sp12_h_r_06(net3545[0:23]),
     .sp12_h_r_07(net3546[0:23]), .sp12_h_r_08(net3547[0:23]),
     .sp12_h_r_09(net3548[0:23]), .sp12_h_l_05(net4033[0:23]),
     .sp4_r_v_b_05(net3550[0:47]), .sp4_r_v_b_06(net3551[0:47]),
     .sp4_r_v_b_07(net3552[0:47]), .sp4_r_v_b_08(net3553[0:47]),
     .sp4_r_v_b_09(net3554[0:47]), .sp4_r_v_b_10(net3555[0:47]),
     .sp4_v_b_10(net4044[0:47]), .sp4_v_b_09(net4043[0:47]),
     .sp4_v_b_08(net4042[0:47]), .sp4_v_b_07(net4041[0:47]),
     .sp4_v_b_06(net4040[0:47]), .sp4_v_b_05(net4039[0:47]),
     .sp4_v_t_16(net3562[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net3565[0:47]),
     .sp4_h_r_12(net3566[0:47]), .sp4_h_r_13(net3567[0:47]),
     .sp4_h_r_14(net3568[0:47]), .sp4_h_r_15(net3569[0:47]),
     .sp4_h_r_16(net3570[0:47]), .sp4_h_l_16(net4059[0:47]),
     .sp4_h_l_15(net4058[0:47]), .sp4_h_l_14(net4057[0:47]),
     .sp4_h_l_13(net4056[0:47]), .sp4_h_l_12(net4055[0:47]),
     .sp4_h_l_11(net4054[0:47]), .tnr_op_16({slf_op_15_33[3],
     slf_op_15_33[2], slf_op_15_33[1], slf_op_15_33[0],
     slf_op_15_33[3], slf_op_15_33[2], slf_op_15_33[1],
     slf_op_15_33[0]}), .tnl_op_16({slf_op_13_33[3], slf_op_13_33[2],
     slf_op_13_33[1], slf_op_13_33[0], slf_op_13_33[3],
     slf_op_13_33[2], slf_op_13_33[1], slf_op_13_33[0]}),
     .lft_op_16(net2169[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net4076[0:7]), .slf_op_14(net4075[0:7]),
     .slf_op_13(net4078[0:7]), .slf_op_12(net4077[0:7]),
     .slf_op_11(net4079[0:7]), .rgt_op_14(net3586[0:7]),
     .rgt_op_15(net3587[0:7]), .rgt_op_12(net3588[0:7]),
     .rgt_op_13(net3589[0:7]), .rgt_op_11(net3590[0:7]),
     .sp4_v_b_16(net4086[0:47]), .sp4_v_b_14(net4089[0:47]),
     .sp4_v_b_15(net4087[0:47]), .sp4_v_b_13(net4088[0:47]),
     .sp4_v_b_11(net4091[0:47]), .sp4_v_b_12(net4090[0:47]),
     .sp4_r_v_b_16(net3597[0:47]), .sp4_r_v_b_15(net3598[0:47]),
     .sp4_r_v_b_13(net3599[0:47]), .sp4_r_v_b_14(net3600[0:47]),
     .sp4_r_v_b_12(net3601[0:47]), .sp4_r_v_b_11(net3602[0:47]),
     .sp12_h_l_16(net4098[0:23]), .sp12_h_l_15(net4100[0:23]),
     .sp12_h_l_14(net4099[0:23]), .sp12_h_l_13(net4102[0:23]),
     .sp12_h_l_12(net4101[0:23]), .sp12_h_l_11(net4103[0:23]),
     .sp12_h_r_16(net3609[0:23]), .sp12_h_r_14(net3610[0:23]),
     .sp12_h_r_15(net3611[0:23]), .sp12_h_r_12(net3612[0:23]),
     .sp12_h_r_13(net3613[0:23]), .sp12_h_r_11(net3614[0:23]),
     .lft_op_14(net3749[0:7]), .lft_op_15(net3750[0:7]),
     .lft_op_12(net3751[0:7]), .lft_op_11(net3753[0:7]),
     .lft_op_13(net3752[0:7]));
array_LT1x16top I_it_12_top ( .glb_netwk(net3647[0:7]),
     .sp12_v_t_16(net3620[0:23]), .rgt_op_16(net2169[0:7]),
     .top_op_16({slf_op_12_33[3], slf_op_12_33[2], slf_op_12_33[1],
     slf_op_12_33[0], slf_op_12_33[3], slf_op_12_33[2],
     slf_op_12_33[1], slf_op_12_33[0]}), .rgt_op_03(net3623[0:7]),
     .slf_op_02(net2647[0:7]), .rgt_op_02(net3625[0:7]),
     .rgt_op_01(slf_op_13_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2818[0:7]), .lft_op_03(net2808[0:7]),
     .lft_op_02(net2810[0:7]), .lft_op_01(slf_op_11_17[7:0]),
     .rgt_op_04(net3633[0:7]), .carry_in(carry_in_12_17),
     .bnl_op_01(bnl_op_12_17[7:0]), .slf_op_04(net2655[0:7]),
     .slf_op_03(net2645[0:7]), .slf_op_01(slf_op_12_17[7:0]),
     .sp4_h_l_04(net2676[0:47]), .carry_out(net3640),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_12_17[23:0]),
     .sp12_h_r_04(net3643[0:23]), .sp12_h_r_03(net3644[0:23]),
     .sp12_h_r_02(net3645[0:23]), .sp12_h_r_01(net3646[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2643[0:7]),
     .sp4_v_b_01(sp4_v_b_12_17[47:0]), .sp4_r_v_b_04(net3650[0:47]),
     .sp4_r_v_b_03(net3651[0:47]), .sp4_r_v_b_02(net3652[0:47]),
     .sp4_r_v_b_01(sp4_v_b_13_17[47:0]), .sp4_h_r_04(net3654[0:47]),
     .sp4_h_r_03(net3655[0:47]), .sp4_h_r_02(net3656[0:47]),
     .sp4_h_r_01(net3657[0:47]), .sp4_h_l_03(net2677[0:47]),
     .sp4_h_l_02(net2678[0:47]), .sp4_h_l_01(net2679[0:47]),
     .bl(bl[653:600]), .bot_op_01(bot_op_12_17[7:0]),
     .sp12_h_l_01(net2668[0:23]), .sp12_h_l_02(net2667[0:23]),
     .sp12_h_l_03(net2666[0:23]), .sp12_h_l_04(net2665[0:23]),
     .sp4_v_b_04(net2672[0:47]), .sp4_v_b_03(net2673[0:47]),
     .sp4_v_b_02(net2674[0:47]), .bnr_op_01(bnr_op_12_17[7:0]),
     .sp4_h_l_05(net2704[0:47]), .sp4_h_l_06(net2703[0:47]),
     .sp4_h_l_07(net2702[0:47]), .sp4_h_l_08(net2701[0:47]),
     .sp4_h_l_09(net2700[0:47]), .sp4_h_l_10(net2699[0:47]),
     .sp4_h_r_10(net3677[0:47]), .sp4_h_r_09(net3678[0:47]),
     .sp4_h_r_08(net3679[0:47]), .sp4_h_r_07(net3680[0:47]),
     .sp4_h_r_06(net3681[0:47]), .sp4_h_r_05(net3682[0:47]),
     .slf_op_05(net2716[0:7]), .slf_op_06(net2715[0:7]),
     .slf_op_07(net2714[0:7]), .slf_op_08(net2713[0:7]),
     .slf_op_09(net2712[0:7]), .slf_op_10(net2711[0:7]),
     .rgt_op_10(net3689[0:7]), .rgt_op_09(net3690[0:7]),
     .rgt_op_08(net3691[0:7]), .rgt_op_07(net3692[0:7]),
     .rgt_op_06(net3693[0:7]), .rgt_op_05(net3694[0:7]),
     .lft_op_10(net2874[0:7]), .lft_op_09(net2875[0:7]),
     .lft_op_08(net2876[0:7]), .lft_op_07(net2877[0:7]),
     .lft_op_06(net2878[0:7]), .lft_op_05(net2879[0:7]),
     .sp12_h_l_10(net2724[0:23]), .sp12_h_r_10(net3702[0:23]),
     .sp12_h_l_09(net2733[0:23]), .sp12_h_l_08(net2732[0:23]),
     .sp12_h_l_07(net2731[0:23]), .sp12_h_l_06(net2730[0:23]),
     .sp12_h_r_05(net3707[0:23]), .sp12_h_r_06(net3708[0:23]),
     .sp12_h_r_07(net3709[0:23]), .sp12_h_r_08(net3710[0:23]),
     .sp12_h_r_09(net3711[0:23]), .sp12_h_l_05(net2729[0:23]),
     .sp4_r_v_b_05(net3713[0:47]), .sp4_r_v_b_06(net3714[0:47]),
     .sp4_r_v_b_07(net3715[0:47]), .sp4_r_v_b_08(net3716[0:47]),
     .sp4_r_v_b_09(net3717[0:47]), .sp4_r_v_b_10(net3718[0:47]),
     .sp4_v_b_10(net2740[0:47]), .sp4_v_b_09(net2739[0:47]),
     .sp4_v_b_08(net2738[0:47]), .sp4_v_b_07(net2737[0:47]),
     .sp4_v_b_06(net2736[0:47]), .sp4_v_b_05(net2735[0:47]),
     .sp4_v_t_16(net3725[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net3728[0:47]),
     .sp4_h_r_12(net3729[0:47]), .sp4_h_r_13(net3730[0:47]),
     .sp4_h_r_14(net3731[0:47]), .sp4_h_r_15(net3732[0:47]),
     .sp4_h_r_16(net3733[0:47]), .sp4_h_l_16(net2755[0:47]),
     .sp4_h_l_15(net2754[0:47]), .sp4_h_l_14(net2753[0:47]),
     .sp4_h_l_13(net2752[0:47]), .sp4_h_l_12(net2751[0:47]),
     .sp4_h_l_11(net2750[0:47]), .tnr_op_16({slf_op_13_33[3],
     slf_op_13_33[2], slf_op_13_33[1], slf_op_13_33[0],
     slf_op_13_33[3], slf_op_13_33[2], slf_op_13_33[1],
     slf_op_13_33[0]}), .tnl_op_16({slf_op_11_33[3], slf_op_11_33[2],
     slf_op_11_33[1], slf_op_11_33[0], slf_op_11_33[3],
     slf_op_11_33[2], slf_op_11_33[1], slf_op_11_33[0]}),
     .lft_op_16(net2167[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net2772[0:7]), .slf_op_14(net2771[0:7]),
     .slf_op_13(net2774[0:7]), .slf_op_12(net2773[0:7]),
     .slf_op_11(net2775[0:7]), .rgt_op_14(net3749[0:7]),
     .rgt_op_15(net3750[0:7]), .rgt_op_12(net3751[0:7]),
     .rgt_op_13(net3752[0:7]), .rgt_op_11(net3753[0:7]),
     .sp4_v_b_16(net2782[0:47]), .sp4_v_b_14(net2785[0:47]),
     .sp4_v_b_15(net2783[0:47]), .sp4_v_b_13(net2784[0:47]),
     .sp4_v_b_11(net2787[0:47]), .sp4_v_b_12(net2786[0:47]),
     .sp4_r_v_b_16(net3760[0:47]), .sp4_r_v_b_15(net3761[0:47]),
     .sp4_r_v_b_13(net3762[0:47]), .sp4_r_v_b_14(net3763[0:47]),
     .sp4_r_v_b_12(net3764[0:47]), .sp4_r_v_b_11(net3765[0:47]),
     .sp12_h_l_16(net2794[0:23]), .sp12_h_l_15(net2796[0:23]),
     .sp12_h_l_14(net2795[0:23]), .sp12_h_l_13(net2798[0:23]),
     .sp12_h_l_12(net2797[0:23]), .sp12_h_l_11(net2799[0:23]),
     .sp12_h_r_16(net3772[0:23]), .sp12_h_r_14(net3773[0:23]),
     .sp12_h_r_15(net3774[0:23]), .sp12_h_r_12(net3775[0:23]),
     .sp12_h_r_13(net3776[0:23]), .sp12_h_r_11(net3777[0:23]),
     .lft_op_14(net2934[0:7]), .lft_op_15(net2935[0:7]),
     .lft_op_12(net2936[0:7]), .lft_op_11(net2938[0:7]),
     .lft_op_13(net2937[0:7]));
array_LT1x16top I_it_07_top ( .glb_netwk(net3810[0:7]),
     .sp12_v_t_16(net3783[0:23]), .rgt_op_16(net2164[0:7]),
     .top_op_16({slf_op_07_33[3], slf_op_07_33[2], slf_op_07_33[1],
     slf_op_07_33[0], slf_op_07_33[3], slf_op_07_33[2],
     slf_op_07_33[1], slf_op_07_33[0]}), .rgt_op_03(net3786[0:7]),
     .slf_op_02(net3136[0:7]), .rgt_op_02(net3788[0:7]),
     .rgt_op_01(slf_op_08_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2492[0:7]), .lft_op_03(net2482[0:7]),
     .lft_op_02(net2484[0:7]), .lft_op_01(slf_op_06_17[7:0]),
     .rgt_op_04(net3796[0:7]), .carry_in(carry_in_07_17),
     .bnl_op_01(bnl_op_07_17[7:0]), .slf_op_04(net3144[0:7]),
     .slf_op_03(net3134[0:7]), .slf_op_01(slf_op_07_17[7:0]),
     .sp4_h_l_04(net3165[0:47]), .carry_out(net3803),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_07_17[23:0]),
     .sp12_h_r_04(net3806[0:23]), .sp12_h_r_03(net3807[0:23]),
     .sp12_h_r_02(net3808[0:23]), .sp12_h_r_01(net3809[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2163[0:7]),
     .sp4_v_b_01(sp4_v_b_07_17[47:0]), .sp4_r_v_b_04(net3813[0:47]),
     .sp4_r_v_b_03(net3814[0:47]), .sp4_r_v_b_02(net3815[0:47]),
     .sp4_r_v_b_01(sp4_v_b_08_17[47:0]), .sp4_h_r_04(net3817[0:47]),
     .sp4_h_r_03(net3818[0:47]), .sp4_h_r_02(net3819[0:47]),
     .sp4_h_r_01(net3820[0:47]), .sp4_h_l_03(net3166[0:47]),
     .sp4_h_l_02(net3167[0:47]), .sp4_h_l_01(net3168[0:47]),
     .bl(bl[395:342]), .bot_op_01(bot_op_07_17[7:0]),
     .sp12_h_l_01(net3157[0:23]), .sp12_h_l_02(net3156[0:23]),
     .sp12_h_l_03(net3155[0:23]), .sp12_h_l_04(net3154[0:23]),
     .sp4_v_b_04(net3161[0:47]), .sp4_v_b_03(net3162[0:47]),
     .sp4_v_b_02(net3163[0:47]), .bnr_op_01(bnr_op_07_17[7:0]),
     .sp4_h_l_05(net3193[0:47]), .sp4_h_l_06(net3192[0:47]),
     .sp4_h_l_07(net3191[0:47]), .sp4_h_l_08(net3190[0:47]),
     .sp4_h_l_09(net3189[0:47]), .sp4_h_l_10(net3188[0:47]),
     .sp4_h_r_10(net3840[0:47]), .sp4_h_r_09(net3841[0:47]),
     .sp4_h_r_08(net3842[0:47]), .sp4_h_r_07(net3843[0:47]),
     .sp4_h_r_06(net3844[0:47]), .sp4_h_r_05(net3845[0:47]),
     .slf_op_05(net3205[0:7]), .slf_op_06(net3204[0:7]),
     .slf_op_07(net3203[0:7]), .slf_op_08(net3202[0:7]),
     .slf_op_09(net3201[0:7]), .slf_op_10(net3200[0:7]),
     .rgt_op_10(net3852[0:7]), .rgt_op_09(net3853[0:7]),
     .rgt_op_08(net3854[0:7]), .rgt_op_07(net3855[0:7]),
     .rgt_op_06(net3856[0:7]), .rgt_op_05(net3857[0:7]),
     .lft_op_10(net2548[0:7]), .lft_op_09(net2549[0:7]),
     .lft_op_08(net2550[0:7]), .lft_op_07(net2551[0:7]),
     .lft_op_06(net2552[0:7]), .lft_op_05(net2553[0:7]),
     .sp12_h_l_10(net3213[0:23]), .sp12_h_r_10(net3865[0:23]),
     .sp12_h_l_09(net3222[0:23]), .sp12_h_l_08(net3221[0:23]),
     .sp12_h_l_07(net3220[0:23]), .sp12_h_l_06(net3219[0:23]),
     .sp12_h_r_05(net3870[0:23]), .sp12_h_r_06(net3871[0:23]),
     .sp12_h_r_07(net3872[0:23]), .sp12_h_r_08(net3873[0:23]),
     .sp12_h_r_09(net3874[0:23]), .sp12_h_l_05(net3218[0:23]),
     .sp4_r_v_b_05(net3876[0:47]), .sp4_r_v_b_06(net3877[0:47]),
     .sp4_r_v_b_07(net3878[0:47]), .sp4_r_v_b_08(net3879[0:47]),
     .sp4_r_v_b_09(net3880[0:47]), .sp4_r_v_b_10(net3881[0:47]),
     .sp4_v_b_10(net3229[0:47]), .sp4_v_b_09(net3228[0:47]),
     .sp4_v_b_08(net3227[0:47]), .sp4_v_b_07(net3226[0:47]),
     .sp4_v_b_06(net3225[0:47]), .sp4_v_b_05(net3224[0:47]),
     .sp4_v_t_16(net3888[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net3891[0:47]),
     .sp4_h_r_12(net3892[0:47]), .sp4_h_r_13(net3893[0:47]),
     .sp4_h_r_14(net3894[0:47]), .sp4_h_r_15(net3895[0:47]),
     .sp4_h_r_16(net3896[0:47]), .sp4_h_l_16(net3244[0:47]),
     .sp4_h_l_15(net3243[0:47]), .sp4_h_l_14(net3242[0:47]),
     .sp4_h_l_13(net3241[0:47]), .sp4_h_l_12(net3240[0:47]),
     .sp4_h_l_11(net3239[0:47]), .tnr_op_16({slf_op_08_33[3],
     slf_op_08_33[2], slf_op_08_33[1], slf_op_08_33[0],
     slf_op_08_33[3], slf_op_08_33[2], slf_op_08_33[1],
     slf_op_08_33[0]}), .tnl_op_16({slf_op_06_33[3], slf_op_06_33[2],
     slf_op_06_33[1], slf_op_06_33[0], slf_op_06_33[3],
     slf_op_06_33[2], slf_op_06_33[1], slf_op_06_33[0]}),
     .lft_op_16(net2162[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net3261[0:7]), .slf_op_14(net3260[0:7]),
     .slf_op_13(net3263[0:7]), .slf_op_12(net3262[0:7]),
     .slf_op_11(net3264[0:7]), .rgt_op_14(net3912[0:7]),
     .rgt_op_15(net3913[0:7]), .rgt_op_12(net3914[0:7]),
     .rgt_op_13(net3915[0:7]), .rgt_op_11(net3916[0:7]),
     .sp4_v_b_16(net3271[0:47]), .sp4_v_b_14(net3274[0:47]),
     .sp4_v_b_15(net3272[0:47]), .sp4_v_b_13(net3273[0:47]),
     .sp4_v_b_11(net3276[0:47]), .sp4_v_b_12(net3275[0:47]),
     .sp4_r_v_b_16(net3923[0:47]), .sp4_r_v_b_15(net3924[0:47]),
     .sp4_r_v_b_13(net3925[0:47]), .sp4_r_v_b_14(net3926[0:47]),
     .sp4_r_v_b_12(net3927[0:47]), .sp4_r_v_b_11(net3928[0:47]),
     .sp12_h_l_16(net3283[0:23]), .sp12_h_l_15(net3285[0:23]),
     .sp12_h_l_14(net3284[0:23]), .sp12_h_l_13(net3287[0:23]),
     .sp12_h_l_12(net3286[0:23]), .sp12_h_l_11(net3288[0:23]),
     .sp12_h_r_16(net3935[0:23]), .sp12_h_r_14(net3936[0:23]),
     .sp12_h_r_15(net3937[0:23]), .sp12_h_r_12(net3938[0:23]),
     .sp12_h_r_13(net3939[0:23]), .sp12_h_r_11(net3940[0:23]),
     .lft_op_14(net2608[0:7]), .lft_op_15(net2609[0:7]),
     .lft_op_12(net2610[0:7]), .lft_op_11(net2612[0:7]),
     .lft_op_13(net2611[0:7]));
array_LT1x16top I_it_13_top ( .glb_netwk(net3973[0:7]),
     .sp12_v_t_16(net3946[0:23]), .rgt_op_16(net2188[0:7]),
     .top_op_16({slf_op_13_33[3], slf_op_13_33[2], slf_op_13_33[1],
     slf_op_13_33[0], slf_op_13_33[3], slf_op_13_33[2],
     slf_op_13_33[1], slf_op_13_33[0]}), .rgt_op_03(net3949[0:7]),
     .slf_op_02(net3625[0:7]), .rgt_op_02(net3951[0:7]),
     .rgt_op_01(slf_op_14_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2655[0:7]), .lft_op_03(net2645[0:7]),
     .lft_op_02(net2647[0:7]), .lft_op_01(slf_op_12_17[7:0]),
     .rgt_op_04(net3959[0:7]), .carry_in(carry_in_13_17),
     .bnl_op_01(bnl_op_13_17[7:0]), .slf_op_04(net3633[0:7]),
     .slf_op_03(net3623[0:7]), .slf_op_01(slf_op_13_17[7:0]),
     .sp4_h_l_04(net3654[0:47]), .carry_out(net3966),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_13_17[23:0]),
     .sp12_h_r_04(net3969[0:23]), .sp12_h_r_03(net3970[0:23]),
     .sp12_h_r_02(net3971[0:23]), .sp12_h_r_01(net3972[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2169[0:7]),
     .sp4_v_b_01(sp4_v_b_13_17[47:0]), .sp4_r_v_b_04(net3976[0:47]),
     .sp4_r_v_b_03(net3977[0:47]), .sp4_r_v_b_02(net3978[0:47]),
     .sp4_r_v_b_01(sp4_v_b_14_17[47:0]), .sp4_h_r_04(net3980[0:47]),
     .sp4_h_r_03(net3981[0:47]), .sp4_h_r_02(net3982[0:47]),
     .sp4_h_r_01(net3983[0:47]), .sp4_h_l_03(net3655[0:47]),
     .sp4_h_l_02(net3656[0:47]), .sp4_h_l_01(net3657[0:47]),
     .bl(bl[707:654]), .bot_op_01(bot_op_13_17[7:0]),
     .sp12_h_l_01(net3646[0:23]), .sp12_h_l_02(net3645[0:23]),
     .sp12_h_l_03(net3644[0:23]), .sp12_h_l_04(net3643[0:23]),
     .sp4_v_b_04(net3650[0:47]), .sp4_v_b_03(net3651[0:47]),
     .sp4_v_b_02(net3652[0:47]), .bnr_op_01(bnr_op_13_17[7:0]),
     .sp4_h_l_05(net3682[0:47]), .sp4_h_l_06(net3681[0:47]),
     .sp4_h_l_07(net3680[0:47]), .sp4_h_l_08(net3679[0:47]),
     .sp4_h_l_09(net3678[0:47]), .sp4_h_l_10(net3677[0:47]),
     .sp4_h_r_10(net4003[0:47]), .sp4_h_r_09(net4004[0:47]),
     .sp4_h_r_08(net4005[0:47]), .sp4_h_r_07(net4006[0:47]),
     .sp4_h_r_06(net4007[0:47]), .sp4_h_r_05(net4008[0:47]),
     .slf_op_05(net3694[0:7]), .slf_op_06(net3693[0:7]),
     .slf_op_07(net3692[0:7]), .slf_op_08(net3691[0:7]),
     .slf_op_09(net3690[0:7]), .slf_op_10(net3689[0:7]),
     .rgt_op_10(net4015[0:7]), .rgt_op_09(net4016[0:7]),
     .rgt_op_08(net4017[0:7]), .rgt_op_07(net4018[0:7]),
     .rgt_op_06(net4019[0:7]), .rgt_op_05(net4020[0:7]),
     .lft_op_10(net2711[0:7]), .lft_op_09(net2712[0:7]),
     .lft_op_08(net2713[0:7]), .lft_op_07(net2714[0:7]),
     .lft_op_06(net2715[0:7]), .lft_op_05(net2716[0:7]),
     .sp12_h_l_10(net3702[0:23]), .sp12_h_r_10(net4028[0:23]),
     .sp12_h_l_09(net3711[0:23]), .sp12_h_l_08(net3710[0:23]),
     .sp12_h_l_07(net3709[0:23]), .sp12_h_l_06(net3708[0:23]),
     .sp12_h_r_05(net4033[0:23]), .sp12_h_r_06(net4034[0:23]),
     .sp12_h_r_07(net4035[0:23]), .sp12_h_r_08(net4036[0:23]),
     .sp12_h_r_09(net4037[0:23]), .sp12_h_l_05(net3707[0:23]),
     .sp4_r_v_b_05(net4039[0:47]), .sp4_r_v_b_06(net4040[0:47]),
     .sp4_r_v_b_07(net4041[0:47]), .sp4_r_v_b_08(net4042[0:47]),
     .sp4_r_v_b_09(net4043[0:47]), .sp4_r_v_b_10(net4044[0:47]),
     .sp4_v_b_10(net3718[0:47]), .sp4_v_b_09(net3717[0:47]),
     .sp4_v_b_08(net3716[0:47]), .sp4_v_b_07(net3715[0:47]),
     .sp4_v_b_06(net3714[0:47]), .sp4_v_b_05(net3713[0:47]),
     .sp4_v_t_16(net4051[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net4054[0:47]),
     .sp4_h_r_12(net4055[0:47]), .sp4_h_r_13(net4056[0:47]),
     .sp4_h_r_14(net4057[0:47]), .sp4_h_r_15(net4058[0:47]),
     .sp4_h_r_16(net4059[0:47]), .sp4_h_l_16(net3733[0:47]),
     .sp4_h_l_15(net3732[0:47]), .sp4_h_l_14(net3731[0:47]),
     .sp4_h_l_13(net3730[0:47]), .sp4_h_l_12(net3729[0:47]),
     .sp4_h_l_11(net3728[0:47]), .tnr_op_16({slf_op_14_33[3],
     slf_op_14_33[2], slf_op_14_33[1], slf_op_14_33[0],
     slf_op_14_33[3], slf_op_14_33[2], slf_op_14_33[1],
     slf_op_14_33[0]}), .tnl_op_16({slf_op_12_33[3], slf_op_12_33[2],
     slf_op_12_33[1], slf_op_12_33[0], slf_op_12_33[3],
     slf_op_12_33[2], slf_op_12_33[1], slf_op_12_33[0]}),
     .lft_op_16(net2643[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net3750[0:7]), .slf_op_14(net3749[0:7]),
     .slf_op_13(net3752[0:7]), .slf_op_12(net3751[0:7]),
     .slf_op_11(net3753[0:7]), .rgt_op_14(net4075[0:7]),
     .rgt_op_15(net4076[0:7]), .rgt_op_12(net4077[0:7]),
     .rgt_op_13(net4078[0:7]), .rgt_op_11(net4079[0:7]),
     .sp4_v_b_16(net3760[0:47]), .sp4_v_b_14(net3763[0:47]),
     .sp4_v_b_15(net3761[0:47]), .sp4_v_b_13(net3762[0:47]),
     .sp4_v_b_11(net3765[0:47]), .sp4_v_b_12(net3764[0:47]),
     .sp4_r_v_b_16(net4086[0:47]), .sp4_r_v_b_15(net4087[0:47]),
     .sp4_r_v_b_13(net4088[0:47]), .sp4_r_v_b_14(net4089[0:47]),
     .sp4_r_v_b_12(net4090[0:47]), .sp4_r_v_b_11(net4091[0:47]),
     .sp12_h_l_16(net3772[0:23]), .sp12_h_l_15(net3774[0:23]),
     .sp12_h_l_14(net3773[0:23]), .sp12_h_l_13(net3776[0:23]),
     .sp12_h_l_12(net3775[0:23]), .sp12_h_l_11(net3777[0:23]),
     .sp12_h_r_16(net4098[0:23]), .sp12_h_r_14(net4099[0:23]),
     .sp12_h_r_15(net4100[0:23]), .sp12_h_r_12(net4101[0:23]),
     .sp12_h_r_13(net4102[0:23]), .sp12_h_r_11(net4103[0:23]),
     .lft_op_14(net2771[0:7]), .lft_op_15(net2772[0:7]),
     .lft_op_12(net2773[0:7]), .lft_op_11(net2775[0:7]),
     .lft_op_13(net2774[0:7]));
array_LT1x16top I_it_09_top ( .glb_netwk(net4136[0:7]),
     .sp12_v_t_16(net4109[0:23]), .rgt_op_16(net2184[0:7]),
     .top_op_16({slf_op_09_33[3], slf_op_09_33[2], slf_op_09_33[1],
     slf_op_09_33[0], slf_op_09_33[3], slf_op_09_33[2],
     slf_op_09_33[1], slf_op_09_33[0]}), .rgt_op_03(net4112[0:7]),
     .slf_op_02(net2259[0:7]), .rgt_op_02(net4114[0:7]),
     .rgt_op_01(slf_op_10_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3796[0:7]), .lft_op_03(net3786[0:7]),
     .lft_op_02(net3788[0:7]), .lft_op_01(slf_op_08_17[7:0]),
     .rgt_op_04(net4122[0:7]), .carry_in(carry_in_09_17),
     .bnl_op_01(bnl_op_09_17[7:0]), .slf_op_04(net2257[0:7]),
     .slf_op_03(net2260[0:7]), .slf_op_01(slf_op_09_17[7:0]),
     .sp4_h_l_04(net2248[0:47]), .carry_out(net4129),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_09_17[23:0]),
     .sp12_h_r_04(net4132[0:23]), .sp12_h_r_03(net4133[0:23]),
     .sp12_h_r_02(net4134[0:23]), .sp12_h_r_01(net4135[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2316[0:7]),
     .sp4_v_b_01(sp4_v_b_09_17[47:0]), .sp4_r_v_b_04(net4139[0:47]),
     .sp4_r_v_b_03(net4140[0:47]), .sp4_r_v_b_02(net4141[0:47]),
     .sp4_r_v_b_01(sp4_v_b_10_17[47:0]), .sp4_h_r_04(net4143[0:47]),
     .sp4_h_r_03(net4144[0:47]), .sp4_h_r_02(net4145[0:47]),
     .sp4_h_r_01(net4146[0:47]), .sp4_h_l_03(net2247[0:47]),
     .sp4_h_l_02(net2246[0:47]), .sp4_h_l_01(net2245[0:47]),
     .bl(bl[491:438]), .bot_op_01(bot_op_09_17[7:0]),
     .sp12_h_l_01(net2282[0:23]), .sp12_h_l_02(net2280[0:23]),
     .sp12_h_l_03(net2349[0:23]), .sp12_h_l_04(net2279[0:23]),
     .sp4_v_b_04(net2320[0:47]), .sp4_v_b_03(net2322[0:47]),
     .sp4_v_b_02(net2324[0:47]), .bnr_op_01(bnr_op_09_17[7:0]),
     .sp4_h_l_05(net2238[0:47]), .sp4_h_l_06(net2240[0:47]),
     .sp4_h_l_07(net2292[0:47]), .sp4_h_l_08(net2291[0:47]),
     .sp4_h_l_09(net2290[0:47]), .sp4_h_l_10(net2289[0:47]),
     .sp4_h_r_10(net4166[0:47]), .sp4_h_r_09(net4167[0:47]),
     .sp4_h_r_08(net4168[0:47]), .sp4_h_r_07(net4169[0:47]),
     .sp4_h_r_06(net4170[0:47]), .sp4_h_r_05(net4171[0:47]),
     .slf_op_05(net2251[0:7]), .slf_op_06(net2250[0:7]),
     .slf_op_07(net2267[0:7]), .slf_op_08(net2266[0:7]),
     .slf_op_09(net2265[0:7]), .slf_op_10(net2268[0:7]),
     .rgt_op_10(net4178[0:7]), .rgt_op_09(net4179[0:7]),
     .rgt_op_08(net4180[0:7]), .rgt_op_07(net4181[0:7]),
     .rgt_op_06(net4182[0:7]), .rgt_op_05(net4183[0:7]),
     .lft_op_10(net3852[0:7]), .lft_op_09(net3853[0:7]),
     .lft_op_08(net3854[0:7]), .lft_op_07(net3855[0:7]),
     .lft_op_06(net3856[0:7]), .lft_op_05(net3857[0:7]),
     .sp12_h_l_10(net2281[0:23]), .sp12_h_r_10(net4191[0:23]),
     .sp12_h_l_09(net2351[0:23]), .sp12_h_l_08(net2353[0:23]),
     .sp12_h_l_07(net2342[0:23]), .sp12_h_l_06(net2356[0:23]),
     .sp12_h_r_05(net4196[0:23]), .sp12_h_r_06(net4197[0:23]),
     .sp12_h_r_07(net4198[0:23]), .sp12_h_r_08(net4199[0:23]),
     .sp12_h_r_09(net4200[0:23]), .sp12_h_l_05(net2354[0:23]),
     .sp4_r_v_b_05(net4202[0:47]), .sp4_r_v_b_06(net4203[0:47]),
     .sp4_r_v_b_07(net4204[0:47]), .sp4_r_v_b_08(net4205[0:47]),
     .sp4_r_v_b_09(net4206[0:47]), .sp4_r_v_b_10(net4207[0:47]),
     .sp4_v_b_10(net2285[0:47]), .sp4_v_b_09(net2286[0:47]),
     .sp4_v_b_08(net2287[0:47]), .sp4_v_b_07(net2288[0:47]),
     .sp4_v_b_06(net2319[0:47]), .sp4_v_b_05(net2315[0:47]),
     .sp4_v_t_16(net4214[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net4217[0:47]),
     .sp4_h_r_12(net4218[0:47]), .sp4_h_r_13(net4219[0:47]),
     .sp4_h_r_14(net4220[0:47]), .sp4_h_r_15(net4221[0:47]),
     .sp4_h_r_16(net4222[0:47]), .sp4_h_l_16(net2337[0:47]),
     .sp4_h_l_15(net2335[0:47]), .sp4_h_l_14(net2338[0:47]),
     .sp4_h_l_13(net2340[0:47]), .sp4_h_l_12(net2343[0:47]),
     .sp4_h_l_11(net2346[0:47]), .tnr_op_16({slf_op_10_33[3],
     slf_op_10_33[2], slf_op_10_33[1], slf_op_10_33[0],
     slf_op_10_33[3], slf_op_10_33[2], slf_op_10_33[1],
     slf_op_10_33[0]}), .tnl_op_16({slf_op_08_33[3], slf_op_08_33[2],
     slf_op_08_33[1], slf_op_08_33[0], slf_op_08_33[3],
     slf_op_08_33[2], slf_op_08_33[1], slf_op_08_33[0]}),
     .lft_op_16(net2164[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net2317[0:7]), .slf_op_14(net2333[0:7]),
     .slf_op_13(net2332[0:7]), .slf_op_12(net2331[0:7]),
     .slf_op_11(net2330[0:7]), .rgt_op_14(net4238[0:7]),
     .rgt_op_15(net4239[0:7]), .rgt_op_12(net4240[0:7]),
     .rgt_op_13(net4241[0:7]), .rgt_op_11(net4242[0:7]),
     .sp4_v_b_16(net2224[0:47]), .sp4_v_b_14(net2222[0:47]),
     .sp4_v_b_15(net2223[0:47]), .sp4_v_b_13(net2218[0:47]),
     .sp4_v_b_11(net2215[0:47]), .sp4_v_b_12(net2213[0:47]),
     .sp4_r_v_b_16(net4249[0:47]), .sp4_r_v_b_15(net4250[0:47]),
     .sp4_r_v_b_13(net4251[0:47]), .sp4_r_v_b_14(net4252[0:47]),
     .sp4_r_v_b_12(net4253[0:47]), .sp4_r_v_b_11(net4254[0:47]),
     .sp12_h_l_16(net2231[0:23]), .sp12_h_l_15(net2229[0:23]),
     .sp12_h_l_14(net2235[0:23]), .sp12_h_l_13(net2226[0:23]),
     .sp12_h_l_12(net2228[0:23]), .sp12_h_l_11(net2236[0:23]),
     .sp12_h_r_16(net4261[0:23]), .sp12_h_r_14(net4262[0:23]),
     .sp12_h_r_15(net4263[0:23]), .sp12_h_r_12(net4264[0:23]),
     .sp12_h_r_13(net4265[0:23]), .sp12_h_r_11(net4266[0:23]),
     .lft_op_14(net3912[0:7]), .lft_op_15(net3913[0:7]),
     .lft_op_12(net3914[0:7]), .lft_op_11(net3916[0:7]),
     .lft_op_13(net3915[0:7]));
array_LT1x16top I_lt_02_top ( .glb_netwk(net4299[0:7]),
     .sp12_v_t_16(net4272[0:23]), .rgt_op_16(net2177[0:7]),
     .top_op_16({slf_op_02_33[3], slf_op_02_33[2], slf_op_02_33[1],
     slf_op_02_33[0], slf_op_02_33[3], slf_op_02_33[2],
     slf_op_02_33[1], slf_op_02_33[0]}), .rgt_op_03(net4275[0:7]),
     .slf_op_02(net4440[0:7]), .rgt_op_02(net4277[0:7]),
     .rgt_op_01(slf_op_03_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net2436[0:7]), .lft_op_03(net2437[0:7]),
     .lft_op_02(net2438[0:7]), .lft_op_01(slf_op_01_17[7:0]),
     .rgt_op_04(net4285[0:7]), .carry_in(carry_in_02_17),
     .bnl_op_01(bnl_op_02_17[7:0]), .slf_op_04(net4448[0:7]),
     .slf_op_03(net4438[0:7]), .slf_op_01(slf_op_02_17[7:0]),
     .sp4_h_l_04(net4469[0:47]), .carry_out(net4292),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_02_17[23:0]),
     .sp12_h_r_04(net4295[0:23]), .sp12_h_r_03(net4296[0:23]),
     .sp12_h_r_02(net4297[0:23]), .sp12_h_r_01(net4298[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net4436[0:7]),
     .sp4_v_b_01(sp4_v_b_02_17[47:0]), .sp4_r_v_b_04(net4302[0:47]),
     .sp4_r_v_b_03(net4303[0:47]), .sp4_r_v_b_02(net4304[0:47]),
     .sp4_r_v_b_01(sp4_v_b_03_17[47:0]), .sp4_h_r_04(net4306[0:47]),
     .sp4_h_r_03(net4307[0:47]), .sp4_h_r_02(net4308[0:47]),
     .sp4_h_r_01(net4309[0:47]), .sp4_h_l_03(net4470[0:47]),
     .sp4_h_l_02(net4471[0:47]), .sp4_h_l_01(net4472[0:47]),
     .bl(bl[125:72]), .bot_op_01(bot_op_02_17[7:0]),
     .sp12_h_l_01(net4461[0:23]), .sp12_h_l_02(net4460[0:23]),
     .sp12_h_l_03(net4459[0:23]), .sp12_h_l_04(net4458[0:23]),
     .sp4_v_b_04(net4465[0:47]), .sp4_v_b_03(net4466[0:47]),
     .sp4_v_b_02(net4467[0:47]), .bnr_op_01(bnr_op_02_17[7:0]),
     .sp4_h_l_05(net4497[0:47]), .sp4_h_l_06(net4496[0:47]),
     .sp4_h_l_07(net4495[0:47]), .sp4_h_l_08(net4494[0:47]),
     .sp4_h_l_09(net4493[0:47]), .sp4_h_l_10(net4492[0:47]),
     .sp4_h_r_10(net4329[0:47]), .sp4_h_r_09(net4330[0:47]),
     .sp4_h_r_08(net4331[0:47]), .sp4_h_r_07(net4332[0:47]),
     .sp4_h_r_06(net4333[0:47]), .sp4_h_r_05(net4334[0:47]),
     .slf_op_05(net4509[0:7]), .slf_op_06(net4508[0:7]),
     .slf_op_07(net4507[0:7]), .slf_op_08(net4506[0:7]),
     .slf_op_09(net4505[0:7]), .slf_op_10(net4504[0:7]),
     .rgt_op_10(net4341[0:7]), .rgt_op_09(net4342[0:7]),
     .rgt_op_08(net4343[0:7]), .rgt_op_07(net4344[0:7]),
     .rgt_op_06(net4345[0:7]), .rgt_op_05(net4346[0:7]),
     .lft_op_10(net2397[0:7]), .lft_op_09(net2398[0:7]),
     .lft_op_08(net2399[0:7]), .lft_op_07(net2400[0:7]),
     .lft_op_06(net2434[0:7]), .lft_op_05(net2435[0:7]),
     .sp12_h_l_10(net4517[0:23]), .sp12_h_r_10(net4354[0:23]),
     .sp12_h_l_09(net4526[0:23]), .sp12_h_l_08(net4525[0:23]),
     .sp12_h_l_07(net4524[0:23]), .sp12_h_l_06(net4523[0:23]),
     .sp12_h_r_05(net4359[0:23]), .sp12_h_r_06(net4360[0:23]),
     .sp12_h_r_07(net4361[0:23]), .sp12_h_r_08(net4362[0:23]),
     .sp12_h_r_09(net4363[0:23]), .sp12_h_l_05(net4522[0:23]),
     .sp4_r_v_b_05(net4365[0:47]), .sp4_r_v_b_06(net4366[0:47]),
     .sp4_r_v_b_07(net4367[0:47]), .sp4_r_v_b_08(net4368[0:47]),
     .sp4_r_v_b_09(net4369[0:47]), .sp4_r_v_b_10(net4370[0:47]),
     .sp4_v_b_10(net4533[0:47]), .sp4_v_b_09(net4532[0:47]),
     .sp4_v_b_08(net4531[0:47]), .sp4_v_b_07(net4530[0:47]),
     .sp4_v_b_06(net4529[0:47]), .sp4_v_b_05(net4528[0:47]),
     .sp4_v_t_16(net4377[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net4380[0:47]),
     .sp4_h_r_12(net4381[0:47]), .sp4_h_r_13(net4382[0:47]),
     .sp4_h_r_14(net4383[0:47]), .sp4_h_r_15(net4384[0:47]),
     .sp4_h_r_16(net4385[0:47]), .sp4_h_l_16(net4548[0:47]),
     .sp4_h_l_15(net4547[0:47]), .sp4_h_l_14(net4546[0:47]),
     .sp4_h_l_13(net4545[0:47]), .sp4_h_l_12(net4544[0:47]),
     .sp4_h_l_11(net4543[0:47]), .tnr_op_16({slf_op_03_33[3],
     slf_op_03_33[2], slf_op_03_33[1], slf_op_03_33[0],
     slf_op_03_33[3], slf_op_03_33[2], slf_op_03_33[1],
     slf_op_03_33[0]}), .tnl_op_16({slf_op_01_33[3], slf_op_01_33[2],
     slf_op_01_33[1], slf_op_01_33[0], slf_op_01_33[3],
     slf_op_01_33[2], slf_op_01_33[1], slf_op_01_33[0]}),
     .lft_op_16(net2175[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net4565[0:7]), .slf_op_14(net4564[0:7]),
     .slf_op_13(net4567[0:7]), .slf_op_12(net4566[0:7]),
     .slf_op_11(net4568[0:7]), .rgt_op_14(net4401[0:7]),
     .rgt_op_15(net4402[0:7]), .rgt_op_12(net4403[0:7]),
     .rgt_op_13(net4404[0:7]), .rgt_op_11(net4405[0:7]),
     .sp4_v_b_16(net4575[0:47]), .sp4_v_b_14(net4578[0:47]),
     .sp4_v_b_15(net4576[0:47]), .sp4_v_b_13(net4577[0:47]),
     .sp4_v_b_11(net4580[0:47]), .sp4_v_b_12(net4579[0:47]),
     .sp4_r_v_b_16(net4412[0:47]), .sp4_r_v_b_15(net4413[0:47]),
     .sp4_r_v_b_13(net4414[0:47]), .sp4_r_v_b_14(net4415[0:47]),
     .sp4_r_v_b_12(net4416[0:47]), .sp4_r_v_b_11(net4417[0:47]),
     .sp12_h_l_16(net4587[0:23]), .sp12_h_l_15(net4589[0:23]),
     .sp12_h_l_14(net4588[0:23]), .sp12_h_l_13(net4591[0:23]),
     .sp12_h_l_12(net4590[0:23]), .sp12_h_l_11(net4592[0:23]),
     .sp12_h_r_16(net4424[0:23]), .sp12_h_r_14(net4425[0:23]),
     .sp12_h_r_15(net4426[0:23]), .sp12_h_r_12(net4427[0:23]),
     .sp12_h_r_13(net4428[0:23]), .sp12_h_r_11(net4429[0:23]),
     .lft_op_14(net2393[0:7]), .lft_op_15(net2433[0:7]),
     .lft_op_12(net2395[0:7]), .lft_op_11(net2396[0:7]),
     .lft_op_13(net2394[0:7]));
array_LT1x16top I_lt_01_top ( .glb_netwk(net4462[0:7]),
     .sp12_v_t_16(net4435[0:23]), .rgt_op_16(net4436[0:7]),
     .top_op_16({slf_op_01_33[3], slf_op_01_33[2], slf_op_01_33[1],
     slf_op_01_33[0], slf_op_01_33[3], slf_op_01_33[2],
     slf_op_01_33[1], slf_op_01_33[0]}), .rgt_op_03(net4438[0:7]),
     .slf_op_02(net2438[0:7]), .rgt_op_02(net4440[0:7]),
     .rgt_op_01(slf_op_02_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04({slf_op_00_20[3], slf_op_00_20[2], slf_op_00_20[1],
     slf_op_00_20[0], slf_op_00_20[3], slf_op_00_20[2],
     slf_op_00_20[1], slf_op_00_20[0]}), .lft_op_03({slf_op_00_19[3],
     slf_op_00_19[2], slf_op_00_19[1], slf_op_00_19[0],
     slf_op_00_19[3], slf_op_00_19[2], slf_op_00_19[1],
     slf_op_00_19[0]}), .lft_op_02({slf_op_00_18[3], slf_op_00_18[2],
     slf_op_00_18[1], slf_op_00_18[0], slf_op_00_18[3],
     slf_op_00_18[2], slf_op_00_18[1], slf_op_00_18[0]}),
     .lft_op_01({slf_op_00_17[3], slf_op_00_17[2], slf_op_00_17[1],
     slf_op_00_17[0], slf_op_00_17[3], slf_op_00_17[2],
     slf_op_00_17[1], slf_op_00_17[0]}), .rgt_op_04(net4448[0:7]),
     .carry_in(carry_in_01_17), .bnl_op_01(bnl_op_01_17[7:0]),
     .slf_op_04(net2436[0:7]), .slf_op_03(net2437[0:7]),
     .slf_op_01(slf_op_01_17[7:0]), .sp4_h_l_04(net2431[0:47]),
     .carry_out(net4455), .vdd_cntl(vdd_cntl_l[255:0]),
     .sp12_v_b__01(sp12_v_b_01_17[23:0]), .sp12_h_r_04(net4458[0:23]),
     .sp12_h_r_03(net4459[0:23]), .sp12_h_r_02(net4460[0:23]),
     .sp12_h_r_01(net4461[0:23]), .glb_netwk_col(clk_tree_drv[7:0]),
     .slf_op_16(net2175[0:7]), .sp4_v_b_01(sp4_v_b_01_17[47:0]),
     .sp4_r_v_b_04(net4465[0:47]), .sp4_r_v_b_03(net4466[0:47]),
     .sp4_r_v_b_02(net4467[0:47]), .sp4_r_v_b_01(sp4_v_b_02_17[47:0]),
     .sp4_h_r_04(net4469[0:47]), .sp4_h_r_03(net4470[0:47]),
     .sp4_h_r_02(net4471[0:47]), .sp4_h_r_01(net4472[0:47]),
     .sp4_h_l_03(net2430[0:47]), .sp4_h_l_02(net2429[0:47]),
     .sp4_h_l_01(net2428[0:47]), .bl(bl[71:18]),
     .bot_op_01(bot_op_01_17[7:0]), .sp12_h_l_01(net2460[0:23]),
     .sp12_h_l_02(net2458[0:23]), .sp12_h_l_03(net2459[0:23]),
     .sp12_h_l_04(net2457[0:23]), .sp4_v_b_04(net4482[0:47]),
     .sp4_v_b_03(net4483[0:47]), .sp4_v_b_02(net4484[0:47]),
     .bnr_op_01(bnr_op_01_17[7:0]), .sp4_h_l_05(net2440[0:47]),
     .sp4_h_l_06(net2441[0:47]), .sp4_h_l_07(net2402[0:47]),
     .sp4_h_l_08(net2413[0:47]), .sp4_h_l_09(net2412[0:47]),
     .sp4_h_l_10(net2401[0:47]), .sp4_h_r_10(net4492[0:47]),
     .sp4_h_r_09(net4493[0:47]), .sp4_h_r_08(net4494[0:47]),
     .sp4_h_r_07(net4495[0:47]), .sp4_h_r_06(net4496[0:47]),
     .sp4_h_r_05(net4497[0:47]), .slf_op_05(net2435[0:7]),
     .slf_op_06(net2434[0:7]), .slf_op_07(net2400[0:7]),
     .slf_op_08(net2399[0:7]), .slf_op_09(net2398[0:7]),
     .slf_op_10(net2397[0:7]), .rgt_op_10(net4504[0:7]),
     .rgt_op_09(net4505[0:7]), .rgt_op_08(net4506[0:7]),
     .rgt_op_07(net4507[0:7]), .rgt_op_06(net4508[0:7]),
     .rgt_op_05(net4509[0:7]), .lft_op_10({slf_op_00_26[3],
     slf_op_00_26[2], slf_op_00_26[1], slf_op_00_26[0],
     slf_op_00_26[3], slf_op_00_26[2], slf_op_00_26[1],
     slf_op_00_26[0]}), .lft_op_09({slf_op_00_25[3], slf_op_00_25[2],
     slf_op_00_25[1], slf_op_00_25[0], slf_op_00_25[3],
     slf_op_00_25[2], slf_op_00_25[1], slf_op_00_25[0]}),
     .lft_op_08({slf_op_00_24[3], slf_op_00_24[2], slf_op_00_24[1],
     slf_op_00_24[0], slf_op_00_24[3], slf_op_00_24[2],
     slf_op_00_24[1], slf_op_00_24[0]}), .lft_op_07({slf_op_00_23[3],
     slf_op_00_23[2], slf_op_00_23[1], slf_op_00_23[0],
     slf_op_00_23[3], slf_op_00_23[2], slf_op_00_23[1],
     slf_op_00_23[0]}), .lft_op_06({slf_op_00_22[3], slf_op_00_22[2],
     slf_op_00_22[1], slf_op_00_22[0], slf_op_00_22[3],
     slf_op_00_22[2], slf_op_00_22[1], slf_op_00_22[0]}),
     .lft_op_05({slf_op_00_21[3], slf_op_00_21[2], slf_op_00_21[1],
     slf_op_00_21[0], slf_op_00_21[3], slf_op_00_21[2],
     slf_op_00_21[1], slf_op_00_21[0]}), .sp12_h_l_10(net2451[0:23]),
     .sp12_h_r_10(net4517[0:23]), .sp12_h_l_09(net2452[0:23]),
     .sp12_h_l_08(net2453[0:23]), .sp12_h_l_07(net2454[0:23]),
     .sp12_h_l_06(net2455[0:23]), .sp12_h_r_05(net4522[0:23]),
     .sp12_h_r_06(net4523[0:23]), .sp12_h_r_07(net4524[0:23]),
     .sp12_h_r_08(net4525[0:23]), .sp12_h_r_09(net4526[0:23]),
     .sp12_h_l_05(net2456[0:23]), .sp4_r_v_b_05(net4528[0:47]),
     .sp4_r_v_b_06(net4529[0:47]), .sp4_r_v_b_07(net4530[0:47]),
     .sp4_r_v_b_08(net4531[0:47]), .sp4_r_v_b_09(net4532[0:47]),
     .sp4_r_v_b_10(net4533[0:47]), .sp4_v_b_10(net4534[0:47]),
     .sp4_v_b_09(net4535[0:47]), .sp4_v_b_08(net4536[0:47]),
     .sp4_v_b_07(net4537[0:47]), .sp4_v_b_06(net4538[0:47]),
     .sp4_v_b_05(net4539[0:47]), .sp4_v_t_16(net4540[0:47]),
     .pgate(pgate_l[255:0]), .reset_b(reset_l[255:0]),
     .sp4_h_r_11(net4543[0:47]), .sp4_h_r_12(net4544[0:47]),
     .sp4_h_r_13(net4545[0:47]), .sp4_h_r_14(net4546[0:47]),
     .sp4_h_r_15(net4547[0:47]), .sp4_h_r_16(net4548[0:47]),
     .sp4_h_l_16(net2418[0:47]), .sp4_h_l_15(net2419[0:47]),
     .sp4_h_l_14(net2424[0:47]), .sp4_h_l_13(net2425[0:47]),
     .sp4_h_l_12(net2426[0:47]), .sp4_h_l_11(net2427[0:47]),
     .tnr_op_16({slf_op_02_33[3], slf_op_02_33[2], slf_op_02_33[1],
     slf_op_02_33[0], slf_op_02_33[3], slf_op_02_33[2],
     slf_op_02_33[1], slf_op_02_33[0]}), .tnl_op_16({tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .lft_op_16({slf_op_00_32[3], slf_op_00_32[2], slf_op_00_32[1],
     slf_op_00_32[0], slf_op_00_32[3], slf_op_00_32[2],
     slf_op_00_32[1], slf_op_00_32[0]}), .wl(wl_l[255:0]),
     .slf_op_15(net2433[0:7]), .slf_op_14(net2393[0:7]),
     .slf_op_13(net2394[0:7]), .slf_op_12(net2395[0:7]),
     .slf_op_11(net2396[0:7]), .rgt_op_14(net4564[0:7]),
     .rgt_op_15(net4565[0:7]), .rgt_op_12(net4566[0:7]),
     .rgt_op_13(net4567[0:7]), .rgt_op_11(net4568[0:7]),
     .sp4_v_b_16(net4569[0:47]), .sp4_v_b_14(net4570[0:47]),
     .sp4_v_b_15(net4571[0:47]), .sp4_v_b_13(net4572[0:47]),
     .sp4_v_b_11(net4573[0:47]), .sp4_v_b_12(net4574[0:47]),
     .sp4_r_v_b_16(net4575[0:47]), .sp4_r_v_b_15(net4576[0:47]),
     .sp4_r_v_b_13(net4577[0:47]), .sp4_r_v_b_14(net4578[0:47]),
     .sp4_r_v_b_12(net4579[0:47]), .sp4_r_v_b_11(net4580[0:47]),
     .sp12_h_l_16(net2445[0:23]), .sp12_h_l_15(net2446[0:23]),
     .sp12_h_l_14(net2447[0:23]), .sp12_h_l_13(net2448[0:23]),
     .sp12_h_l_12(net2449[0:23]), .sp12_h_l_11(net2450[0:23]),
     .sp12_h_r_16(net4587[0:23]), .sp12_h_r_14(net4588[0:23]),
     .sp12_h_r_15(net4589[0:23]), .sp12_h_r_12(net4590[0:23]),
     .sp12_h_r_13(net4591[0:23]), .sp12_h_r_11(net4592[0:23]),
     .lft_op_14({slf_op_00_30[3], slf_op_00_30[2], slf_op_00_30[1],
     slf_op_00_30[0], slf_op_00_30[3], slf_op_00_30[2],
     slf_op_00_30[1], slf_op_00_30[0]}), .lft_op_15({slf_op_00_31[3],
     slf_op_00_31[2], slf_op_00_31[1], slf_op_00_31[0],
     slf_op_00_31[3], slf_op_00_31[2], slf_op_00_31[1],
     slf_op_00_31[0]}), .lft_op_12({slf_op_00_28[3], slf_op_00_28[2],
     slf_op_00_28[1], slf_op_00_28[0], slf_op_00_28[3],
     slf_op_00_28[2], slf_op_00_28[1], slf_op_00_28[0]}),
     .lft_op_11({slf_op_00_27[3], slf_op_00_27[2], slf_op_00_27[1],
     slf_op_00_27[0], slf_op_00_27[3], slf_op_00_27[2],
     slf_op_00_27[1], slf_op_00_27[0]}), .lft_op_13({slf_op_00_29[3],
     slf_op_00_29[2], slf_op_00_29[1], slf_op_00_29[0],
     slf_op_00_29[3], slf_op_00_29[2], slf_op_00_29[1],
     slf_op_00_29[0]}));
array_LT1x16top I_it_16_top ( .glb_netwk(net4625[0:7]),
     .sp12_v_t_16(net4598[0:23]), .rgt_op_16(rgt_op_16_32[7:0]),
     .top_op_16({slf_op_16_33[3], slf_op_16_33[2], slf_op_16_33[1],
     slf_op_16_33[0], slf_op_16_33[3], slf_op_16_33[2],
     slf_op_16_33[1], slf_op_16_33[0]}), .rgt_op_03(rgt_op_16_19[7:0]),
     .slf_op_02(slf_op_16_18[7:0]), .rgt_op_02(rgt_op_16_18[7:0]),
     .rgt_op_01(rgt_op_16_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net3470[0:7]), .lft_op_03(net3460[0:7]),
     .lft_op_02(net3462[0:7]), .lft_op_01(slf_op_15_17[7:0]),
     .rgt_op_04(rgt_op_16_20[7:0]), .carry_in(carry_in_16_17),
     .bnl_op_01(bnl_op_16_17[7:0]), .slf_op_04(slf_op_16_20[7:0]),
     .slf_op_03(slf_op_16_19[7:0]), .slf_op_01(slf_op_16_17[7:0]),
     .sp4_h_l_04(net3002[0:47]), .carry_out(net4618),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_16_17[23:0]),
     .sp12_h_r_04(sp12_h_r_16_20[23:0]),
     .sp12_h_r_03(sp12_h_r_16_19[23:0]),
     .sp12_h_r_02(sp12_h_r_16_18[23:0]),
     .sp12_h_r_01(sp12_h_r_16_17[23:0]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(slf_op_16_32[7:0]),
     .sp4_v_b_01(sp4_v_b_16_17[47:0]),
     .sp4_r_v_b_04(sp4_r_v_b_16_20[47:0]),
     .sp4_r_v_b_03(sp4_r_v_b_16_19[47:0]),
     .sp4_r_v_b_02(sp4_r_v_b_16_18[47:0]),
     .sp4_r_v_b_01(sp4_r_v_b_16_17[47:0]),
     .sp4_h_r_04(sp4_h_r_16_20[47:0]),
     .sp4_h_r_03(sp4_h_r_16_19[47:0]),
     .sp4_h_r_02(sp4_h_r_16_18[47:0]),
     .sp4_h_r_01(sp4_h_r_16_17[47:0]), .sp4_h_l_03(net3003[0:47]),
     .sp4_h_l_02(net3004[0:47]), .sp4_h_l_01(net3005[0:47]),
     .bl(bl[869:816]), .bot_op_01(bot_op_16_17[7:0]),
     .sp12_h_l_01(net2994[0:23]), .sp12_h_l_02(net2993[0:23]),
     .sp12_h_l_03(net2992[0:23]), .sp12_h_l_04(net2991[0:23]),
     .sp4_v_b_04(net2998[0:47]), .sp4_v_b_03(net2999[0:47]),
     .sp4_v_b_02(net3000[0:47]), .bnr_op_01(bnr_op_16_17[7:0]),
     .sp4_h_l_05(net3030[0:47]), .sp4_h_l_06(net3029[0:47]),
     .sp4_h_l_07(net3028[0:47]), .sp4_h_l_08(net3027[0:47]),
     .sp4_h_l_09(net3026[0:47]), .sp4_h_l_10(net3025[0:47]),
     .sp4_h_r_10(sp4_h_r_16_26[47:0]),
     .sp4_h_r_09(sp4_h_r_16_25[47:0]),
     .sp4_h_r_08(sp4_h_r_16_24[47:0]),
     .sp4_h_r_07(sp4_h_r_16_23[47:0]),
     .sp4_h_r_06(sp4_h_r_16_22[47:0]),
     .sp4_h_r_05(sp4_h_r_16_21[47:0]), .slf_op_05(slf_op_16_21[7:0]),
     .slf_op_06(slf_op_16_22[7:0]), .slf_op_07(slf_op_16_23[7:0]),
     .slf_op_08(slf_op_16_24[7:0]), .slf_op_09(slf_op_16_25[7:0]),
     .slf_op_10(slf_op_16_26[7:0]), .rgt_op_10(rgt_op_16_26[7:0]),
     .rgt_op_09(rgt_op_16_25[7:0]), .rgt_op_08(rgt_op_16_24[7:0]),
     .rgt_op_07(rgt_op_16_23[7:0]), .rgt_op_06(rgt_op_16_22[7:0]),
     .rgt_op_05(rgt_op_16_21[7:0]), .lft_op_10(net3526[0:7]),
     .lft_op_09(net3527[0:7]), .lft_op_08(net3528[0:7]),
     .lft_op_07(net3529[0:7]), .lft_op_06(net3530[0:7]),
     .lft_op_05(net3531[0:7]), .sp12_h_l_10(net3050[0:23]),
     .sp12_h_r_10(sp12_h_r_16_26[23:0]), .sp12_h_l_09(net3059[0:23]),
     .sp12_h_l_08(net3058[0:23]), .sp12_h_l_07(net3057[0:23]),
     .sp12_h_l_06(net3056[0:23]), .sp12_h_r_05(sp12_h_r_16_21[23:0]),
     .sp12_h_r_06(sp12_h_r_16_22[23:0]),
     .sp12_h_r_07(sp12_h_r_16_23[23:0]),
     .sp12_h_r_08(sp12_h_r_16_24[23:0]),
     .sp12_h_r_09(sp12_h_r_16_25[23:0]), .sp12_h_l_05(net3055[0:23]),
     .sp4_r_v_b_05(sp4_r_v_b_16_21[47:0]),
     .sp4_r_v_b_06(sp4_r_v_b_16_22[47:0]),
     .sp4_r_v_b_07(sp4_r_v_b_16_23[47:0]),
     .sp4_r_v_b_08(sp4_r_v_b_16_24[47:0]),
     .sp4_r_v_b_09(sp4_r_v_b_16_25[47:0]),
     .sp4_r_v_b_10(sp4_r_v_b_16_26[47:0]), .sp4_v_b_10(net3066[0:47]),
     .sp4_v_b_09(net3065[0:47]), .sp4_v_b_08(net3064[0:47]),
     .sp4_v_b_07(net3063[0:47]), .sp4_v_b_06(net3062[0:47]),
     .sp4_v_b_05(net3061[0:47]), .sp4_v_t_16(net4703[0:47]),
     .pgate(pgate_l[255:0]), .reset_b(reset_l[255:0]),
     .sp4_h_r_11(sp4_h_r_16_27[47:0]),
     .sp4_h_r_12(sp4_h_r_16_28[47:0]),
     .sp4_h_r_13(sp4_h_r_16_29[47:0]),
     .sp4_h_r_14(sp4_h_r_16_30[47:0]),
     .sp4_h_r_15(sp4_h_r_16_31[47:0]),
     .sp4_h_r_16(sp4_h_r_16_32[47:0]), .sp4_h_l_16(net3081[0:47]),
     .sp4_h_l_15(net3080[0:47]), .sp4_h_l_14(net3079[0:47]),
     .sp4_h_l_13(net3078[0:47]), .sp4_h_l_12(net3077[0:47]),
     .sp4_h_l_11(net3076[0:47]), .tnr_op_16({tnr_op_16_32[3],
     tnr_op_16_32[2], tnr_op_16_32[1], tnr_op_16_32[0],
     tnr_op_16_32[3], tnr_op_16_32[2], tnr_op_16_32[1],
     tnr_op_16_32[0]}), .tnl_op_16({slf_op_15_33[3], slf_op_15_33[2],
     slf_op_15_33[1], slf_op_15_33[0], slf_op_15_33[3],
     slf_op_15_33[2], slf_op_15_33[1], slf_op_15_33[0]}),
     .lft_op_16(net3458[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(slf_op_16_31[7:0]), .slf_op_14(slf_op_16_30[7:0]),
     .slf_op_13(slf_op_16_29[7:0]), .slf_op_12(slf_op_16_28[7:0]),
     .slf_op_11(slf_op_16_27[7:0]), .rgt_op_14(rgt_op_16_30[7:0]),
     .rgt_op_15(rgt_op_16_31[7:0]), .rgt_op_12(rgt_op_16_28[7:0]),
     .rgt_op_13(rgt_op_16_29[7:0]), .rgt_op_11(rgt_op_16_27[7:0]),
     .sp4_v_b_16(net3108[0:47]), .sp4_v_b_14(net3111[0:47]),
     .sp4_v_b_15(net3109[0:47]), .sp4_v_b_13(net3110[0:47]),
     .sp4_v_b_11(net3113[0:47]), .sp4_v_b_12(net3112[0:47]),
     .sp4_r_v_b_16(sp4_r_v_b_16_32[47:0]),
     .sp4_r_v_b_15(sp4_r_v_b_16_31[47:0]),
     .sp4_r_v_b_13(sp4_r_v_b_16_29[47:0]),
     .sp4_r_v_b_14(sp4_r_v_b_16_30[47:0]),
     .sp4_r_v_b_12(sp4_r_v_b_16_28[47:0]),
     .sp4_r_v_b_11(sp4_r_v_b_16_27[47:0]), .sp12_h_l_16(net3120[0:23]),
     .sp12_h_l_15(net3122[0:23]), .sp12_h_l_14(net3121[0:23]),
     .sp12_h_l_13(net3124[0:23]), .sp12_h_l_12(net3123[0:23]),
     .sp12_h_l_11(net3125[0:23]), .sp12_h_r_16(sp12_h_r_16_32[23:0]),
     .sp12_h_r_14(sp12_h_r_16_30[23:0]),
     .sp12_h_r_15(sp12_h_r_16_31[23:0]),
     .sp12_h_r_12(sp12_h_r_16_28[23:0]),
     .sp12_h_r_13(sp12_h_r_16_29[23:0]),
     .sp12_h_r_11(sp12_h_r_16_27[23:0]), .lft_op_14(net3586[0:7]),
     .lft_op_15(net3587[0:7]), .lft_op_12(net3588[0:7]),
     .lft_op_11(net3590[0:7]), .lft_op_13(net3589[0:7]));
array_LT1x16top I_it_04_top ( .glb_netwk(net4788[0:7]),
     .sp12_v_t_16(net4761[0:23]), .rgt_op_16(net2179[0:7]),
     .top_op_16({slf_op_04_33[3], slf_op_04_33[2], slf_op_04_33[1],
     slf_op_04_33[0], slf_op_04_33[3], slf_op_04_33[2],
     slf_op_04_33[1], slf_op_04_33[0]}), .rgt_op_03(net4764[0:7]),
     .slf_op_02(net3299[0:7]), .rgt_op_02(net4766[0:7]),
     .rgt_op_01(slf_op_05_17[7:0]), .purst(purst), .prog(prog),
     .lft_op_04(net4285[0:7]), .lft_op_03(net4275[0:7]),
     .lft_op_02(net4277[0:7]), .lft_op_01(slf_op_03_17[7:0]),
     .rgt_op_04(net4774[0:7]), .carry_in(carry_in_04_17),
     .bnl_op_01(bnl_op_04_17[7:0]), .slf_op_04(net3307[0:7]),
     .slf_op_03(net3297[0:7]), .slf_op_01(slf_op_04_17[7:0]),
     .sp4_h_l_04(net3328[0:47]), .carry_out(net4781),
     .vdd_cntl(vdd_cntl_l[255:0]), .sp12_v_b__01(sp12_v_b_04_17[23:0]),
     .sp12_h_r_04(net4784[0:23]), .sp12_h_r_03(net4785[0:23]),
     .sp12_h_r_02(net4786[0:23]), .sp12_h_r_01(net4787[0:23]),
     .glb_netwk_col(clk_tree_drv[7:0]), .slf_op_16(net2160[0:7]),
     .sp4_v_b_01(sp4_v_b_04_17[47:0]), .sp4_r_v_b_04(net4791[0:47]),
     .sp4_r_v_b_03(net4792[0:47]), .sp4_r_v_b_02(net4793[0:47]),
     .sp4_r_v_b_01(sp4_v_b_05_17[47:0]), .sp4_h_r_04(net4795[0:47]),
     .sp4_h_r_03(net4796[0:47]), .sp4_h_r_02(net4797[0:47]),
     .sp4_h_r_01(net4798[0:47]), .sp4_h_l_03(net3329[0:47]),
     .sp4_h_l_02(net3330[0:47]), .sp4_h_l_01(net3331[0:47]),
     .bl(bl[233:180]), .bot_op_01(bot_op_04_17[7:0]),
     .sp12_h_l_01(net3320[0:23]), .sp12_h_l_02(net3319[0:23]),
     .sp12_h_l_03(net3318[0:23]), .sp12_h_l_04(net3317[0:23]),
     .sp4_v_b_04(net3324[0:47]), .sp4_v_b_03(net3325[0:47]),
     .sp4_v_b_02(net3326[0:47]), .bnr_op_01(bnr_op_04_17[7:0]),
     .sp4_h_l_05(net3356[0:47]), .sp4_h_l_06(net3355[0:47]),
     .sp4_h_l_07(net3354[0:47]), .sp4_h_l_08(net3353[0:47]),
     .sp4_h_l_09(net3352[0:47]), .sp4_h_l_10(net3351[0:47]),
     .sp4_h_r_10(net4818[0:47]), .sp4_h_r_09(net4819[0:47]),
     .sp4_h_r_08(net4820[0:47]), .sp4_h_r_07(net4821[0:47]),
     .sp4_h_r_06(net4822[0:47]), .sp4_h_r_05(net4823[0:47]),
     .slf_op_05(net3368[0:7]), .slf_op_06(net3367[0:7]),
     .slf_op_07(net3366[0:7]), .slf_op_08(net3365[0:7]),
     .slf_op_09(net3364[0:7]), .slf_op_10(net3363[0:7]),
     .rgt_op_10(net4830[0:7]), .rgt_op_09(net4831[0:7]),
     .rgt_op_08(net4832[0:7]), .rgt_op_07(net4833[0:7]),
     .rgt_op_06(net4834[0:7]), .rgt_op_05(net4835[0:7]),
     .lft_op_10(net4341[0:7]), .lft_op_09(net4342[0:7]),
     .lft_op_08(net4343[0:7]), .lft_op_07(net4344[0:7]),
     .lft_op_06(net4345[0:7]), .lft_op_05(net4346[0:7]),
     .sp12_h_l_10(net3376[0:23]), .sp12_h_r_10(net4843[0:23]),
     .sp12_h_l_09(net3385[0:23]), .sp12_h_l_08(net3384[0:23]),
     .sp12_h_l_07(net3383[0:23]), .sp12_h_l_06(net3382[0:23]),
     .sp12_h_r_05(net4848[0:23]), .sp12_h_r_06(net4849[0:23]),
     .sp12_h_r_07(net4850[0:23]), .sp12_h_r_08(net4851[0:23]),
     .sp12_h_r_09(net4852[0:23]), .sp12_h_l_05(net3381[0:23]),
     .sp4_r_v_b_05(net4854[0:47]), .sp4_r_v_b_06(net4855[0:47]),
     .sp4_r_v_b_07(net4856[0:47]), .sp4_r_v_b_08(net4857[0:47]),
     .sp4_r_v_b_09(net4858[0:47]), .sp4_r_v_b_10(net4859[0:47]),
     .sp4_v_b_10(net3392[0:47]), .sp4_v_b_09(net3391[0:47]),
     .sp4_v_b_08(net3390[0:47]), .sp4_v_b_07(net3389[0:47]),
     .sp4_v_b_06(net3388[0:47]), .sp4_v_b_05(net3387[0:47]),
     .sp4_v_t_16(net4866[0:47]), .pgate(pgate_l[255:0]),
     .reset_b(reset_l[255:0]), .sp4_h_r_11(net4869[0:47]),
     .sp4_h_r_12(net4870[0:47]), .sp4_h_r_13(net4871[0:47]),
     .sp4_h_r_14(net4872[0:47]), .sp4_h_r_15(net4873[0:47]),
     .sp4_h_r_16(net4874[0:47]), .sp4_h_l_16(net3407[0:47]),
     .sp4_h_l_15(net3406[0:47]), .sp4_h_l_14(net3405[0:47]),
     .sp4_h_l_13(net3404[0:47]), .sp4_h_l_12(net3403[0:47]),
     .sp4_h_l_11(net3402[0:47]), .tnr_op_16({slf_op_05_33[3],
     slf_op_05_33[2], slf_op_05_33[1], slf_op_05_33[0],
     slf_op_05_33[3], slf_op_05_33[2], slf_op_05_33[1],
     slf_op_05_33[0]}), .tnl_op_16({slf_op_03_33[3], slf_op_03_33[2],
     slf_op_03_33[1], slf_op_03_33[0], slf_op_03_33[3],
     slf_op_03_33[2], slf_op_03_33[1], slf_op_03_33[0]}),
     .lft_op_16(net2177[0:7]), .wl(wl_l[255:0]),
     .slf_op_15(net3424[0:7]), .slf_op_14(net3423[0:7]),
     .slf_op_13(net3426[0:7]), .slf_op_12(net3425[0:7]),
     .slf_op_11(net3427[0:7]), .rgt_op_14(net4890[0:7]),
     .rgt_op_15(net4891[0:7]), .rgt_op_12(net4892[0:7]),
     .rgt_op_13(net4893[0:7]), .rgt_op_11(net4894[0:7]),
     .sp4_v_b_16(net3434[0:47]), .sp4_v_b_14(net3437[0:47]),
     .sp4_v_b_15(net3435[0:47]), .sp4_v_b_13(net3436[0:47]),
     .sp4_v_b_11(net3439[0:47]), .sp4_v_b_12(net3438[0:47]),
     .sp4_r_v_b_16(net4901[0:47]), .sp4_r_v_b_15(net4902[0:47]),
     .sp4_r_v_b_13(net4903[0:47]), .sp4_r_v_b_14(net4904[0:47]),
     .sp4_r_v_b_12(net4905[0:47]), .sp4_r_v_b_11(net4906[0:47]),
     .sp12_h_l_16(net3446[0:23]), .sp12_h_l_15(net3448[0:23]),
     .sp12_h_l_14(net3447[0:23]), .sp12_h_l_13(net3450[0:23]),
     .sp12_h_l_12(net3449[0:23]), .sp12_h_l_11(net3451[0:23]),
     .sp12_h_r_16(net4913[0:23]), .sp12_h_r_14(net4914[0:23]),
     .sp12_h_r_15(net4915[0:23]), .sp12_h_r_12(net4916[0:23]),
     .sp12_h_r_13(net4917[0:23]), .sp12_h_r_11(net4918[0:23]),
     .lft_op_14(net4401[0:7]), .lft_op_15(net4402[0:7]),
     .lft_op_12(net4403[0:7]), .lft_op_11(net4405[0:7]),
     .lft_op_13(net4404[0:7]));
bram_bufferx4 I332 ( .in(net02116), .out(ceb_o));
bram_bufferx4 I283 ( .in(net2066), .out(bs_en_o));
bram_bufferx4 I287 ( .in(net2047), .out(r_o));
bram_bufferx4 I288 ( .in(net4938), .out(shift_o));
bram_bufferx4 I289 ( .in(net4940), .out(mode_o));
bram_bufferx4 I286 ( .in(net2043), .out(update_o));
bram_bufferx4 I284 ( .in(net2049), .out(hiz_b_o));

endmodule
// Library - leafcell, Cell - bram_bufferx16_2inv, View - schematic
// LAST TIME SAVED: Aug  4 12:31:20 2007
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module bram_bufferx16_2inv ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(in), .Y(net6));

endmodule
// Library - leafcell, Cell - bram_hbuffer_1xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:50:36 2007
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module bram_hbuffer_1xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;
output [1:0]  bm_sdi_o;
output [1:0]  bm_banksel_o;
output [1:0]  bm_sdo_o;

input [1:0]  bm_sdo_i;
input [1:0]  bm_banksel_i;
input [1:0]  bm_sdi_i;
input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_icg, View - schematic
// LAST TIME SAVED: Jun 25 14:02:00 2007
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module bram_icg ( clkout, clk, en );
output  clkout;

input  clk, en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I193 ( .A(net027), .Y(net014), .B(c));
inv_tri_2_hvt I7 ( .Tb(cn), .T(c), .A(net027), .Y(net023));
inv_tri_2_hvt I5 ( .Tb(c), .T(cn), .A(en), .Y(net023));
inv_hvt I391 ( .A(net014), .Y(clkout));
inv_hvt I6 ( .A(net023), .Y(net027));
inv_hvt I4 ( .A(cn), .Y(c));
inv_hvt I3 ( .A(clk), .Y(cn));

endmodule
// Library - misc, Cell - ml_osc_logic, View - schematic
// LAST TIME SAVED: Aug 28 08:48:45 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_osc_logic ( sel_trim, clkin, smc_osc_fsel, smc_oscen );

input  clkin, smc_oscen;

output [3:0]  sel_trim;

input [1:0]  smc_osc_fsel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [1:2]  in_sel;



tiehi I280 ( .tiehi(net058));
ml_dff I174 ( .R(reset_ff), .D(net050), .CLK(clkin_buf_b), .QN(net150),
     .Q(net172));
ml_dff I238 ( .R(reset_ff), .D(net050), .CLK(clkin_buf), .QN(net154),
     .Q(net177));
ml_dff I244 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf),
     .QN(net155), .Q(net182));
ml_dff I245 ( .R(reset_ff), .D(smc_osc_fsel[1]), .CLK(clkin_buf_b),
     .QN(net153), .Q(net187));
ml_dff I242 ( .R(reset_ff), .D(net048), .CLK(clkin_buf_b), .QN(net191),
     .Q(net192));
ml_dff I243 ( .R(reset_ff), .D(net048), .CLK(clkin_buf), .QN(net152),
     .Q(net197));
ml_mux2_hvt I279 ( .in1(net182), .in0(net187), .out(sel_trim[0]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I277 ( .in1(net057), .in0(net061), .out(sel_trim[2]),
     .sel(clkin_buf_delay));
ml_mux2_hvt I278 ( .in1(net052), .in0(net054), .out(sel_trim[1]),
     .sel(clkin_buf_delay));
nor2_hvt I256 ( .A(smc_osc_fsel[1]), .B(smc_osc_fsel[0]),
     .Y(in_sel[2]));
inv_hvt I263 ( .A(clkin_buf), .Y(net065));
inv_hvt I252 ( .A(smc_oscen), .Y(reset_ff));
inv_hvt I264 ( .A(net065), .Y(net063));
inv_hvt I253 ( .A(clkin_buf_b), .Y(clkin_buf));
inv_hvt I254 ( .A(clkin), .Y(clkin_buf_b));
inv_hvt I255 ( .A(smc_osc_fsel[1]), .Y(in_sel[1]));
inv_hvt I266 ( .A(net063), .Y(net059));
inv_hvt I265 ( .A(net059), .Y(net0143));
inv_hvt I274 ( .A(net177), .Y(net057));
inv_hvt I273 ( .A(net172), .Y(net061));
inv_hvt I275 ( .A(net192), .Y(net054));
inv_hvt I276 ( .A(net197), .Y(net052));
inv_hvt I261 ( .A(in_sel[2]), .Y(net050));
inv_hvt I267 ( .A(net0143), .Y(net0144));
inv_hvt I262 ( .A(in_sel[1]), .Y(net048));
inv_hvt I268 ( .A(net0144), .Y(net0145));
inv_hvt I269 ( .A(net0142), .Y(clkin_buf_delay));
inv_hvt I270 ( .A(net0145), .Y(net0142));
inv_hvt I176 ( .A(net058), .Y(sel_trim[3]));

endmodule
// Library - leafcell, Cell - bram_hbuffer_dff_2xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:02:56 2007
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module bram_hbuffer_dff_2xbank ( bm_banksel_o, bm_init_o,
     bm_rcapmux_en_o, bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o,
     bm_sdo_o, bm_sreb_o, bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i,
     bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i,
     bm_sdi_i, bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclkrw_o, bm_sreb_o, bm_sweb_o,
     bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [3:0]  bm_sdi_o;
output [3:0]  bm_banksel_o;
output [1:0]  bm_sclk_o;
output [7:0]  bm_sa_o;
output [3:0]  bm_sdo_o;

input [7:0]  bm_sa_i;
input [3:0]  bm_sdo_i;
input [3:0]  bm_banksel_i;
input [3:0]  bm_sdi_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net102;

wire  [0:3]  net103;



tielo I23 ( .tielo(net057));
bram_icg I47 ( .en(net74), .clk(bm_sclk_i), .clkout(net61));
bram_icg I19 ( .en(net72), .clk(bm_sclk_i), .clkout(net64));
bram_bufferx16_2inv I16_3_ ( .in(net103[0]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I16_2_ ( .in(net103[1]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I16_1_ ( .in(net103[2]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I16_0_ ( .in(net103[3]), .out(bm_sdo_o[0]));
bram_bufferx4 I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx4 I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx4 I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx4 I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx4 I22 ( .in(net64), .out(bm_sclk_o[1]));
bram_bufferx4 I5 ( .in(bm_wdummymux_en_i), .out(bm_wdummymux_en_o));
bram_bufferx4 I13_3_ ( .in(bm_banksel_i[3]), .out(bm_banksel_o[3]));
bram_bufferx4 I13_2_ ( .in(bm_banksel_i[2]), .out(bm_banksel_o[2]));
bram_bufferx4 I13_1_ ( .in(bm_banksel_i[1]), .out(bm_banksel_o[1]));
bram_bufferx4 I13_0_ ( .in(bm_banksel_i[0]), .out(bm_banksel_o[0]));
bram_bufferx4 I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx4 I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx4 I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx4 I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx4 I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx4 I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx4 I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx4 I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx4 I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx4 I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx4 I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx4 I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx4 I18 ( .in(net61), .out(bm_sclk_o[0]));
bram_bufferx4 I11 ( .in(bm_sreb_i), .out(bm_sreb_o));
leafcell_ml_dff_schematic I48_3_ ( .R(net057), .D(bm_sdo_i[3]),
     .CLK(bm_sclk_i), .QN(net102[0]), .Q(net103[0]));
leafcell_ml_dff_schematic I48_2_ ( .R(net057), .D(bm_sdo_i[2]),
     .CLK(bm_sclk_i), .QN(net102[1]), .Q(net103[1]));
leafcell_ml_dff_schematic I48_1_ ( .R(net057), .D(bm_sdo_i[1]),
     .CLK(bm_sclk_i), .QN(net102[2]), .Q(net103[2]));
leafcell_ml_dff_schematic I48_0_ ( .R(net057), .D(bm_sdo_i[0]),
     .CLK(bm_sclk_i), .QN(net102[3]), .Q(net103[3]));
nor2_hvt I20 ( .A(bm_banksel_i[2]), .B(bm_banksel_i[3]), .Y(net67));
nor2_hvt I49 ( .A(bm_banksel_i[0]), .B(bm_banksel_i[1]), .Y(net70));
inv_hvt I21 ( .A(net67), .Y(net72));
inv_hvt I17 ( .A(net70), .Y(net74));

endmodule
// Library - leafcell, Cell - bram_hbuffer_2xbank, View - schematic
// LAST TIME SAVED: Aug  4 13:01:06 2007
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module bram_hbuffer_2xbank ( bm_banksel_o, bm_init_o, bm_rcapmux_en_o,
     bm_sa_o, bm_sclk_o, bm_sclkrw_o, bm_sdi_o, bm_sdo_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o, bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sdo_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i );
output  bm_init_o, bm_rcapmux_en_o, bm_sclk_o, bm_sclkrw_o, bm_sreb_o,
     bm_sweb_o, bm_wdummymux_en_o;

input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i;

output [7:0]  bm_sa_o;
output [3:0]  bm_sdi_o;
output [3:0]  bm_sdo_o;
output [3:0]  bm_banksel_o;

input [3:0]  bm_sdi_i;
input [3:0]  bm_banksel_i;
input [3:0]  bm_sdo_i;
input [7:0]  bm_sa_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



bram_bufferx16_2inv I6_3_ ( .in(bm_sdi_i[3]), .out(bm_sdi_o[3]));
bram_bufferx16_2inv I6_2_ ( .in(bm_sdi_i[2]), .out(bm_sdi_o[2]));
bram_bufferx16_2inv I6_1_ ( .in(bm_sdi_i[1]), .out(bm_sdi_o[1]));
bram_bufferx16_2inv I6_0_ ( .in(bm_sdi_i[0]), .out(bm_sdi_o[0]));
bram_bufferx16_2inv I5 ( .in(bm_wdummymux_en_i),
     .out(bm_wdummymux_en_o));
bram_bufferx16_2inv I2_3_ ( .in(bm_sdo_i[3]), .out(bm_sdo_o[3]));
bram_bufferx16_2inv I2_2_ ( .in(bm_sdo_i[2]), .out(bm_sdo_o[2]));
bram_bufferx16_2inv I2_1_ ( .in(bm_sdo_i[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I2_0_ ( .in(bm_sdo_i[0]), .out(bm_sdo_o[0]));
bram_bufferx16_2inv I13_3_ ( .in(bm_banksel_i[3]),
     .out(bm_banksel_o[3]));
bram_bufferx16_2inv I13_2_ ( .in(bm_banksel_i[2]),
     .out(bm_banksel_o[2]));
bram_bufferx16_2inv I13_1_ ( .in(bm_banksel_i[1]),
     .out(bm_banksel_o[1]));
bram_bufferx16_2inv I13_0_ ( .in(bm_banksel_i[0]),
     .out(bm_banksel_o[0]));
bram_bufferx16_2inv I12 ( .in(bm_sclk_i), .out(bm_sclk_o));
bram_bufferx16_2inv I9 ( .in(bm_sweb_i), .out(bm_sweb_o));
bram_bufferx16_2inv I0 ( .in(bm_sclkrw_i), .out(bm_sclkrw_o));
bram_bufferx16_2inv I7 ( .in(bm_rcapmux_en_i), .out(bm_rcapmux_en_o));
bram_bufferx16_2inv I8 ( .in(bm_init_i), .out(bm_init_o));
bram_bufferx16_2inv I10_7_ ( .in(bm_sa_i[7]), .out(bm_sa_o[7]));
bram_bufferx16_2inv I10_6_ ( .in(bm_sa_i[6]), .out(bm_sa_o[6]));
bram_bufferx16_2inv I10_5_ ( .in(bm_sa_i[5]), .out(bm_sa_o[5]));
bram_bufferx16_2inv I10_4_ ( .in(bm_sa_i[4]), .out(bm_sa_o[4]));
bram_bufferx16_2inv I10_3_ ( .in(bm_sa_i[3]), .out(bm_sa_o[3]));
bram_bufferx16_2inv I10_2_ ( .in(bm_sa_i[2]), .out(bm_sa_o[2]));
bram_bufferx16_2inv I10_1_ ( .in(bm_sa_i[1]), .out(bm_sa_o[1]));
bram_bufferx16_2inv I10_0_ ( .in(bm_sa_i[0]), .out(bm_sa_o[0]));
bram_bufferx16_2inv I11 ( .in(bm_sreb_i), .out(bm_sreb_o));

endmodule
// Library - leafcell, Cell - bram_bufferx2e, View - schematic
// LAST TIME SAVED: Jun 25 13:54:30 2007
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module bram_bufferx2e ( out, en, in );
output  out;

input  en, in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I391 ( .A(net7), .Y(out));
nand2_hvt I193 ( .A(en), .Y(net7), .B(in));

endmodule
// Library - leafcell, Cell - bram_bank_logic_bot, View - schematic
// LAST TIME SAVED: Aug 31 18:48:17 2007
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module bram_bank_logic_bot ( bm_sclkrw_o, bm_sdo_o, bm_sweb_o,
     bm_banksel_i, bm_sclk_i, bm_sclkrw_i, bm_sdo_i, bm_sweb_i );

input  bm_sclk_i, bm_sclkrw_i, bm_sweb_i;

output [1:0]  bm_sweb_o;
output [1:0]  bm_sdo_o;
output [1:0]  bm_sclkrw_o;

input [1:0]  bm_banksel_i;
input [1:0]  bm_sdo_i;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:1]  net25;

wire  [1:0]  net26;



bram_bufferx16_2inv I51_1_ ( .in(net26[1]), .out(bm_sdo_o[1]));
bram_bufferx16_2inv I51_0_ ( .in(net26[0]), .out(bm_sdo_o[0]));
leafcell_ml_dff_schematic I52_1_ ( .R(net020), .D(bm_sdo_i[1]),
     .CLK(bm_sclk_i), .QN(net25[0]), .Q(net26[1]));
leafcell_ml_dff_schematic I52_0_ ( .R(net020), .D(bm_sdo_i[0]),
     .CLK(bm_sclk_i), .QN(net25[1]), .Q(net26[0]));
bram_bufferx2e I54_1_ ( .in(bm_sweb_i), .en(bm_banksel_i[1]),
     .out(bm_sweb_o[1]));
bram_bufferx2e I54_0_ ( .in(bm_sweb_i), .en(bm_banksel_i[0]),
     .out(bm_sweb_o[0]));
bram_bufferx2e I48_1_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[1]),
     .out(bm_sclkrw_o[1]));
bram_bufferx2e I48_0_ ( .in(bm_sclkrw_i), .en(bm_banksel_i[0]),
     .out(bm_sclkrw_o[0]));
tielo I55 ( .tielo(net020));

endmodule
// Library - leafcell, Cell - quad_x4_ice8, View - schematic
// LAST TIME SAVED: Oct 16 14:41:17 2008
// NETLIST TIME: Nov 14 16:17:20 2008
`timescale 1ns / 1ns 

module quad_x4_ice8 ( bm_sdo_o, cf_b, cf_l, cf_r, cf_t,
     fabric_out_32_00, fabric_out_33_01, fabric_out_33_02, padeb_b,
     padeb_l, padeb_r, padeb_t, pado_b, pado_l, pado_r, pado_t,
     sdo_pad, spi_ss_in_b, spi_ss_in_l, spi_ss_in_r, bl_bot, bl_top,
     bm_banksel_i, bm_init_i, bm_rcapmux_en_i, bm_sa_i, bm_sclk_i,
     bm_sclkrw_i, bm_sdi_i, bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i,
     bs_en, ceb, end_of_startup_bot_r, end_of_startup_l,
     end_of_startup_r, end_of_startup_top, hiz_b, mode, padin_b,
     padin_l, padin_r, padin_t, pgate_l, pgate_r, prog, purst, r,
     reset_b_l, reset_b_r, sdi_pad, shift, spieb_b, spioeb_l, spiout_b,
     spiout_l, spiout_r, tclk, tiegnd, tievdd, update, vdd_cntl_l,
     vdd_cntl_r, wl_l, wl_r );
output  fabric_out_32_00, fabric_out_33_01, fabric_out_33_02, sdo_pad;


input  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en, ceb, hiz_b, mode, prog,
     purst, r, sdi_pad, shift, tclk, tiegnd, tievdd, update;

output [3:0]  bm_sdo_o;
output [767:0]  cf_r;
output [767:0]  cf_b;
output [63:0]  spi_ss_in_r;
output [767:0]  cf_t;
output [59:0]  padeb_t;
output [56:0]  padeb_b;
output [49:0]  pado_l;
output [63:32]  spi_ss_in_b;
output [59:0]  pado_t;
output [54:0]  pado_r;
output [54:0]  padeb_r;
output [49:0]  padeb_l;
output [31:0]  spi_ss_in_l;
output [56:0]  pado_b;
output [767:0]  cf_l;

inout [1743:0]  bl_bot;
inout [1743:0]  bl_top;

input [31:0]  spiout_r;
input [3:0]  bm_banksel_i;
input [3:0]  bm_sdi_i;
input [31:0]  spiout_l;
input [59:0]  padin_t;
input [543:0]  reset_b_l;
input [56:0]  padin_b;
input [543:0]  pgate_r;
input [543:0]  wl_l;
input [31:16]  end_of_startup_bot_r;
input [7:0]  bm_sa_i;
input [54:0]  padin_r;
input [31:0]  end_of_startup_l;
input [543:0]  wl_r;
input [63:32]  spiout_b;
input [49:0]  padin_l;
input [543:0]  pgate_l;
input [31:0]  end_of_startup_top;
input [543:0]  vdd_cntl_r;
input [543:0]  vdd_cntl_l;
input [63:32]  spieb_b;
input [31:0]  spioeb_l;
input [543:0]  reset_b_r;
input [31:0]  end_of_startup_r;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:23]  net1207;

wire  [0:7]  net1647;

wire  [0:23]  net1202;

wire  [0:23]  net1203;

wire  [0:7]  net1105;

wire  [0:47]  net2038;

wire  [0:7]  net1589;

wire  [0:47]  net01772;

wire  [0:23]  net1600;

wire  [0:7]  net1648;

wire  [0:7]  net1652;

wire  [0:47]  net2071;

wire  [0:7]  net1897;

wire  [0:23]  net1606;

wire  [0:7]  net1108;

wire  [0:47]  net1233;

wire  [0:23]  net2010;

wire  [0:23]  net2001;

wire  [0:3]  net1835;

wire  [0:47]  net2033;

wire  [0:7]  net1941;

wire  [0:7]  net1462;

wire  [0:7]  net1946;

wire  [0:7]  net1656;

wire  [0:23]  net2021;

wire  [0:7]  net1162;

wire  [0:7]  net1942;

wire  [0:7]  net1868;

wire  [0:47]  net1634;

wire  [0:47]  net01767;

wire  [0:7]  net1161;

wire  [0:7]  net1156;

wire  [0:47]  net01760;

wire  [0:7]  net1587;

wire  [0:47]  net01764;

wire  [0:47]  net01769;

wire  [0:47]  net01763;

wire  [0:47]  net01762;

wire  [3:0]  slf_op_00_16;

wire  [7:0]  n_slf_op_01_17;

wire  [7:0]  bm_sa_b1_o;

wire  [0:47]  net1236;

wire  [7:0]  n_slf_op_16_23;

wire  [1:0]  bm_sdi_b0_o;

wire  [1:0]  bm_sclkrw_b0_o;

wire  [1:0]  bm_sweb_b2_o;

wire  [0:7]  net1909;

wire  [0:23]  net1199;

wire  [3:0]  bm_bank30_banksel_o;

wire  [1:0]  bm_sweb_b0_o;

wire  [7:0]  n_slf_op_16_17;

wire  [1:0]  bm_sclkrw_b2_o;

wire  [3:0]  bm_bank30_sdi_o;

wire  [1:0]  bm_bank10_banksel_o;

wire  [3:0]  bm_bank30_sdo_i;

wire  [0:23]  net2014;

wire  [1:0]  bm_sdi_b2_o;

wire  [1:0]  bm_bank30_sclk_o;

wire  [0:7]  net1958;

wire  [0:7]  net1586;

wire  [0:47]  net2076;

wire  [0:7]  net1860;

wire  [0:47]  net2032;

wire  [0:47]  net2066;

wire  [0:15]  net1243;

wire  [0:7]  net1107;

wire  [0:47]  net2061;

wire  [0:47]  net1237;

wire  [0:47]  net1241;

wire  [0:47]  net2037;

wire  [0:7]  net1098;

wire  [0:47]  net2055;

wire  [0:7]  net1899;

wire  [0:47]  net01765;

wire  [0:7]  net1904;

wire  [0:47]  net1632;

wire  [0:7]  net1110;

wire  [0:23]  net2020;

wire  [0:7]  net1152;

wire  [0:23]  net2015;

wire  [7:0]  glb_net;

wire  [0:7]  net1901;

wire  [0:23]  net1613;

wire  [0:7]  net1654;

wire  [0:47]  net1640;

wire  [0:47]  net2053;

wire  [0:47]  net01770;

wire  [0:7]  net1106;

wire  [0:23]  net2004;

wire  [0:1]  net1925;

wire  [0:7]  net1936;

wire  [0:7]  net1952;

wire  [0:7]  net1943;

wire  [0:23]  net1205;

wire  [0:47]  net2048;

wire  [0:7]  net1956;

wire  [0:3]  net1777;

wire  [0:47]  net2046;

wire  [0:7]  net1944;

wire  [0:7]  net1104;

wire  [0:23]  net1608;

wire  [0:47]  net1644;

wire  [0:47]  net1238;

wire  [0:7]  net1594;

wire  [0:7]  net1959;

wire  [0:23]  net2023;

wire  [0:47]  net01771;

wire  [0:47]  net2069;

wire  [0:47]  net1239;

wire  [0:47]  net1228;

wire  [0:23]  net1200;

wire  [0:47]  net2064;

wire  [0:7]  net1163;

wire  [0:23]  net1198;

wire  [0:23]  net2030;

wire  [0:47]  net1756;

wire  [0:7]  net1903;

wire  [0:7]  net1588;

wire  [0:7]  net1649;

wire  [0:47]  net2042;

wire  [0:23]  net2007;

wire  [0:23]  net2026;

wire  [0:47]  net2056;

wire  [0:23]  net2013;

wire  [0:7]  net1955;

wire  [0:47]  net2045;

wire  [0:7]  net1962;

wire  [0:7]  net1593;

wire  [0:1]  net1293;

wire  [0:7]  net1898;

wire  [0:3]  net1920;

wire  [0:7]  net2083;

wire  [0:47]  net01774;

wire  [0:1]  net936;

wire  [0:7]  net1657;

wire  [0:47]  net1639;

wire  [0:7]  net1907;

wire  [0:7]  net1099;

wire  [0:47]  net1232;

wire  [0:7]  net1164;

wire  [0:7]  net1940;

wire  [0:7]  net1650;

wire  [0:23]  net1603;

wire  [0:23]  net2025;

wire  [0:7]  net1859;

wire  [0:23]  net2024;

wire  [0:47]  net2078;

wire  [0:7]  net1775;

wire  [0:23]  net2005;

wire  [0:47]  net2052;

wire  [0:47]  net1642;

wire  [0:47]  net1231;

wire  [0:23]  net2012;

wire  [0:7]  net1951;

wire  [0:47]  net1229;

wire  [0:47]  net2058;

wire  [0:47]  net2039;

wire  [0:47]  net1645;

wire  [0:47]  net1636;

wire  [0:7]  net1865;

wire  [0:3]  net1038;

wire  [0:47]  net2065;

wire  [0:47]  net2041;

wire  [0:47]  net01761;

wire  [0:7]  net1900;

wire  [0:47]  net2074;

wire  [0:7]  net1103;

wire  [0:7]  net1934;

wire  [0:47]  net1242;

wire  [0:47]  net2073;

wire  [0:7]  net1871;

wire  [0:7]  net1933;

wire  [0:1]  net935;

wire  [0:23]  net1999;

wire  [0:7]  net1896;

wire  [0:47]  net2040;

wire  [0:23]  net1605;

wire  [0:47]  net01773;

wire  [0:47]  net1599;

wire  [0:47]  net1637;

wire  [0:7]  net1662;

wire  [0:7]  net1862;

wire  [0:3]  net975;

wire  [0:47]  net2034;

wire  [0:47]  net2050;

wire  [0:47]  net2060;

wire  [0:47]  net2044;

wire  [0:7]  net1591;

wire  [0:7]  net1872;

wire  [0:47]  net2067;

wire  [0:7]  net1863;

wire  [0:7]  net1935;

wire  [0:7]  net1100;

wire  [0:23]  net1211;

wire  [0:23]  net2027;

wire  [0:1]  net1990;

wire  [0:7]  net1905;

wire  [0:23]  net1601;

wire  [0:47]  net2062;

wire  [0:47]  net1641;

wire  [0:7]  net1213;

wire  [0:7]  net1101;

wire  [0:47]  net2077;

wire  [0:47]  net2068;

wire  [0:23]  net1206;

wire  [0:47]  net1633;

wire  [0:7]  net1954;

wire  [0:7]  net1755;

wire  [0:7]  net1160;

wire  [0:47]  net1128;

wire  [0:7]  net1908;

wire  [0:7]  net1658;

wire  [0:47]  net1635;

wire  [0:47]  net2075;

wire  [0:7]  net1158;

wire  [0:7]  net1928;

wire  [0:47]  net2035;

wire  [0:7]  net1102;

wire  [0:7]  net1938;

wire  [0:7]  net1653;

wire  [0:7]  net1157;

wire  [0:7]  net1659;

wire  [0:47]  net1234;

wire  [0:47]  net1235;

wire  [0:23]  net1168;

wire  [0:7]  net1861;

wire  [0:7]  net1592;

wire  [0:23]  net1609;

wire  [0:7]  net1660;

wire  [0:23]  net2022;

wire  [3:0]  slf_op_33_16;

wire  [0:7]  net1651;

wire  [0:23]  net1612;

wire  [0:23]  net1208;

wire  [0:47]  net2051;

wire  [0:47]  net2070;

wire  [0:7]  net1945;

wire  [0:23]  net1204;

wire  [0:7]  net920;

wire  [0:7]  net942;

wire  [0:7]  net1159;

wire  [0:47]  net2059;

wire  [0:7]  net1961;

wire  [0:7]  net1949;

wire  [0:7]  net1902;

wire  [0:23]  net2003;

wire  [0:23]  net2017;

wire  [0:7]  net1244;

wire  [0:47]  net1638;

wire  [0:1]  net1926;

wire  [0:23]  net1210;

wire  [0:7]  net1153;

wire  [0:47]  net2079;

wire  [0:7]  net1994;

wire  [3:0]  slf_op_00_17;

wire  [0:23]  net2009;

wire  [0:23]  net1607;

wire  [0:7]  net1939;

wire  [0:1]  net1310;

wire  [0:7]  net1271;

wire  [0:23]  net2028;

wire  [0:15]  net2047;

wire  [0:7]  net1597;

wire  [0:7]  net1109;

wire  [0:47]  net2031;

wire  [0:15]  net1577;

wire  [0:47]  net2043;

wire  [0:23]  net2018;

wire  [3:0]  slf_op_33_17;

wire  [0:3]  net974;

wire  [0:47]  net2036;

wire  [0:47]  net1643;

wire  [0:23]  net1602;

wire  [0:47]  net2057;

wire  [0:47]  net2049;

wire  [0:7]  net1585;

wire  [0:7]  net1596;

wire  [0:1]  net1290;

wire  [0:7]  net1950;

wire  [0:23]  net1610;

wire  [0:7]  net1864;

wire  [0:47]  net2054;

wire  [0:7]  net1262;

wire  [0:23]  net2002;

wire  [0:7]  net1576;

wire  [0:7]  net1646;

wire  [0:47]  net01768;

wire  [0:7]  net1590;

wire  [0:7]  net1937;

wire  [0:23]  net2000;

wire  [0:7]  net1165;

wire  [0:23]  net1212;

wire  [0:7]  net1314;

wire  [0:23]  net1201;

wire  [0:7]  net962;

wire  [0:7]  net1155;

wire  [0:47]  net2063;

wire  [0:1]  net918;

wire  [0:7]  net1953;

wire  [0:7]  net1275;

wire  [0:7]  net1869;

wire  [0:47]  net2072;

wire  [0:23]  net1209;

wire  [0:7]  net1957;

wire  [0:23]  net1614;

wire  [0:7]  net1906;

wire  [0:7]  net1867;

wire  [0:23]  net2011;

wire  [0:7]  net1960;

wire  [0:1]  net1007;

wire  [0:23]  net2029;

wire  [0:47]  net1230;

wire  [0:7]  net1948;

wire  [0:7]  net1870;

wire  [0:7]  net1947;

wire  [0:23]  net1615;

wire  [0:47]  net01766;

wire  [0:1]  net1922;

wire  [0:7]  net1595;

wire  [0:23]  net2019;

wire  [0:7]  net1866;

wire  [0:23]  net1604;

wire  [0:23]  net2008;

wire  [0:3]  net979;

wire  [0:15]  net1837;

wire  [0:23]  net2006;

wire  [0:23]  net2016;

wire  [0:47]  net1240;

wire  [0:23]  net1611;



clk_mux2to1x48k I_glb_ck_tree_bot ( .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[271:270]), .bl(bl_bot[873:870]),
     .min3({padin_193, fabric_out_33_16}), .min2({padin_80,
     fabric_out_00_16}), .min1({padin_27, fabric_out_17_33}),
     .min0({padin_135, fabric_out_17_00}), .wl_l(wl_l[271:270]),
     .reset_l(reset_b_l[271:270]), .pgate_l(pgate_l[271:270]),
     .gnet({glb_net[7], glb_net[6], glb_net[1], glb_net[0]}),
     .pgate_r(pgate_r[271:270]), .wl_r(wl_r[271:270]),
     .reset_r(reset_b_r[271:270]), .vdd_cntl_r(vdd_cntl_r[271:270]));
clk_mux2to1x48k I_glb_ck_tree_top ( .prog(prog),
     .vdd_cntl_l(vdd_cntl_l[273:272]), .bl(bl_top[873:870]),
     .min3({padin_136, fabric_out_16_00}), .min2({padin_26,
     fabric_out_16_33}), .min1({padin_81, fabric_out_00_17}),
     .min0({padin_192, fabric_out_33_17}), .wl_l(wl_l[273:272]),
     .reset_l(reset_b_l[273:272]), .pgate_l(pgate_l[273:272]),
     .gnet(glb_net[5:2]), .pgate_r(pgate_r[273:272]),
     .wl_r(wl_r[273:272]), .reset_r(reset_b_r[273:272]),
     .vdd_cntl_r(vdd_cntl_r[273:272]));
cram_row270col4 I_mem270bot ( .bl(bl_bot[873:870]),
     .pgate_l(pgate_l[269:0]), .pgate_r(pgate_r[269:0]),
     .reset_l(reset_b_l[269:0]), .reset_r(reset_b_r[269:0]),
     .vdd_cntl_l(vdd_cntl_l[269:0]), .vdd_cntl_r(vdd_cntl_r[269:0]),
     .wl_l(wl_l[269:0]), .wl_r(wl_r[269:0]));
cram_row270col4 I_mem270top ( .bl(bl_top[873:870]),
     .pgate_l(pgate_l[543:274]), .pgate_r(pgate_r[543:274]),
     .reset_l(reset_b_l[543:274]), .reset_r(reset_b_r[543:274]),
     .vdd_cntl_l(vdd_cntl_l[543:274]),
     .vdd_cntl_r(vdd_cntl_r[543:274]), .wl_l(wl_l[543:274]),
     .wl_r(wl_r[543:274]));
quad_bl_ice8 I_quad_bl_ice8 ( .tnr_op_00_16(n_slf_op_01_17[7:0]),
     .ceb_i(net0901), .ceb_o(net0902), .padin_80(padin_80),
     .padin_b(padin_b[29:0]), .padeb_b(padeb_b[29:0]),
     .pado_b(pado_b[29:0]), .fabric_out_00_15(hold_lbank),
     .pado_l(pado_l[23:0]), .padin_l(padin_l[23:0]),
     .padeb_l(padeb_l[23:0]), .fabric_out_00_16(fabric_out_00_16),
     .fabric_out_16_00(fabric_out_16_00), .padin_27(padin_27),
     .slf_op_16_00(net1835[0:3]), .slf_op_00_16(slf_op_00_16[3:0]),
     .sp4_h_r_16_00(net1837[0:15]), .spi_ss_in_l(spi_ss_in_l[31:0]),
     .spioeb_l(spioeb_l[31:0]), .spiout_l(spiout_l[31:0]),
     .update_i(net1841), .top_op_16_16(n_slf_op_16_17[7:0]),
     .top_op_15_16(net1859[0:7]), .top_op_14_16(net1860[0:7]),
     .top_op_13_16(net1861[0:7]), .top_op_12_16(net1862[0:7]),
     .top_op_11_16(net1863[0:7]), .top_op_10_16(net1864[0:7]),
     .top_op_09_16(net1865[0:7]), .top_op_08_16(net1866[0:7]),
     .top_op_07_16(net1867[0:7]), .top_op_06_16(net1868[0:7]),
     .top_op_05_16(net1869[0:7]), .top_op_04_16(net1870[0:7]),
     .top_op_03_16(net1871[0:7]), .top_op_02_16(net1872[0:7]),
     .top_op_01_16(n_slf_op_01_17[7:0]),
     .tnr_op_15_16(n_slf_op_16_17[7:0]), .tnr_op_14_16(net1859[0:7]),
     .tnr_op_13_16(net1860[0:7]), .tnr_op_12_16(net1861[0:7]),
     .tnr_op_11_16(net1862[0:7]), .tnr_op_10_16(net1863[0:7]),
     .tnr_op_09_16(net1864[0:7]), .tnr_op_08_16(net1865[0:7]),
     .tnr_op_07_16(net1866[0:7]), .tnr_op_06_16(net1867[0:7]),
     .tnr_op_05_16(net1868[0:7]), .tnr_op_04_16(net1869[0:7]),
     .tnr_op_03_16(net1870[0:7]), .tnr_op_02_16(net1871[0:7]),
     .tnr_op_01_16(net1872[0:7]), .tnl_op_16_16(net1859[0:7]),
     .tnl_op_15_16(net1860[0:7]), .tnl_op_14_16(net1861[0:7]),
     .tnl_op_13_16(net1862[0:7]), .tnl_op_12_16(net1863[0:7]),
     .tnl_op_11_16(net1864[0:7]), .tnl_op_10_16(net1865[0:7]),
     .tnl_op_09_16(net1866[0:7]), .tnl_op_08_16(net1867[0:7]),
     .tnl_op_07_16(net1868[0:7]), .tnl_op_06_16(net1869[0:7]),
     .tnl_op_05_16(net1870[0:7]), .tnl_op_04_16(net1871[0:7]),
     .tnl_op_03_16(net1872[0:7]), .tnl_op_02_16(n_slf_op_01_17[7:0]),
     .tnl_op_01_16({slf_op_00_17[3], slf_op_00_17[2], slf_op_00_17[1],
     slf_op_00_17[0], slf_op_00_17[3], slf_op_00_17[2],
     slf_op_00_17[1], slf_op_00_17[0]}), .tievdd(tievdd),
     .tiegnd(tiegnd), .tclk_i(net1892), .shift_i(net1893),
     .sdi(net1894), .rgt_op_16_16(net1775[0:7]),
     .rgt_op_16_14(net1896[0:7]), .rgt_op_16_13(net1897[0:7]),
     .rgt_op_16_12(net1898[0:7]), .rgt_op_16_11(net1899[0:7]),
     .rgt_op_16_10(net1900[0:7]), .rgt_op_16_09(net1901[0:7]),
     .rgt_op_16_08(net1902[0:7]), .rgt_op_16_07(net1903[0:7]),
     .rgt_op_16_06(net1904[0:7]), .rgt_op_16_05(net1905[0:7]),
     .rgt_op_16_04(net1906[0:7]), .rgt_op_16_03(net1907[0:7]),
     .rgt_op_16_02(net1908[0:7]), .rgt_op_16_01(net1909[0:7]),
     .r_i(net1910), .purst(purst), .prog(prog), .mode_i(net1913),
     .hold_l_b(hold_lbank), .hold_b_l(hold_bbank), .hiz_b_i(net1916),
     .glb_in(glb_net[7:0]),
     .end_of_startup_lft_b(end_of_startup_l[15:0]), .bs_en_i(net1919),
     .bnr_op_16_01(net1920[0:3]), .bm_wdummymux_en_i(net1921),
     .bm_sweb_i(net1922[0:1]), .bm_sreb_i(net1923),
     .bm_sdo_i({bm_sdo_b1_o, bm_sdi_b0_o[0]}), .bm_sdi_i(net1925[0:1]),
     .bm_sclkrw_i(net1926[0:1]), .bm_sclk_i(net1927),
     .bm_sa_i(net1928[0:7]), .bm_rcapmux_en_i(net1929),
     .bm_init_i(net1930), .update_o(net1931), .tclk_o(net1932),
     .slf_op_16_16(net1933[0:7]), .slf_op_16_15(net1934[0:7]),
     .slf_op_16_14(net1935[0:7]), .slf_op_16_13(net1936[0:7]),
     .slf_op_16_12(net1937[0:7]), .slf_op_16_11(net1938[0:7]),
     .slf_op_16_10(net1939[0:7]), .slf_op_16_09(net1940[0:7]),
     .slf_op_16_08(net1941[0:7]), .slf_op_16_07(net1942[0:7]),
     .slf_op_16_06(net1943[0:7]), .slf_op_16_05(net1944[0:7]),
     .slf_op_16_04(net1945[0:7]), .slf_op_16_03(net1946[0:7]),
     .slf_op_16_02(net1947[0:7]), .slf_op_16_01(net1948[0:7]),
     .slf_op_15_16(net1949[0:7]), .slf_op_14_16(net1950[0:7]),
     .slf_op_13_16(net1951[0:7]), .slf_op_12_16(net1952[0:7]),
     .slf_op_11_16(net1953[0:7]), .slf_op_10_16(net1954[0:7]),
     .slf_op_09_16(net1955[0:7]), .slf_op_08_16(net1956[0:7]),
     .slf_op_07_16(net1957[0:7]), .slf_op_06_16(net1958[0:7]),
     .slf_op_05_16(net1959[0:7]), .slf_op_04_16(net1960[0:7]),
     .slf_op_03_16(net1961[0:7]), .slf_op_02_16(net1962[0:7]),
     .slf_op_01_16(net1576[0:7]), .shift_o(net1964), .sdo(net1965),
     .r_o(net1966), .mode_o(net1967), .hiz_b_o(net1968),
     .cf_l(cf_l[383:0]), .cf_b(cf_b[383:0]), .carry_out_16_16(net1971),
     .carry_out_15_16(net1972), .carry_out_14_16(net1973),
     .carry_out_13_16(net1974), .carry_out_12_16(net1975),
     .carry_out_11_16(net1976), .carry_out_10_16(net1977),
     .carry_out_09_16(net1978), .carry_out_07_16(net1979),
     .carry_out_06_16(net1980), .carry_out_05_16(net1981),
     .carry_out_04_16(net1982), .carry_out_03_16(net1983),
     .carry_out_02_16(net1984), .carry_out_01_16(net1985),
     .bs_en_o(net1986), .bm_wdummymux_en_o(net1987),
     .bm_sweb_o(bm_sweb_b0_o[1:0]), .bm_sreb_o(net1989),
     .bm_sdo_o(net1990[0:1]), .bm_sdi_o(bm_sdi_b0_o[1:0]),
     .bm_sclkrw_o(bm_sclkrw_b0_o[1:0]), .bm_sclk_o(net1993),
     .bm_sa_o(net1994[0:7]), .bm_rcapmux_en_o(net1995),
     .bm_init_o(net1996), .wl_l(wl_l[271:0]),
     .vdd_cntl_l(vdd_cntl_l[271:0]), .sp12_v_t_16_16(net1999[0:23]),
     .sp12_v_t_15_16(net2000[0:23]), .sp12_v_t_14_16(net2001[0:23]),
     .sp12_v_t_13_16(net2002[0:23]), .sp12_v_t_12_16(net2003[0:23]),
     .sp12_v_t_11_16(net2004[0:23]), .sp12_v_t_10_16(net2005[0:23]),
     .sp12_v_t_09_16(net2006[0:23]), .sp12_v_t_08_16(net2007[0:23]),
     .sp12_v_t_07_16(net2008[0:23]), .sp12_v_t_06_16(net2009[0:23]),
     .sp12_v_t_05_16(net2010[0:23]), .sp12_v_t_04_16(net2011[0:23]),
     .sp12_v_t_03_16(net2012[0:23]), .sp12_v_t_02_16(net2013[0:23]),
     .sp12_v_t_01_16(net2014[0:23]), .sp12_h_r_16_16(net2015[0:23]),
     .sp12_h_r_16_15(net2016[0:23]), .sp12_h_r_16_14(net2017[0:23]),
     .sp12_h_r_16_13(net2018[0:23]), .sp12_h_r_16_12(net2019[0:23]),
     .sp12_h_r_16_11(net2020[0:23]), .sp12_h_r_16_10(net2021[0:23]),
     .sp12_h_r_16_09(net2022[0:23]), .sp12_h_r_16_08(net2023[0:23]),
     .sp12_h_r_16_07(net2024[0:23]), .sp12_h_r_16_06(net2025[0:23]),
     .sp12_h_r_16_05(net2026[0:23]), .sp12_h_r_16_04(net2027[0:23]),
     .sp12_h_r_16_03(net2028[0:23]), .sp12_h_r_16_02(net2029[0:23]),
     .sp12_h_r_16_01(net2030[0:23]), .sp4_v_t_16_16(net2046[0:47]),
     .sp4_v_t_15_16(net2045[0:47]), .sp4_v_t_14_16(net2044[0:47]),
     .sp4_v_t_13_16(net2043[0:47]), .sp4_v_t_12_16(net2042[0:47]),
     .sp4_v_t_11_16(net2041[0:47]), .sp4_v_t_10_16(net2040[0:47]),
     .sp4_v_t_09_16(net2039[0:47]), .sp4_v_t_08_16(net2038[0:47]),
     .sp4_v_t_07_16(net2037[0:47]), .sp4_v_t_06_16(net2036[0:47]),
     .sp4_v_t_05_16(net2035[0:47]), .sp4_v_t_04_16(net2034[0:47]),
     .sp4_v_t_03_16(net2033[0:47]), .sp4_v_t_02_16(net2032[0:47]),
     .sp4_v_t_01_16(net2031[0:47]), .sp4_v_t_00_16(net2047[0:15]),
     .sp4_r_v_b_16_16(net2048[0:47]), .sp4_r_v_b_16_15(net2049[0:47]),
     .sp4_r_v_b_16_14(net2050[0:47]), .sp4_r_v_b_16_13(net2051[0:47]),
     .sp4_r_v_b_16_12(net2052[0:47]), .sp4_r_v_b_16_11(net2053[0:47]),
     .sp4_r_v_b_16_10(net2054[0:47]), .sp4_r_v_b_16_09(net2055[0:47]),
     .sp4_r_v_b_16_08(net2056[0:47]), .sp4_r_v_b_16_07(net2057[0:47]),
     .sp4_r_v_b_16_06(net2058[0:47]), .sp4_r_v_b_16_05(net2059[0:47]),
     .sp4_r_v_b_16_04(net2060[0:47]), .sp4_r_v_b_16_03(net2061[0:47]),
     .sp4_r_v_b_16_02(net2062[0:47]), .sp4_r_v_b_16_01(net2063[0:47]),
     .sp4_h_r_16_16(net2064[0:47]), .sp4_h_r_16_15(net2065[0:47]),
     .sp4_h_r_16_14(net2066[0:47]), .sp4_h_r_16_13(net2067[0:47]),
     .sp4_h_r_16_12(net2068[0:47]), .sp4_h_r_16_11(net2069[0:47]),
     .sp4_h_r_16_10(net2070[0:47]), .sp4_h_r_16_09(net2071[0:47]),
     .sp4_h_r_16_08(net2072[0:47]), .sp4_h_r_16_07(net2073[0:47]),
     .sp4_h_r_16_06(net2074[0:47]), .sp4_h_r_16_05(net2075[0:47]),
     .sp4_h_r_16_04(net2076[0:47]), .sp4_h_r_16_03(net2077[0:47]),
     .sp4_h_r_16_02(net2078[0:47]), .sp4_h_r_16_01(net2079[0:47]),
     .reset_l(reset_b_l[271:0]), .pgate_l(pgate_l[271:0]),
     .bl(bl_bot[869:0]), .rgt_op_16_15(net2083[0:7]),
     .tnr_op_16_16(net1244[0:7]));
quad_br_ice8 I_quad_br_ice8 ( .ceb_o(net01437), .ceb_mi(ceb),
     .ceb_i(net0902),
     .end_of_startup_bot_r(end_of_startup_bot_r[31:16]),
     .end_of_startup_rgt_b(end_of_startup_r[15:0]),
     .spiout_b(spiout_b[63:32]), .spioeb_b(spieb_b[63:32]),
     .spi_ss_in_b(spi_ss_in_b[63:32]), .padin_81(padin_81),
     .fabric_out_18_00(hold_bbank), .padin_b(padin_b[56:30]),
     .padeb_b(padeb_b[56:30]), .pado_b(pado_b[56:30]),
     .pado_r(pado_r[27:0]), .padin_r(padin_r[27:0]),
     .padeb_r(padeb_r[27:0]), .fabric_out_33_16(fabric_out_33_16),
     .fabric_out_33_01(fabric_out_33_01),
     .fabric_out_33_02(fabric_out_33_02),
     .fabric_out_32_00(fabric_out_32_00),
     .fabric_out_17_00(fabric_out_17_00), .padin_135(padin_135),
     .bm_sdo_i({bm_sdo_b3_o, bm_sdi_b2_o[0]}),
     .slf_op_17_00(net1920[0:3]), .slf_op_33_16(slf_op_33_16[3:0]),
     .spi_ss_in_r(spi_ss_in_r[31:0]), .spiout_r(spiout_r[31:0]),
     .spioeb_r({tievdd, tievdd, tievdd, tievdd, tiegnd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd}), .sp4_v_b_17_16(net2048[0:47]),
     .sp4_v_b_17_15(net2049[0:47]), .sp4_v_b_17_14(net2050[0:47]),
     .sp4_v_b_17_13(net2051[0:47]), .sp4_v_b_17_12(net2052[0:47]),
     .sp4_v_b_17_11(net2053[0:47]), .sp4_v_b_17_10(net2054[0:47]),
     .sp4_v_b_17_09(net2055[0:47]), .sp4_v_b_17_08(net2056[0:47]),
     .sp4_v_b_17_07(net2057[0:47]), .sp4_v_b_17_06(net2058[0:47]),
     .sp4_v_b_17_05(net2059[0:47]), .sp4_v_b_17_04(net2060[0:47]),
     .sp4_v_b_17_03(net2061[0:47]), .sp4_v_b_17_02(net2062[0:47]),
     .sp4_v_b_17_01(net2063[0:47]), .mode_mi(mode),
     .carry_out_17_16(net1082), .top_op_32_16(net1110[0:7]),
     .top_op_31_16(net1109[0:7]), .top_op_30_16(net1108[0:7]),
     .top_op_29_16(net1107[0:7]), .top_op_28_16(net1106[0:7]),
     .top_op_27_16(net1105[0:7]), .top_op_26_16(net1104[0:7]),
     .top_op_25_16(net1103[0:7]), .top_op_24_16(net1102[0:7]),
     .top_op_23_16(net1101[0:7]), .top_op_22_16(net1100[0:7]),
     .top_op_21_16(net1099[0:7]), .top_op_20_16(net1098[0:7]),
     .top_op_19_16(net1275[0:7]), .top_op_18_16(net1213[0:7]),
     .tnr_op_19_16(net1098[0:7]), .tnr_op_20_16(net1099[0:7]),
     .tnr_op_21_16(net1100[0:7]), .tnr_op_22_16(net1101[0:7]),
     .tnr_op_23_16(net1102[0:7]), .tnr_op_24_16(net1103[0:7]),
     .tnr_op_25_16(net1104[0:7]), .tnr_op_26_16(net1105[0:7]),
     .tnr_op_27_16(net1106[0:7]), .tnr_op_28_16(net1107[0:7]),
     .tnr_op_29_16(net1108[0:7]), .tnr_op_30_16(net1109[0:7]),
     .tnr_op_31_16(net1110[0:7]), .tnr_op_32_16({slf_op_33_17[3],
     slf_op_33_17[2], slf_op_33_17[1], slf_op_33_17[0],
     slf_op_33_17[3], slf_op_33_17[2], slf_op_33_17[1],
     slf_op_33_17[0]}), .tnl_op_18_16(net1244[0:7]),
     .tnl_op_19_16(net1213[0:7]), .tnl_op_20_16(net1275[0:7]),
     .tnl_op_21_16(net1098[0:7]), .tnl_op_22_16(net1099[0:7]),
     .tnl_op_23_16(net1100[0:7]), .tnl_op_24_16(net1101[0:7]),
     .tnl_op_25_16(net1102[0:7]), .tnl_op_26_16(net1103[0:7]),
     .tnl_op_27_16(net1104[0:7]), .tnl_op_28_16(net1105[0:7]),
     .tnl_op_29_16(net1106[0:7]), .tnl_op_30_16(net1107[0:7]),
     .tnl_op_31_16(net1108[0:7]), .tnl_op_32_16(net1109[0:7]),
     .tnl_op_33_16(net1110[0:7]), .sp4_v_t_17_16(net1128[0:47]),
     .hold_r_b(hold_rbank), .lft_op_17_13(net1936[0:7]),
     .lft_op_17_14(net1935[0:7]), .lft_op_17_11(net1938[0:7]),
     .lft_op_17_10(net1939[0:7]), .lft_op_17_08(net1941[0:7]),
     .lft_op_17_04(net1945[0:7]), .lft_op_17_09(net1940[0:7]),
     .lft_op_17_07(net1942[0:7]), .lft_op_17_06(net1943[0:7]),
     .lft_op_17_05(net1944[0:7]), .lft_op_17_03(net1946[0:7]),
     .lft_op_17_02(net1947[0:7]), .lft_op_17_01(net1948[0:7]),
     .sdi_pad(sdi_pad), .shift_mi(shift), .sdo_pad(sdo_pad),
     .hold_b_r(hold_bbank), .hiz_b_mi(hiz_b), .update_mi(update),
     .r_mi(r), .tclk_mi(tclk), .bs_en_mi(bs_en),
     .slf_op_19_16(net1152[0:7]), .slf_op_18_16(net1153[0:7]),
     .sp12_h_l_17_15(net2016[0:23]), .slf_op_28_16(net1155[0:7]),
     .slf_op_27_16(net1156[0:7]), .slf_op_26_16(net1157[0:7]),
     .slf_op_25_16(net1158[0:7]), .slf_op_24_16(net1159[0:7]),
     .slf_op_23_16(net1160[0:7]), .slf_op_22_16(net1161[0:7]),
     .slf_op_21_16(net1162[0:7]), .slf_op_31_16(net1163[0:7]),
     .slf_op_30_16(net1164[0:7]), .slf_op_29_16(net1165[0:7]),
     .bnl_op_17_01(net1835[0:3]), .sp4_h_l_17_16(net2064[0:47]),
     .sp12_v_t_17_16(net1168[0:23]), .carry_out_31_16(net1169),
     .carry_out_30_16(net1170), .carry_out_29_16(net1171),
     .carry_out_28_16(net1172), .carry_out_27_16(net1173),
     .carry_out_26_16(net1174), .carry_out_24_16(net1175),
     .carry_out_23_16(net1176), .carry_out_22_16(net1177),
     .carry_out_21_16(net1178), .carry_out_20_16(net1179),
     .carry_out_19_16(net1180), .carry_out_18_16(net1181),
     .slf_op_17_01(net1909[0:7]), .slf_op_17_02(net1908[0:7]),
     .slf_op_17_03(net1907[0:7]), .slf_op_17_04(net1906[0:7]),
     .slf_op_17_05(net1905[0:7]), .slf_op_17_06(net1904[0:7]),
     .slf_op_17_07(net1903[0:7]), .slf_op_17_08(net1902[0:7]),
     .slf_op_17_09(net1901[0:7]), .slf_op_17_10(net1900[0:7]),
     .slf_op_17_11(net1899[0:7]), .slf_op_17_12(net1898[0:7]),
     .slf_op_17_13(net1897[0:7]), .slf_op_17_14(net1896[0:7]),
     .slf_op_17_15(net2083[0:7]), .cf_r(cf_r[383:0]),
     .sp12_v_t_18_16(net1198[0:23]), .sp12_v_t_19_16(net1199[0:23]),
     .sp12_v_t_20_16(net1200[0:23]), .sp12_v_t_22_16(net1201[0:23]),
     .sp12_v_t_21_16(net1202[0:23]), .sp12_v_t_23_16(net1203[0:23]),
     .sp12_v_t_24_16(net1204[0:23]), .sp12_v_t_25_16(net1205[0:23]),
     .sp12_v_t_26_16(net1206[0:23]), .sp12_v_t_27_16(net1207[0:23]),
     .sp12_v_t_28_16(net1208[0:23]), .sp12_v_t_29_16(net1209[0:23]),
     .sp12_v_t_30_16(net1210[0:23]), .sp12_v_t_31_16(net1211[0:23]),
     .sp12_v_t_32_16(net1212[0:23]), .tnr_op_17_16(net1213[0:7]),
     .sp12_h_l_17_13(net2018[0:23]), .sp12_h_l_17_11(net2020[0:23]),
     .sp12_h_l_17_10(net2021[0:23]), .sp12_h_l_17_12(net2019[0:23]),
     .sp12_h_l_17_08(net2023[0:23]), .sp12_h_l_17_07(net2024[0:23]),
     .sp12_h_l_17_09(net2022[0:23]), .sp12_h_l_17_06(net2025[0:23]),
     .sp12_h_l_17_04(net2027[0:23]), .sp12_h_l_17_02(net2029[0:23]),
     .sp12_h_l_17_05(net2026[0:23]), .sp12_h_l_17_03(net2028[0:23]),
     .sp12_h_l_17_16(net2015[0:23]), .sp12_h_l_17_01(net2030[0:23]),
     .sp4_v_t_18_16(net1228[0:47]), .sp4_v_t_19_16(net1229[0:47]),
     .sp4_v_t_20_16(net1230[0:47]), .sp4_v_t_21_16(net1231[0:47]),
     .sp4_v_t_22_16(net1232[0:47]), .sp4_v_t_23_16(net1233[0:47]),
     .sp4_v_t_24_16(net1234[0:47]), .sp4_v_t_25_16(net1235[0:47]),
     .sp4_v_t_26_16(net1236[0:47]), .sp4_v_t_27_16(net1237[0:47]),
     .sp4_v_t_28_16(net1238[0:47]), .sp4_v_t_29_16(net1239[0:47]),
     .sp4_v_t_30_16(net1240[0:47]), .sp4_v_t_31_16(net1241[0:47]),
     .sp4_v_t_32_16(net1242[0:47]), .sp4_v_t_33_16(net1243[0:15]),
     .top_op_17_16(net1244[0:7]), .sp12_h_l_17_14(net2017[0:23]),
     .sp4_h_l_17_14(net2066[0:47]), .sp4_h_l_17_13(net2067[0:47]),
     .sp4_h_l_17_12(net2068[0:47]), .sp4_h_l_17_11(net2069[0:47]),
     .sp4_h_l_17_10(net2070[0:47]), .sp4_h_l_17_09(net2071[0:47]),
     .sp4_h_l_17_08(net2072[0:47]), .sp4_h_l_17_07(net2073[0:47]),
     .sp4_h_l_17_06(net2074[0:47]), .sp4_h_l_17_05(net2075[0:47]),
     .sp4_h_l_17_04(net2076[0:47]), .sp4_h_l_17_03(net2077[0:47]),
     .sp4_h_l_17_02(net2078[0:47]), .slf_op_17_16(net1775[0:7]),
     .tnl_op_17_16(n_slf_op_16_17[7:0]), .sp4_h_l_17_01(net2079[0:47]),
     .slf_op_20_16(net1262[0:7]), .vdd_cntl_r(vdd_cntl_r[271:0]),
     .lft_op_17_12(net1937[0:7]), .wl_r(wl_r[271:0]),
     .bl(bl_bot[1743:874]), .reset_r(reset_b_r[271:0]),
     .pgate_r(pgate_r[271:0]), .lft_op_17_15(net1934[0:7]),
     .lft_op_17_16(net1933[0:7]), .slf_op_32_16(net1271[0:7]),
     .carry_out_32_16(net1272), .sp4_h_l_17_00(net1837[0:15]),
     .sp4_h_l_17_15(net2065[0:47]), .tnr_op_18_16(net1275[0:7]),
     .update_i(net1931), .tiegnd(tiegnd), .tclk_i(net1932),
     .shift_i(net1964), .sdi(net1965), .r_i(net1966), .purst(purst),
     .prog(prog), .mode_i(net1967), .hiz_b_i(net1968),
     .glb_in(glb_net[7:0]), .bs_en_i(net1986),
     .bm_wdummymux_en_i(net946), .bm_sweb_i(net1290[0:1]),
     .bm_sreb_i(net939), .bm_sdi_i(bm_bank30_sdi_o[3:2]),
     .bm_sclkrw_i(net1293[0:1]), .bm_sclk_i(bm_bank30_sclk_o[1]),
     .bm_sa_i(net942[0:7]), .bm_rcapmux_en_i(net945),
     .bm_init_i(net943), .update_o(net1298), .tclk_o(net1299),
     .shift_o(net1300), .sdo(net1301), .r_o(net1302), .mode_o(net1303),
     .hiz_b_o(net1304), .cf_b(cf_b[767:384]), .bs_en_o(net1306),
     .bm_wdummymux_en_o(net1307), .bm_sweb_o(bm_sweb_b2_o[1:0]),
     .bm_sreb_o(net1309), .bm_sdo_o(net1310[0:1]),
     .bm_sdi_o(bm_sdi_b2_o[1:0]), .bm_sclkrw_o(bm_sclkrw_b2_o[1:0]),
     .bm_sclk_o(net1313), .bm_sa_o(net1314[0:7]),
     .bm_rcapmux_en_o(net1315), .bm_init_o(net1316));
quad_tr_ice8 I_quad_tr_ice8 ( .slf_op_17_33(net1038[0:3]),
     .sp4_v_b_17_32(net01760[0:47]), .sp4_v_b_17_31(net01761[0:47]),
     .sp4_v_b_17_30(net01762[0:47]), .sp4_v_b_17_29(net01763[0:47]),
     .sp4_v_b_17_28(net01764[0:47]), .sp4_v_b_17_27(net01765[0:47]),
     .sp4_v_b_17_26(net01766[0:47]), .sp4_v_b_17_25(net01767[0:47]),
     .sp4_v_b_17_24(net01768[0:47]), .sp4_v_b_17_23(net01769[0:47]),
     .sp4_v_b_17_22(net01770[0:47]), .sp4_v_b_17_21(net01771[0:47]),
     .sp4_v_b_17_20(net01772[0:47]), .sp4_v_b_17_19(net01773[0:47]),
     .sp4_v_b_17_18(net01774[0:47]), .ceb_i(net01437),
     .ceb_o(net01682),
     .end_of_startup_top_r(end_of_startup_top[31:16]),
     .fabric_out_33_18(hold_rbank), .pado_t(pado_t[59:30]),
     .padeb_t(padeb_t[59:30]), .padin_t(padin_t[59:30]),
     .pado_r(pado_r[54:28]), .padin_r(padin_r[54:28]),
     .padeb_r(padeb_r[54:28]), .fabric_out_17_33(fabric_out_17_33),
     .fabric_out_33_17(fabric_out_33_17), .padin_136(padin_136),
     .padin_192(padin_192), .bm_sdo_i(net1459),
     .slf_op_33_17(slf_op_33_17[3:0]), .sp4_h_l_17_33(net1577[0:15]),
     .cf_t(cf_t[767:384]), .carry_in_27_17(net1173),
     .carry_in_29_17(net1171), .carry_in_30_17(net1170),
     .carry_in_31_17(net1169), .carry_in_32_17(net1272),
     .carry_in_23_17(net1176), .carry_in_18_17(net1181),
     .carry_in_19_17(net1180), .carry_in_20_17(net1179),
     .carry_in_21_17(net1178), .carry_in_22_17(net1177),
     .bot_op_17_17(net1775[0:7]), .bot_op_18_17(net1153[0:7]),
     .bnr_op_32_17({slf_op_33_16[3], slf_op_33_16[2], slf_op_33_16[1],
     slf_op_33_16[0], slf_op_33_16[3], slf_op_33_16[2],
     slf_op_33_16[1], slf_op_33_16[0]}), .bnr_op_31_17(net1271[0:7]),
     .bnr_op_30_17(net1163[0:7]), .bnr_op_29_17(net1164[0:7]),
     .bnr_op_28_17(net1165[0:7]), .bnr_op_27_17(net1155[0:7]),
     .bnr_op_26_17(net1156[0:7]), .bnr_op_25_17(net1157[0:7]),
     .bnr_op_24_17(net1158[0:7]), .bnr_op_23_17(net1159[0:7]),
     .bnr_op_22_17(net1160[0:7]), .bnr_op_21_17(net1161[0:7]),
     .bnr_op_20_17(net1162[0:7]), .bnr_op_19_17(net1262[0:7]),
     .bnr_op_18_17(net1152[0:7]), .bnr_op_17_17(net1153[0:7]),
     .slf_op_27_17(net1105[0:7]), .sp12_v_b_32_17(net1212[0:23]),
     .sp12_v_b_31_17(net1211[0:23]), .sp12_v_b_30_17(net1210[0:23]),
     .sp12_v_b_29_17(net1209[0:23]), .sp12_v_b_28_17(net1208[0:23]),
     .sp12_v_b_27_17(net1207[0:23]), .sp12_v_b_26_17(net1206[0:23]),
     .sp12_v_b_25_17(net1205[0:23]), .sp12_v_b_24_17(net1204[0:23]),
     .sp12_v_b_23_17(net1203[0:23]), .sp12_v_b_22_17(net1201[0:23]),
     .sp12_v_b_21_17(net1202[0:23]), .sp12_v_b_20_17(net1200[0:23]),
     .sp12_v_b_19_17(net1199[0:23]), .sp12_v_b_18_17(net1198[0:23]),
     .sp12_v_b_17_17(net1168[0:23]), .tievdd(tievdd), .tiegnd(tiegnd),
     .sp4_h_l_17_29(net1634[0:47]), .sp4_h_l_17_30(net1633[0:47]),
     .sp4_h_l_17_27(net1636[0:47]), .sp4_h_l_17_26(net1637[0:47]),
     .sp4_h_l_17_24(net1639[0:47]), .sp4_h_l_17_20(net1643[0:47]),
     .sp4_h_l_17_25(net1638[0:47]), .sp4_h_l_17_23(net1640[0:47]),
     .sp4_h_l_17_22(net1641[0:47]), .sp4_h_l_17_21(net1642[0:47]),
     .sp4_h_l_17_19(net1644[0:47]), .sp4_h_l_17_18(net1645[0:47]),
     .sp4_h_l_17_17(net1599[0:47]), .purst(purst), .prog(prog),
     .glb_in(glb_net[7:0]),
     .end_of_startup_lft_b(end_of_startup_r[31:16]),
     .bm_sreb_i(net1309), .bm_sdi_i(bm_sdi_b2_o[1]),
     .bm_sclkrw_i(bm_sclkrw_b2_o[1]), .bm_sclk_i(net1313),
     .bm_sa_i(net1314[0:7]), .bm_rcapmux_en_i(net1315),
     .bm_init_i(net1316), .update_o(net1785), .tclk_o(net1788),
     .sdi(net1301), .sp4_v_b_32_17(net1242[0:47]),
     .sp4_v_b_31_17(net1241[0:47]), .slf_op_17_30(net1662[0:7]),
     .sp4_v_b_30_17(net1240[0:47]), .sp4_v_b_29_17(net1239[0:47]),
     .sp4_v_b_28_17(net1238[0:47]), .sp4_v_b_27_17(net1237[0:47]),
     .sp4_v_b_26_17(net1236[0:47]), .sp4_v_b_25_17(net1235[0:47]),
     .sp4_v_b_24_17(net1234[0:47]), .sp4_v_b_23_17(net1233[0:47]),
     .sp4_v_b_22_17(net1232[0:47]), .sp4_v_b_21_17(net1231[0:47]),
     .sp4_v_b_20_17(net1230[0:47]), .sp4_v_b_19_17(net1229[0:47]),
     .sp4_v_b_18_17(net1228[0:47]), .shift_o(net1789),
     .shift_i(net1300), .hold_t_r(hold_tbank), .r_o(net1791),
     .update_i(net1298), .mode_i(net1303), .tnl_op_17_32(net1777[0:3]),
     .sdo(net1790), .mode_o(net1794), .hiz_b_i(net1304),
     .hiz_b_o(net1795), .bs_en_i(net1306), .r_i(net1302),
     .spi_ss_in_b_r(spi_ss_in_r[63:32]),
     .sp12_h_l_17_32(net1600[0:23]), .bot_op_26_17(net1157[0:7]),
     .bot_op_27_17(net1156[0:7]), .bot_op_28_17(net1155[0:7]),
     .bot_op_29_17(net1165[0:7]), .bot_op_30_17(net1164[0:7]),
     .bot_op_31_17(net1163[0:7]), .bot_op_32_17(net1271[0:7]),
     .sp4_v_b_33_17(net1243[0:15]), .bot_op_24_17(net1159[0:7]),
     .bot_op_19_17(net1152[0:7]), .bot_op_20_17(net1262[0:7]),
     .bot_op_21_17(net1162[0:7]), .bot_op_22_17(net1161[0:7]),
     .bot_op_23_17(net1160[0:7]), .bs_en_o(net1797), .tclk_i(net1299),
     .bm_sweb_o(net1456), .bm_sreb_o(net1457), .bm_sdo_o(bm_sdo_b3_o),
     .bm_sdi_o(net1459), .bm_sclkrw_o(net1460), .bm_sclk_o(net1461),
     .bm_sa_o(net1462[0:7]), .bm_rcapmux_en_o(net1463),
     .bm_init_o(net1464), .lft_op_17_17(n_slf_op_16_17[7:0]),
     .lft_op_17_18(net1660[0:7]), .lft_op_17_19(net1659[0:7]),
     .lft_op_17_20(net1658[0:7]), .lft_op_17_21(net1657[0:7]),
     .lft_op_17_22(net1656[0:7]), .lft_op_17_23(n_slf_op_16_23[7:0]),
     .lft_op_17_24(net1654[0:7]), .lft_op_17_25(net1653[0:7]),
     .lft_op_17_26(net1652[0:7]), .lft_op_17_27(net1651[0:7]),
     .lft_op_17_28(net1650[0:7]), .lft_op_17_29(net1649[0:7]),
     .lft_op_17_30(net1648[0:7]), .lft_op_17_31(net1647[0:7]),
     .cf_r(cf_r[767:384]), .sp4_v_b_17_17(net1128[0:47]),
     .bnl_op_33_17(net1271[0:7]), .bnl_op_32_17(net1163[0:7]),
     .bnl_op_31_17(net1164[0:7]), .bnl_op_30_17(net1165[0:7]),
     .bnl_op_29_17(net1155[0:7]), .bnl_op_28_17(net1156[0:7]),
     .bnl_op_27_17(net1157[0:7]), .bnl_op_26_17(net1158[0:7]),
     .bnl_op_25_17(net1159[0:7]), .bnl_op_24_17(net1160[0:7]),
     .bnl_op_23_17(net1161[0:7]), .bnl_op_22_17(net1162[0:7]),
     .bnl_op_21_17(net1262[0:7]), .bnl_op_20_17(net1152[0:7]),
     .bnl_op_19_17(net1153[0:7]), .slf_op_17_28(net1587[0:7]),
     .slf_op_17_26(net1589[0:7]), .slf_op_17_25(net1590[0:7]),
     .slf_op_17_27(net1588[0:7]), .slf_op_17_23(net1592[0:7]),
     .slf_op_17_22(net1593[0:7]), .slf_op_17_24(net1591[0:7]),
     .slf_op_17_21(net1594[0:7]), .slf_op_17_19(net1596[0:7]),
     .slf_op_17_20(net1595[0:7]), .slf_op_17_18(net1597[0:7]),
     .slf_op_17_31(net1585[0:7]), .slf_op_21_17(net1099[0:7]),
     .slf_op_20_17(net1098[0:7]), .slf_op_19_17(net1275[0:7]),
     .slf_op_18_17(net1213[0:7]), .slf_op_31_17(net1109[0:7]),
     .slf_op_30_17(net1108[0:7]), .slf_op_29_17(net1107[0:7]),
     .slf_op_28_17(net1106[0:7]), .slf_op_32_17(net1110[0:7]),
     .slf_op_26_17(net1104[0:7]), .slf_op_25_17(net1103[0:7]),
     .slf_op_24_17(net1102[0:7]), .slf_op_23_17(net1101[0:7]),
     .slf_op_17_17(net1244[0:7]), .slf_op_22_17(net1100[0:7]),
     .carry_in_24_17(net1175), .carry_in_26_17(net1174),
     .slf_op_17_32(net1755[0:7]), .slf_op_17_29(net1586[0:7]),
     .sp12_h_l_17_30(net1602[0:23]), .sp12_h_l_17_29(net1603[0:23]),
     .sp12_h_l_17_28(net1604[0:23]), .sp12_h_l_17_27(net1605[0:23]),
     .sp12_h_l_17_26(net1606[0:23]), .sp12_h_l_17_25(net1607[0:23]),
     .sp12_h_l_17_24(net1608[0:23]), .sp12_h_l_17_23(net1609[0:23]),
     .sp12_h_l_17_22(net1610[0:23]), .sp12_h_l_17_21(net1611[0:23]),
     .sp12_h_l_17_20(net1612[0:23]), .sp12_h_l_17_19(net1613[0:23]),
     .sp12_h_l_17_18(net1614[0:23]), .lft_op_17_32(net1646[0:7]),
     .sp12_h_l_17_17(net1615[0:23]), .vdd_cntl_r(vdd_cntl_r[543:272]),
     .carry_in_17_17(net1082), .sp4_h_l_17_28(net1635[0:47]),
     .wl_r(wl_r[543:272]), .bm_wdummymux_en_o(net1548),
     .bm_wdummymux_en_i(net1307), .bm_sweb_i(bm_sweb_b2_o[1]),
     .carry_in_28_17(net1172), .bnl_op_17_17(net1933[0:7]),
     .bl(bl_top[1743:874]), .reset_r(reset_b_r[543:272]),
     .pgate_r(pgate_r[543:272]), .sp4_h_l_17_31(net1632[0:47]),
     .sp4_h_l_17_32(net1756[0:47]), .bnl_op_18_17(net1775[0:7]),
     .bot_op_25_17(net1158[0:7]), .sp12_h_l_17_31(net1601[0:23]),
     .hold_r_t(hold_rbank));
quad_tl_ice8 I_quad_tl_ice8 ( .ceb_i(net01682), .ceb_o(net0901),
     .tnr_op_16_32(net1038[0:3]),
     .end_of_startup_top_l(end_of_startup_top[15:0]),
     .padin_l_t(padin_l[49:24]), .padeb_l_t(padeb_l[49:24]),
     .pado_l_t(pado_l[49:24]), .fabric_out_15_33(hold_tbank),
     .pado_t_l(pado_t[29:0]), .padeb_t_l(padeb_t[29:0]),
     .padin_t_l(padin_t[29:0]), .fabric_out_16_33(fabric_out_16_33),
     .fabric_out_00_17(fabric_out_00_17), .padin_26(padin_26),
     .padin_193(padin_193), .bm_sdo_o(bm_sdo_b1_o),
     .slf_op_00_17(slf_op_00_17[3:0]), .bnr_op_00_17(net1576[0:7]),
     .sp4_h_r_16_33(net1577[0:15]), .cf_t(cf_t[383:0]),
     .hold_l_t(hold_lbank), .hold_t_l(hold_tbank),
     .bnr_op_08_17(net1955[0:7]), .rgt_op_16_31(net1585[0:7]),
     .rgt_op_16_29(net1586[0:7]), .rgt_op_16_28(net1587[0:7]),
     .rgt_op_16_27(net1588[0:7]), .rgt_op_16_26(net1589[0:7]),
     .rgt_op_16_25(net1590[0:7]), .rgt_op_16_24(net1591[0:7]),
     .rgt_op_16_23(net1592[0:7]), .rgt_op_16_22(net1593[0:7]),
     .rgt_op_16_21(net1594[0:7]), .rgt_op_16_20(net1595[0:7]),
     .rgt_op_16_19(net1596[0:7]), .rgt_op_16_18(net1597[0:7]),
     .rgt_op_16_17(net1244[0:7]), .sp4_h_r_16_17(net1599[0:47]),
     .sp12_h_r_16_32(net1600[0:23]), .sp12_h_r_16_31(net1601[0:23]),
     .sp12_h_r_16_30(net1602[0:23]), .sp12_h_r_16_29(net1603[0:23]),
     .sp12_h_r_16_28(net1604[0:23]), .sp12_h_r_16_27(net1605[0:23]),
     .sp12_h_r_16_26(net1606[0:23]), .sp12_h_r_16_25(net1607[0:23]),
     .sp12_h_r_16_24(net1608[0:23]), .sp12_h_r_16_23(net1609[0:23]),
     .sp12_h_r_16_22(net1610[0:23]), .sp12_h_r_16_21(net1611[0:23]),
     .sp12_h_r_16_20(net1612[0:23]), .sp12_h_r_16_19(net1613[0:23]),
     .sp12_h_r_16_18(net1614[0:23]), .sp12_h_r_16_17(net1615[0:23]),
     .sp4_r_v_b_16_32(net01760[0:47]),
     .sp4_r_v_b_16_31(net01761[0:47]),
     .sp4_r_v_b_16_30(net01762[0:47]),
     .sp4_r_v_b_16_29(net01763[0:47]),
     .sp4_r_v_b_16_28(net01764[0:47]),
     .sp4_r_v_b_16_27(net01765[0:47]),
     .sp4_r_v_b_16_26(net01766[0:47]),
     .sp4_r_v_b_16_25(net01767[0:47]),
     .sp4_r_v_b_16_24(net01768[0:47]),
     .sp4_r_v_b_16_23(net01769[0:47]),
     .sp4_r_v_b_16_22(net01770[0:47]),
     .sp4_r_v_b_16_21(net01771[0:47]),
     .sp4_r_v_b_16_20(net01772[0:47]),
     .sp4_r_v_b_16_19(net01773[0:47]),
     .sp4_r_v_b_16_18(net01774[0:47]), .sp4_r_v_b_16_17(net1128[0:47]),
     .sp4_h_r_16_31(net1632[0:47]), .sp4_h_r_16_30(net1633[0:47]),
     .sp4_h_r_16_29(net1634[0:47]), .sp4_h_r_16_28(net1635[0:47]),
     .sp4_h_r_16_27(net1636[0:47]), .sp4_h_r_16_26(net1637[0:47]),
     .sp4_h_r_16_25(net1638[0:47]), .sp4_h_r_16_24(net1639[0:47]),
     .sp4_h_r_16_23(net1640[0:47]), .sp4_h_r_16_22(net1641[0:47]),
     .sp4_h_r_16_21(net1642[0:47]), .sp4_h_r_16_20(net1643[0:47]),
     .sp4_h_r_16_19(net1644[0:47]), .sp4_h_r_16_18(net1645[0:47]),
     .slf_op_16_32(net1646[0:7]), .slf_op_16_31(net1647[0:7]),
     .slf_op_16_30(net1648[0:7]), .slf_op_16_29(net1649[0:7]),
     .slf_op_16_28(net1650[0:7]), .slf_op_16_27(net1651[0:7]),
     .slf_op_16_26(net1652[0:7]), .slf_op_16_25(net1653[0:7]),
     .slf_op_16_24(net1654[0:7]), .slf_op_16_23(n_slf_op_16_23[7:0]),
     .slf_op_16_22(net1656[0:7]), .slf_op_16_21(net1657[0:7]),
     .slf_op_16_20(net1658[0:7]), .slf_op_16_19(net1659[0:7]),
     .slf_op_16_18(net1660[0:7]), .slf_op_16_17(n_slf_op_16_17[7:0]),
     .rgt_op_16_30(net1662[0:7]), .bnr_op_07_17(net1956[0:7]),
     .bnr_op_06_17(net1957[0:7]), .sp4_v_b_15_17(net2045[0:47]),
     .sp4_v_b_16_17(net2046[0:47]), .bnl_op_01_17({slf_op_00_16[3],
     slf_op_00_16[2], slf_op_00_16[1], slf_op_00_16[0],
     slf_op_00_16[3], slf_op_00_16[2], slf_op_00_16[1],
     slf_op_00_16[0]}), .bnl_op_02_17(net1576[0:7]),
     .bnl_op_03_17(net1962[0:7]), .bnl_op_04_17(net1961[0:7]),
     .bnl_op_05_17(net1960[0:7]), .bnl_op_06_17(net1959[0:7]),
     .bnl_op_07_17(net1958[0:7]), .bnl_op_08_17(net1957[0:7]),
     .bnl_op_09_17(net1956[0:7]), .bnl_op_10_17(net1955[0:7]),
     .bnl_op_11_17(net1954[0:7]), .bnl_op_12_17(net1953[0:7]),
     .bnl_op_13_17(net1952[0:7]), .bnl_op_14_17(net1951[0:7]),
     .bnl_op_15_17(net1950[0:7]), .bnl_op_16_17(net1949[0:7]),
     .bnr_op_09_17(net1954[0:7]), .bnr_op_10_17(net1953[0:7]),
     .bnr_op_11_17(net1952[0:7]), .bnr_op_12_17(net1951[0:7]),
     .bnr_op_13_17(net1950[0:7]), .bnr_op_14_17(net1949[0:7]),
     .bnr_op_15_17(net1933[0:7]), .sp4_v_b_00_17(net2047[0:15]),
     .sp4_v_b_01_17(net2031[0:47]), .sp4_v_b_02_17(net2032[0:47]),
     .sp4_v_b_03_17(net2033[0:47]), .sp4_v_b_04_17(net2034[0:47]),
     .sp4_v_b_05_17(net2035[0:47]), .sp4_v_b_06_17(net2036[0:47]),
     .sp4_v_b_07_17(net2037[0:47]), .sp4_v_b_08_17(net2038[0:47]),
     .sp4_v_b_09_17(net2039[0:47]), .sp4_v_b_10_17(net2040[0:47]),
     .sp4_v_b_11_17(net2041[0:47]), .sp4_v_b_12_17(net2042[0:47]),
     .sp4_v_b_13_17(net2043[0:47]), .sp4_v_b_14_17(net2044[0:47]),
     .bnr_op_05_17(net1958[0:7]), .bnr_op_04_17(net1959[0:7]),
     .bnr_op_03_17(net1960[0:7]), .bnr_op_02_17(net1961[0:7]),
     .bnr_op_01_17(net1962[0:7]), .slf_op_15_17(net1859[0:7]),
     .slf_op_14_17(net1860[0:7]), .slf_op_13_17(net1861[0:7]),
     .slf_op_12_17(net1862[0:7]), .slf_op_11_17(net1863[0:7]),
     .slf_op_10_17(net1864[0:7]), .slf_op_09_17(net1865[0:7]),
     .slf_op_08_17(net1866[0:7]), .slf_op_07_17(net1867[0:7]),
     .slf_op_06_17(net1868[0:7]), .slf_op_05_17(net1869[0:7]),
     .slf_op_04_17(net1870[0:7]), .slf_op_03_17(net1871[0:7]),
     .slf_op_02_17(net1872[0:7]), .slf_op_01_17(n_slf_op_01_17[7:0]),
     .sp12_v_b_15_17(net2000[0:23]), .sp12_v_b_14_17(net2001[0:23]),
     .sp12_v_b_13_17(net2002[0:23]), .sp12_v_b_12_17(net2003[0:23]),
     .sp12_v_b_11_17(net2004[0:23]), .sp12_v_b_10_17(net2005[0:23]),
     .sp12_v_b_09_17(net2006[0:23]), .sp12_v_b_08_17(net2007[0:23]),
     .sp12_v_b_07_17(net2008[0:23]), .sp12_v_b_06_17(net2009[0:23]),
     .sp12_v_b_05_17(net2010[0:23]), .sp12_v_b_04_17(net2011[0:23]),
     .sp12_v_b_03_17(net2012[0:23]), .sp12_v_b_02_17(net2013[0:23]),
     .sp12_v_b_01_17(net2014[0:23]), .bot_op_15_17(net1949[0:7]),
     .bot_op_14_17(net1950[0:7]), .bot_op_13_17(net1951[0:7]),
     .bot_op_12_17(net1952[0:7]), .bot_op_11_17(net1953[0:7]),
     .bot_op_10_17(net1954[0:7]), .bot_op_09_17(net1955[0:7]),
     .bot_op_08_17(net1956[0:7]), .bot_op_07_17(net1957[0:7]),
     .bot_op_06_17(net1958[0:7]), .bot_op_05_17(net1959[0:7]),
     .bot_op_04_17(net1960[0:7]), .bot_op_03_17(net1961[0:7]),
     .bot_op_02_17(net1962[0:7]), .bot_op_01_17(net1576[0:7]),
     .rgt_op_16_32(net1755[0:7]), .sp4_h_r_16_32(net1756[0:47]),
     .carry_in_16_17(net1971), .carry_in_15_17(net1972),
     .carry_in_14_17(net1973), .carry_in_13_17(net1974),
     .carry_in_12_17(net1975), .carry_in_11_17(net1976),
     .carry_in_10_17(net1977), .carry_in_09_17(net1978),
     .carry_in_07_17(net1979), .carry_in_06_17(net1980),
     .carry_in_01_17(net1985), .carry_in_02_17(net1984),
     .carry_in_03_17(net1983), .carry_in_04_17(net1982),
     .carry_in_05_17(net1981),
     .end_of_startup_lft_t(end_of_startup_l[31:16]),
     .bot_op_16_17(net1933[0:7]), .sp12_v_b_16_17(net1999[0:23]),
     .bnr_op_16_17(net1775[0:7]), .slf_op_16_33(net1777[0:3]),
     .bm_sclkrw_o(bm_sclkrw_b1_o), .bm_sdi_o(bm_sdo_b1_i),
     .bm_sweb_o(bm_sweb_b1_o), .bm_sdo_i(bm_sdo_b1_i),
     .bm_sclkrw_i(bm_sclkrw_b0_o[1]), .bm_sdi_i(bm_sdi_b0_o[1]),
     .bm_sweb_i(bm_sweb_b0_o[1]), .update_i(net1785), .tievdd(tievdd),
     .tiegnd(tiegnd), .tclk_i(net1788), .shift_i(net1789),
     .sdi(net1790), .r_i(net1791), .purst(purst), .prog(prog),
     .mode_i(net1794), .hiz_b_i(net1795), .glb_in(glb_net[7:0]),
     .bs_en_i(net1797), .bm_wdummymux_en_i(net1987),
     .bm_sreb_i(net1989), .bm_sclk_i(net1993), .bm_sa_i(net1994[0:7]),
     .bm_rcapmux_en_i(net1995), .bm_init_i(net1996),
     .update_o(net1841), .tclk_o(net1892), .shift_o(net1893),
     .sdo(net1894), .r_o(net1910), .mode_o(net1913), .hiz_b_o(net1916),
     .cf_l(cf_l[767:384]), .bs_en_o(net1919),
     .bm_wdummymux_en_o(bm_wdummymux_en_b1_o),
     .bm_sreb_o(bm_sreb_b1_o), .bm_sclk_o(bm_sclk_b1_o),
     .bm_sa_o(bm_sa_b1_o[7:0]), .bm_rcapmux_en_o(bm_rcapmux_en_b1_o),
     .bm_init_o(bm_init_b1_o), .wl_l(wl_l[543:272]),
     .vdd_cntl_l(vdd_cntl_l[543:272]), .reset_l(reset_b_l[543:272]),
     .pgate_l(pgate_l[543:272]), .bl(bl_top[869:0]));
bram_hbuffer_1xbank I2 ( .bm_wdummymux_en_o(net1921),
     .bm_sweb_i(net916), .bm_sreb_i(net917), .bm_sdi_i(net918[0:1]),
     .bm_sclk_i(net919), .bm_sa_i(net920[0:7]), .bm_init_i(net921),
     .bm_banksel_o(bm_bank10_banksel_o[1:0]), .bm_rcapmux_en_i(net923),
     .bm_wdummymux_en_i(net924), .bm_sweb_o(net1006),
     .bm_sreb_o(net1923), .bm_sdi_o(net1925[0:1]), .bm_sclk_o(net1927),
     .bm_sa_o(net1928[0:7]), .bm_init_o(net1930),
     .bm_rcapmux_en_o(net1929), .bm_sclkrw_i(net932),
     .bm_sclkrw_o(net1005), .bm_sdo_i(net1007[0:1]),
     .bm_banksel_i(net935[0:1]), .bm_sdo_o(net936[0:1]));
bram_hbuffer_1xbank I17 ( .bm_wdummymux_en_o(net924),
     .bm_sweb_i(net938), .bm_sreb_i(net939),
     .bm_sdi_i(bm_bank30_sdi_o[1:0]), .bm_sclk_i(bm_bank30_sclk_o[0]),
     .bm_sa_i(net942[0:7]), .bm_init_i(net943),
     .bm_banksel_o(net935[0:1]), .bm_rcapmux_en_i(net945),
     .bm_wdummymux_en_i(net946), .bm_sweb_o(net916),
     .bm_sreb_o(net917), .bm_sdi_o(net918[0:1]), .bm_sclk_o(net919),
     .bm_sa_o(net920[0:7]), .bm_init_o(net921),
     .bm_rcapmux_en_o(net923), .bm_sclkrw_i(net954),
     .bm_sclkrw_o(net932), .bm_sdo_i(net936[0:1]),
     .bm_banksel_i(bm_bank30_banksel_o[1:0]),
     .bm_sdo_o(bm_bank30_sdo_i[1:0]));
bram_hbuffer_dff_2xbank I24 ( .bm_sweb_i(net959), .bm_sreb_i(net960),
     .bm_sclk_i(net961), .bm_sa_i(net962[0:7]), .bm_init_i(net963),
     .bm_banksel_o(bm_bank30_banksel_o[3:0]), .bm_rcapmux_en_i(net965),
     .bm_wdummymux_en_i(net966), .bm_sweb_o(net938),
     .bm_sreb_o(net939), .bm_sclk_o(bm_bank30_sclk_o[1:0]),
     .bm_sa_o(net942[0:7]), .bm_init_o(net943), .bm_sclkrw_i(net972),
     .bm_sclkrw_o(net954), .bm_sdi_i(net974[0:3]),
     .bm_sdo_o(net975[0:3]), .bm_sdi_o(bm_bank30_sdi_o[3:0]),
     .bm_rcapmux_en_o(net945), .bm_wdummymux_en_o(net946),
     .bm_banksel_i(net979[0:3]), .bm_sdo_i(bm_bank30_sdo_i[3:0]));
bram_hbuffer_2xbank I20 ( .bm_wdummymux_en_o(net966),
     .bm_sweb_i(bm_sweb_i), .bm_sreb_i(bm_sreb_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_init_i(bm_init_i), .bm_banksel_o(net979[0:3]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_o(net959),
     .bm_sreb_o(net960), .bm_sclk_o(net961), .bm_sa_o(net962[0:7]),
     .bm_init_o(net963), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclkrw_o(net972), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sdo_o(bm_sdo_o[3:0]), .bm_sdi_o(net974[0:3]),
     .bm_rcapmux_en_o(net965), .bm_banksel_i(bm_banksel_i[3:0]),
     .bm_sdo_i(net975[0:3]));
bram_bank_logic_bot I10 ( .bm_sdo_i(net1990[0:1]), .bm_sclk_i(net1927),
     .bm_sclkrw_i(net1005), .bm_sweb_i(net1006),
     .bm_sdo_o(net1007[0:1]), .bm_sweb_o(net1922[0:1]),
     .bm_sclkrw_o(net1926[0:1]),
     .bm_banksel_i(bm_bank10_banksel_o[1:0]));
bram_bank_logic_bot I21 ( .bm_sdo_i(net1310[0:1]),
     .bm_sclk_i(bm_bank30_sclk_o[1]), .bm_sclkrw_i(net954),
     .bm_sweb_i(net938), .bm_sdo_o(bm_bank30_sdo_i[3:2]),
     .bm_sweb_o(net1290[0:1]), .bm_sclkrw_o(net1293[0:1]),
     .bm_banksel_i(bm_bank30_banksel_o[3:2]));

endmodule
// Library - chip, Cell - chip_ice8f, View - schematic
// LAST TIME SAVED: Jun  6 17:34:55 2008
// NETLIST TIME: Nov 14 16:17:21 2008
`timescale 1ns / 1ns 

module chip_ice8f ( tdo, VREFSSTL, cdone, uio_bbank, uio_lbank,
     uio_rbank, uio_tbank, vpp, creset_b, tck, tdi, tms, trstb );

output  tdo;

inout  VREFSSTL, cdone, vpp;

input  creset_b, tck, tdi, tms, trstb;

inout [59:0]  uio_tbank;
inout [56:0]  uio_bbank;
inout [49:0]  uio_lbank;
inout [54:0]  uio_rbank;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [49:0]  in_lbank;

wire  [54:0]  out_rbank;

wire  [7:0]  bm_sa_i;

wire  [543:0]  pgate_r;

wire  [543:0]  wl_r;

wire  [0:31]  net190;

wire  [3:0]  bm_sdi_i;

wire  [59:0]  in_tbank;

wire  [543:0]  wl_l;

wire  [3:0]  bm_sdo_o;

wire  [543:0]  vdd_cntl_r;

wire  [59:0]  out_tbank;

wire  [7:1]  psdo;

wire  [767:0]  cf_rbank;

wire  [59:0]  oen_tbank;

wire  [767:0]  cf_bbank;

wire  [56:0]  padin_b;

wire  [1743:0]  bl_top;

wire  [49:0]  out_lbank;

wire  [54:0]  oeb_rbank;

wire  [56:0]  padeb_b;

wire  [63:32]  spi_ss_in_bbank;

wire  [1743:0]  bl_bot;

wire  [3:0]  bm_banksel_i;

wire  [543:0]  reset_l;

wire  [49:0]  oen_lbank;

wire  [63:0]  spi_ss_in_r;

wire  [543:0]  vdd_cntl_l;

wire  [56:0]  pado_b;

wire  [767:0]  cf_tbank;

wire  [543:0]  reset_r;

wire  [767:0]  cf_lbank;

wire  [543:0]  pgate_l;

wire  [54:0]  in_rbank;

wire  [3:0]  last_rsr;



ring_route8k_f Iring_route ( .tiegnd(tiegnd), .tievdd(tievdd),
     .vpp(vpp), .ceb0(ceb), .cf_lbank({cf_lbank[736], cf_lbank[735],
     cf_lbank[734], cf_lbank[733], cf_lbank[732], cf_lbank[731],
     cf_lbank[730], cf_lbank[729], cf_lbank[728], cf_lbank[727],
     cf_lbank[726], cf_lbank[725], cf_lbank[724], cf_lbank[723],
     cf_lbank[722], cf_lbank[721], cf_lbank[720], cf_lbank[710],
     cf_lbank[709], cf_lbank[708], cf_lbank[707], cf_lbank[706],
     cf_lbank[705], cf_lbank[704], cf_lbank[703], cf_lbank[702],
     cf_lbank[701], cf_lbank[700], cf_lbank[699], cf_lbank[698],
     cf_lbank[697], cf_lbank[696], cf_lbank[662], cf_lbank[661],
     cf_lbank[660], cf_lbank[659], cf_lbank[658], cf_lbank[657],
     cf_lbank[656], cf_lbank[655], cf_lbank[654], cf_lbank[653],
     cf_lbank[652], cf_lbank[651], cf_lbank[650], cf_lbank[649],
     cf_lbank[648], cf_lbank[638], cf_lbank[637], cf_lbank[636],
     cf_lbank[635], cf_lbank[634], cf_lbank[633], cf_lbank[632],
     cf_lbank[631], cf_lbank[630], cf_lbank[629], cf_lbank[628],
     cf_lbank[627], cf_lbank[626], cf_lbank[625], cf_lbank[624],
     cf_lbank[590], cf_lbank[589], cf_lbank[588], cf_lbank[587],
     cf_lbank[586], cf_lbank[585], cf_lbank[584], cf_lbank[583],
     cf_lbank[582], cf_lbank[581], cf_lbank[580], cf_lbank[579],
     cf_lbank[578], cf_lbank[577], cf_lbank[576], cf_lbank[566],
     cf_lbank[565], cf_lbank[564], cf_lbank[563], cf_lbank[562],
     cf_lbank[561], cf_lbank[560], cf_lbank[559], cf_lbank[558],
     cf_lbank[557], cf_lbank[556], cf_lbank[555], cf_lbank[554],
     cf_lbank[553], cf_lbank[552], cf_lbank[542], cf_lbank[541],
     cf_lbank[540], cf_lbank[539], cf_lbank[538], cf_lbank[537],
     cf_lbank[536], cf_lbank[535], cf_lbank[534], cf_lbank[533],
     cf_lbank[532], cf_lbank[531], cf_lbank[530], cf_lbank[529],
     cf_lbank[528], cf_lbank[518], cf_lbank[517], cf_lbank[516],
     cf_lbank[515], cf_lbank[514], cf_lbank[513], cf_lbank[512],
     cf_lbank[511], cf_lbank[510], cf_lbank[509], cf_lbank[508],
     cf_lbank[507], cf_lbank[506], cf_lbank[505], cf_lbank[504],
     cf_lbank[494], cf_lbank[493], cf_lbank[492], cf_lbank[491],
     cf_lbank[490], cf_lbank[489], cf_lbank[488], cf_lbank[487],
     cf_lbank[486], cf_lbank[485], cf_lbank[484], cf_lbank[483],
     cf_lbank[482], cf_lbank[481], cf_lbank[480], cf_lbank[470],
     cf_lbank[469], cf_lbank[468], cf_lbank[467], cf_lbank[466],
     cf_lbank[465], cf_lbank[464], cf_lbank[463], cf_lbank[462],
     cf_lbank[461], cf_lbank[460], cf_lbank[459], cf_lbank[458],
     cf_lbank[457], cf_lbank[456], cf_lbank[446], cf_lbank[445],
     cf_lbank[444], cf_lbank[443], cf_lbank[442], cf_lbank[441],
     cf_lbank[440], cf_lbank[439], cf_lbank[438], cf_lbank[437],
     cf_lbank[436], cf_lbank[435], cf_lbank[434], cf_lbank[433],
     cf_lbank[432], cf_lbank[422], cf_lbank[421], cf_lbank[420],
     cf_lbank[419], cf_lbank[418], cf_lbank[417], cf_lbank[416],
     cf_lbank[415], cf_lbank[414], cf_lbank[413], cf_lbank[412],
     cf_lbank[411], cf_lbank[410], cf_lbank[409], cf_lbank[408],
     cf_lbank[398], cf_lbank[397], cf_lbank[396], cf_lbank[395],
     cf_lbank[394], cf_lbank[393], cf_lbank[392], cf_lbank[391],
     cf_lbank[390], cf_lbank[389], cf_lbank[388], cf_lbank[387],
     cf_lbank[386], cf_lbank[385], cf_lbank[384], cf_lbank[374],
     cf_lbank[373], cf_lbank[372], cf_lbank[371], cf_lbank[370],
     cf_lbank[369], cf_lbank[368], cf_lbank[367], cf_lbank[366],
     cf_lbank[365], cf_lbank[364], cf_lbank[363], cf_lbank[362],
     cf_lbank[361], cf_lbank[360], cf_lbank[326], cf_lbank[325],
     cf_lbank[324], cf_lbank[323], cf_lbank[322], cf_lbank[321],
     cf_lbank[320], cf_lbank[319], cf_lbank[318], cf_lbank[317],
     cf_lbank[316], cf_lbank[315], cf_lbank[314], cf_lbank[313],
     cf_lbank[312], cf_lbank[302], cf_lbank[301], cf_lbank[300],
     cf_lbank[299], cf_lbank[298], cf_lbank[297], cf_lbank[296],
     cf_lbank[295], cf_lbank[294], cf_lbank[293], cf_lbank[292],
     cf_lbank[291], cf_lbank[290], cf_lbank[289], cf_lbank[288],
     cf_lbank[278], cf_lbank[277], cf_lbank[276], cf_lbank[275],
     cf_lbank[274], cf_lbank[273], cf_lbank[272], cf_lbank[271],
     cf_lbank[270], cf_lbank[269], cf_lbank[268], cf_lbank[267],
     cf_lbank[266], cf_lbank[265], cf_lbank[264], cf_lbank[254],
     cf_lbank[253], cf_lbank[252], cf_lbank[251], cf_lbank[250],
     cf_lbank[249], cf_lbank[248], cf_lbank[247], cf_lbank[246],
     cf_lbank[245], cf_lbank[244], cf_lbank[243], cf_lbank[242],
     cf_lbank[241], cf_lbank[240], cf_lbank[230], cf_lbank[229],
     cf_lbank[228], cf_lbank[227], cf_lbank[226], cf_lbank[225],
     cf_lbank[224], cf_lbank[223], cf_lbank[222], cf_lbank[221],
     cf_lbank[220], cf_lbank[219], cf_lbank[218], cf_lbank[217],
     cf_lbank[216], cf_lbank[206], cf_lbank[205], cf_lbank[204],
     cf_lbank[203], cf_lbank[202], cf_lbank[201], cf_lbank[200],
     cf_lbank[199], cf_lbank[198], cf_lbank[197], cf_lbank[196],
     cf_lbank[195], cf_lbank[194], cf_lbank[193], cf_lbank[192],
     cf_lbank[182], cf_lbank[181], cf_lbank[180], cf_lbank[179],
     cf_lbank[178], cf_lbank[177], cf_lbank[176], cf_lbank[175],
     cf_lbank[174], cf_lbank[173], cf_lbank[172], cf_lbank[171],
     cf_lbank[170], cf_lbank[169], cf_lbank[168], cf_lbank[158],
     cf_lbank[157], cf_lbank[156], cf_lbank[155], cf_lbank[154],
     cf_lbank[153], cf_lbank[152], cf_lbank[151], cf_lbank[150],
     cf_lbank[149], cf_lbank[148], cf_lbank[147], cf_lbank[146],
     cf_lbank[145], cf_lbank[144], cf_lbank[134], cf_lbank[133],
     cf_lbank[132], cf_lbank[131], cf_lbank[130], cf_lbank[129],
     cf_lbank[128], cf_lbank[127], cf_lbank[126], cf_lbank[125],
     cf_lbank[124], cf_lbank[123], cf_lbank[122], cf_lbank[121],
     cf_lbank[120], cf_lbank[86], cf_lbank[85], cf_lbank[84],
     cf_lbank[83], cf_lbank[82], cf_lbank[81], cf_lbank[80],
     cf_lbank[79], cf_lbank[78], cf_lbank[77], cf_lbank[76],
     cf_lbank[75], cf_lbank[74], cf_lbank[73], cf_lbank[72],
     cf_lbank[62], cf_lbank[61], cf_lbank[60], cf_lbank[59],
     cf_lbank[58], cf_lbank[57], cf_lbank[56], cf_lbank[55],
     cf_lbank[54], cf_lbank[53], cf_lbank[52], cf_lbank[51],
     cf_lbank[50], cf_lbank[49], cf_lbank[48]}),
     .cf_r_ext(cf_rbank[450:449]), .cf_rbank({cf_rbank[720],
     cf_rbank[706], cf_rbank[696], cf_rbank[682], cf_rbank[672],
     cf_rbank[658], cf_rbank[648], cf_rbank[634], cf_rbank[624],
     cf_rbank[610], cf_rbank[600], cf_rbank[586], cf_rbank[576],
     cf_rbank[562], cf_rbank[552], cf_rbank[538], cf_rbank[528],
     cf_rbank[514], cf_rbank[504], cf_rbank[490], cf_rbank[480],
     cf_rbank[466], cf_rbank[456], cf_rbank[442], cf_rbank[432],
     cf_rbank[394], cf_rbank[384], cf_rbank[370], cf_rbank[360],
     cf_rbank[346], cf_rbank[336], cf_rbank[322], cf_rbank[312],
     cf_rbank[298], cf_rbank[288], cf_rbank[274], cf_rbank[264],
     cf_rbank[250], cf_rbank[240], cf_rbank[226], cf_rbank[216],
     cf_rbank[202], cf_rbank[192], cf_rbank[178], cf_rbank[168],
     cf_rbank[154], cf_rbank[144], cf_rbank[130], cf_rbank[120],
     cf_rbank[106], cf_rbank[96], cf_rbank[82], cf_rbank[72],
     cf_rbank[58], cf_rbank[48]}), .oen_bbank(padeb_b[56:0]),
     .cf_bbank({cf_bbank[730], cf_bbank[720], cf_bbank[706],
     cf_bbank[696], cf_bbank[682], cf_bbank[672], cf_bbank[648],
     cf_bbank[634], cf_bbank[624], cf_bbank[610], cf_bbank[600],
     cf_bbank[586], cf_bbank[576], cf_bbank[562], cf_bbank[552],
     cf_bbank[538], cf_bbank[528], cf_bbank[514], cf_bbank[504],
     cf_bbank[490], cf_bbank[480], cf_bbank[466], cf_bbank[456],
     cf_bbank[442], cf_bbank[432], cf_bbank[394], cf_bbank[384],
     cf_bbank[370], cf_bbank[360], cf_bbank[346], cf_bbank[336],
     cf_bbank[322], cf_bbank[312], cf_bbank[298], cf_bbank[288],
     cf_bbank[274], cf_bbank[264], cf_bbank[250], cf_bbank[240],
     cf_bbank[226], cf_bbank[216], cf_bbank[202], cf_bbank[192],
     cf_bbank[178], cf_bbank[168], cf_bbank[154], cf_bbank[144],
     cf_bbank[130], cf_bbank[120], cf_bbank[106], cf_bbank[96],
     cf_bbank[82], cf_bbank[72], cf_bbank[58], cf_bbank[48],
     cf_bbank[34], cf_bbank[24]}),
     .spi_ss_in_bbank(spi_ss_in_bbank[61:56]), .j_tck(j_tck),
     .fabric_out_32_00(fabric_out_32_00),
     .fabric_out_33_02(fabric_out_33_02),
     .fabric_out_33_01(fabric_out_33_01),
     .en_8bconfig_b(en_8bconfig_b), .trstb(trstb), .tms(tms),
     .tdi(tdi), .tck(tck), .spi_ss_in_r(spi_ss_in_r[11:5]),
     .out_tbank(out_tbank[59:0]), .out_rbank(out_rbank[54:0]),
     .out_lbank(out_lbank[49:0]), .out_bbank(pado_b[56:0]),
     .oen_tbank(oen_tbank[59:0]), .oen_rbank(oeb_rbank[54:0]),
     .oen_lbank(oen_lbank[49:0]), .fromsdo(fromsdo),
     .creset_b(creset_b), .bm_sdo_o(bm_sdo_o[3:0]),
     .VREFSSTL(VREFSSTL), .wl_r(wl_r[543:0]), .wl_l(wl_l[543:0]),
     .vdd_cntl_r(vdd_cntl_r[543:0]), .vdd_cntl_l(vdd_cntl_l[543:0]),
     .update0(net163), .tdo(tdo), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .spi_clk_out(spi_clk_out), .shift0(net165),
     .reset_r(reset_r[543:0]), .reset_l(reset_l[543:0]),
     .psdo(psdo[7:1]), .pgate_r(pgate_r[543:0]),
     .pgate_l(pgate_l[543:0]), .mode0(net170), .md_spi_b(md_spi_b),
     .last_rsr(last_rsr[3:0]),
     .jtag_rowtest_mode_rowu3_b(jtag_rowtest_mode_rowu3_b),
     .jtag_rowtest_mode_rowu2_b(jtag_rowtest_mode_rowu2_b),
     .jtag_rowtest_mode_rowu1_b(jtag_rowtest_mode_rowu1_b),
     .jtag_rowtest_mode_rowu0_b(jtag_rowtest_mode_rowu0_b),
     .j_tdi(net166), .in_tbank(in_tbank[59:0]),
     .in_rbank(in_rbank[54:0]), .in_lbank(in_lbank[49:0]),
     .in_bbank(padin_b[56:0]), .hiz_b0(net171), .gsr(gsr),
     .gint_hz(gint_hz), .end_of_startup(end_of_startup),
     .bs_en0(net172), .bm_wdummymux_en_i(bm_wdummymux_en_i),
     .bm_sweb_i(bm_sweb_i), .bm_sreb_i(bm_sreb_i),
     .bm_sdi_i(bm_sdi_i[3:0]), .bm_sclkrw_i(bm_sclkrw_i),
     .bm_sclk_i(bm_sclk_i), .bm_sa_i(bm_sa_i[7:0]),
     .bm_rcapmux_en_i(bm_rcapmux_en_i), .bm_init_i(bm_init_i),
     .bm_banksel_i(bm_banksel_i[3:0]), .uio_tbank(uio_tbank[59:0]),
     .uio_rbank(uio_rbank[54:0]), .uio_lbank(uio_lbank[49:0]),
     .uio_bbank(uio_bbank[56:0]), .cdone(cdone),
     .bl_top(bl_top[1743:0]), .bl_bot(bl_bot[1743:0]),
     .cf_tbank({cf_tbank[730], cf_tbank[720], cf_tbank[706],
     cf_tbank[696], cf_tbank[682], cf_tbank[672], cf_tbank[658],
     cf_tbank[648], cf_tbank[634], cf_tbank[624], cf_tbank[610],
     cf_tbank[600], cf_tbank[586], cf_tbank[576], cf_tbank[562],
     cf_tbank[552], cf_tbank[538], cf_tbank[528], cf_tbank[514],
     cf_tbank[504], cf_tbank[490], cf_tbank[480], cf_tbank[466],
     cf_tbank[456], cf_tbank[442], cf_tbank[432], cf_tbank[418],
     cf_tbank[408], cf_tbank[394], cf_tbank[384], cf_tbank[370],
     cf_tbank[360], cf_tbank[322], cf_tbank[312], cf_tbank[298],
     cf_tbank[288], cf_tbank[274], cf_tbank[264], cf_tbank[250],
     cf_tbank[240], cf_tbank[226], cf_tbank[216], cf_tbank[202],
     cf_tbank[192], cf_tbank[178], cf_tbank[168], cf_tbank[154],
     cf_tbank[144], cf_tbank[130], cf_tbank[120], cf_tbank[106],
     cf_tbank[96], cf_tbank[82], cf_tbank[72], cf_tbank[58],
     cf_tbank[48], cf_tbank[34], cf_tbank[24], cf_tbank[10],
     cf_tbank[0]}));
quad_x4_ice8 Iquad_x4 ( .ceb(ceb), .end_of_startup_bot_r({tievdd,
     end_of_startup, end_of_startup, end_of_startup, en_8bconfig_b,
     en_8bconfig_b, en_8bconfig_b, en_8bconfig_b, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .spi_ss_in_r(spi_ss_in_r[63:0]), .end_of_startup_r({tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     jtag_rowtest_mode_rowu3_b, jtag_rowtest_mode_rowu2_b, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     en_8bconfig_b, en_8bconfig_b, en_8bconfig_b, en_8bconfig_b,
     tievdd, tievdd}), .spiout_b({tiegnd, tiegnd, spi_ss_out_b,
     spi_clk_out, tiegnd, spi_sdo, tiegnd, tiegnd, tiegnd, psdo[2],
     psdo[3], psdo[4], psdo[5], psdo[6], psdo[7], tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .spi_ss_in_l(net190[0:31]), .spiout_r({tiegnd, last_rsr[3],
     last_rsr[2], tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, psdo[1], tiegnd, tiegnd, tiegnd, tiegnd}),
     .spi_ss_in_b(spi_ss_in_bbank[63:32]), .spiout_l({tiegnd,
     last_rsr[1], tiegnd, tiegnd, last_rsr[0], tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd}),
     .spioeb_l({tievdd, tiegnd, tievdd, tievdd, tiegnd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd}), .end_of_startup_top({tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd}), .spieb_b({tievdd, tievdd,
     md_spi_b, md_spi_b, tievdd, spi_sdo_oe_b, tievdd, tievdd, tievdd,
     tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tiegnd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .fabric_out_33_01(fabric_out_33_01),
     .fabric_out_32_00(fabric_out_32_00),
     .fabric_out_33_02(fabric_out_33_02), .bl_bot(bl_bot[1743:0]),
     .padin_b(padin_b[56:0]), .padeb_b(padeb_b[56:0]),
     .cf_b(cf_bbank[767:0]), .pado_b(pado_b[56:0]),
     .pgate_r(pgate_r[543:0]), .reset_b_r(reset_r[543:0]),
     .vdd_cntl_r(vdd_cntl_r[543:0]), .wl_r(wl_r[543:0]),
     .padeb_r(oeb_rbank[54:0]), .pado_r(out_rbank[54:0]),
     .cf_r(cf_rbank[767:0]), .padin_r(in_rbank[54:0]),
     .cf_l(cf_lbank[767:0]), .bl_top(bl_top[1743:0]),
     .pado_t(out_tbank[59:0]), .padeb_t(oen_tbank[59:0]),
     .padin_t(in_tbank[59:0]), .cf_t(cf_tbank[767:0]),
     .end_of_startup_l({tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, jtag_rowtest_mode_rowu1_b, tievdd,
     jtag_rowtest_mode_rowu0_b, tievdd, tievdd, tievdd, tievdd, tievdd,
     tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd, tievdd}),
     .pado_l(out_lbank[49:0]), .padin_l(in_lbank[49:0]),
     .reset_b_l(reset_l[543:0]), .vdd_cntl_l(vdd_cntl_l[543:0]),
     .wl_l(wl_l[543:0]), .padeb_l(oen_lbank[49:0]),
     .pgate_l(pgate_l[543:0]), .update(net163), .tclk(j_tck),
     .shift(net165), .sdi_pad(net166), .r(gsr), .purst(gsr),
     .prog(gint_hz), .mode(net170), .hiz_b(net171), .bs_en(net172),
     .bm_wdummymux_en_i(bm_wdummymux_en_i), .bm_sweb_i(bm_sweb_i),
     .bm_sreb_i(bm_sreb_i), .bm_sdi_i(bm_sdi_i[3:0]),
     .bm_sclkrw_i(bm_sclkrw_i), .bm_sclk_i(bm_sclk_i),
     .bm_sa_i(bm_sa_i[7:0]), .bm_rcapmux_en_i(bm_rcapmux_en_i),
     .bm_init_i(bm_init_i), .bm_banksel_i(bm_banksel_i[3:0]),
     .sdo_pad(fromsdo), .bm_sdo_o(bm_sdo_o[3:0]), .tievdd(tievdd),
     .tiegnd(tiegnd));
tielo4x I469 ( .tielo(tiegnd));
tiehi4x I468 ( .tiehi(tievdd));

endmodule
// Library - misc, Cell - ml_osc, View - schematic
// LAST TIME SAVED: Sep 30 17:24:55 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_osc ( clk_out, smc_osc_fsel, smc_oscen );
output  clk_out;

input  smc_oscen;

input [1:0]  smc_osc_fsel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:0]  sel_trim;



tielo I272 ( .tielo(net0104));
tielo I273 ( .tielo(net0188));
tiehi I275 ( .tiehi(net0205));
tiehi I219 ( .tiehi(net0106));
ml_osc_stage I254 ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_b_buf), .out(out_bot), .sel_trim(sel_trim[3:0]));
ml_osc_stage I255 ( .pbias(pbias), .oscen_b(oscen_b),
     .clkin(clkby2_buf), .out(out_top), .sel_trim(sel_trim[3:0]));
ml_osc_logic Iosc_logic ( .sel_trim(sel_trim[3:0]),
     .smc_oscen(smc_oscen), .smc_osc_fsel(smc_osc_fsel[1:0]),
     .clkin(clk_out));
ml_dff I174 ( .R(oscen_b), .D(clkby2_b), .CLK(clk_dffin),
     .QN(clkby2_b), .Q(clkby2));
nor3_hvt I256 ( .B(net079), .Y(net075), .A(net079), .C(net079));
nor3_hvt I218 ( .B(net083), .Y(net079), .A(net083), .C(net083));
nor3_hvt I217 ( .B(net0106), .Y(net083), .A(net0106), .C(net0106));
nand3_hvt I224 ( .Y(net088), .B(net0106), .C(net0106), .A(net0106));
nand3_hvt I230 ( .Y(net092), .B(net088), .C(net088), .A(net088));
nand3_hvt I231 ( .Y(net096), .B(net092), .C(net092), .A(net092));
rppolywo_m  R18 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net362), .PLUS(net356), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net356), .PLUS(pbias), .BULK(gnd_));
rppolywo_m  R7 ( .BULK(gnd_), .MINUS(net383), .PLUS(net366));
rppolywo_m  R2 ( .MINUS(net366), .PLUS(net362), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net437), .PLUS(net437), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net437), .PLUS(net383), .BULK(gnd_));
nand2_hvt I175 ( .A(out_bot), .Y(clk_dffin), .B(out_top));
inv_hvt I222 ( .A(clkby2), .Y(clkby2_b_buf));
inv_hvt I220 ( .A(clkby2_b), .Y(clkby2_buf));
inv_hvt I176 ( .A(clkby2_b), .Y(clk_out));
inv_hvt I248 ( .A(net0104), .Y(net0226));
inv_hvt I198 ( .A(smc_oscen), .Y(oscen_b));
nch_hvt  M45 ( .D(gnd_), .B(gnd_), .G(net0188), .S(gnd_));
nch_hvt  MN31 ( .D(net437), .B(gnd_), .G(smc_oscen), .S(gnd_));
nch_hvt  MN44 ( .D(pbias), .B(gnd_), .G(net0104), .S(net371));
pch_hvt  MP77 ( .D(net371), .B(vdd_), .G(net0226), .S(pbias));
pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(net0205), .S(vdd_));
pch_hvt  MP37 ( .D(pbias), .B(vdd_), .G(pbias), .S(vdd_));
pch_hvt  MP41 ( .D(pbias), .B(vdd_), .G(smc_oscen), .S(vdd_));

endmodule
// Library - misc, Cell - ml_osc_top, View - schematic
// LAST TIME SAVED: Oct 14 15:44:25 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_osc_top ( cnt_podt_out, smc_clk, crst_b, por_b, smc_osc_fsel,
     smc_oscoff_b, smc_podt_off, smc_podt_rst );
output  cnt_podt_out, smc_clk;

input  crst_b, por_b, smc_oscoff_b, smc_podt_off, smc_podt_rst;

input [1:0]  smc_osc_fsel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [10:0]  q_b;

wire  [10:0]  q;



tiehi I179 ( .tiehi(net076));
nor2_hvt I256 ( .A(rst_osc_b), .B(smc_oscoff_b), .Y(net066));
nor2_hvt I266 ( .A(clk_out), .B(smc_podt_off), .Y(net078));
nor2_hvt I257 ( .A(disable_osc), .B(net066), .Y(smc_oscen));
nor2_hvt I264 ( .A(smc_podt_rst), .B(net090), .Y(net054));
nor2_hvt I252 ( .A(cnt_rst), .B(smc_oscoff_b), .Y(net0124));
nand2_hvt I227 ( .A(smc_off_b), .B(rst_osc_b), .Y(disable_osc));
nand2_hvt I270 ( .A(crst_b), .Y(net064), .B(por_b));
ml_dff I230 ( .R(cnt_rst), .D(net076), .CLK(q_b[10]), .QN(net067),
     .Q(net063));
ml_dff I243 ( .R(rst_off_latch), .D(net0174), .CLK(clk_out_b),
     .QN(smc_off_b), .Q(net0152));
ml_dff I228_10_ ( .R(cnt_rst), .D(q_b[10]), .CLK(q[9]), .QN(q_b[10]),
     .Q(q[10]));
ml_dff I228_9_ ( .R(cnt_rst), .D(q_b[9]), .CLK(q[8]), .QN(q_b[9]),
     .Q(q[9]));
ml_dff I228_8_ ( .R(cnt_rst), .D(q_b[8]), .CLK(q[7]), .QN(q_b[8]),
     .Q(q[8]));
ml_dff I228_7_ ( .R(cnt_rst), .D(q_b[7]), .CLK(q[6]), .QN(q_b[7]),
     .Q(q[7]));
ml_dff I228_6_ ( .R(cnt_rst), .D(q_b[6]), .CLK(q[5]), .QN(q_b[6]),
     .Q(q[6]));
ml_dff I228_5_ ( .R(cnt_rst), .D(q_b[5]), .CLK(q[4]), .QN(q_b[5]),
     .Q(q[5]));
ml_dff I228_4_ ( .R(cnt_rst), .D(q_b[4]), .CLK(q[3]), .QN(q_b[4]),
     .Q(q[4]));
ml_dff I228_3_ ( .R(cnt_rst), .D(q_b[3]), .CLK(q[2]), .QN(q_b[3]),
     .Q(q[3]));
ml_dff I228_2_ ( .R(cnt_rst), .D(q_b[2]), .CLK(q[1]), .QN(q_b[2]),
     .Q(q[2]));
ml_dff I228_1_ ( .R(cnt_rst), .D(q_b[1]), .CLK(q[0]), .QN(q_b[1]),
     .Q(q[1]));
ml_dff I228_0_ ( .R(cnt_rst), .D(q_b[0]), .CLK(clk_in), .QN(q_b[0]),
     .Q(q[0]));
inv_hvt I233 ( .A(clk_out), .Y(clk_out_b));
inv_hvt I271 ( .A(net064), .Y(rst_osc_b));
inv_hvt I267 ( .A(net078), .Y(clk_in));
inv_hvt I262 ( .A(net067), .Y(cnt_podt_out));
inv_hvt I244 ( .A(smc_oscoff_b), .Y(net0174));
inv_hvt I265 ( .A(net054), .Y(cnt_rst));
inv_hvt I229 ( .A(rst_osc_b), .Y(net090));
inv_hvt I253 ( .A(net0124), .Y(rst_off_latch));
inv_hvt I232 ( .A(clk_out_b), .Y(smc_clk));
ml_osc Iml_osc ( .smc_osc_fsel(smc_osc_fsel[1:0]), .clk_out(clk_out),
     .smc_oscen(smc_oscen));

endmodule
// Library - leafcell, Cell - bram_bufferx16, View - schematic
// LAST TIME SAVED: Jun 25 13:49:31 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module bram_bufferx16 ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I0 ( .A(net07), .Y(net09));
inv_hvt I2 ( .A(in), .Y(net07));
inv_hvt I4 ( .A(net6), .Y(out));
inv_hvt I3 ( .A(net09), .Y(net6));

endmodule
// Library - xpmem, Cell - ml_cram_logic, View - schematic
// LAST TIME SAVED: Sep 28 20:58:40 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_cram_logic ( cram_pgateoff, cram_prec, cram_pullup_b,
     cram_rst, cram_vddoff, cram_wl_en, cram_write, smc_clk_out, por,
     smc_clk, smc_read, smc_rprec, smc_rpull_b, smc_rrst_pullwlen,
     smc_rwl_en, smc_seq_rst, smc_wcram_rst, smc_write, smc_wset_prec,
     smc_wset_precgnd, smc_wwlwrt_dis, smc_wwlwrt_en );
output  cram_pgateoff, cram_prec, cram_pullup_b, cram_rst, cram_vddoff,
     cram_wl_en, cram_write, smc_clk_out;

input  por, smc_clk, smc_read, smc_rprec, smc_rpull_b,
     smc_rrst_pullwlen, smc_rwl_en, smc_seq_rst, smc_wcram_rst,
     smc_write, smc_wset_prec, smc_wset_precgnd, smc_wwlwrt_dis,
     smc_wwlwrt_en;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I213 ( .A(net208), .Y(net177), .B(net248));
inv_hvt I370 ( .A(net273), .Y(rst_rpull_rwl));
inv_hvt I373 ( .A(cram_rst), .Y(net257));
inv_hvt I346 ( .A(net315), .Y(net220));
inv_hvt I263 ( .A(net269), .Y(net218));
inv_hvt I266 ( .A(cram_write_int), .Y(net216));
inv_hvt I286 ( .A(net359), .Y(net299));
inv_hvt I422 ( .A(smc_rwl_en), .Y(net212));
inv_hvt I323 ( .A(net282), .Y(net210));
inv_hvt I378 ( .A(net276), .Y(net248));
inv_hvt I333 ( .A(net279), .Y(net208));
inv_hvt I324 ( .A(net210), .Y(cram_pgateoff));
inv_hvt I403 ( .A(net285), .Y(net204));
inv_hvt I292 ( .A(net200), .Y(cram_prec));
inv_hvt I267 ( .A(net303), .Y(net200));
inv_hvt I224 ( .A(net291), .Y(reset_logic));
inv_hvt I401 ( .A(net294), .Y(net196));
inv_hvt I381 ( .A(net309), .Y(net194));
inv_hvt I268 ( .A(net257), .Y(net253));
inv_hvt I293 ( .A(net236), .Y(cram_vddoff));
inv_hvt I269 ( .A(net255), .Y(net251));
inv_hvt I330 ( .A(net265), .Y(net190));
inv_hvt I374 ( .A(net253), .Y(net255));
inv_hvt I294 ( .A(cram_rst_int_b), .Y(cram_rst));
inv_hvt I375 ( .A(net252), .Y(cram_rst_dly));
inv_hvt I421 ( .A(net394), .Y(net186));
inv_hvt I249 ( .A(net262), .Y(net184));
inv_hvt I250 ( .A(net184), .Y(cram_pullup_b));
inv_hvt I359 ( .A(net179), .Y(net180));
inv_hvt I376 ( .A(net251), .Y(net252));
inv_hvt I336 ( .A(smc_clk), .Y(sm_clk_b));
inv_hvt I367 ( .A(net306), .Y(dis_pgatewrt));
inv_hvt I281 ( .A(net399), .Y(net226));
inv_hvt I399 ( .A(net300), .Y(net240));
inv_hvt I290 ( .A(net218), .Y(cram_wl_en));
inv_hvt I425 ( .A(net299), .Y(net262));
inv_hvt I337 ( .A(sm_clk_b), .Y(smc_clk_out));
inv_hvt I256 ( .A(net379), .Y(cram_write_int));
inv_hvt I291 ( .A(net216), .Y(cram_write));
inv_hvt I415 ( .A(net312), .Y(net260));
inv_hvt I312 ( .A(net177), .Y(net228));
inv_hvt I270 ( .A(net228), .Y(net236));
inv_hvt I271 ( .A(net226), .Y(cram_rst_int_b));
mux2_hvt I161 ( .in1(cram_write_int), .in0(net186), .out(net269),
     .sel(net208));
mux2_hvt I295 ( .in1(net194), .in0(net220), .out(net265),
     .sel(net208));
nor2_hvt I402 ( .A(net283), .B(smc_wset_precgnd), .Y(net285));
nor2_hvt I329 ( .A(net190), .B(smc_seq_rst), .Y(net303));
nor2_hvt I398 ( .A(smc_rpull_b), .B(net299), .Y(net300));
nor2_hvt I393 ( .A(cram_rst_dly), .B(reset_logic), .Y(net179));
nor2_hvt I364 ( .A(net389), .B(smc_seq_rst), .Y(net282));
nor2_hvt I400 ( .A(net292), .B(smc_wset_prec), .Y(net294));
nor2_hvt I366 ( .A(reset_logic), .B(net370), .Y(net306));
nor2_hvt I223 ( .A(net318), .B(por), .Y(net291));
nor2_hvt I390 ( .A(smc_write), .B(smc_seq_rst), .Y(net279));
nor2_hvt I392 ( .A(net283), .B(cram_rst), .Y(net276));
nor2_hvt I389 ( .A(net375), .B(reset_logic), .Y(net273));
nor2_hvt I385 ( .A(smc_rprec), .B(net287), .Y(net315));
nor2_hvt I414 ( .A(net310), .B(smc_wwlwrt_en), .Y(net312));
nor2_hvt I391 ( .A(net292), .B(cram_rst), .Y(net309));
nor3_hvt I220 ( .B(net322), .Y(net326), .A(net322), .C(net322));
nor3_hvt I217 ( .B(net401), .Y(net330), .A(net401), .C(net401));
nor3_hvt I386 ( .B(smc_seq_rst), .Y(net318), .A(smc_write),
     .C(smc_read));
nor3_hvt I218 ( .B(net330), .Y(net322), .A(net330), .C(net330));
nor3_hvt I387 ( .B(smc_rwl_en), .Y(net287), .A(net315),
     .C(reset_logic));
nand3_hvt I230 ( .Y(net348), .B(net344), .C(net344), .A(net344));
nand3_hvt I231 ( .Y(net352), .B(net348), .C(net348), .A(net348));
nand3_hvt I426 ( .Y(net344), .B(net401), .C(net401), .A(net401));
ml_dff_schematic I411 ( .R(reset_logic), .D(smc_wwlwrt_dis),
     .CLK(smc_clk), .QN(net369), .Q(net370));
ml_dff_schematic I408 ( .R(rst_rpull_rwl), .D(net401), .CLK(net212),
     .QN(net394), .Q(net395));
ml_dff_schematic I405 ( .R(dis_pgatewrt), .D(net401),
     .CLK(cram_rst_int_b), .QN(net389), .Q(net390));
ml_dff_schematic I412 ( .R(net180), .D(net196), .CLK(smc_clk_out),
     .QN(net337), .Q(net292));
ml_dff_schematic I410 ( .R(dis_pgatewrt), .D(net260),
     .CLK(smc_clk_out), .QN(net379), .Q(net310));
ml_dff_schematic I108 ( .R(reset_logic), .D(smc_rrst_pullwlen),
     .CLK(smc_clk_out), .QN(net343), .Q(net375));
ml_dff_schematic I413 ( .R(net180), .D(net204), .CLK(smc_clk_out),
     .QN(net333), .Q(net283));
ml_dff_schematic I407 ( .R(rst_rpull_rwl), .D(net240),
     .CLK(smc_clk_out), .QN(net359), .Q(net360));
ml_dff_schematic I406 ( .R(reset_logic), .D(smc_wcram_rst),
     .CLK(smc_clk_out), .QN(net399), .Q(net400));
tiehi I427 ( .tiehi(net401));

endmodule
// Library - chip, Cell - CHIP_route_right_ice8f, View - schematic
// LAST TIME SAVED: Sep 24 09:02:30 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module CHIP_route_right_ice8f ( bm_banksel_i, bm_init_i,
     bm_rcapmux_en_i, bm_sa_i, bm_sclk_i, bm_sclkrw_i, bm_sdi_i,
     bm_sreb_i, bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bldld, cm_banksel_bltrd1_3_,
     cm_clk_blbrd, cm_clk_bltrd1, cm_sdi_u0, cm_sdi_u1, cm_sdi_u2d,
     cm_sdi_u3d2, core_por_b0, core_por_b1, core_por_b_rowu2,
     core_por_b_rowu3, core_por_bb, cram_pgateoff, cram_prec,
     cram_prec_bltrd1, cram_pullup_b, cram_pullup_b_bltrd1, cram_rst,
     cram_vddoff, cram_wl_en, cram_write, cram_write_bltrd1,
     data_muxsel1_blbrd, data_muxsel1_bltrd1, data_muxsel_blbrd,
     data_muxsel_bltrd1, .en_8bcibfig_b_bltrd1(en_8bconfig_b_bltrd1),
     en_8bconfig_b, en_8bconfig_b_blbrd, end_of_startup, gint_hz, gsr,
     hiz_b0, j_rst_b, j_tck, j_tdi, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, last_rsr, md_spi_b, mode0,
     nvcm_spi_sdi, nvcm_spi_ss_b, pgate_r, psdo, reset_b_r, row_test0,
     rst_b, sdo_enable, shift0, smc_load_nvcm_bstream, smc_row_inc,
     smc_rsr_rst, smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1,
     smc_write0, spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out_b,
     totdopad, update0, vdd_cntl_r, wl_r, bm_sdo_o, bp0, cdone_in,
     cf_r, cm_sdo_u0d1, cm_sdo_u1d3, cm_sdo_u2d1, cm_sdo_u3,
     crst_filterout, fabric_out_32_00, fabric_out_33_01,
     fabric_out_33_02, fromsdo, idcode_msb20bits, last_rsr3,
     monitor_celld4, nvcm_boot, nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo,
     nvcm_spi_sdo_oe_b, smc_core_por_bottom1, smc_core_por_bottom2,
     spi_ss_in_bbank, spi_ss_in_r, tck_pad, tdi_pad, tms_pad, trst_pad,
     vddio_rightbank );
output  bm_init_i, bm_rcapmux_en_i, bm_sclk_i, bm_sclkrw_i, bm_sreb_i,
     bm_sweb_i, bm_wdummymux_en_i, bs_en0, cdone_out, ceb0,
     cm_banksel_blbrd_2_, cm_banksel_bltrd1_3_, cm_clk_blbrd,
     cm_clk_bltrd1, core_por_b0, core_por_b1, core_por_b_rowu2,
     core_por_b_rowu3, core_por_bb, cram_pgateoff, cram_prec,
     cram_prec_bltrd1, cram_pullup_b, cram_pullup_b_bltrd1, cram_rst,
     cram_vddoff, cram_wl_en, cram_write, cram_write_bltrd1,
     data_muxsel1_blbrd, data_muxsel1_bltrd1, data_muxsel_blbrd,
     data_muxsel_bltrd1, en_8bconfig_b_bltrd1, en_8bconfig_b,
     en_8bconfig_b_blbrd, end_of_startup, gint_hz, gsr, hiz_b0,
     j_rst_b, j_tck, j_tdi, jtag_rowtest_mode_rowu2_b,
     jtag_rowtest_mode_rowu3_b, md_spi_b, mode0, nvcm_spi_sdi,
     nvcm_spi_ss_b, row_test0, rst_b, sdo_enable, shift0,
     smc_load_nvcm_bstream, smc_row_inc, smc_rsr_rst,
     smc_wdis_dclk_blbrd, smc_wdis_dclk_bltrd1, smc_write0,
     spi_clk_out, spi_sdo, spi_sdo_oe_b, spi_ss_out_b, totdopad,
     update0;

input  bp0, cdone_in, crst_filterout, fabric_out_32_00,
     fabric_out_33_01, fabric_out_33_02, fromsdo, last_rsr3, nvcm_boot,
     nvcm_rdy, nvcm_relextspi, nvcm_spi_sdo, nvcm_spi_sdo_oe_b,
     smc_core_por_bottom1, smc_core_por_bottom2, tck_pad, tdi_pad,
     tms_pad, trst_pad, vddio_rightbank;

output [3:0]  bm_sdi_i;
output [1:0]  cm_sdi_u1;
output [1:0]  cm_banksel_bldld;
output [1:0]  cm_sdi_u0;
output [7:1]  psdo;
output [7:0]  bm_sa_i;
output [543:0]  wl_r;
output [1:0]  cm_sdi_u3d2;
output [1:0]  cm_sdi_u2d;
output [3:0]  bm_banksel_i;
output [1:0]  last_rsr;
output [543:0]  vdd_cntl_r;
output [543:0]  pgate_r;
output [543:0]  reset_b_r;

input [3:0]  bm_sdo_o;
input [7:1]  spi_ss_in_r;
input [19:0]  idcode_msb20bits;
input [1:0]  cm_sdo_u1d3;
input [1:0]  monitor_celld4;
input [1:0]  cm_sdo_u3;
input [1:0]  cm_sdo_u0d1;
input [4:0]  spi_ss_in_bbank;
input [1:0]  cf_r;
input [1:0]  cm_sdo_u2d1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [3:3]  cm_banksel_bltrd;

wire  [1:0]  smc_osco_fsel;

wire  [0:1]  net0206;

wire  [1:0]  u1_in;

wire  [0:1]  net0207;

wire  [1:0]  u0_in;

wire  [1:0]  cm_sdi_u3d0;

wire  [3:3]  cm_banksel_bltrd0;

wire  [1:0]  cm_sdo_u3d;

wire  [3:3]  monitor_celld1;

wire  [1:0]  cm_sdi_u3;

wire  [3:3]  monitor_celld2;

wire  [3:2]  monitor_celldd;

wire  [1:0]  cm_sdo_u3d1;

wire  [1:0]  dff_out_top;

wire  [1:0]  dff_out_bot;

wire  [2:3]  monitor_celld;

wire  [1:0]  cm_sdo_u3dd;

wire  [3:0]  cm_banksel;

wire  [1:0]  cm_sdi_u2;

wire  [1:0]  cm_sdi_u3d;

wire  [1:0]  cm_sdo_u3d0;

wire  [7:1]  spi_ss_in_rd;



tielo I474_1_ ( .tielo(net0207[0]));
tielo I474_0_ ( .tielo(net0207[1]));
tielo I475_1_ ( .tielo(net0206[0]));
tielo I475_0_ ( .tielo(net0206[1]));
sg_dffbuf_modified I286_1_ ( .r(net0207[0]), .d(cm_sdo_u3d[1]),
     .clk(net507), .dffout(dff_out_top[1]));
sg_dffbuf_modified I286_0_ ( .r(net0207[1]), .d(cm_sdo_u3d[0]),
     .clk(net507), .dffout(dff_out_top[0]));
sg_dffbuf_modified I453_1_ ( .r(net0206[0]), .d(cm_sdo_u3dd[1]),
     .clk(net509), .dffout(dff_out_bot[1]));
sg_dffbuf_modified I453_0_ ( .r(net0206[1]), .d(cm_sdo_u3dd[0]),
     .clk(net509), .dffout(dff_out_bot[0]));
// smc_and_jtag_ice8f I_smc_and_jtag (
smc_and_jtag I_smc_and_jtag (
     .idcode_msb20bits(idcode_msb20bits[19:0]),
     .nvcm_spi_sdo_oe_b(nvcm_spi_sdo_oe_b),
     .nvcm_spi_sdo(nvcm_spi_sdo), .nvcm_relextspi(nvcm_relextspi),
     .nvcm_rdy(nvcm_rdy), .nvcm_boot(nvcm_boot), .bp0(bp0),
     .smc_load_nvcm_bstream(smc_load_nvcm_bstream), .rst_b(rst_b),
     .nvcm_spi_ss_b(nvcm_spi_ss_b), .nvcm_spi_sdi(nvcm_spi_sdi),
     .j_shift0(shift0), .j_ceb0(ceb0), .warmboot_sel({fabric_out_33_02,
     fabric_out_33_01}), .trst_pad(trst_pad), .tms_pad(tms_pad),
     .tdi_pad(tdi_pad), .tck_pad(tck_pad),
     .spi_ss_in_b(spi_ss_in_bbank[4]), .spi_sdi(spi_ss_in_bbank[2]),
     .spi_clk_in(spi_ss_in_bbank[3]), .psdi(spi_ss_in_rd[7:1]),
     .por_b(smc_por_b0), .osc_clk(osc_clk), .creset_b(crst_filterout),
     .coldboot_sel(spi_ss_in_bbank[1:0]), .cnt_podt_out(cnt_podt_out),
     .cm_sdo_u3(cm_sdo_u3d1[1:0]), .cm_sdo_u2(cm_sdo_u2d1[1:0]),
     .cm_sdo_u1(cm_sdo_u1d3[1:0]), .cm_sdo_u0(cm_sdo_u0d1[1:0]),
     .cm_monitor_cell({monitor_celldd[3:2], monitor_celld4[1:0]}),
     .cm_last_rsr(last_rsr3), .cdone_in(cdone_in),
     .bschain_sdo(fromsdo), .boot(fabric_out_32_00),
     .bm_bank_sdo(bm_sdo_o[3:0]), .tdo_pad(totdopad),
     .tdo_oe_pad(sdo_enable), .spi_ss_out_b(spi_ss_out_b),
     .spi_sdo_oe_b(spi_sdo_oe_b), .spi_sdo(spi_sdo),
     .spi_clk_out(spi_clk_out), .smc_wwlwrt_en(smc_wwlwrt_en),
     .smc_wwlwrt_dis(smc_wwlwrt_dis),
     .smc_wset_precgnd(smc_wset_precgnd),
     .smc_wset_prec(smc_wset_prec), .smc_write(smc_write0),
     .smc_wdis_dclk(smc_wdis_dclk), .smc_wcram_rst(smc_wcram_rst),
     .smc_seq_rst(smc_seq_rst), .smc_rwl_en(smc_rwl_en),
     .smc_rsr_rst(net257), .smc_rrst_pullwlen(smc_rrst_pullwlen),
     .smc_rpull_b(smc_rpull_b), .smc_rprec(smc_rprec),
     .smc_row_inc(net261), .cm_clk(cm_clk), .smc_read(net263),
     .smc_podt_rst(smc_podt_rst), .smc_podt_off(smc_podt_off),
     .smc_oscoff_b(smc_oscoff_b), .smc_osc_fsel(smc_osco_fsel[1:0]),
     .psdo(psdo[7:1]), .md_spi_b(md_spi_b), .j_upd_dr(update0),
     .j_tdi(j_tdi), .j_tck(j_tck), .j_sft_dr(shiftfromsmc),
     .j_rst_b(j_rst_b), .j_row_test(row_test0), .j_mode(mode0),
     .j_hiz_b(hiz_b0), .gsr(gsr), .gint_hz(gint_hz),
     .end_of_startup(end_of_startup), .en_8bconfig_b(en_8bconfig_b),
     .data_muxsel1(data_muxsel1), .data_muxsel(data_muxsel),
     .cm_sdi_u3(cm_sdi_u3[1:0]), .cm_sdi_u2(cm_sdi_u2[1:0]),
     .cm_sdi_u1(u1_in[1:0]), .cm_sdi_u0(u0_in[1:0]),
     .cm_banksel(cm_banksel[3:0]), .cdone_out(cdone_out),
     .bs_en(bs_en0), .bm_wdummymux_en(bm_wdummymux_en_i),
     .bm_sreb(bm_sreb_i), .bm_sclkrw(bm_sclkrw_i),
     .bm_sa(bm_sa_i[7:0]), .bm_rcapmux_en(bm_rcapmux_en_i),
     .bm_init(bm_init_i), .bm_clk(bm_sclk_i),
     .bm_banksel(bm_banksel_i[3:0]), .bm_bank_sdi(bm_sdi_i[3:0]),
     .bm_sweb(bm_sweb_i));
ml_rowdrv_bank10k Irowur ( .vddctrl({vdd_cntl_r[272], vdd_cntl_r[273],
     vdd_cntl_r[274], vdd_cntl_r[275], vdd_cntl_r[276],
     vdd_cntl_r[277], vdd_cntl_r[278], vdd_cntl_r[279],
     vdd_cntl_r[280], vdd_cntl_r[281], vdd_cntl_r[282],
     vdd_cntl_r[283], vdd_cntl_r[284], vdd_cntl_r[285],
     vdd_cntl_r[286], vdd_cntl_r[287], vdd_cntl_r[288],
     vdd_cntl_r[289], vdd_cntl_r[290], vdd_cntl_r[291],
     vdd_cntl_r[292], vdd_cntl_r[293], vdd_cntl_r[294],
     vdd_cntl_r[295], vdd_cntl_r[296], vdd_cntl_r[297],
     vdd_cntl_r[298], vdd_cntl_r[299], vdd_cntl_r[300],
     vdd_cntl_r[301], vdd_cntl_r[302], vdd_cntl_r[303],
     vdd_cntl_r[304], vdd_cntl_r[305], vdd_cntl_r[306],
     vdd_cntl_r[307], vdd_cntl_r[308], vdd_cntl_r[309],
     vdd_cntl_r[310], vdd_cntl_r[311], vdd_cntl_r[312],
     vdd_cntl_r[313], vdd_cntl_r[314], vdd_cntl_r[315],
     vdd_cntl_r[316], vdd_cntl_r[317], vdd_cntl_r[318],
     vdd_cntl_r[319], vdd_cntl_r[320], vdd_cntl_r[321],
     vdd_cntl_r[322], vdd_cntl_r[323], vdd_cntl_r[324],
     vdd_cntl_r[325], vdd_cntl_r[326], vdd_cntl_r[327],
     vdd_cntl_r[328], vdd_cntl_r[329], vdd_cntl_r[330],
     vdd_cntl_r[331], vdd_cntl_r[332], vdd_cntl_r[333],
     vdd_cntl_r[334], vdd_cntl_r[335], vdd_cntl_r[336],
     vdd_cntl_r[337], vdd_cntl_r[338], vdd_cntl_r[339],
     vdd_cntl_r[340], vdd_cntl_r[341], vdd_cntl_r[342],
     vdd_cntl_r[343], vdd_cntl_r[344], vdd_cntl_r[345],
     vdd_cntl_r[346], vdd_cntl_r[347], vdd_cntl_r[348],
     vdd_cntl_r[349], vdd_cntl_r[350], vdd_cntl_r[351],
     vdd_cntl_r[352], vdd_cntl_r[353], vdd_cntl_r[354],
     vdd_cntl_r[355], vdd_cntl_r[356], vdd_cntl_r[357],
     vdd_cntl_r[358], vdd_cntl_r[359], vdd_cntl_r[360],
     vdd_cntl_r[361], vdd_cntl_r[362], vdd_cntl_r[363],
     vdd_cntl_r[364], vdd_cntl_r[365], vdd_cntl_r[366],
     vdd_cntl_r[367], vdd_cntl_r[368], vdd_cntl_r[369],
     vdd_cntl_r[370], vdd_cntl_r[371], vdd_cntl_r[372],
     vdd_cntl_r[373], vdd_cntl_r[374], vdd_cntl_r[375],
     vdd_cntl_r[376], vdd_cntl_r[377], vdd_cntl_r[378],
     vdd_cntl_r[379], vdd_cntl_r[380], vdd_cntl_r[381],
     vdd_cntl_r[382], vdd_cntl_r[383], vdd_cntl_r[384],
     vdd_cntl_r[385], vdd_cntl_r[386], vdd_cntl_r[387],
     vdd_cntl_r[388], vdd_cntl_r[389], vdd_cntl_r[390],
     vdd_cntl_r[391], vdd_cntl_r[392], vdd_cntl_r[393],
     vdd_cntl_r[394], vdd_cntl_r[395], vdd_cntl_r[396],
     vdd_cntl_r[397], vdd_cntl_r[398], vdd_cntl_r[399],
     vdd_cntl_r[400], vdd_cntl_r[401], vdd_cntl_r[402],
     vdd_cntl_r[403], vdd_cntl_r[404], vdd_cntl_r[405],
     vdd_cntl_r[406], vdd_cntl_r[407], vdd_cntl_r[408],
     vdd_cntl_r[409], vdd_cntl_r[410], vdd_cntl_r[411],
     vdd_cntl_r[412], vdd_cntl_r[413], vdd_cntl_r[414],
     vdd_cntl_r[415], vdd_cntl_r[416], vdd_cntl_r[417],
     vdd_cntl_r[418], vdd_cntl_r[419], vdd_cntl_r[420],
     vdd_cntl_r[421], vdd_cntl_r[422], vdd_cntl_r[423],
     vdd_cntl_r[424], vdd_cntl_r[425], vdd_cntl_r[426],
     vdd_cntl_r[427], vdd_cntl_r[428], vdd_cntl_r[429],
     vdd_cntl_r[430], vdd_cntl_r[431], vdd_cntl_r[432],
     vdd_cntl_r[433], vdd_cntl_r[434], vdd_cntl_r[435],
     vdd_cntl_r[436], vdd_cntl_r[437], vdd_cntl_r[438],
     vdd_cntl_r[439], vdd_cntl_r[440], vdd_cntl_r[441],
     vdd_cntl_r[442], vdd_cntl_r[443], vdd_cntl_r[444],
     vdd_cntl_r[445], vdd_cntl_r[446], vdd_cntl_r[447],
     vdd_cntl_r[448], vdd_cntl_r[449], vdd_cntl_r[450],
     vdd_cntl_r[451], vdd_cntl_r[452], vdd_cntl_r[453],
     vdd_cntl_r[454], vdd_cntl_r[455], vdd_cntl_r[456],
     vdd_cntl_r[457], vdd_cntl_r[458], vdd_cntl_r[459],
     vdd_cntl_r[460], vdd_cntl_r[461], vdd_cntl_r[462],
     vdd_cntl_r[463], vdd_cntl_r[464], vdd_cntl_r[465],
     vdd_cntl_r[466], vdd_cntl_r[467], vdd_cntl_r[468],
     vdd_cntl_r[469], vdd_cntl_r[470], vdd_cntl_r[471],
     vdd_cntl_r[472], vdd_cntl_r[473], vdd_cntl_r[474],
     vdd_cntl_r[475], vdd_cntl_r[476], vdd_cntl_r[477],
     vdd_cntl_r[478], vdd_cntl_r[479], vdd_cntl_r[480],
     vdd_cntl_r[481], vdd_cntl_r[482], vdd_cntl_r[483],
     vdd_cntl_r[484], vdd_cntl_r[485], vdd_cntl_r[486],
     vdd_cntl_r[487], vdd_cntl_r[488], vdd_cntl_r[489],
     vdd_cntl_r[490], vdd_cntl_r[491], vdd_cntl_r[492],
     vdd_cntl_r[493], vdd_cntl_r[494], vdd_cntl_r[495],
     vdd_cntl_r[496], vdd_cntl_r[497], vdd_cntl_r[498],
     vdd_cntl_r[499], vdd_cntl_r[500], vdd_cntl_r[501],
     vdd_cntl_r[502], vdd_cntl_r[503], vdd_cntl_r[504],
     vdd_cntl_r[505], vdd_cntl_r[506], vdd_cntl_r[507],
     vdd_cntl_r[508], vdd_cntl_r[509], vdd_cntl_r[510],
     vdd_cntl_r[511], vdd_cntl_r[512], vdd_cntl_r[513],
     vdd_cntl_r[514], vdd_cntl_r[515], vdd_cntl_r[516],
     vdd_cntl_r[517], vdd_cntl_r[518], vdd_cntl_r[519],
     vdd_cntl_r[520], vdd_cntl_r[521], vdd_cntl_r[522],
     vdd_cntl_r[523], vdd_cntl_r[524], vdd_cntl_r[525],
     vdd_cntl_r[526], vdd_cntl_r[527], vdd_cntl_r[528],
     vdd_cntl_r[529], vdd_cntl_r[530], vdd_cntl_r[531],
     vdd_cntl_r[532], vdd_cntl_r[533], vdd_cntl_r[534],
     vdd_cntl_r[535], vdd_cntl_r[536], vdd_cntl_r[537],
     vdd_cntl_r[538], vdd_cntl_r[539], vdd_cntl_r[540],
     vdd_cntl_r[541], vdd_cntl_r[542], vdd_cntl_r[543]}),
     .pgate({pgate_r[272], pgate_r[273], pgate_r[274], pgate_r[275],
     pgate_r[276], pgate_r[277], pgate_r[278], pgate_r[279],
     pgate_r[280], pgate_r[281], pgate_r[282], pgate_r[283],
     pgate_r[284], pgate_r[285], pgate_r[286], pgate_r[287],
     pgate_r[288], pgate_r[289], pgate_r[290], pgate_r[291],
     pgate_r[292], pgate_r[293], pgate_r[294], pgate_r[295],
     pgate_r[296], pgate_r[297], pgate_r[298], pgate_r[299],
     pgate_r[300], pgate_r[301], pgate_r[302], pgate_r[303],
     pgate_r[304], pgate_r[305], pgate_r[306], pgate_r[307],
     pgate_r[308], pgate_r[309], pgate_r[310], pgate_r[311],
     pgate_r[312], pgate_r[313], pgate_r[314], pgate_r[315],
     pgate_r[316], pgate_r[317], pgate_r[318], pgate_r[319],
     pgate_r[320], pgate_r[321], pgate_r[322], pgate_r[323],
     pgate_r[324], pgate_r[325], pgate_r[326], pgate_r[327],
     pgate_r[328], pgate_r[329], pgate_r[330], pgate_r[331],
     pgate_r[332], pgate_r[333], pgate_r[334], pgate_r[335],
     pgate_r[336], pgate_r[337], pgate_r[338], pgate_r[339],
     pgate_r[340], pgate_r[341], pgate_r[342], pgate_r[343],
     pgate_r[344], pgate_r[345], pgate_r[346], pgate_r[347],
     pgate_r[348], pgate_r[349], pgate_r[350], pgate_r[351],
     pgate_r[352], pgate_r[353], pgate_r[354], pgate_r[355],
     pgate_r[356], pgate_r[357], pgate_r[358], pgate_r[359],
     pgate_r[360], pgate_r[361], pgate_r[362], pgate_r[363],
     pgate_r[364], pgate_r[365], pgate_r[366], pgate_r[367],
     pgate_r[368], pgate_r[369], pgate_r[370], pgate_r[371],
     pgate_r[372], pgate_r[373], pgate_r[374], pgate_r[375],
     pgate_r[376], pgate_r[377], pgate_r[378], pgate_r[379],
     pgate_r[380], pgate_r[381], pgate_r[382], pgate_r[383],
     pgate_r[384], pgate_r[385], pgate_r[386], pgate_r[387],
     pgate_r[388], pgate_r[389], pgate_r[390], pgate_r[391],
     pgate_r[392], pgate_r[393], pgate_r[394], pgate_r[395],
     pgate_r[396], pgate_r[397], pgate_r[398], pgate_r[399],
     pgate_r[400], pgate_r[401], pgate_r[402], pgate_r[403],
     pgate_r[404], pgate_r[405], pgate_r[406], pgate_r[407],
     pgate_r[408], pgate_r[409], pgate_r[410], pgate_r[411],
     pgate_r[412], pgate_r[413], pgate_r[414], pgate_r[415],
     pgate_r[416], pgate_r[417], pgate_r[418], pgate_r[419],
     pgate_r[420], pgate_r[421], pgate_r[422], pgate_r[423],
     pgate_r[424], pgate_r[425], pgate_r[426], pgate_r[427],
     pgate_r[428], pgate_r[429], pgate_r[430], pgate_r[431],
     pgate_r[432], pgate_r[433], pgate_r[434], pgate_r[435],
     pgate_r[436], pgate_r[437], pgate_r[438], pgate_r[439],
     pgate_r[440], pgate_r[441], pgate_r[442], pgate_r[443],
     pgate_r[444], pgate_r[445], pgate_r[446], pgate_r[447],
     pgate_r[448], pgate_r[449], pgate_r[450], pgate_r[451],
     pgate_r[452], pgate_r[453], pgate_r[454], pgate_r[455],
     pgate_r[456], pgate_r[457], pgate_r[458], pgate_r[459],
     pgate_r[460], pgate_r[461], pgate_r[462], pgate_r[463],
     pgate_r[464], pgate_r[465], pgate_r[466], pgate_r[467],
     pgate_r[468], pgate_r[469], pgate_r[470], pgate_r[471],
     pgate_r[472], pgate_r[473], pgate_r[474], pgate_r[475],
     pgate_r[476], pgate_r[477], pgate_r[478], pgate_r[479],
     pgate_r[480], pgate_r[481], pgate_r[482], pgate_r[483],
     pgate_r[484], pgate_r[485], pgate_r[486], pgate_r[487],
     pgate_r[488], pgate_r[489], pgate_r[490], pgate_r[491],
     pgate_r[492], pgate_r[493], pgate_r[494], pgate_r[495],
     pgate_r[496], pgate_r[497], pgate_r[498], pgate_r[499],
     pgate_r[500], pgate_r[501], pgate_r[502], pgate_r[503],
     pgate_r[504], pgate_r[505], pgate_r[506], pgate_r[507],
     pgate_r[508], pgate_r[509], pgate_r[510], pgate_r[511],
     pgate_r[512], pgate_r[513], pgate_r[514], pgate_r[515],
     pgate_r[516], pgate_r[517], pgate_r[518], pgate_r[519],
     pgate_r[520], pgate_r[521], pgate_r[522], pgate_r[523],
     pgate_r[524], pgate_r[525], pgate_r[526], pgate_r[527],
     pgate_r[528], pgate_r[529], pgate_r[530], pgate_r[531],
     pgate_r[532], pgate_r[533], pgate_r[534], pgate_r[535],
     pgate_r[536], pgate_r[537], pgate_r[538], pgate_r[539],
     pgate_r[540], pgate_r[541], pgate_r[542], pgate_r[543]}),
     .reset({reset_b_r[272], reset_b_r[273], reset_b_r[274],
     reset_b_r[275], reset_b_r[276], reset_b_r[277], reset_b_r[278],
     reset_b_r[279], reset_b_r[280], reset_b_r[281], reset_b_r[282],
     reset_b_r[283], reset_b_r[284], reset_b_r[285], reset_b_r[286],
     reset_b_r[287], reset_b_r[288], reset_b_r[289], reset_b_r[290],
     reset_b_r[291], reset_b_r[292], reset_b_r[293], reset_b_r[294],
     reset_b_r[295], reset_b_r[296], reset_b_r[297], reset_b_r[298],
     reset_b_r[299], reset_b_r[300], reset_b_r[301], reset_b_r[302],
     reset_b_r[303], reset_b_r[304], reset_b_r[305], reset_b_r[306],
     reset_b_r[307], reset_b_r[308], reset_b_r[309], reset_b_r[310],
     reset_b_r[311], reset_b_r[312], reset_b_r[313], reset_b_r[314],
     reset_b_r[315], reset_b_r[316], reset_b_r[317], reset_b_r[318],
     reset_b_r[319], reset_b_r[320], reset_b_r[321], reset_b_r[322],
     reset_b_r[323], reset_b_r[324], reset_b_r[325], reset_b_r[326],
     reset_b_r[327], reset_b_r[328], reset_b_r[329], reset_b_r[330],
     reset_b_r[331], reset_b_r[332], reset_b_r[333], reset_b_r[334],
     reset_b_r[335], reset_b_r[336], reset_b_r[337], reset_b_r[338],
     reset_b_r[339], reset_b_r[340], reset_b_r[341], reset_b_r[342],
     reset_b_r[343], reset_b_r[344], reset_b_r[345], reset_b_r[346],
     reset_b_r[347], reset_b_r[348], reset_b_r[349], reset_b_r[350],
     reset_b_r[351], reset_b_r[352], reset_b_r[353], reset_b_r[354],
     reset_b_r[355], reset_b_r[356], reset_b_r[357], reset_b_r[358],
     reset_b_r[359], reset_b_r[360], reset_b_r[361], reset_b_r[362],
     reset_b_r[363], reset_b_r[364], reset_b_r[365], reset_b_r[366],
     reset_b_r[367], reset_b_r[368], reset_b_r[369], reset_b_r[370],
     reset_b_r[371], reset_b_r[372], reset_b_r[373], reset_b_r[374],
     reset_b_r[375], reset_b_r[376], reset_b_r[377], reset_b_r[378],
     reset_b_r[379], reset_b_r[380], reset_b_r[381], reset_b_r[382],
     reset_b_r[383], reset_b_r[384], reset_b_r[385], reset_b_r[386],
     reset_b_r[387], reset_b_r[388], reset_b_r[389], reset_b_r[390],
     reset_b_r[391], reset_b_r[392], reset_b_r[393], reset_b_r[394],
     reset_b_r[395], reset_b_r[396], reset_b_r[397], reset_b_r[398],
     reset_b_r[399], reset_b_r[400], reset_b_r[401], reset_b_r[402],
     reset_b_r[403], reset_b_r[404], reset_b_r[405], reset_b_r[406],
     reset_b_r[407], reset_b_r[408], reset_b_r[409], reset_b_r[410],
     reset_b_r[411], reset_b_r[412], reset_b_r[413], reset_b_r[414],
     reset_b_r[415], reset_b_r[416], reset_b_r[417], reset_b_r[418],
     reset_b_r[419], reset_b_r[420], reset_b_r[421], reset_b_r[422],
     reset_b_r[423], reset_b_r[424], reset_b_r[425], reset_b_r[426],
     reset_b_r[427], reset_b_r[428], reset_b_r[429], reset_b_r[430],
     reset_b_r[431], reset_b_r[432], reset_b_r[433], reset_b_r[434],
     reset_b_r[435], reset_b_r[436], reset_b_r[437], reset_b_r[438],
     reset_b_r[439], reset_b_r[440], reset_b_r[441], reset_b_r[442],
     reset_b_r[443], reset_b_r[444], reset_b_r[445], reset_b_r[446],
     reset_b_r[447], reset_b_r[448], reset_b_r[449], reset_b_r[450],
     reset_b_r[451], reset_b_r[452], reset_b_r[453], reset_b_r[454],
     reset_b_r[455], reset_b_r[456], reset_b_r[457], reset_b_r[458],
     reset_b_r[459], reset_b_r[460], reset_b_r[461], reset_b_r[462],
     reset_b_r[463], reset_b_r[464], reset_b_r[465], reset_b_r[466],
     reset_b_r[467], reset_b_r[468], reset_b_r[469], reset_b_r[470],
     reset_b_r[471], reset_b_r[472], reset_b_r[473], reset_b_r[474],
     reset_b_r[475], reset_b_r[476], reset_b_r[477], reset_b_r[478],
     reset_b_r[479], reset_b_r[480], reset_b_r[481], reset_b_r[482],
     reset_b_r[483], reset_b_r[484], reset_b_r[485], reset_b_r[486],
     reset_b_r[487], reset_b_r[488], reset_b_r[489], reset_b_r[490],
     reset_b_r[491], reset_b_r[492], reset_b_r[493], reset_b_r[494],
     reset_b_r[495], reset_b_r[496], reset_b_r[497], reset_b_r[498],
     reset_b_r[499], reset_b_r[500], reset_b_r[501], reset_b_r[502],
     reset_b_r[503], reset_b_r[504], reset_b_r[505], reset_b_r[506],
     reset_b_r[507], reset_b_r[508], reset_b_r[509], reset_b_r[510],
     reset_b_r[511], reset_b_r[512], reset_b_r[513], reset_b_r[514],
     reset_b_r[515], reset_b_r[516], reset_b_r[517], reset_b_r[518],
     reset_b_r[519], reset_b_r[520], reset_b_r[521], reset_b_r[522],
     reset_b_r[523], reset_b_r[524], reset_b_r[525], reset_b_r[526],
     reset_b_r[527], reset_b_r[528], reset_b_r[529], reset_b_r[530],
     reset_b_r[531], reset_b_r[532], reset_b_r[533], reset_b_r[534],
     reset_b_r[535], reset_b_r[536], reset_b_r[537], reset_b_r[538],
     reset_b_r[539], reset_b_r[540], reset_b_r[541], reset_b_r[542],
     reset_b_r[543]}), .wl({wl_r[272], wl_r[273], wl_r[274], wl_r[275],
     wl_r[276], wl_r[277], wl_r[278], wl_r[279], wl_r[280], wl_r[281],
     wl_r[282], wl_r[283], wl_r[284], wl_r[285], wl_r[286], wl_r[287],
     wl_r[288], wl_r[289], wl_r[290], wl_r[291], wl_r[292], wl_r[293],
     wl_r[294], wl_r[295], wl_r[296], wl_r[297], wl_r[298], wl_r[299],
     wl_r[300], wl_r[301], wl_r[302], wl_r[303], wl_r[304], wl_r[305],
     wl_r[306], wl_r[307], wl_r[308], wl_r[309], wl_r[310], wl_r[311],
     wl_r[312], wl_r[313], wl_r[314], wl_r[315], wl_r[316], wl_r[317],
     wl_r[318], wl_r[319], wl_r[320], wl_r[321], wl_r[322], wl_r[323],
     wl_r[324], wl_r[325], wl_r[326], wl_r[327], wl_r[328], wl_r[329],
     wl_r[330], wl_r[331], wl_r[332], wl_r[333], wl_r[334], wl_r[335],
     wl_r[336], wl_r[337], wl_r[338], wl_r[339], wl_r[340], wl_r[341],
     wl_r[342], wl_r[343], wl_r[344], wl_r[345], wl_r[346], wl_r[347],
     wl_r[348], wl_r[349], wl_r[350], wl_r[351], wl_r[352], wl_r[353],
     wl_r[354], wl_r[355], wl_r[356], wl_r[357], wl_r[358], wl_r[359],
     wl_r[360], wl_r[361], wl_r[362], wl_r[363], wl_r[364], wl_r[365],
     wl_r[366], wl_r[367], wl_r[368], wl_r[369], wl_r[370], wl_r[371],
     wl_r[372], wl_r[373], wl_r[374], wl_r[375], wl_r[376], wl_r[377],
     wl_r[378], wl_r[379], wl_r[380], wl_r[381], wl_r[382], wl_r[383],
     wl_r[384], wl_r[385], wl_r[386], wl_r[387], wl_r[388], wl_r[389],
     wl_r[390], wl_r[391], wl_r[392], wl_r[393], wl_r[394], wl_r[395],
     wl_r[396], wl_r[397], wl_r[398], wl_r[399], wl_r[400], wl_r[401],
     wl_r[402], wl_r[403], wl_r[404], wl_r[405], wl_r[406], wl_r[407],
     wl_r[408], wl_r[409], wl_r[410], wl_r[411], wl_r[412], wl_r[413],
     wl_r[414], wl_r[415], wl_r[416], wl_r[417], wl_r[418], wl_r[419],
     wl_r[420], wl_r[421], wl_r[422], wl_r[423], wl_r[424], wl_r[425],
     wl_r[426], wl_r[427], wl_r[428], wl_r[429], wl_r[430], wl_r[431],
     wl_r[432], wl_r[433], wl_r[434], wl_r[435], wl_r[436], wl_r[437],
     wl_r[438], wl_r[439], wl_r[440], wl_r[441], wl_r[442], wl_r[443],
     wl_r[444], wl_r[445], wl_r[446], wl_r[447], wl_r[448], wl_r[449],
     wl_r[450], wl_r[451], wl_r[452], wl_r[453], wl_r[454], wl_r[455],
     wl_r[456], wl_r[457], wl_r[458], wl_r[459], wl_r[460], wl_r[461],
     wl_r[462], wl_r[463], wl_r[464], wl_r[465], wl_r[466], wl_r[467],
     wl_r[468], wl_r[469], wl_r[470], wl_r[471], wl_r[472], wl_r[473],
     wl_r[474], wl_r[475], wl_r[476], wl_r[477], wl_r[478], wl_r[479],
     wl_r[480], wl_r[481], wl_r[482], wl_r[483], wl_r[484], wl_r[485],
     wl_r[486], wl_r[487], wl_r[488], wl_r[489], wl_r[490], wl_r[491],
     wl_r[492], wl_r[493], wl_r[494], wl_r[495], wl_r[496], wl_r[497],
     wl_r[498], wl_r[499], wl_r[500], wl_r[501], wl_r[502], wl_r[503],
     wl_r[504], wl_r[505], wl_r[506], wl_r[507], wl_r[508], wl_r[509],
     wl_r[510], wl_r[511], wl_r[512], wl_r[513], wl_r[514], wl_r[515],
     wl_r[516], wl_r[517], wl_r[518], wl_r[519], wl_r[520], wl_r[521],
     wl_r[522], wl_r[523], wl_r[524], wl_r[525], wl_r[526], wl_r[527],
     wl_r[528], wl_r[529], wl_r[530], wl_r[531], wl_r[532], wl_r[533],
     wl_r[534], wl_r[535], wl_r[536], wl_r[537], wl_r[538], wl_r[539],
     wl_r[540], wl_r[541], wl_r[542], wl_r[543]}),
     .smc_write(smc_write_rowu3), .smc_rsr_inc(smc_row_inc_rowu3),
     .rsr_rst(smc_rsr_rst_rowu3), .por_rst(core_por_b_rowu3),
     .cram_wl_en(cram_wl_en_rowu3), .cram_vddoff(cram_vddoff_rowu3),
     .cram_rst(cram_rst_rowu3), .cram_pgateoff(cram_pgateoff_rowu3),
     .banksel(cm_banksel_bltrd0[3]), .last_rsr(last_rsr[1]),
     .trst_b(j_rst_b_rowu3), .jtag_rowtest_rst(row_test_rowu3),
     .jtag_clk(tck_pad_rowu3),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu3_b));
ml_rowdrv_bank10k Irowlr ( .vddctrl(vdd_cntl_r[271:0]),
     .pgate(pgate_r[271:0]), .reset(reset_b_r[271:0]),
     .wl(wl_r[271:0]), .smc_write(smc_write_rowu2),
     .smc_rsr_inc(smc_row_inc_rowu2), .rsr_rst(smc_rsr_rst_rowu2),
     .por_rst(core_por_b_rowu2), .cram_wl_en(cram_wl_en_rowu2),
     .cram_vddoff(cram_vddoff_rowu2), .cram_rst(cram_rst_rowu2),
     .cram_pgateoff(cram_pgateoff_rowu2),
     .banksel(cm_banksel_blbrd_2_), .last_rsr(last_rsr[0]),
     .trst_b(j_rst_b_rowu2), .jtag_rowtest_rst(row_test_rowu2),
     .jtag_clk(tck_pad_rowu2),
     .jtag_rowtest_mode_b(jtag_rowtest_mode_rowu2_b));
SMC_CORE_POR_right I450 ( .vddio_rightbank(vddio_rightbank),
     .smc_por_b(smc_por_b0), .core_por_b(core_por_b0),
     .smc_core_por_bottom1(smc_core_por_bottom1),
     .smc_core_por_bottom2(smc_core_por_bottom2));
sg_bufx10 I460_1_ ( .in(cm_banksel[1]), .out(cm_banksel_bldld[1]));
sg_bufx10 I460_0_ ( .in(cm_banksel[0]), .out(cm_banksel_bldld[0]));
sg_bufx10 I307 ( .in(cram_pgateoff), .out(cram_pgateoffr0));
sg_bufx10 I208 ( .in(cm_banksel[3]), .out(cm_banksel_bltrd[3]));
sg_bufx10 I308 ( .in(cram_rst), .out(cram_rstr0));
sg_bufx10 I309 ( .in(cram_vddoff), .out(cram_vddoffr0));
sg_bufx10 I310 ( .in(cram_wl_en), .out(cram_wl_enr0));
sg_bufx10 I311 ( .in(smc_row_inc), .out(smc_row_incr0));
sg_bufx10 I151 ( .in(cram_prec), .out(cram_prec_blbrd));
sg_bufx10 I312 ( .in(smc_write0), .out(smc_writer0));
sg_bufx10 I315 ( .in(cram_pgateoffr0), .out(cram_pgateoffr1));
sg_bufx10 I201 ( .in(cm_banksel_bltrd[3]), .out(cm_banksel_bltrd0[3]));
sg_bufx10 I157 ( .in(smc_wdis_dclk), .out(smc_wdis_dclk_blbrd));
sg_bufx10 I431 ( .in(monitor_celld[3]), .out(monitor_celld1[3]));
sg_bufx10 I282_1_ ( .in(cm_sdi_u3d[1]), .out(cm_sdi_u3d0[1]));
sg_bufx10 I282_0_ ( .in(cm_sdi_u3d[0]), .out(cm_sdi_u3d0[0]));
sg_bufx10 I320 ( .in(smc_writer0), .out(smc_writer1));
sg_bufx10 I322 ( .in(tck_padr0), .out(tck_padr1));
sg_bufx10 I317 ( .in(cram_vddoffr0), .out(cram_vddoffr1));
sg_bufx10 I432 ( .in(cf_r[0]), .out(monitor_celld[2]));
sg_bufx10 I323 ( .in(row_test1), .out(row_testr1));
sg_bufx10 I455_1_ ( .in(dff_out_bot[1]), .out(cm_sdo_u3d0[1]));
sg_bufx10 I455_0_ ( .in(dff_out_bot[0]), .out(cm_sdo_u3d0[0]));
sg_bufx10 I207 ( .in(en_8bconfig_b_blbrd), .out(en_8bconfig_b_bltrd0));
sg_bufx10 I434_1_ ( .in(monitor_celld2[3]), .out(monitor_celldd[3]));
sg_bufx10 I434_0_ ( .in(monitor_celld[2]), .out(monitor_celldd[2]));
sg_bufx10 I210 ( .in(cram_write_bltrd0), .out(cram_write_bltrd1));
sg_bufx10 I205 ( .in(data_muxsel_blbrd), .out(data_muxsel_bltrd0));
sg_bufx10 I206 ( .in(cram_write_blbrd), .out(cram_write_bltrd0));
sg_bufx10 I153 ( .in(data_muxsel), .out(data_muxsel_blbrd));
sg_bufx10 I458_1_ ( .in(u0_in[1]), .out(cm_sdi_u0[1]));
sg_bufx10 I458_0_ ( .in(u0_in[0]), .out(cm_sdi_u0[0]));
sg_bufx10 I433 ( .in(monitor_celld1[3]), .out(monitor_celld2[3]));
sg_bufx10 I152 ( .in(cram_write), .out(cram_write_blbrd));
sg_bufx10 I304 ( .in(j_tck), .out(tck_padr0));
sg_bufx10 I319 ( .in(smc_row_incr0), .out(smc_row_incr1));
sg_bufx10 I457 ( .in(net257), .out(smc_rsr_rst));
sg_bufx10 I454_1_ ( .in(dff_out_top[1]), .out(cm_sdo_u3dd[1]));
sg_bufx10 I454_0_ ( .in(dff_out_top[0]), .out(cm_sdo_u3dd[0]));
sg_bufx10 I198 ( .in(cram_pullup_b), .out(cram_pullup_b_bldrd));
sg_bufx10 I156 ( .in(smc_clk_out), .out(cm_clk_blbrd));
sg_bufx10 I150 ( .in(cm_banksel[2]), .out(cm_banksel_blbrd_2_));
sg_bufx10 I288_1_ ( .in(cm_sdo_u3d0[1]), .out(cm_sdo_u3d1[1]));
sg_bufx10 I288_0_ ( .in(cm_sdo_u3d0[0]), .out(cm_sdo_u3d1[0]));
sg_bufx10 I155 ( .in(en_8bconfig_b), .out(en_8bconfig_b_blbrd));
sg_bufx10 I115_1_ ( .in(cm_sdi_u2[1]), .out(cm_sdi_u2d[1]));
sg_bufx10 I115_0_ ( .in(cm_sdi_u2[0]), .out(cm_sdi_u2d[0]));
sg_bufx10 I116_1_ ( .in(cm_sdi_u3[1]), .out(cm_sdi_u3d[1]));
sg_bufx10 I116_0_ ( .in(cm_sdi_u3[0]), .out(cm_sdi_u3d[0]));
sg_bufx10 I154 ( .in(data_muxsel1), .out(data_muxsel1_blbrd));
sg_bufx10 I324 ( .in(smc_rsr_rstr0), .out(smc_rsr_rstr1));
sg_bufx10 I202 ( .in(cm_clk_blbrd), .out(cm_clk_bltrd0));
sg_bufx10 I459_1_ ( .in(u1_in[1]), .out(cm_sdi_u1[1]));
sg_bufx10 I459_0_ ( .in(u1_in[0]), .out(cm_sdi_u1[0]));
sg_bufx10 I203 ( .in(data_muxsel1_blbrd), .out(data_muxsel1_bltrd0));
sg_bufx10 I325 ( .in(core_por_bbr0), .out(core_por_b_rowu3));
sg_bufx10 I456 ( .in(net261), .out(smc_row_inc));
sg_bufx10 I215 ( .in(cm_banksel_bltrd0[3]),
     .out(cm_banksel_bltrd1_3_));
sg_bufx10 I443 ( .in(j_rst_br0), .out(j_rst_br1));
sg_bufx10 I306 ( .in(row_test0), .out(row_test1));
sg_bufx10 I212 ( .in(smc_wdis_dclk_bltrd0),
     .out(smc_wdis_dclk_bltrd1));
sg_bufx10 I209 ( .in(en_8bconfig_b_bltrd0),
     .out(en_8bconfig_b_bltrd1));
sg_bufx10 I213 ( .in(data_muxsel1_bltrd0), .out(data_muxsel1_bltrd1));
sg_bufx10 I204 ( .in(smc_wdis_dclk_blbrd), .out(smc_wdis_dclk_bltrd0));
sg_bufx10 I200 ( .in(cram_prec_blbrd), .out(cram_prec_bltrd0));
sg_bufx10 I199 ( .in(cram_pullup_b_bldrd), .out(cram_pullup_b_bltrd0));
sg_bufx10 I211 ( .in(data_muxsel_bltrd0), .out(data_muxsel_bltrd1));
sg_bufx10 I217 ( .in(cram_pullup_b_bltrd0),
     .out(cram_pullup_b_bltrd1));
sg_bufx10 I440 ( .in(j_rst_b), .out(j_rst_br0));
sg_bufx10 I214 ( .in(cm_clk_bltrd0), .out(cm_clk_bltrd1));
sg_bufx10 I216 ( .in(cram_prec_bltrd0), .out(cram_prec_bltrd1));
sg_bufx10 I305 ( .in(smc_rsr_rst), .out(smc_rsr_rstr0));
sg_bufx10 I285_1_ ( .in(cm_sdo_u3[1]), .out(cm_sdo_u3d[1]));
sg_bufx10 I285_0_ ( .in(cm_sdo_u3[0]), .out(cm_sdo_u3d[0]));
sg_bufx10 I318 ( .in(cram_wl_enr0), .out(cram_wl_enr1));
sg_bufx10 I283_1_ ( .in(cm_sdi_u3d0[1]), .out(cm_sdi_u3d2[1]));
sg_bufx10 I283_0_ ( .in(cm_sdi_u3d0[0]), .out(cm_sdi_u3d2[0]));
sg_bufx10 I314 ( .in(core_por_bb), .out(core_por_bbr0));
sg_bufx10 I316 ( .in(cram_rstr0), .out(cram_rstr1));
sg_bufx10 I430 ( .in(cf_r[1]), .out(monitor_celld[3]));
inv_hvt I136 ( .A(core_por_b0), .Y(core_por_bb));
ml_osc_top Iml_osc ( .smc_podt_rst(smc_podt_rst),
     .smc_podt_off(smc_podt_off), .smc_oscoff_b(smc_oscoff_b),
     .smc_osc_fsel(smc_osco_fsel[1:0]), .por_b(core_por_b0),
     .crst_b(crst_filterout), .smc_clk(osc_clk),
     .cnt_podt_out(cnt_podt_out));
bram_bufferx16 I407 ( .in(cram_wl_enr0), .out(cram_wl_en_rowu2));
bram_bufferx16 I416 ( .in(cram_rstr1), .out(cram_rst_rowu3));
bram_bufferx16 I185 ( .in(core_por_b0), .out(core_por_b1));
bram_bufferx16 I442 ( .in(j_rst_br1), .out(j_rst_b_rowu3));
bram_bufferx16 I441 ( .in(j_rst_br0), .out(j_rst_b_rowu2));
bram_bufferx16 I409 ( .in(smc_writer0), .out(smc_write_rowu2));
bram_bufferx16 I287 ( .in(cm_clk_bltrd0), .out(net507));
bram_bufferx16 I452 ( .in(smc_clk_out), .out(net509));
bram_bufferx16 I451_6_ ( .in(spi_ss_in_r[7]), .out(spi_ss_in_rd[7]));
bram_bufferx16 I451_5_ ( .in(spi_ss_in_r[6]), .out(spi_ss_in_rd[6]));
bram_bufferx16 I451_4_ ( .in(spi_ss_in_r[5]), .out(spi_ss_in_rd[5]));
bram_bufferx16 I451_3_ ( .in(spi_ss_in_r[4]), .out(spi_ss_in_rd[4]));
bram_bufferx16 I451_2_ ( .in(spi_ss_in_r[3]), .out(spi_ss_in_rd[3]));
bram_bufferx16 I451_1_ ( .in(spi_ss_in_r[2]), .out(spi_ss_in_rd[2]));
bram_bufferx16 I451_0_ ( .in(spi_ss_in_r[1]), .out(spi_ss_in_rd[1]));
bram_bufferx16 I402 ( .in(smc_rsr_rstr0), .out(smc_rsr_rst_rowu2));
bram_bufferx16 I410 ( .in(core_por_bbr0), .out(core_por_b_rowu2));
bram_bufferx16 I406 ( .in(cram_vddoffr0), .out(cram_vddoff_rowu2));
bram_bufferx16 I405 ( .in(cram_rstr0), .out(cram_rst_rowu2));
bram_bufferx16 I401 ( .in(tck_padr0), .out(tck_pad_rowu2));
bram_bufferx16 I403 ( .in(row_test1), .out(row_test_rowu2));
bram_bufferx16 I420 ( .in(tck_padr1), .out(tck_pad_rowu3));
bram_bufferx16 I418 ( .in(row_testr1), .out(row_test_rowu3));
bram_bufferx16 I408 ( .in(smc_row_incr0), .out(smc_row_inc_rowu2));
bram_bufferx16 I404 ( .in(cram_pgateoffr0), .out(cram_pgateoff_rowu2));
bram_bufferx16 I412 ( .in(smc_writer1), .out(smc_write_rowu3));
bram_bufferx16 I414 ( .in(cram_wl_enr1), .out(cram_wl_en_rowu3));
bram_bufferx16 I413 ( .in(smc_row_incr1), .out(smc_row_inc_rowu3));
bram_bufferx16 I417 ( .in(cram_pgateoffr1), .out(cram_pgateoff_rowu3));
bram_bufferx16 I419 ( .in(smc_rsr_rstr1), .out(smc_rsr_rst_rowu3));
bram_bufferx16 I415 ( .in(cram_vddoffr1), .out(cram_vddoff_rowu3));
ml_cram_logic Iml_cram_logic ( .smc_wwlwrt_en(smc_wwlwrt_en),
     .smc_wset_precgnd(smc_wset_precgnd), .smc_write(smc_write0),
     .cram_pgateoff(cram_pgateoff), .smc_wcram_rst(smc_wcram_rst),
     .smc_rwl_en(smc_rwl_en), .smc_rrst_pullwlen(smc_rrst_pullwlen),
     .smc_rpull_b(smc_rpull_b), .smc_rprec(smc_rprec),
     .smc_read(net263), .smc_clk(cm_clk), .por(core_por_bb),
     .cram_write(cram_write), .cram_wl_en(cram_wl_en),
     .cram_rst(cram_rst), .cram_pullup_b(cram_pullup_b),
     .cram_prec(cram_prec), .cram_vddoff(cram_vddoff),
     .smc_seq_rst(smc_seq_rst), .smc_clk_out(smc_clk_out),
     .smc_wwlwrt_dis(smc_wwlwrt_dis), .smc_wset_prec(smc_wset_prec));

endmodule
// Library - NVCM, Cell - ml_lshv_6v_hold, View - schematic
// LAST TIME SAVED: Dec 20 11:32:52 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_lshv_6v_hold ( out_b_hv, out_hv, in_hv, sel_25, sel_b_25,
     vddp_tieh );
output  out_b_hv, out_hv;

inout  in_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M2 ( .D(out_b_hv), .B(net129), .G(sel_25), .S(net129));
pch_25  M5 ( .D(out_hv), .B(net121), .G(sel_b_25), .S(net121));
pch_25  M7 ( .D(net129), .B(in_hv), .G(out_hv), .S(in_hv));
pch_25  M6 ( .D(net121), .B(in_hv), .G(out_b_hv), .S(in_hv));
nch_25  M12 ( .D(out_hv), .B(GND_), .G(vddp_tieh), .S(net132));
nch_25  M15 ( .D(net132), .B(GND_), .G(sel_b_25), .S(gnd_));
nch_25  M10 ( .D(out_b_hv), .B(GND_), .G(vddp_tieh), .S(net140));
nch_25  M14 ( .D(net140), .B(GND_), .G(sel_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_hv_inv, View - schematic
// LAST TIME SAVED: Jan 21 18:15:24 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_hv_inv ( out_b_hv, in_hv, sel_25, sel_hv, vddp_tieh );
output  out_b_hv;

inout  in_hv;

input  sel_25, sel_hv, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M16 ( .D(net86), .B(in_hv), .G(sel_hv), .S(in_hv));
pch_25  M39 ( .D(out_b_hv), .B(net86), .G(sel_25), .S(net86));
nch_25  M29 ( .D(net89), .B(gnd_), .G(sel_25), .S(gnd_));
nch_25  M21 ( .D(out_b_hv), .B(gnd_), .G(vddp_tieh), .S(net89));

endmodule
// Library - io, Cell - PVSS3DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:17:04 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module PVSS3DGZ ( VSS );
input  VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_hv_ls_inv, View - schematic
// LAST TIME SAVED: Jan  8 14:11:13 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_hv_ls_inv ( in_hv, out_b_hv, sel_25, sel_b_25, vddp_tieh );
inout  in_hv, out_b_hv;

input  sel_25, sel_b_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_lshv_6v_hold Ishv_6v_hold ( .vddp_tieh(vddp_tieh), .out_b_hv(net61),
     .in_hv(in_hv), .sel_b_25(sel_b_25), .sel_25(sel_25),
     .out_hv(sel_hv));
ml_hv_inv Ihv_inv ( .vddp_tieh(vddp_tieh), .out_b_hv(out_b_hv),
     .sel_25(sel_25), .in_hv(in_hv), .sel_hv(sel_hv));

endmodule
// Library - tsmcN65lo, Cell - nand3_25, View - schematic
// LAST TIME SAVED: Mar 29 20:19:50 2006
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nand3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(net21), .B(Gb), .G(C), .S(G));
nch_25  M2 ( .D(net25), .B(Gb), .G(B), .S(net21));
nch_25  NM1 ( .D(Y), .B(Gb), .G(A), .S(net25));
pch_25  PM1 ( .D(Y), .B(Pb), .G(A), .S(P));
pch_25  M1 ( .D(Y), .B(Pb), .G(C), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(P));

endmodule
// Library - tsmcN65lo, Cell - nor3_25, View - schematic
// LAST TIME SAVED: Mar 29 20:26:16 2006
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nor3_25 ( Y, A, B, C, G, Gb, P, Pb );
output  Y;

input  A, B, C, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M2 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  M3 ( .D(Y), .B(Gb), .G(C), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  M1 ( .D(Y), .B(Pb), .G(C), .S(net16));
pch_25  PM1 ( .D(net12), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(net16), .B(Pb), .G(B), .S(net12));

endmodule
// Library - NVCM, Cell - ml_ls_vdd2vdd25, View - schematic
// LAST TIME SAVED: Apr  4 14:26:57 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ls_vdd2vdd25 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(out_vddio_b), .B(sup), .G(in), .S(net29));
pch_25  M13 ( .D(out_vddio), .B(sup), .G(in_b), .S(net33));
pch_25  M4 ( .D(net29), .B(sup), .G(out_vddio), .S(sup));
pch_25  M6 ( .D(net33), .B(sup), .G(out_vddio_b), .S(sup));
nch_25  M9 ( .D(out_vddio), .B(gnd_), .G(in_b), .S(gnd_));
nch_25  M7 ( .D(out_vddio_b), .B(gnd_), .G(in), .S(gnd_));

endmodule
// Library - tsmcN65lo, Cell - inv_25, View - schematic
// LAST TIME SAVED: Mar 29 20:14:12 2006
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module inv_25 ( OUT, G, Gb, IN, P, Pb );
output  OUT;

input  G, Gb, IN, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  NM1 ( .D(OUT), .B(Gb), .G(IN), .S(G));
pch_25  PM1 ( .D(OUT), .B(Pb), .G(IN), .S(P));

endmodule
// Library - sbtlibn65lp, Cell - vdd_tielow, View - schematic
// LAST TIME SAVED: May  8 16:23:59 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module vdd_tielow ( gnd_tiel );
inout  gnd_tiel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(gnd_tiel), .B(GND_), .G(net9), .S(gnd_));
pch_hvt  M3 ( .D(net9), .B(vdd_), .G(net9), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_chip_spare, View - schematic
// LAST TIME SAVED: Sep 11 18:02:11 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_chip_spare (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M14 ( .D(net96), .B(net85), .G(net286), .S(net85));
pch_25  M5 ( .D(net85), .B(net123), .G(net114), .S(net123));
pch_25  M3 ( .D(net108), .B(net89), .G(net316), .S(net89));
pch_25  M2 ( .D(net89), .B(net126), .G(net119), .S(net126));
nch_25  M7 ( .D(net100), .B(GND_), .G(net286), .S(gnd_));
nch_25  M1 ( .D(net96), .B(GND_), .G(net121), .S(net100));
nch_25  M6 ( .D(net104), .B(GND_), .G(net316), .S(gnd_));
nch_25  M4 ( .D(net108), .B(GND_), .G(net121), .S(net104));
ml_hv_ls_inv I132 ( .sel_b_25(net316), .sel_25(net405),
     .out_b_hv(net119), .in_hv(net126), .vddp_tieh(net121));
ml_hv_ls_inv Iml_hv_ls_inv_vppt ( .sel_b_25(net286), .sel_25(net404),
     .out_b_hv(net114), .in_hv(net123), .vddp_tieh(net121));
rppolywo_m  R8 ( .MINUS(vddp_), .PLUS(net123), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(vddp_), .PLUS(net126), .BULK(gnd_));
nand3_25 I257 ( .B(net0373), .A(net0373), .Y(net0397), .C(net0373),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I256 ( .B(net0381), .A(net0381), .Y(net0373), .C(net0381),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I255 ( .B(net215), .A(net215), .Y(net0381), .C(net215),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I248 ( .B(net0397), .A(net0397), .Y(net0405), .C(net0397),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I247 ( .B(net0405), .A(net0405), .Y(net0413), .C(net0405),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I245 ( .B(net0413), .A(net0413), .Y(net0421), .C(net0413),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I244 ( .B(net0421), .A(net0421), .Y(net0453), .C(net0421),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I231 ( .B(net0453), .A(net0453), .Y(net0445), .C(net0453),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I233 ( .B(net0437), .A(net0437), .Y(net0429), .C(net0437),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I234 ( .B(net0429), .A(net0429), .Y(net0595), .C(net0429),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I232 ( .B(net0445), .A(net0445), .Y(net0437), .C(net0445),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nor3_25 I215 ( .B(net0460), .A(net0460), .C(net0460), .Y(net0594),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I214 ( .B(net0468), .A(net0468), .C(net0468), .Y(net0460),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I212 ( .B(net0476), .A(net0476), .C(net0476), .Y(net0468),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I211 ( .B(net160), .A(net160), .C(net160), .Y(net0492),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I209 ( .B(net0500), .A(net0500), .C(net0500), .Y(net0476),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I42 ( .B(net191), .A(net191), .C(net191), .Y(net160), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I78 ( .B(net199), .A(net199), .C(net199), .Y(net191), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I83 ( .B(net207), .A(net207), .C(net207), .Y(net199), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I84 ( .B(net215), .A(net215), .C(net215), .Y(net207), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I210 ( .B(net0492), .A(net0492), .C(net0492), .Y(net0500),
     .G(gnd_), .Gb(gnd_), .Pb(vddp_), .P(vddp_));
inv_hvt I120 ( .A(net253), .Y(net249));
inv_hvt I119 ( .A(net231), .Y(net253));
inv_hvt I118 ( .A(net231), .Y(net258));
inv_hvt I117 ( .A(net258), .Y(net254));
inv_hvt I319 ( .A(net263), .Y(net259));
inv_hvt I323 ( .A(net231), .Y(net263));
inv_hvt I57 ( .A(net231), .Y(net268));
inv_hvt I58 ( .A(net268), .Y(net264));
ml_ls_vdd2vdd25 I122 ( .in(net249), .sup(vddp_), .out_vddio_b(net291),
     .out_vddio(net252), .in_b(net253));
ml_ls_vdd2vdd25 I121 ( .in(net254), .sup(vddp_), .out_vddio_b(net297),
     .out_vddio(net257), .in_b(net258));
ml_ls_vdd2vdd25 I335 ( .in(net259), .sup(vddp_), .out_vddio_b(net303),
     .out_vddio(net262), .in_b(net263));
ml_ls_vdd2vdd25 I56 ( .in(net264), .sup(vddp_), .out_vddio_b(net309),
     .out_vddio(net267), .in_b(net268));
inv_25 I126 ( .IN(net291), .OUT(net271), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I125 ( .IN(net297), .OUT(net272), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I139 ( .IN(net405), .OUT(net316), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(net404), .OUT(net286), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I384 ( .IN(net303), .OUT(net274), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I54 ( .IN(net309), .OUT(net273), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nand3_hvt I185 ( .Y(net0665), .B(net0661), .C(net0661), .A(net0661));
nand3_hvt I186 ( .Y(net0661), .B(net0657), .C(net0657), .A(net0657));
nand3_hvt I187 ( .Y(net0657), .B(net0653), .C(net0653), .A(net0653));
nand3_hvt I188 ( .Y(net0653), .B(net0649), .C(net0649), .A(net0649));
nand3_hvt I183 ( .Y(net0649), .B(net281), .C(net281), .A(net281));
nand3_hvt I246 ( .Y(net328), .B(net324), .C(net324), .A(net324));
nand3_hvt I61 ( .Y(net332), .B(net328), .C(net328), .A(net328));
nand3_hvt I62 ( .Y(net336), .B(net332), .C(net332), .A(net332));
nand3_hvt I63 ( .Y(net340), .B(net336), .C(net336), .A(net336));
nand3_hvt I64 ( .Y(net360), .B(net340), .C(net340), .A(net340));
nand3_hvt I104 ( .Y(net281), .B(net344), .C(net344), .A(net344));
nand3_hvt I105 ( .Y(net344), .B(net348), .C(net348), .A(net348));
nand3_hvt I106 ( .Y(net348), .B(net352), .C(net352), .A(net352));
nand3_hvt I107 ( .Y(net352), .B(net356), .C(net356), .A(net356));
nand3_hvt I108 ( .Y(net356), .B(net360), .C(net360), .A(net360));
nand3_hvt I184 ( .Y(net0596), .B(net0665), .C(net0665), .A(net0665));
nor3_hvt I177 ( .B(net0732), .Y(net0728), .A(net0732), .C(net0732));
nor3_hvt I178 ( .B(net0728), .Y(net0724), .A(net0728), .C(net0728));
nor3_hvt I179 ( .B(net0724), .Y(net0720), .A(net0724), .C(net0724));
nor3_hvt I180 ( .B(net0720), .Y(net0716), .A(net0720), .C(net0720));
nor3_hvt I181 ( .B(net0716), .Y(net0712), .A(net0716), .C(net0716));
nor3_hvt I182 ( .B(net0712), .Y(net0597), .A(net0712), .C(net0712));
nor3_hvt I65 ( .B(net363), .Y(net383), .A(net363), .C(net363));
nor3_hvt I70 ( .B(net367), .Y(net363), .A(net367), .C(net367));
nor3_hvt I71 ( .B(net371), .Y(net367), .A(net371), .C(net371));
nor3_hvt I72 ( .B(net375), .Y(net371), .A(net375), .C(net375));
nor3_hvt I73 ( .B(net379), .Y(net375), .A(net379), .C(net379));
nor3_hvt I99 ( .B(net383), .Y(net387), .A(net383), .C(net383));
nor3_hvt I100 ( .B(net387), .Y(net391), .A(net387), .C(net387));
nor3_hvt I101 ( .B(net391), .Y(net395), .A(net391), .C(net391));
nor3_hvt I102 ( .B(net395), .Y(net399), .A(net395), .C(net395));
nor3_hvt I103 ( .B(net399), .Y(net0732), .A(net399), .C(net399));
vddp_tiehigh I140 ( .vddp_tieh(net121));
vdd_tielow I154 ( .gnd_tiel(net405));
vdd_tielow I155 ( .gnd_tiel(net404));
vdd_tielow I153 ( .gnd_tiel(net231));
vdd_tielow I146 ( .gnd_tiel(net215));
vdd_tielow I145 ( .gnd_tiel(net324));
vdd_tielow I144 ( .gnd_tiel(net379));

endmodule
// Library - NVCM, Cell - ml_chip_buf, View - schematic
// LAST TIME SAVED: Feb 26 16:35:06 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_chip_buf ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I131 ( .A(in), .Y(net120));
inv_hvt I45 ( .A(net120), .Y(out));

endmodule
// Library - NVCM, Cell - ml_chip_buf_top_8f, View - schematic
// LAST TIME SAVED: Sep  3 10:26:28 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_chip_buf_top_8f ( fsm_blkadd_b_buf, fsm_blkadd_buf,
     fsm_coladd_buf, fsm_din_buf, fsm_gwlbdis_buf, fsm_lshven_buf,
     fsm_multibl_read_buf, fsm_nv_bstream_buf, fsm_nv_rri_trim_buf,
     fsm_nv_rrow_buf, fsm_nv_sisi_ui_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmhv_buf, fsm_pgmien_buf, fsm_pgmvfy_buf,
     fsm_rd_buf, fsm_rowadd_buf, fsm_rst_b_buf, fsm_sample_buf,
     fsm_tm_rd_mode_buf, fsm_tm_testdec_buf, fsm_tm_trow_buf,
     fsm_trim_ipp_buf, fsm_trim_rrefpgm_buf, fsm_trim_rrefrd_buf,
     fsm_trim_vbg_buf, fsm_vpgmwl_buf, fsm_vpxaset_buf, fsm_wgnden_buf,
     fsm_wpen_buf, fsm_wren_buf, fsm_ymuxdis_buf, nv_dataout_buf,
     tm_allbank_sel_buf, tm_allbl_h_buf, tm_allbl_l_buf,
     tm_allwl_h_buf, tm_allwl_l_buf, tm_dma_buf, tm_tcol_buf,
     tm_testdec_wr_buf, fsm_blkadd, fsm_blkadd_b, fsm_coladd, fsm_din,
     fsm_gwlbdis, fsm_lshven, fsm_multibl_read, fsm_nv_bstream,
     fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm,
     fsm_pgmdisc, fsm_pgmhv, fsm_pgmien, fsm_pgmvfy, fsm_rd,
     fsm_rowadd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_ipp, fsm_trim_rrefpgm, fsm_trim_rrefrd,
     fsm_trim_vbg, fsm_vpgmwl, fsm_vpxaset, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, nv_dataout, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr
     );
output  fsm_din_buf, fsm_gwlbdis_buf, fsm_lshven_buf,
     fsm_multibl_read_buf, fsm_nv_bstream_buf, fsm_nv_rri_trim_buf,
     fsm_nv_rrow_buf, fsm_nv_sisi_ui_buf, fsm_nvcmen_buf, fsm_pgm_buf,
     fsm_pgmdisc_buf, fsm_pgmhv_buf, fsm_pgmien_buf, fsm_pgmvfy_buf,
     fsm_rd_buf, fsm_rst_b_buf, fsm_sample_buf, fsm_tm_rd_mode_buf,
     fsm_tm_testdec_buf, fsm_tm_trow_buf, fsm_vpxaset_buf,
     fsm_wgnden_buf, fsm_wpen_buf, fsm_wren_buf, fsm_ymuxdis_buf,
     tm_allbank_sel_buf, tm_allbl_h_buf, tm_allbl_l_buf,
     tm_allwl_h_buf, tm_allwl_l_buf, tm_dma_buf, tm_tcol_buf,
     tm_testdec_wr_buf;

input  fsm_din, fsm_gwlbdis, fsm_lshven, fsm_multibl_read,
     fsm_nv_bstream, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmdisc, fsm_pgmhv, fsm_pgmien,
     fsm_pgmvfy, fsm_rd, fsm_rst_b, fsm_sample, fsm_tm_rd_mode,
     fsm_tm_testdec, fsm_tm_trow, fsm_vpxaset, fsm_wgnden, fsm_wpen,
     fsm_wren, fsm_ymuxdis, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [3:0]  fsm_blkadd_b_buf;
output [3:0]  fsm_trim_ipp_buf;
output [2:0]  fsm_vpgmwl_buf;
output [3:0]  fsm_blkadd_buf;
output [2:0]  fsm_trim_rrefrd_buf;
output [3:0]  nv_dataout_buf;
output [9:0]  fsm_coladd_buf;
output [7:0]  fsm_rowadd_buf;
output [3:0]  fsm_trim_vbg_buf;
output [2:0]  fsm_trim_rrefpgm_buf;

input [7:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_trim_ipp;
input [3:0]  nv_dataout;
input [2:0]  fsm_trim_rrefpgm;
input [9:0]  fsm_coladd;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_vpgmwl;
input [3:0]  fsm_trim_vbg;
input [3:0]  fsm_blkadd_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:3]  net188;



mux2_hvt I134 ( .in1(net0182), .in0(net0182), .out(net0281),
     .sel(gnd_in));
mux2_hvt I206 ( .in1(gnd_in), .in0(gnd_in), .out(net0190),
     .sel(gnd_in));
mux2_hvt I132 ( .in1(net0190), .in0(net0190), .out(net0186),
     .sel(gnd_in));
mux2_hvt I133 ( .in1(net0186), .in0(net0186), .out(net0182),
     .sel(gnd_in));
vdd_tielow I135 ( .gnd_tiel(gnd_in));
vdd_tielow I145 ( .gnd_tiel(net0280));
vdd_tielow I144 ( .gnd_tiel(net0223));
nor3_hvt I125 ( .B(net0239), .Y(net0219), .A(net0239), .C(net0239));
nor3_hvt I126 ( .B(net0235), .Y(net0239), .A(net0235), .C(net0235));
nor3_hvt I127 ( .B(net0231), .Y(net0235), .A(net0231), .C(net0231));
nor3_hvt I128 ( .B(net0227), .Y(net0231), .A(net0227), .C(net0227));
nor3_hvt I129 ( .B(net0223), .Y(net0227), .A(net0223), .C(net0223));
nor3_hvt I99 ( .B(net0219), .Y(net0215), .A(net0219), .C(net0219));
nor3_hvt I100 ( .B(net0215), .Y(net0211), .A(net0215), .C(net0215));
nor3_hvt I101 ( .B(net0211), .Y(net0207), .A(net0211), .C(net0211));
nor3_hvt I130 ( .B(net0207), .Y(net0203), .A(net0207), .C(net0207));
nor3_hvt I103 ( .B(net0203), .Y(net0282), .A(net0203), .C(net0203));
nand3_hvt I246 ( .Y(net0276), .B(net0280), .C(net0280), .A(net0280));
nand3_hvt I61 ( .Y(net0272), .B(net0276), .C(net0276), .A(net0276));
nand3_hvt I62 ( .Y(net0268), .B(net0272), .C(net0272), .A(net0272));
nand3_hvt I123 ( .Y(net0264), .B(net0268), .C(net0268), .A(net0268));
nand3_hvt I124 ( .Y(net0244), .B(net0264), .C(net0264), .A(net0264));
nand3_hvt I104 ( .Y(net0283), .B(net0260), .C(net0260), .A(net0260));
nand3_hvt I105 ( .Y(net0260), .B(net0256), .C(net0256), .A(net0256));
nand3_hvt I106 ( .Y(net0256), .B(net0252), .C(net0252), .A(net0252));
nand3_hvt I107 ( .Y(net0252), .B(net0248), .C(net0248), .A(net0248));
nand3_hvt I108 ( .Y(net0248), .B(net0244), .C(net0244), .A(net0244));
vdd_tiehigh I117 ( .vdd_tieh(vdd_spare));
ml_chip_buf I120_3_ ( .in(vdd_spare), .out(net188[0]));
ml_chip_buf I120_2_ ( .in(vdd_spare), .out(net188[1]));
ml_chip_buf I120_1_ ( .in(vdd_spare), .out(net188[2]));
ml_chip_buf I120_0_ ( .in(vdd_spare), .out(net188[3]));
ml_chip_buf I118 ( .in(tm_allbank_sel), .out(tm_allbank_sel_buf));
ml_chip_buf I102_3_ ( .in(nv_dataout[3]), .out(nv_dataout_buf[3]));
ml_chip_buf I102_2_ ( .in(nv_dataout[2]), .out(nv_dataout_buf[2]));
ml_chip_buf I102_1_ ( .in(nv_dataout[1]), .out(nv_dataout_buf[1]));
ml_chip_buf I102_0_ ( .in(nv_dataout[0]), .out(nv_dataout_buf[0]));
ml_chip_buf I95_3_ ( .in(fsm_trim_ipp[3]), .out(fsm_trim_ipp_buf[3]));
ml_chip_buf I95_2_ ( .in(fsm_trim_ipp[2]), .out(fsm_trim_ipp_buf[2]));
ml_chip_buf I95_1_ ( .in(fsm_trim_ipp[1]), .out(fsm_trim_ipp_buf[1]));
ml_chip_buf I95_0_ ( .in(fsm_trim_ipp[0]), .out(fsm_trim_ipp_buf[0]));
ml_chip_buf I94 ( .in(fsm_wren), .out(fsm_wren_buf));
ml_chip_buf I93 ( .in(fsm_pgmhv), .out(fsm_pgmhv_buf));
ml_chip_buf I87 ( .in(fsm_ymuxdis), .out(fsm_ymuxdis_buf));
ml_chip_buf I86 ( .in(tm_allbl_h), .out(tm_allbl_h_buf));
ml_chip_buf I85 ( .in(tm_allbl_l), .out(tm_allbl_l_buf));
ml_chip_buf I84 ( .in(tm_tcol), .out(tm_tcol_buf));
ml_chip_buf I83 ( .in(tm_allwl_l), .out(tm_allwl_l_buf));
ml_chip_buf I82 ( .in(tm_allwl_h), .out(tm_allwl_h_buf));
ml_chip_buf I81 ( .in(fsm_nv_rrow), .out(fsm_nv_rrow_buf));
ml_chip_buf I80 ( .in(tm_testdec_wr), .out(tm_testdec_wr_buf));
ml_chip_buf I89 ( .in(fsm_tm_trow), .out(fsm_tm_trow_buf));
ml_chip_buf I88 ( .in(fsm_gwlbdis), .out(fsm_gwlbdis_buf));
ml_chip_buf I91 ( .in(fsm_nv_bstream), .out(fsm_nv_bstream_buf));
ml_chip_buf I90 ( .in(tm_dma), .out(tm_dma_buf));
ml_chip_buf I92 ( .in(fsm_din), .out(fsm_din_buf));
ml_chip_buf I79_2_ ( .in(fsm_trim_rrefrd[2]),
     .out(fsm_trim_rrefrd_buf[2]));
ml_chip_buf I79_1_ ( .in(fsm_trim_rrefrd[1]),
     .out(fsm_trim_rrefrd_buf[1]));
ml_chip_buf I79_0_ ( .in(fsm_trim_rrefrd[0]),
     .out(fsm_trim_rrefrd_buf[0]));
ml_chip_buf I78 ( .in(fsm_vpxaset), .out(fsm_vpxaset_buf));
ml_chip_buf I77 ( .in(fsm_wpen), .out(fsm_wpen_buf));
ml_chip_buf I76_2_ ( .in(fsm_trim_rrefpgm[2]),
     .out(fsm_trim_rrefpgm_buf[2]));
ml_chip_buf I76_1_ ( .in(fsm_trim_rrefpgm[1]),
     .out(fsm_trim_rrefpgm_buf[1]));
ml_chip_buf I76_0_ ( .in(fsm_trim_rrefpgm[0]),
     .out(fsm_trim_rrefpgm_buf[0]));
ml_chip_buf I75 ( .in(fsm_sample), .out(fsm_sample_buf));
ml_chip_buf I74 ( .in(fsm_tm_testdec), .out(fsm_tm_testdec_buf));
ml_chip_buf I73_7_ ( .in(fsm_rowadd[7]), .out(fsm_rowadd_buf[7]));
ml_chip_buf I73_6_ ( .in(fsm_rowadd[6]), .out(fsm_rowadd_buf[6]));
ml_chip_buf I73_5_ ( .in(fsm_rowadd[5]), .out(fsm_rowadd_buf[5]));
ml_chip_buf I73_4_ ( .in(fsm_rowadd[4]), .out(fsm_rowadd_buf[4]));
ml_chip_buf I73_3_ ( .in(fsm_rowadd[3]), .out(fsm_rowadd_buf[3]));
ml_chip_buf I73_2_ ( .in(fsm_rowadd[2]), .out(fsm_rowadd_buf[2]));
ml_chip_buf I73_1_ ( .in(fsm_rowadd[1]), .out(fsm_rowadd_buf[1]));
ml_chip_buf I73_0_ ( .in(fsm_rowadd[0]), .out(fsm_rowadd_buf[0]));
ml_chip_buf I72 ( .in(fsm_tm_rd_mode), .out(fsm_tm_rd_mode_buf));
ml_chip_buf I71 ( .in(fsm_pgmien), .out(fsm_pgmien_buf));
ml_chip_buf I70 ( .in(fsm_rd), .out(fsm_rd_buf));
ml_chip_buf I69 ( .in(fsm_rst_b), .out(fsm_rst_b_buf));
ml_chip_buf I68 ( .in(fsm_nv_rri_trim), .out(fsm_nv_rri_trim_buf));
ml_chip_buf I63 ( .in(fsm_multibl_read), .out(fsm_multibl_read_buf));
ml_chip_buf I50_2_ ( .in(fsm_vpgmwl[2]), .out(fsm_vpgmwl_buf[2]));
ml_chip_buf I50_1_ ( .in(fsm_vpgmwl[1]), .out(fsm_vpgmwl_buf[1]));
ml_chip_buf I50_0_ ( .in(fsm_vpgmwl[0]), .out(fsm_vpgmwl_buf[0]));
ml_chip_buf I56 ( .in(fsm_wgnden), .out(fsm_wgnden_buf));
ml_chip_buf I49_3_ ( .in(fsm_trim_vbg[3]), .out(fsm_trim_vbg_buf[3]));
ml_chip_buf I49_2_ ( .in(fsm_trim_vbg[2]), .out(fsm_trim_vbg_buf[2]));
ml_chip_buf I49_1_ ( .in(fsm_trim_vbg[1]), .out(fsm_trim_vbg_buf[1]));
ml_chip_buf I49_0_ ( .in(fsm_trim_vbg[0]), .out(fsm_trim_vbg_buf[0]));
ml_chip_buf I51 ( .in(fsm_lshven), .out(fsm_lshven_buf));
ml_chip_buf I53 ( .in(fsm_nvcmen), .out(fsm_nvcmen_buf));
ml_chip_buf I54 ( .in(fsm_pgmdisc), .out(fsm_pgmdisc_buf));
ml_chip_buf I57 ( .in(fsm_pgmvfy), .out(fsm_pgmvfy_buf));
ml_chip_buf I55 ( .in(fsm_pgm), .out(fsm_pgm_buf));
ml_chip_buf I65_3_ ( .in(fsm_blkadd_b[3]), .out(fsm_blkadd_b_buf[3]));
ml_chip_buf I65_2_ ( .in(fsm_blkadd_b[2]), .out(fsm_blkadd_b_buf[2]));
ml_chip_buf I65_1_ ( .in(fsm_blkadd_b[1]), .out(fsm_blkadd_b_buf[1]));
ml_chip_buf I65_0_ ( .in(fsm_blkadd_b[0]), .out(fsm_blkadd_b_buf[0]));
ml_chip_buf I64_3_ ( .in(fsm_blkadd[3]), .out(fsm_blkadd_buf[3]));
ml_chip_buf I64_2_ ( .in(fsm_blkadd[2]), .out(fsm_blkadd_buf[2]));
ml_chip_buf I64_1_ ( .in(fsm_blkadd[1]), .out(fsm_blkadd_buf[1]));
ml_chip_buf I64_0_ ( .in(fsm_blkadd[0]), .out(fsm_blkadd_buf[0]));
ml_chip_buf I66_9_ ( .in(fsm_coladd[9]), .out(fsm_coladd_buf[9]));
ml_chip_buf I66_8_ ( .in(fsm_coladd[8]), .out(fsm_coladd_buf[8]));
ml_chip_buf I66_7_ ( .in(fsm_coladd[7]), .out(fsm_coladd_buf[7]));
ml_chip_buf I66_6_ ( .in(fsm_coladd[6]), .out(fsm_coladd_buf[6]));
ml_chip_buf I66_5_ ( .in(fsm_coladd[5]), .out(fsm_coladd_buf[5]));
ml_chip_buf I66_4_ ( .in(fsm_coladd[4]), .out(fsm_coladd_buf[4]));
ml_chip_buf I66_3_ ( .in(fsm_coladd[3]), .out(fsm_coladd_buf[3]));
ml_chip_buf I66_2_ ( .in(fsm_coladd[2]), .out(fsm_coladd_buf[2]));
ml_chip_buf I66_1_ ( .in(fsm_coladd[1]), .out(fsm_coladd_buf[1]));
ml_chip_buf I66_0_ ( .in(fsm_coladd[0]), .out(fsm_coladd_buf[0]));
ml_chip_buf I67 ( .in(fsm_nv_sisi_ui), .out(fsm_nv_sisi_ui_buf));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_spare_right, View - schematic
// LAST TIME SAVED: Sep 23 13:32:35 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_ctrl_spare_right (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:9]  net0260;



vdd_tielow I141_9_ ( .gnd_tiel(net0260[0]));
vdd_tielow I141_8_ ( .gnd_tiel(net0260[1]));
vdd_tielow I141_7_ ( .gnd_tiel(net0260[2]));
vdd_tielow I141_6_ ( .gnd_tiel(net0260[3]));
vdd_tielow I141_5_ ( .gnd_tiel(net0260[4]));
vdd_tielow I141_4_ ( .gnd_tiel(net0260[5]));
vdd_tielow I141_3_ ( .gnd_tiel(net0260[6]));
vdd_tielow I141_2_ ( .gnd_tiel(net0260[7]));
vdd_tielow I141_1_ ( .gnd_tiel(net0260[8]));
vdd_tielow I141_0_ ( .gnd_tiel(net0260[9]));
rppolywo_m  R1 ( .MINUS(net0257), .PLUS(net0280), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net302), .PLUS(net0283), .BULK(gnd_));
rppolywo_m  R2 ( .MINUS(net0254), .PLUS(net0277), .BULK(gnd_));
rppolywo_m  R5 ( .MINUS(net0249), .PLUS(net0268), .BULK(gnd_));
rppolywo_m  R6 ( .MINUS(net0246), .PLUS(net0265), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(net0245), .PLUS(net0262), .BULK(gnd_));

endmodule
// Library - io, Cell - PVDD1DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:14:35 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module PVDD1DGZ ( VDD );
input  VDD;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_core_ctrl_spare_left, View - schematic
// LAST TIME SAVED: Sep 17 13:53:07 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_ctrl_spare_left (  );supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nmoscap_25  C7 ( .MINUS(GND_), .PLUS(vddp_));
pch_25  M14 ( .D(net96), .B(net85), .G(net286), .S(net85));
pch_25  M5 ( .D(net85), .B(net123), .G(net114), .S(net123));
pch_25  M3 ( .D(net108), .B(net89), .G(net316), .S(net89));
pch_25  M2 ( .D(net89), .B(net126), .G(net119), .S(net126));
nch_25  M7 ( .D(net100), .B(GND_), .G(net286), .S(gnd_));
nch_25  M1 ( .D(net96), .B(GND_), .G(net121), .S(net100));
nch_25  M6 ( .D(net104), .B(GND_), .G(net316), .S(gnd_));
nch_25  M4 ( .D(net108), .B(GND_), .G(net121), .S(net104));
ml_hv_ls_inv I132 ( .sel_b_25(net316), .sel_25(net405),
     .out_b_hv(net119), .in_hv(net126), .vddp_tieh(net121));
ml_hv_ls_inv Iml_hv_ls_inv_vppt ( .sel_b_25(net286), .sel_25(net404),
     .out_b_hv(net114), .in_hv(net123), .vddp_tieh(net121));
rppolywo_m  R8 ( .MINUS(vddp_), .PLUS(net123), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(vddp_), .PLUS(net126), .BULK(gnd_));
rppolywo_m  R10 ( .MINUS(net0388), .PLUS(net0385), .BULK(gnd_));
rppolywo_m  R11 ( .MINUS(net0379), .PLUS(net0382), .BULK(gnd_));
rppolywo_m  R13 ( .MINUS(net0370), .PLUS(net0376), .BULK(gnd_));
rppolywo_m  R14 ( .MINUS(net0376), .PLUS(gnd_), .BULK(gnd_));
rppolywo_m  R15 ( .MINUS(net0367), .PLUS(net0370), .BULK(gnd_));
rppolywo_m  R16 ( .MINUS(net0382), .PLUS(net0367), .BULK(gnd_));
rppolywo_m  R9 ( .MINUS(gnd_), .PLUS(net0388), .BULK(gnd_));
rppolywo_m  R12 ( .MINUS(net0385), .PLUS(net0379), .BULK(gnd_));
nand3_25 I96 ( .B(net160), .A(net160), .Y(net168), .C(net160),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I45 ( .B(net168), .A(net168), .Y(net176), .C(net168),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I48 ( .B(net176), .A(net176), .Y(net184), .C(net176),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nand3_25 I53 ( .B(net184), .A(net184), .Y(net284), .C(net184),
     .P(vddp_), .Pb(vddp_), .Gb(gnd_), .G(gnd_));
nor3_25 I42 ( .B(net191), .A(net191), .C(net191), .Y(net160), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I78 ( .B(net199), .A(net199), .C(net199), .Y(net191), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I83 ( .B(net207), .A(net207), .C(net207), .Y(net199), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
nor3_25 I84 ( .B(net215), .A(net215), .C(net215), .Y(net207), .G(gnd_),
     .Gb(gnd_), .Pb(vddp_), .P(vddp_));
inv_hvt I120 ( .A(net253), .Y(net249));
inv_hvt I119 ( .A(net231), .Y(net253));
inv_hvt I118 ( .A(net231), .Y(net258));
inv_hvt I117 ( .A(net258), .Y(net254));
inv_hvt I319 ( .A(net263), .Y(net259));
inv_hvt I323 ( .A(net231), .Y(net263));
inv_hvt I57 ( .A(net231), .Y(net268));
inv_hvt I58 ( .A(net268), .Y(net264));
ml_ls_vdd2vdd25 I122 ( .in(net249), .sup(vddp_), .out_vddio_b(net291),
     .out_vddio(net252), .in_b(net253));
ml_ls_vdd2vdd25 I121 ( .in(net254), .sup(vddp_), .out_vddio_b(net297),
     .out_vddio(net257), .in_b(net258));
ml_ls_vdd2vdd25 I335 ( .in(net259), .sup(vddp_), .out_vddio_b(net303),
     .out_vddio(net262), .in_b(net263));
ml_ls_vdd2vdd25 I56 ( .in(net264), .sup(vddp_), .out_vddio_b(net309),
     .out_vddio(net267), .in_b(net268));
inv_25 I126 ( .IN(net291), .OUT(net271), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I125 ( .IN(net297), .OUT(net272), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I139 ( .IN(net405), .OUT(net316), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I114 ( .IN(net404), .OUT(net286), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I384 ( .IN(net303), .OUT(net274), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I54 ( .IN(net309), .OUT(net273), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nand3_hvt I246 ( .Y(net328), .B(net324), .C(net324), .A(net324));
nand3_hvt I61 ( .Y(net332), .B(net328), .C(net328), .A(net328));
nand3_hvt I62 ( .Y(net336), .B(net332), .C(net332), .A(net332));
nand3_hvt I63 ( .Y(net340), .B(net336), .C(net336), .A(net336));
nand3_hvt I64 ( .Y(net360), .B(net340), .C(net340), .A(net340));
nor3_hvt I65 ( .B(net363), .Y(net282), .A(net363), .C(net363));
nor3_hvt I70 ( .B(net367), .Y(net363), .A(net367), .C(net367));
nor3_hvt I71 ( .B(net371), .Y(net367), .A(net371), .C(net371));
nor3_hvt I72 ( .B(net375), .Y(net371), .A(net375), .C(net375));
nor3_hvt I73 ( .B(net379), .Y(net375), .A(net379), .C(net379));
vddp_tiehigh I140 ( .vddp_tieh(net121));
vdd_tielow I154 ( .gnd_tiel(net405));
vdd_tielow I155 ( .gnd_tiel(net404));
vdd_tielow I153 ( .gnd_tiel(net231));
vdd_tielow I146 ( .gnd_tiel(net215));
vdd_tielow I145 ( .gnd_tiel(net324));
vdd_tielow I144 ( .gnd_tiel(net379));

endmodule
// Library - sbtlibn65lp, Cell - ml_mux2_25, View - schematic
// LAST TIME SAVED: Aug  6 15:48:57 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_mux2_25 ( out_25, in_a_25, in_b_25, sel_a_25 );
output  out_25;

input  in_a_25, in_b_25, sel_a_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M10 ( .D(in_b_25), .B(vddp_), .G(sel_a_25), .S(out_25));
pch_25  M13 ( .D(in_a_25), .B(vddp_), .G(EN_B_25), .S(out_25));
nch_25  M14 ( .D(in_a_25), .B(GND_), .G(sel_a_25), .S(out_25));
nch_25  M12 ( .D(in_b_25), .B(GND_), .G(EN_B_25), .S(out_25));
inv_25 I156 ( .IN(sel_a_25), .OUT(EN_B_25), .P(vddp_), .Pb(vddp_),
     .G(GND_), .Gb(GND_));

endmodule
// Library - sbtlibn65lp, Cell - oai21x2_sup_25, View - schematic
// LAST TIME SAVED: Dec 18 17:40:05 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module oai21x2_sup_25 ( Y, A0, A1, B0, ysup_25 );
output  Y;

input  A0, A1, B0, ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(gnd_), .G(A0), .S(net024));
nch_25  M6 ( .D(Y), .B(gnd_), .G(A1), .S(net024));
nch_25  M7 ( .D(net024), .B(gnd_), .G(B0), .S(gnd_));
pch_25  M4 ( .D(Y), .B(ysup_25), .G(A0), .S(net017));
pch_25  M0 ( .D(net017), .B(ysup_25), .G(A1), .S(ysup_25));
pch_25  M5 ( .D(Y), .B(ysup_25), .G(B0), .S(ysup_25));

endmodule
// Library - tsmcN65lo, Cell - nor2_25, View - schematic
// LAST TIME SAVED: Mar 29 20:24:25 2006
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nor2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(Y), .B(Gb), .G(A), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(B), .S(G));
pch_25  PM1 ( .D(net15), .B(Pb), .G(A), .S(P));
pch_25  M0 ( .D(Y), .B(Pb), .G(B), .S(net15));

endmodule
// Library - NVCM, Cell - ml_ls_vdd25_nor2, View - schematic
// LAST TIME SAVED: Jan 12 15:33:21 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ls_vdd25_nor2 ( out_vddio, out_vddio_b, sup, in, in_b );
output  out_vddio, out_vddio_b;

inout  sup;

input  in, in_b;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_25 I79 ( .A(in), .Y(out_vddio_b), .Gb(gnd_), .G(gnd_), .Pb(sup),
     .P(sup), .B(out_vddio));
nor2_25 I151 ( .A(out_vddio_b), .Y(out_vddio), .Gb(gnd_), .G(gnd_),
     .Pb(sup), .P(sup), .B(in_b));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yptest, View - schematic
// LAST TIME SAVED: Feb 26 14:41:48 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yptest ( yp_test_25, yp_test_b_25, yp_test,
     yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25, ysup_25 );
output  yp_test_25, yp_test_b_25;

input  yp_test, yp_test_b_high_b_ysup_25, yp_test_b_low_ysup_25,
     ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



oai21x2_sup_25 I180 ( .A1(yp_test_b_low_ysup_25), .Y(yp_test_b_25),
     .A0(net37), .B0(yp_test_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(yp_test), .sup(ysup_25),
     .out_vddio_b(net028), .out_vddio(net37), .in_b(net40));
inv_hvt I181 ( .A(yp_test), .Y(net40));
inv_25 I182 ( .IN(net028), .OUT(yp_test_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yp3, View - schematic
// LAST TIME SAVED: Feb 26 14:41:31 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp3 ( yp3_25, yp3_b_25, yp3_b_high_b_ysup_25,
     yp3_b_low_ysup_25, yp3_sel, ysup_25 );
output  yp3_25, yp3_b_25;

input  yp3_b_high_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_hvt I201 ( .A(yp3_sel), .Y(net075));
inv_hvt I101 ( .A(net075), .Y(net070));
oai21x2_sup_25 I202 ( .A1(yp3_b_low_ysup_25), .Y(yp3_b_25),
     .A0(net069), .B0(yp3_b_high_b_ysup_25), .ysup_25(ysup_25));
ml_ls_vdd25_nor2 I192 ( .in(net070), .sup(ysup_25),
     .out_vddio_b(yp3_25_b), .out_vddio(net069), .in_b(net075));
inv_25 I204 ( .IN(yp3_25_b), .OUT(yp3_25), .P(ysup_25), .Pb(ysup_25),
     .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_yp21, View - schematic
// LAST TIME SAVED: Feb 26 14:41:20 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_yp21 ( yp21, yp21_b_25, yp21_b_low_b, yp21_sel,
     ysup_25 );
output  yp21, yp21_b_25;

input  yp21_b_low_b, yp21_sel, ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nand2_hvt I206 ( .A(yp21_sel_b), .Y(net50), .B(yp21_b_low_b));
inv_hvt I207 ( .A(net50), .Y(net68));
inv_hvt I208 ( .A(yp21_sel), .Y(yp21_sel_b));
inv_hvt I209 ( .A(yp21_sel_b), .Y(yp21));
ml_ls_vdd25_nor2 I194 ( .in(net68), .sup(ysup_25),
     .out_vddio_b(yp21_b_25_b), .out_vddio(net72), .in_b(net50));
inv_25 I213 ( .IN(yp21_b_25_b), .OUT(yp21_b_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));

endmodule
// Library - NVCM, Cell - ml_ymux_vblinhi_pgm_drv, View - schematic
// LAST TIME SAVED: Apr  8 10:44:07 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_vblinhi_pgm_drv ( vblinhi_pgm_25, ysup_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25 );
inout  vblinhi_pgm_25, ysup_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_na25  M13 ( .D(vdd_), .B(GND_), .G(en_blinhi_pgm_b_ysup_25),
     .S(vblinhi_pgm_25));
pch_25  M5 ( .D(net10), .B(ysup_25), .G(en_blinhi_pgm_b_ysup_25),
     .S(ysup_25));
pch_25  M0 ( .D(net10), .B(vblinhi_pgm_25), .G(en_blinhi_pgm_b),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_ctrl_8f, View - schematic
// LAST TIME SAVED: Jul 16 15:24:32 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_ctrl_8f ( yp1, yp1_b_25, yp2, yp2_b_25, yp3_25,
     yp3_b_25, yp_test_25, yp_test_b_25, vblinhi_pgm_25,
     en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b, yp1_sel,
     yp2_b_low_b, yp2_sel, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp3_sel, yp_test,
     yp_test_b_high_b, yp_test_b_low_b, ysup_25 );

inout  vblinhi_pgm_25;

input  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, yp1_b_low_b,
     yp2_b_low_b, yp3_b_high_even_b_ysup_25, yp3_b_high_odd_b_ysup_25,
     yp3_b_low_ysup_25, yp_test_b_high_b, yp_test_b_low_b, ysup_25;

output [7:0]  yp2;
output [10:0]  yp1;
output [1:0]  yp_test_b_25;
output [7:0]  yp3_25;
output [10:0]  yp1_b_25;
output [1:0]  yp_test_25;
output [7:0]  yp3_b_25;
output [7:0]  yp2_b_25;

input [7:0]  yp3_sel;
input [7:0]  yp2_sel;
input [1:0]  yp_test;
input [10:0]  yp1_sel;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_1_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1]), .yp_test(yp_test[1]),
     .yp_test_25(yp_test_25[1]));
ml_ymux_ctrl_yptest Iml_ymux_ctrl_yptest_0_ (
     .yp_test_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp_test_b_low_ysup_25(yp3_b_low_ysup_25), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[0]), .yp_test(yp_test[0]),
     .yp_test_25(yp_test_25[0]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_7_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[7]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[7]), .yp3_25(yp3_25[7]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_6_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[6]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[6]), .yp3_25(yp3_25[6]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_5_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[5]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[5]), .yp3_25(yp3_25[5]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_4_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[4]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[4]), .yp3_25(yp3_25[4]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_3_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[3]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[3]), .yp3_25(yp3_25[3]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_2_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[2]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[2]), .yp3_25(yp3_25[2]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_1_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[1]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[1]), .yp3_25(yp3_25[1]));
ml_ymux_ctrl_yp3 Iml_ymux_ctrl_yp3_0_ (
     .yp3_b_high_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25), .yp3_sel(yp3_sel[0]),
     .ysup_25(ysup_25), .yp3_b_25(yp3_b_25[0]), .yp3_25(yp3_25[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_7_ ( .yp21_sel(yp2_sel[7]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[7]), .yp21(yp2[7]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_6_ ( .yp21_sel(yp2_sel[6]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[6]), .yp21(yp2[6]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_5_ ( .yp21_sel(yp2_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[5]), .yp21(yp2[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_4_ ( .yp21_sel(yp2_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[4]), .yp21(yp2[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_3_ ( .yp21_sel(yp2_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[3]), .yp21(yp2[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_2_ ( .yp21_sel(yp2_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[2]), .yp21(yp2[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_1_ ( .yp21_sel(yp2_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[1]), .yp21(yp2[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp2_0_ ( .yp21_sel(yp2_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp2_b_low_b),
     .yp21_b_25(yp2_b_25[0]), .yp21(yp2[0]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_10_ ( .yp21_sel(yp1_sel[10]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[10]), .yp21(yp1[10]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_9_ ( .yp21_sel(yp1_sel[9]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[9]), .yp21(yp1[9]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_8_ ( .yp21_sel(yp1_sel[8]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[8]), .yp21(yp1[8]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_7_ ( .yp21_sel(yp1_sel[7]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[7]), .yp21(yp1[7]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_6_ ( .yp21_sel(yp1_sel[6]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[6]), .yp21(yp1[6]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_5_ ( .yp21_sel(yp1_sel[5]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[5]), .yp21(yp1[5]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_4_ ( .yp21_sel(yp1_sel[4]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[4]), .yp21(yp1[4]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_3_ ( .yp21_sel(yp1_sel[3]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[3]), .yp21(yp1[3]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_2_ ( .yp21_sel(yp1_sel[2]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[2]), .yp21(yp1[2]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_1_ ( .yp21_sel(yp1_sel[1]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[1]), .yp21(yp1[1]));
ml_ymux_ctrl_yp21 Iml_ymux_ctrl_yp1_0_ ( .yp21_sel(yp1_sel[0]),
     .ysup_25(ysup_25), .yp21_b_low_b(yp1_b_low_b),
     .yp21_b_25(yp1_b_25[0]), .yp21(yp1[0]));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_1_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_vblinhi_pgm_drv Iml_ymux_vblinhi_pgm_drv_0_ (
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_ysup_25),
     .ysup_25(ysup_25), .en_blinhi_pgm_b(en_blinhi_pgm_b),
     .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - io, Cell - PVDD2POC, View - schematic
// LAST TIME SAVED: Jul 28 17:15:17 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module PVDD2POC ( VDDPST );
input  VDDPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_pump_a_clkdly, View - schematic
// LAST TIME SAVED: Feb 11 09:24:13 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_pump_a_clkdly ( out, in );
output  out;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_hvt  M80 ( .D(vdd_), .B(vdd_), .G(net66), .S(vdd_));
pch_hvt  M0 ( .D(vdd_), .B(vdd_), .G(net62), .S(vdd_));
inv_hvt I206 ( .A(in), .Y(net66));
inv_hvt I204 ( .A(net64), .Y(net62));
inv_hvt I205 ( .A(net66), .Y(net64));
inv_hvt I207 ( .A(net70), .Y(out));
inv_hvt I208 ( .A(net62), .Y(net70));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_logic_8f_sbb, View - schematic
// LAST TIME SAVED: Jul 14 12:21:35 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_8f_sbb ( out_hv_winv, out_hv_woinv, in );
output  out_hv_winv, out_hv_woinv;

input  in;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I140 ( .A(net268), .B(in), .Y(net255));
nor2_hvt I128 ( .A(net264), .B(net270), .Y(net258));
inv_hvt I142 ( .A(net258), .Y(net266));
inv_hvt I134 ( .A(in), .Y(net264));
inv_hvt I143 ( .A(net255), .Y(net262));
ml_pump_a_clkdly I141 ( .in(net262), .out(net270));
ml_pump_a_clkdly I219 ( .in(net266), .out(net268));
ml_ls_vdd2vdd25 I144 ( .in(net266), .sup(vddp_),
     .out_vddio_b(out_hv_winv), .out_vddio(net279), .in_b(net258));
ml_ls_vdd2vdd25 I148 ( .in(net262), .sup(vddp_),
     .out_vddio_b(out_hv_woinv), .out_vddio(net274), .in_b(net255));

endmodule
// Library - sbtlibn65lp, Cell - oai2211x2_hvt, View - schematic
// LAST TIME SAVED: Jul 31 10:31:37 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module oai2211x2_hvt ( Y, A0, A1, B0, B1, C0, D0 );
output  Y;

input  A0, A1, B0, B1, C0, D0;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(net040), .B(GND_), .G(A0), .S(net024));
nch_hvt  M13 ( .D(net044), .B(GND_), .G(D0), .S(net040));
nch_hvt  M11 ( .D(Y), .B(GND_), .G(C0), .S(net044));
nch_hvt  M8 ( .D(net040), .B(GND_), .G(A1), .S(net024));
nch_hvt  M10 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M12 ( .D(Y), .B(VDD_), .G(D0), .S(vdd_));
pch_hvt  M7 ( .D(Y), .B(VDD_), .G(C0), .S(vdd_));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M4 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - sbtlibn65lp, Cell - anor31_hvt, View - schematic
// LAST TIME SAVED: Feb 13 14:15:10 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module anor31_hvt ( Y, A, B, C, D );
output  Y;

input  A, B, C, D;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M1 ( .D(Y), .B(gnd_), .G(A), .S(net23));
nch_hvt  M8 ( .D(net030), .B(gnd_), .G(C), .S(gnd_));
nch_hvt  M6 ( .D(net23), .B(gnd_), .G(B), .S(net030));
nch_hvt  M7 ( .D(Y), .B(gnd_), .G(D), .S(gnd_));
pch_hvt  M5 ( .D(Y), .B(vdd_), .G(D), .S(net35));
pch_hvt  M4 ( .D(net35), .B(vdd_), .G(A), .S(vdd_));
pch_hvt  M3 ( .D(net35), .B(vdd_), .G(B), .S(vdd_));
pch_hvt  M2 ( .D(net35), .B(vdd_), .G(C), .S(vdd_));

endmodule
// Library - sbtlibn65lp, Cell - oai22x2_hvt, View - schematic
// LAST TIME SAVED: Jan 24 13:53:38 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module oai22x2_hvt ( Y, A0, A1, B0, B1 );
output  Y;

input  A0, A1, B0, B1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_hvt  M2 ( .D(Y), .B(GND_), .G(A0), .S(net024));
nch_hvt  M8 ( .D(Y), .B(GND_), .G(A1), .S(net024));
nch_hvt  M10 ( .D(net024), .B(GND_), .G(B1), .S(gnd_));
nch_hvt  M9 ( .D(net024), .B(GND_), .G(B0), .S(gnd_));
pch_hvt  M3 ( .D(net017), .B(VDD_), .G(A1), .S(vdd_));
pch_hvt  M6 ( .D(Y), .B(VDD_), .G(B1), .S(net061));
pch_hvt  M4 ( .D(Y), .B(VDD_), .G(A0), .S(net017));
pch_hvt  M5 ( .D(net061), .B(VDD_), .G(B0), .S(vdd_));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_logic_8f, View - schematic
// LAST TIME SAVED: Jul 31 10:32:24 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_ctrl_logic_8f ( dec_trim, en_blinhi_pgm_b,
     en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa, sa_bl_to_pgm_glb,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25,
     sel_dec_l_25, yp1_sel, yp2_sel, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp3_sel,
     yp21_b_low_b, yp_test, fsm_blkadd, fsm_coladd, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h, fsm_tm_allwl_l,
     fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow, fsm_trim_rrefpgm,
     fsm_trim_rrefrd, fsm_vpxaset, fsm_wpen, fsm_ymuxdis,
     tm_allbank_sel, tm_tcol, ysup_25 );
output  en_blinhi_pgm_b, en_blinhi_pgm_b_ysup_25, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, sel_dec_l_25, yp3_b_high_even_b_ysup_25,
     yp3_b_high_odd_b_ysup_25, yp3_b_low_ysup_25, yp21_b_low_b;

input  fsm_lshven, fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow,
     fsm_nv_sisi_ui, fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy,
     fsm_rd, fsm_tm_allbl_h, fsm_tm_allbl_l, fsm_tm_allwl_h,
     fsm_tm_allwl_l, fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, tm_allbank_sel, tm_tcol,
     ysup_25;

output [7:5]  dec_trim;
output [3:0]  sb25_gnd_25;
output [3:0]  sbhv_high_25;
output [7:0]  yp3_sel;
output [7:0]  yp2_sel;
output [10:0]  yp1_sel;
output [3:0]  sb25_high_25;
output [3:0]  sbhv_gnd_25;
output [1:0]  yp_test;

input [9:0]  fsm_coladd;
input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [3:0]  fsm_blkadd;
input [2:0]  fsm_trim_rrefpgm;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp2_sel_b;

wire  [7:0]  yp3_sel_b;

wire  [7:5]  dec_trim_b;

wire  [2:0]  tdec_b;

wire  [2:0]  tdec;

wire  [3:0]  sb25low_b;

wire  [0:2]  net634;

wire  [1:0]  yp_test_b;

wire  [1:0]  xadd;

wire  [3:0]  sbhvlow_b;

wire  [1:0]  xadd_b;

wire  [10:0]  yp1_sel_b;

wire  [9:0]  yadd_b;

wire  [9:0]  yadd;

wire  [0:3]  net348;



ml_core_ctrl_logic_8f_sbb Isb25_3_ ( .in(sb25low_b[3]),
     .out_hv_woinv(sb25_gnd_25[3]), .out_hv_winv(sb25_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isb25_2_ ( .in(sb25low_b[2]),
     .out_hv_woinv(sb25_gnd_25[2]), .out_hv_winv(sb25_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isb25_1_ ( .in(sb25low_b[1]),
     .out_hv_woinv(sb25_gnd_25[1]), .out_hv_winv(sb25_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isb25_0_ ( .in(sb25low_b[0]),
     .out_hv_woinv(sb25_gnd_25[0]), .out_hv_winv(sb25_high_25[0]));
ml_core_ctrl_logic_8f_sbb Isbhv_3_ ( .in(sbhvlow_b[3]),
     .out_hv_woinv(sbhv_gnd_25[3]), .out_hv_winv(sbhv_high_25[3]));
ml_core_ctrl_logic_8f_sbb Isbhv_2_ ( .in(sbhvlow_b[2]),
     .out_hv_woinv(sbhv_gnd_25[2]), .out_hv_winv(sbhv_high_25[2]));
ml_core_ctrl_logic_8f_sbb Isbhv_1_ ( .in(sbhvlow_b[1]),
     .out_hv_woinv(sbhv_gnd_25[1]), .out_hv_winv(sbhv_high_25[1]));
ml_core_ctrl_logic_8f_sbb Isbhv_0_ ( .in(sbhvlow_b[0]),
     .out_hv_woinv(sbhv_gnd_25[0]), .out_hv_winv(sbhv_high_25[0]));
oai2211x2_hvt I86_3_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net570),
     .Y(yp1_sel_b[3]), .A0(yadd[7]), .B0(vddp_rd_overw), .B1(yadd[6]));
oai2211x2_hvt I86_2_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net570),
     .Y(yp1_sel_b[2]), .A0(yadd[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
oai2211x2_hvt I86_1_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net570),
     .Y(yp1_sel_b[1]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd[6]));
oai2211x2_hvt I86_0_ ( .D0(yadd_b[9]), .C0(yadd_b[8]), .A1(net570),
     .Y(yp1_sel_b[0]), .A0(yadd_b[7]), .B0(vddp_rd_overw),
     .B1(yadd_b[6]));
oai21x2 I36 ( .A1(fsm_pgmvfy), .A0(fsm_rd), .B0(net441),
     .Y(all_blk_sel_b));
vdd_tiehigh I198 ( .vdd_tieh(vdd_tieh));
exor2_hvt I151_3_ ( .A(net348[0]), .Y(sb25low_b[3]), .B(pgm_hvact_b));
exor2_hvt I151_2_ ( .A(net348[1]), .Y(sb25low_b[2]), .B(pgm_hvact_b));
exor2_hvt I151_1_ ( .A(net348[2]), .Y(sb25low_b[1]), .B(pgm_hvact_b));
exor2_hvt I151_0_ ( .A(net348[3]), .Y(sb25low_b[0]), .B(pgm_hvact_b));
anor21_hvt I119_1_ ( .A(fsm_rowadd[1]), .B(x1_desel_b), .Y(xadd_b[1]),
     .C(fsm_tm_trow));
anor21_hvt I119_0_ ( .A(fsm_rowadd[0]), .B(vdd_tieh), .Y(xadd_b[0]),
     .C(fsm_nv_sisi_ui));
anor21_hvt I109 ( .A(pgm_hvact), .B(fsm_tm_allwl_h), .Y(net410),
     .C(nvcmen_buf_b));
ml_ls_vdd2vdd25 I213 ( .in(net0556), .sup(vddp_),
     .out_vddio_b(sel_dec_l_25), .out_vddio(net0540), .in_b(net0397));
nor3_hvt I111 ( .B(fsm_tm_allbl_l), .Y(yp3_b_high_b),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_l));
nor3_hvt I112 ( .C(yp3_b_high_b), .A(nvcmen_buf_b), .B(fsm_tm_allbl_h),
     .Y(net340));
nor3_hvt I57 ( .C(fsm_tm_allbl_h), .A(fsm_tm_allbl_l),
     .B(fsm_tm_testdec), .Y(net344));
anor31_hvt I155_3_ ( .A(ensb25_dec), .D(net411), .B(xadd[1]),
     .Y(net348[0]), .C(xadd[0]));
anor31_hvt I155_2_ ( .A(ensb25_dec), .D(net411), .B(xadd[1]),
     .Y(net348[1]), .C(xadd_b[0]));
anor31_hvt I155_1_ ( .A(ensb25_dec), .D(net411), .B(xadd_b[1]),
     .Y(net348[2]), .C(xadd[0]));
anor31_hvt I155_0_ ( .A(ensb25_dec), .D(net411), .B(xadd_b[1]),
     .Y(net348[3]), .C(xadd_b[0]));
anor31_hvt I121_3_ ( .A(net413), .D(net415), .B(xadd[1]),
     .Y(sbhvlow_b[3]), .C(xadd[0]));
anor31_hvt I121_2_ ( .A(net413), .D(net415), .B(xadd[1]),
     .Y(sbhvlow_b[2]), .C(xadd_b[0]));
anor31_hvt I121_1_ ( .A(net413), .D(net415), .B(xadd_b[1]),
     .Y(sbhvlow_b[1]), .C(xadd[0]));
anor31_hvt I121_0_ ( .A(net413), .D(net415), .B(xadd_b[1]),
     .Y(sbhvlow_b[0]), .C(xadd_b[0]));
anor31_hvt I107 ( .A(fsm_tm_testdec), .D(net340), .B(nvcmen_buf),
     .Y(net358), .C(yadd[0]));
anor31_hvt I108 ( .A(fsm_tm_testdec), .D(net340), .B(nvcmen_buf),
     .Y(net363), .C(yadd_b[0]));
oai22x2_hvt I93 ( .A1(net397), .Y(net366), .A0(net469),
     .B0(fsm_nv_rri_trim), .B1(fsm_nv_sisi_ui));
nand4_hvt I210_10_ ( .D(yadd_b[6]), .A(yadd[9]), .C(yadd[7]),
     .Y(yp1_sel_b[10]), .B(yadd_b[8]));
nand4_hvt I210_9_ ( .D(yadd[6]), .A(yadd[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[9]), .B(yadd_b[8]));
nand4_hvt I210_8_ ( .D(yadd_b[6]), .A(yadd[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[8]), .B(yadd_b[8]));
nand4_hvt I210_7_ ( .D(yadd[6]), .A(yadd_b[9]), .C(yadd[7]),
     .Y(yp1_sel_b[7]), .B(yadd[8]));
nand4_hvt I210_6_ ( .D(yadd_b[6]), .A(yadd_b[9]), .C(yadd[7]),
     .Y(yp1_sel_b[6]), .B(yadd[8]));
nand4_hvt I210_5_ ( .D(yadd[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[5]), .B(yadd[8]));
nand4_hvt I210_4_ ( .D(yadd_b[6]), .A(yadd_b[9]), .C(yadd_b[7]),
     .Y(yp1_sel_b[4]), .B(yadd[8]));
nand4_hvt I122 ( .D(fsm_lshven), .C(pgm_hvact), .A(tm_allwl_l_b),
     .Y(net412), .B(blk_dec));
nand4_hvt I49_7_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[7]), .B(yadd[2]));
nand4_hvt I49_6_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[6]), .B(yadd[2]));
nand4_hvt I49_5_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[5]), .B(yadd[2]));
nand4_hvt I49_4_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[4]), .B(yadd[2]));
nand4_hvt I49_3_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[3]), .B(yadd_b[2]));
nand4_hvt I49_2_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd[1]),
     .Y(yp3_sel_b[2]), .B(yadd_b[2]));
nand4_hvt I49_1_ ( .D(yadd[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[1]), .B(yadd_b[2]));
nand4_hvt I49_0_ ( .D(yadd_b[0]), .A(ymux_en_core), .C(yadd_b[1]),
     .Y(yp3_sel_b[0]), .B(yadd_b[2]));
nand4_hvt I27 ( .D(fsm_blkadd[0]), .Y(blk_dec_b), .B(fsm_blkadd[2]),
     .C(fsm_blkadd[1]), .A(fsm_blkadd[3]));
inv_hvt I207 ( .A(net576), .Y(ref_pgm));
inv_hvt I200 ( .A(fsm_tm_testdec), .Y(net393));
inv_hvt I120_1_ ( .A(xadd_b[1]), .Y(xadd[1]));
inv_hvt I120_0_ ( .A(xadd_b[0]), .Y(xadd[0]));
inv_hvt I181 ( .A(all_blk_sel_b), .Y(net397));
inv_hvt I161 ( .A(net578), .Y(net399));
inv_hvt I158 ( .A(pgm_hvact_b), .Y(pgm_hvact));
inv_hvt I157 ( .A(fsm_pgmvfy), .Y(net405));
inv_hvt I160 ( .A(net410), .Y(net411));
inv_hvt I123 ( .A(net412), .Y(net413));
inv_hvt I125 ( .A(net498), .Y(net415));
inv_hvt I189 ( .A(fsm_nvcmen), .Y(nvcmen_buf_b));
inv_hvt I164 ( .A(net418), .Y(net419));
inv_hvt I224 ( .A(tm_allbank_sel), .Y(tm_pgm_rd_allblk_n));
inv_hvt I131 ( .A(fsm_tm_allwl_l), .Y(tm_allwl_l_b));
inv_hvt I218 ( .A(net0556), .Y(net0397));
inv_hvt I97 ( .A(fsm_multibl_read), .Y(net429));
inv_hvt I94 ( .A(net366), .Y(vddp_rd_overw));
inv_hvt I84 ( .A(nvcmen_buf_b), .Y(nvcmen_buf));
inv_hvt I72_7_ ( .A(yp2_sel_b[7]), .Y(yp2_sel[7]));
inv_hvt I72_6_ ( .A(yp2_sel_b[6]), .Y(yp2_sel[6]));
inv_hvt I72_5_ ( .A(yp2_sel_b[5]), .Y(yp2_sel[5]));
inv_hvt I72_4_ ( .A(yp2_sel_b[4]), .Y(yp2_sel[4]));
inv_hvt I72_3_ ( .A(yp2_sel_b[3]), .Y(yp2_sel[3]));
inv_hvt I72_2_ ( .A(yp2_sel_b[2]), .Y(yp2_sel[2]));
inv_hvt I72_1_ ( .A(yp2_sel_b[1]), .Y(yp2_sel[1]));
inv_hvt I72_0_ ( .A(yp2_sel_b[0]), .Y(yp2_sel[0]));
inv_hvt I66 ( .A(net358), .Y(net627));
inv_hvt I46_9_ ( .A(fsm_coladd[9]), .Y(yadd_b[9]));
inv_hvt I46_8_ ( .A(fsm_coladd[8]), .Y(yadd_b[8]));
inv_hvt I46_7_ ( .A(fsm_coladd[7]), .Y(yadd_b[7]));
inv_hvt I46_6_ ( .A(fsm_coladd[6]), .Y(yadd_b[6]));
inv_hvt I46_5_ ( .A(fsm_coladd[5]), .Y(yadd_b[5]));
inv_hvt I46_4_ ( .A(fsm_coladd[4]), .Y(yadd_b[4]));
inv_hvt I46_3_ ( .A(fsm_coladd[3]), .Y(yadd_b[3]));
inv_hvt I46_2_ ( .A(fsm_coladd[2]), .Y(yadd_b[2]));
inv_hvt I46_1_ ( .A(fsm_coladd[1]), .Y(yadd_b[1]));
inv_hvt I46_0_ ( .A(fsm_coladd[0]), .Y(yadd_b[0]));
inv_hvt I201 ( .A(fsm_tm_rd_mode), .Y(net441));
inv_hvt I25_2_ ( .A(tdec_b[2]), .Y(tdec[2]));
inv_hvt I25_1_ ( .A(tdec_b[1]), .Y(tdec[1]));
inv_hvt I25_0_ ( .A(tdec_b[0]), .Y(tdec[0]));
inv_hvt I24_2_ ( .A(net634[0]), .Y(tdec_b[2]));
inv_hvt I24_1_ ( .A(net634[1]), .Y(tdec_b[1]));
inv_hvt I24_0_ ( .A(net634[2]), .Y(tdec_b[0]));
inv_hvt I38_7_ ( .A(dec_trim_b[7]), .Y(dec_trim[7]));
inv_hvt I38_6_ ( .A(dec_trim_b[6]), .Y(dec_trim[6]));
inv_hvt I38_5_ ( .A(dec_trim_b[5]), .Y(dec_trim[5]));
inv_hvt I40 ( .A(net596), .Y(sa_bl_to_pgm_glb));
inv_hvt I103 ( .A(net519), .Y(en_blinhi_pgm_b));
inv_hvt I47_9_ ( .A(yadd_b[9]), .Y(yadd[9]));
inv_hvt I47_8_ ( .A(yadd_b[8]), .Y(yadd[8]));
inv_hvt I47_7_ ( .A(yadd_b[7]), .Y(yadd[7]));
inv_hvt I47_6_ ( .A(yadd_b[6]), .Y(yadd[6]));
inv_hvt I47_5_ ( .A(yadd_b[5]), .Y(yadd[5]));
inv_hvt I47_4_ ( .A(yadd_b[4]), .Y(yadd[4]));
inv_hvt I47_3_ ( .A(yadd_b[3]), .Y(yadd[3]));
inv_hvt I47_2_ ( .A(yadd_b[2]), .Y(yadd[2]));
inv_hvt I47_1_ ( .A(yadd_b[1]), .Y(yadd[1]));
inv_hvt I47_0_ ( .A(yadd_b[0]), .Y(yadd[0]));
inv_hvt I71 ( .A(net508), .Y(yp21_b_low_b));
inv_hvt I51_7_ ( .A(yp3_sel_b[7]), .Y(yp3_sel[7]));
inv_hvt I51_6_ ( .A(yp3_sel_b[6]), .Y(yp3_sel[6]));
inv_hvt I51_5_ ( .A(yp3_sel_b[5]), .Y(yp3_sel[5]));
inv_hvt I51_4_ ( .A(yp3_sel_b[4]), .Y(yp3_sel[4]));
inv_hvt I51_3_ ( .A(yp3_sel_b[3]), .Y(yp3_sel[3]));
inv_hvt I51_2_ ( .A(yp3_sel_b[2]), .Y(yp3_sel[2]));
inv_hvt I51_1_ ( .A(yp3_sel_b[1]), .Y(yp3_sel[1]));
inv_hvt I51_0_ ( .A(yp3_sel_b[0]), .Y(yp3_sel[0]));
inv_hvt I61 ( .A(net599), .Y(net459));
inv_hvt I69 ( .A(net363), .Y(net617));
inv_hvt I117_1_ ( .A(yp_test_b[1]), .Y(yp_test[1]));
inv_hvt I117_0_ ( .A(yp_test_b[0]), .Y(yp_test[0]));
inv_hvt I185 ( .A(tm_tcol), .Y(net467));
inv_hvt I90 ( .A(net567), .Y(net469));
inv_25 I104 ( .IN(net611), .OUT(en_blinhi_pgm_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net625), .OUT(yp3_b_high_even_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I79 ( .IN(net615), .OUT(yp3_b_high_odd_b_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
inv_25 I77 ( .IN(net620), .OUT(yp3_b_low_ysup_25), .P(ysup_25),
     .Pb(ysup_25), .G(gnd_), .Gb(gnd_));
nand3_hvt I156 ( .Y(pgm_hvact_b), .B(fsm_pgm), .C(net405),
     .A(fsm_lshven));
nand3_hvt I127 ( .Y(net498), .B(pgm_hvact), .C(fsm_tm_allwl_h),
     .A(fsm_lshven));
nand3_hvt I163 ( .C(tm_allwl_l_b), .A(fsm_vpxaset), .Y(net418),
     .B(sa_bl_to_blsa));
nand3_hvt I215 ( .Y(net0502), .B(yp1_sel_b[1]), .C(yp1_sel_b[2]),
     .A(yp1_sel_b[0]));
nand3_hvt I70 ( .C(nvcmen_buf), .A(net593), .Y(net508), .B(net393));
nand3_hvt I37_7_ ( .Y(dec_trim_b[7]), .B(tdec[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I37_6_ ( .Y(dec_trim_b[6]), .B(tdec[1]), .C(tdec_b[0]),
     .A(tdec[2]));
nand3_hvt I37_5_ ( .Y(dec_trim_b[5]), .B(tdec_b[1]), .C(tdec[0]),
     .A(tdec[2]));
nand3_hvt I73_7_ ( .A(yadd[5]), .C(yadd[3]), .Y(yp2_sel_b[7]),
     .B(yadd[4]));
nand3_hvt I73_6_ ( .A(yadd[5]), .C(yadd_b[3]), .Y(yp2_sel_b[6]),
     .B(yadd[4]));
nand3_hvt I73_5_ ( .A(yadd[5]), .C(yadd[3]), .Y(yp2_sel_b[5]),
     .B(yadd_b[4]));
nand3_hvt I73_4_ ( .A(yadd[5]), .C(yadd_b[3]), .Y(yp2_sel_b[4]),
     .B(yadd_b[4]));
nand3_hvt I73_3_ ( .A(yadd_b[5]), .C(yadd[3]), .Y(yp2_sel_b[3]),
     .B(yadd[4]));
nand3_hvt I73_2_ ( .A(yadd_b[5]), .C(yadd_b[3]), .Y(yp2_sel_b[2]),
     .B(yadd[4]));
nand3_hvt I73_1_ ( .A(yadd_b[5]), .C(yadd[3]), .Y(yp2_sel_b[1]),
     .B(yadd_b[4]));
nand3_hvt I73_0_ ( .A(yadd_b[5]), .C(yadd_b[3]), .Y(yp2_sel_b[0]),
     .B(yadd_b[4]));
nor4_hvt I98 ( .B(fsm_tm_allbl_l), .Y(net519), .D(nvcmen_buf_b),
     .A(net581), .C(fsm_tm_allbl_l));
nor4_hvt I52 ( .D(net588), .B(fsm_tm_allbl_h), .Y(ymux_dis_b),
     .A(fsm_tm_allbl_l), .C(fsm_tm_allbl_h));
nor2_hvt I211_10_ ( .A(tm_tcol), .B(yp1_sel_b[10]), .Y(yp1_sel[10]));
nor2_hvt I211_9_ ( .A(tm_tcol), .B(yp1_sel_b[9]), .Y(yp1_sel[9]));
nor2_hvt I211_8_ ( .A(tm_tcol), .B(yp1_sel_b[8]), .Y(yp1_sel[8]));
nor2_hvt I211_7_ ( .A(tm_tcol), .B(yp1_sel_b[7]), .Y(yp1_sel[7]));
nor2_hvt I211_6_ ( .A(tm_tcol), .B(yp1_sel_b[6]), .Y(yp1_sel[6]));
nor2_hvt I211_5_ ( .A(tm_tcol), .B(yp1_sel_b[5]), .Y(yp1_sel[5]));
nor2_hvt I211_4_ ( .A(tm_tcol), .B(yp1_sel_b[4]), .Y(yp1_sel[4]));
nor2_hvt I195 ( .A(fsm_nv_rri_trim), .B(fsm_nv_sisi_ui),
     .Y(x1_desel_b));
nor2_hvt I217 ( .A(net0502), .B(net0594), .Y(net0556));
nor2_hvt I114 ( .A(tm_tcol), .B(net605), .Y(ymux_en_core));
nor2_hvt I186 ( .A(net467), .B(net605), .Y(ymux_test_en));
nor2_hvt I88 ( .A(fsm_tm_rd_mode), .B(fsm_pgmvfy), .Y(net567));
nor2_hvt I96 ( .A(net366), .B(net429), .Y(net570));
nor2_hvt I75_3_ ( .A(yp1_sel_b[3]), .B(tm_tcol), .Y(yp1_sel[3]));
nor2_hvt I75_2_ ( .A(yp1_sel_b[2]), .B(tm_tcol), .Y(yp1_sel[2]));
nor2_hvt I75_1_ ( .A(yp1_sel_b[1]), .B(tm_tcol), .Y(yp1_sel[1]));
nor2_hvt I75_0_ ( .A(yp1_sel_b[0]), .B(tm_tcol), .Y(yp1_sel[0]));
nor2_hvt I206 ( .A(fsm_pgmvfy), .B(fsm_pgm), .Y(net576));
nand2_hvt I221 ( .A(blk_dec_b), .Y(blk_dec), .B(tm_pgm_rd_allblk_n));
nand2_hvt I162 ( .A(blk_dec), .Y(net578), .B(tm_allwl_l_b));
nand2_hvt I101 ( .A(pgm_hvact), .Y(net581), .B(pgm_hvact));
nand2_hvt I35 ( .B(one_blk_sel_b), .Y(sa_bl_to_blsa),
     .A(all_blk_sel_b));
nand2_hvt I216 ( .A(yp1_sel_b[4]), .Y(net0594), .B(yp1_sel_b[3]));
nand2_hvt I53 ( .A(fsm_nvcmen), .B(fsm_lshven), .Y(net588));
nand2_hvt I116_1_ ( .A(yadd[0]), .Y(yp_test_b[1]), .B(ymux_test_en));
nand2_hvt I116_0_ ( .A(yadd_b[0]), .Y(yp_test_b[0]), .B(ymux_test_en));
nand2_hvt I59 ( .A(fsm_lshven), .Y(net593), .B(pgm_hvact));
nand2_hvt I39 ( .A(blk_dec), .Y(net596), .B(fsm_pgmien));
nand2_hvt I60 ( .A(net593), .Y(net599), .B(net344));
nand2_hvt I89 ( .A(fsm_tm_rd_mode), .Y(one_blk_sel_b), .B(blk_dec));
oai21x2_hvt I55 ( .A1(sa_bl_to_blsa), .Y(net605), .A0(blk_dec),
     .B0(ymux_dis_b));
ml_ls_vdd25_nor2 I106 ( .in(net519), .sup(ysup_25),
     .out_vddio_b(net610), .out_vddio(net611), .in_b(en_blinhi_pgm_b));
ml_ls_vdd25_nor2 I68 ( .in(net363), .sup(ysup_25),
     .out_vddio_b(net615), .out_vddio(net616), .in_b(net617));
ml_ls_vdd25_nor2 I192 ( .in(net599), .sup(ysup_25),
     .out_vddio_b(net620), .out_vddio(net621), .in_b(net459));
ml_ls_vdd25_nor2 I65 ( .in(net358), .sup(ysup_25),
     .out_vddio_b(net625), .out_vddio(net626), .in_b(net627));
mux2_hvt I152 ( .in1(net399), .in0(net419), .out(ensb25_dec),
     .sel(pgm_hvact));
mux2_hvt I133_2_ ( .in1(fsm_trim_rrefpgm[2]), .in0(fsm_trim_rrefrd[2]),
     .out(net634[0]), .sel(ref_pgm));
mux2_hvt I133_1_ ( .in1(fsm_trim_rrefpgm[1]), .in0(fsm_trim_rrefrd[1]),
     .out(net634[1]), .sel(ref_pgm));
mux2_hvt I133_0_ ( .in1(fsm_trim_rrefpgm[0]), .in0(fsm_trim_rrefrd[0]),
     .out(net634[2]), .sel(ref_pgm));

endmodule
// Library - NVCM, Cell - ml_core_sa_resbot_m2, View - schematic
// LAST TIME SAVED: Sep 11 10:45:00 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_sa_resbot_m2 ( bl_in, bl_out, div_2r, div_3r, nwell,
     sa_ngate_25, sa_pgate_vpxa );
inout  bl_in, bl_out, div_2r, div_3r, nwell;


input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M4 ( .D(net115), .B(gnd_), .G(sa_ngate_25[4]), .S(bl_out));
nch_25  M3 ( .D(net090), .B(gnd_), .G(sa_ngate_25[3]), .S(net115));
nch_25  M0 ( .D(net086), .B(gnd_), .G(sa_ngate_25[2]), .S(net090));
nch_25  M32 ( .D(net111), .B(gnd_), .G(sa_ngate_25[1]), .S(net086));
pch_25  M5 ( .D(bl_out), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net115));
pch_25  M1 ( .D(net090), .B(nwell), .G(sa_pgate_vpxa[2]), .S(net086));
pch_25  M2 ( .D(net115), .B(nwell), .G(sa_pgate_vpxa[3]), .S(net090));
pch_25  M37 ( .D(net086), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net111));
rppolywo_m  R31 ( .MINUS(net099), .PLUS(div_3r), .BULK(gnd_));
rppolywo_m  R32 ( .MINUS(div_2r), .PLUS(net099), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(div_3r), .PLUS(net111), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net111), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R30 ( .MINUS(net0111), .PLUS(div_2r), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(net0111), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_rock_gwlgnd_nor2, View - schematic
// LAST TIME SAVED: Jan 23 10:17:03 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_rock_gwlgnd_nor2 ( gwl_gnd_25, gwl_b_sup_25, gwl_b_25,
     gwl_b_gnden_25 );
output  gwl_gnd_25;

inout  gwl_b_sup_25;

input  gwl_b_25, gwl_b_gnden_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(net14), .B(GND_), .G(gwl_b_gnden_25), .S(GND_));
nch_25  M0 ( .D(gwl_gnd_25), .B(GND_), .G(gwl_b_25), .S(net14));
pch_25  M2 ( .D(gwl_gnd_25), .B(gwl_b_sup_25), .G(gwl_b_25),
     .S(gwl_b_sup_25));

endmodule
// Library - NVCM, Cell - ml_core_sa_refres, View - schematic
// LAST TIME SAVED: Sep 11 10:40:27 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_sa_refres ( bot, nwell, wp_ref, sa_ngate_25,
     sa_pgate_vpxa );
inout  bot, nwell, wp_ref;


input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M32 ( .D(net44), .B(gnd_), .G(sa_ngate_25[1]), .S(net40));
nch_25  M2 ( .D(net50), .B(gnd_), .G(sa_ngate_25[3]), .S(net084));
nch_25  M6 ( .D(net084), .B(gnd_), .G(sa_ngate_25[4]), .S(bot));
nch_25  M1 ( .D(net40), .B(gnd_), .G(sa_ngate_25[2]), .S(net50));
pch_25  M3 ( .D(net084), .B(nwell), .G(sa_pgate_vpxa[3]), .S(net50));
pch_25  M37 ( .D(net40), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net44));
pch_25  M5 ( .D(bot), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net084));
pch_25  M0 ( .D(net50), .B(nwell), .G(sa_pgate_vpxa[2]), .S(net40));
rppolywo_m  R2 ( .MINUS(net096), .PLUS(net090), .BULK(gnd_));
rppolywo_m  R7 ( .MINUS(bot), .PLUS(net32), .BULK(gnd_));
rppolywo_m  R6 ( .MINUS(net32), .PLUS(net096), .BULK(gnd_));
rppolywo_m  R1 ( .MINUS(net090), .PLUS(net44), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net44), .PLUS(wp_ref), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_resbot, View - schematic
// LAST TIME SAVED: Apr  9 15:18:14 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_sa_resbot ( bl_in, bl_out, div_2r, div_3r, nwell,
     sa_ngate_25, sa_pgate_vpxa );
inout  bl_in, bl_out, div_2r, div_3r, nwell;


input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M4 ( .D(net115), .B(gnd_), .G(sa_ngate_25[4]), .S(bl_out));
nch_25  M3 ( .D(div_2r), .B(gnd_), .G(sa_ngate_25[3]), .S(net115));
nch_25  M0 ( .D(div_3r), .B(gnd_), .G(sa_ngate_25[2]), .S(div_2r));
nch_25  M32 ( .D(net111), .B(gnd_), .G(sa_ngate_25[1]), .S(div_3r));
pch_25  M5 ( .D(bl_out), .B(nwell), .G(sa_pgate_vpxa[4]), .S(net115));
pch_25  M1 ( .D(div_2r), .B(nwell), .G(sa_pgate_vpxa[2]), .S(div_3r));
pch_25  M2 ( .D(net115), .B(nwell), .G(sa_pgate_vpxa[3]), .S(div_2r));
pch_25  M37 ( .D(div_3r), .B(nwell), .G(sa_pgate_vpxa[1]), .S(net111));
rppolywo_m  R31 ( .MINUS(net099), .PLUS(div_3r), .BULK(gnd_));
rppolywo_m  R32 ( .MINUS(div_2r), .PLUS(net099), .BULK(gnd_));
rppolywo_m  R18 ( .MINUS(div_3r), .PLUS(net111), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net111), .PLUS(bl_in), .BULK(gnd_));
rppolywo_m  R30 ( .MINUS(net115), .PLUS(div_2r), .BULK(gnd_));
rppolywo_m  R24 ( .MINUS(bl_out), .PLUS(net115), .BULK(gnd_));

endmodule
// Library - io, Cell - PVDD2DGZ, View - schematic
// LAST TIME SAVED: Jul 28 17:14:57 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module PVDD2DGZ ( VDDPST );
input  VDDPST;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;




endmodule
// Library - NVCM, Cell - ml_rock_lwldrv_wp, View - schematic
// LAST TIME SAVED: Jan 21 10:22:42 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_rock_lwldrv_wp ( wp, ngate_25, gwl_b_25, gwl_gnd_25, gwp_hv,
     s_b_25, s_b_hv );
output  wp;

inout  ngate_25;

input  gwl_b_25, gwl_gnd_25, gwp_hv, s_b_25, s_b_hv;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M6 ( .D(wp), .B(gwp_hv), .G(s_b_hv), .S(gwp_hv));
nch_25  M11 ( .D(net18), .B(GND_), .G(s_b_25), .S(gwl_gnd_25));
nch_25  M12 ( .D(wp), .B(GND_), .G(ngate_25), .S(net18));
nch_25  M10 ( .D(net18), .B(GND_), .G(gwl_b_25), .S(gwl_gnd_25));

endmodule
// Library - sbtlibn65lp, Cell - ml_dff, View - schematic
// LAST TIME SAVED: Aug  3 14:03:13 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module sbtlibn65lp_ml_dff_schematic ( Q, QN, CLK, D, R );
output  Q, QN;

input  CLK, D, R;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nor2_hvt I129 ( .A(net057), .B(R), .Y(net052));
nor2_hvt I125 ( .A(net028), .B(R), .Y(net035));
inv_tri_2_hvt I128 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net028));
inv_tri_2_hvt I130 ( .Tb(clk_buf), .T(clk_b), .A(net052), .Y(net057));
inv_tri_2_hvt I127 ( .Tb(clk_b), .T(clk_buf), .A(net035), .Y(net057));
inv_tri_2_hvt I124 ( .Tb(clk_buf), .T(clk_b), .A(D), .Y(net028));
inv_hvt I146 ( .A(net057), .Y(Q));
inv_hvt I147 ( .A(net052), .Y(QN));
inv_hvt I131 ( .A(CLK), .Y(clk_b));
inv_hvt I132 ( .A(clk_b), .Y(clk_buf));

endmodule
// Library - tsmcN65lo, Cell - nand2_25, View - schematic
// LAST TIME SAVED: Mar 29 20:17:19 2006
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nand2_25 ( Y, A, B, G, Gb, P, Pb );
output  Y;

input  A, B, G, Gb, P, Pb;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .D(net16), .B(Gb), .G(B), .S(G));
nch_25  NM1 ( .D(Y), .B(Gb), .G(A), .S(net16));
pch_25  M2 ( .D(Y), .B(Pb), .G(B), .S(P));
pch_25  PM1 ( .D(Y), .B(Pb), .G(A), .S(P));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp, View - schematic
// LAST TIME SAVED: Jan 21 17:21:12 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp ( out_div, out_ref, in_div, in_ref, sa_bias,
     saen_b_25 );
output  out_div, out_ref;

input  in_div, in_ref, sa_bias, saen_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M4_1_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(net65), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M0 ( .D(out_div), .B(vddp_), .G(in_div), .S(net65));
pch_25  M3 ( .D(out_ref), .B(vddp_), .G(in_ref), .S(net65));
nch_25  M1 ( .D(out_ref), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M2 ( .D(out_div), .B(GND_), .G(out_ref), .S(gnd_));
nch_25  M8 ( .D(out_ref), .B(GND_), .G(saen_b_25), .S(gnd_));
nch_25  M5 ( .D(out_div), .B(GND_), .G(saen_b_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa_comp_top, View - schematic
// LAST TIME SAVED: Jan 21 17:21:37 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_sa_comp_top ( sa_out, in_div, in_ref, saen_25 );
output  sa_out;

input  in_div, in_ref, saen_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I85 ( .IN(saen_25), .OUT(saen_b_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I38 ( .IN(sa_out_b_25), .OUT(net051), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I82 ( .IN(net038), .OUT(sa_out), .P(vdd_), .Pb(vdd_), .G(gnd_),
     .Gb(gnd_));
nand2_25 I80 ( .G(gnd_), .Pb(vdd_), .A(net051), .Y(net038), .P(vdd_),
     .B(saen_25), .Gb(gnd_));
nand2_25 I96 ( .G(gnd_), .Pb(vddp_), .A(out_div2), .Y(sa_out_b_25),
     .P(vddp_), .B(saen_25), .Gb(gnd_));
ml_core_sa_comp Icore_sa_comp0 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref), .in_div(in_div),
     .out_ref(in_ref2), .out_div(in_div2));
ml_core_sa_comp Icore_sa_comp1 ( .saen_b_25(saen_b_25),
     .sa_bias(sa_bias), .in_ref(in_ref2), .in_div(in_div2),
     .out_ref(net73), .out_div(out_div2));
nch_25  M0 ( .D(net039), .B(gnd_), .G(saen_25), .S(gnd_));
pch_25  M43 ( .D(sa_bias), .B(vddp_), .G(saen_25), .S(vddp_));
pch_25  M4_4_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_3_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_2_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_1_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
pch_25  M4_0_ ( .D(sa_bias), .B(vddp_), .G(sa_bias), .S(vddp_));
rppolywo_m  R0 ( .MINUS(net039), .PLUS(net45), .BULK(gnd_));
rppolywo_m  R17 ( .MINUS(net45), .PLUS(sa_bias), .BULK(gnd_));

endmodule
// Library - NVCM, Cell - ml_core_sa, View - schematic
// LAST TIME SAVED: Sep 12 16:00:47 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_sa ( nv_dataout, blsa, vpxa, dec_ok_25, dec_trim,
     fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, tm_testdec_wr );
output  nv_dataout;

inout  blsa, vpxa;

input  dec_ok_25, fsm_rst_b, fsm_sample, fsm_tm_testdec, saen_25,
     saen_b_vpxa, testdec_en_b_25, tm_testdec_wr;

input [4:1]  sa_pgate_vpxa;
input [4:1]  sa_ngate_25;
input [7:5]  dec_trim;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_core_sa_resbot_m2 res_bot_ref_m2 ( .div_2r(dec_ref_2r),
     .div_3r(net0155), .bl_out(net0181), .nwell(nwell),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .bl_in(blsa_ref));
nch  M1 ( .D(net0173), .B(GND_), .G(testdec_b), .S(net0269));
nch  M27 ( .D(net0103), .B(GND_), .G(vdd_tieh), .S(blsa_ref));
vdd_tielow I204 ( .gnd_tiel(gnnd_tlow));
inv_25 I38 ( .IN(testdec_en_b_25), .OUT(dec_gate_25), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
inv_25 I222 ( .IN(dec_ok_25), .OUT(net0114), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I224 ( .IN(net0114), .OUT(net098), .P(vdd_), .Pb(vdd_),
     .G(gnd_), .Gb(gnd_));
nor2_hvt I214 ( .B(high_res_b), .Y(net0132), .A(testdec));
mux2_hvt I206 ( .in1(blsa), .in0(dec_in_3r), .out(in_div),
     .sel(testdec_b));
mux2_hvt I207 ( .in1(dec_ref_2r), .in0(dec_ref_2r), .out(in_ref),
     .sel(testdec_b));
mux2_hvt I219 ( .in1(net098), .in0(sa_out), .out(net0191),
     .sel(tm_testdec_wr));
rppolywo_m  R3 ( .MINUS(net0115), .PLUS(net0112), .BULK(gnd_));
rppolywo_m  R0 ( .MINUS(net0169), .PLUS(net0115), .BULK(gnd_));
ml_rock_gwlgnd_nor2 Iml_rock_gwlgnd_nor2 ( .gwl_b_gnden_25(vdd_tieh),
     .gwl_b_sup_25(vpxa), .gwl_b_25(saen_b_vpxa),
     .gwl_gnd_25(gwl_gnd_25_ref));
inv_hvt I208 ( .A(fsm_tm_testdec), .Y(testdec_b));
inv_hvt I220 ( .A(testdec_b), .Y(testdec));
inv_hvt I213 ( .A(net0132), .Y(net0120));
inv_hvt I215 ( .A(fsm_rst_b), .Y(net131));
inv_hvt I136 ( .A(rd_out_b), .Y(nv_dataout));
nor3_hvt I102 ( .B(dec_trim[6]), .Y(high_res_b), .A(dec_trim[5]),
     .C(dec_trim[7]));
vddp_tiehigh I169 ( .vddp_tieh(vddp_tieh));
vdd_tiehigh I117_2_ ( .vdd_tieh(nwell));
vdd_tiehigh I117_1_ ( .vdd_tieh(nwell));
vdd_tiehigh I117_0_ ( .vdd_tieh(nwell));
vdd_tiehigh I168 ( .vdd_tieh(vdd_tieh));
ml_core_sa_refres Irefres ( .nwell(wp_ref),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .wp_ref(wp_ref), .bot(net0173));
ml_core_sa_resbot res_bot_sen ( .div_2r(net0228), .div_3r(dec_in_3r),
     .bl_out(net0112), .nwell(nwell),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .bl_in(blsa));
ml_rock_lwldrv_wp Irock_lwldrv_wp ( .gwl_gnd_25(gwl_gnd_25_ref),
     .s_b_hv(vddp_tieh), .gwp_hv(vddp_tieh), .gwl_b_25(gnnd_tlow),
     .ngate_25(vpxa), .s_b_25(vpxa), .wp(wp_ref));
sbtlibn65lp_ml_dff_schematic I132 ( .R(net131), .D(net0191),
     .CLK(fsm_sample), .QN(rd_out_b), .Q(net135));
ml_core_sa_comp_top Icore_sa_comp_top ( .saen_25(saen_25),
     .in_ref(in_ref), .in_div(in_div), .sa_out(sa_out));
nch_hvt  M48 ( .D(net0169), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M46 ( .D(net0112), .B(GND_), .G(net0120), .S(gnd_));
nch_hvt  M45 ( .D(net0181), .B(GND_), .G(vdd_tieh), .S(gnd_));
nch_hvt  M47 ( .D(net0115), .B(GND_), .G(dec_trim[5]), .S(gnd_));
nch_hvt  M14 ( .D(net184), .B(GND_), .G(vdd_tieh), .S(net0103));
nch_hvt  M16 ( .D(net208), .B(GND_), .G(vdd_tieh), .S(net184));
nch_25  M21 ( .D(blsa_ref), .B(GND_), .G(saen_b_vpxa), .S(gnd_));
nch_25  M23 ( .D(vdd_), .B(gnd_), .G(dec_gate_25), .S(net0269));
nch_25  M25 ( .D(net0269), .B(GND_), .G(vddp_tieh), .S(net208));

endmodule
// Library - NVCM, Cell - ml_core_sa_top, View - schematic
// LAST TIME SAVED: Apr 18 11:05:06 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_sa_top ( nv_dataout, bl_out, bl_pgm_glb, vpxa,
     dec_ok_25, dec_trim, fsm_rst_b, fsm_sample, fsm_tm_testdec,
     sa_bl_to_blsa, sa_bl_to_pgm_glb, sa_ngate_25, sa_pgate_vpxa,
     saen_25, saen_b_vpxa, testdec_en_b_25, tm_dma, tm_testdec_wr );
output  nv_dataout;

inout  bl_out, bl_pgm_glb, vpxa;

input  dec_ok_25, fsm_rst_b, fsm_sample, fsm_tm_testdec, sa_bl_to_blsa,
     sa_bl_to_pgm_glb, saen_25, saen_b_vpxa, testdec_en_b_25, tm_dma,
     tm_testdec_wr;

input [7:5]  dec_trim;
input [4:1]  sa_ngate_25;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch  M27 ( .D(bl_out), .B(GND_), .G(net81), .S(net71));
inv_hvt I108 ( .A(net063), .Y(net061));
inv_hvt I131 ( .A(tm_dma), .Y(net063));
inv_hvt I101 ( .A(net69), .Y(net77));
inv_hvt I102 ( .A(sa_bl_to_pgm_glb), .Y(net69));
inv_hvt I167 ( .A(sa_bl_to_blsa), .Y(net73));
inv_hvt I96 ( .A(net73), .Y(net81));
pch_hvt  M1 ( .D(bl_pgm_glb), .B(VDD_), .G(net69), .S(bl_out));
pch_hvt  M11 ( .D(VDD_), .B(VDD_), .G(net73), .S(VDD_));
nch_hvt  M2 ( .D(bl_out), .B(GND_), .G(net77), .S(bl_pgm_glb));
nch_hvt  M4 ( .D(net71), .B(GND_), .G(net061), .S(gnd_));
ml_core_sa Iml_core_sa ( .tm_testdec_wr(tm_testdec_wr),
     .testdec_en_b_25(testdec_en_b_25),
     .fsm_tm_testdec(fsm_tm_testdec), .dec_ok_25(dec_ok_25),
     .saen_b_vpxa(saen_b_vpxa), .saen_25(saen_25),
     .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .dec_trim(dec_trim[7:5]),
     .nv_dataout(nv_dataout), .vpxa(vpxa), .blsa(net71));

endmodule
// Library - NVCM, Cell - ml_s_b_hv_sw, View - schematic
// LAST TIME SAVED: May 16 11:29:12 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_s_b_hv_sw ( sbout_hv, ssup_hv, sbout_gnd_25, sbout_high_25,
     vddp_tieh );
inout  sbout_hv, ssup_hv;

input  sbout_gnd_25, sbout_high_25, vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I114 ( .IN(sbout_high_25), .OUT(net62), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
nch_25  M23 ( .D(sbout_hv), .B(GND_), .G(vddp_tieh), .S(net34));
nch_25  M7 ( .D(net34), .B(GND_), .G(sbout_gnd_25), .S(gnd_));
pch_25  M5 ( .D(net46), .B(ssup_hv), .G(sbout_hv_b), .S(ssup_hv));
pch_25  M14 ( .D(sbout_hv), .B(net46), .G(sbout_gnd_25), .S(net46));
ml_hv_ls_inv Iml_hv_ls_inv_vppt ( .vddp_tieh(vddp_tieh),
     .sel_b_25(net62), .sel_25(sbout_high_25), .out_b_hv(sbout_hv_b),
     .in_hv(ssup_hv));

endmodule
// Library - NVCM, Cell - ml_wp_ctrl, View - schematic
// LAST TIME SAVED: Mar  9 16:06:25 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_wp_ctrl ( s_b_25, s_b_hv, sb25sup_25, sbhvsup_hv,
     sb25_gnd_25, sb25_high_25, sbhv_gnd_25, sbhv_high_25 );
inout  sb25sup_25, sbhvsup_hv;


inout [3:0]  s_b_25;
inout [3:0]  s_b_hv;

input [3:0]  sbhv_high_25;
input [3:0]  sb25_gnd_25;
input [3:0]  sbhv_gnd_25;
input [3:0]  sb25_high_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I21_7_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_6_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_5_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_4_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_3_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_2_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_1_ ( .vddp_tieh(vddp_tieh));
vddp_tiehigh I21_0_ ( .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_25_sw_3_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[3]),
     .sbout_hv(s_b_25[3]), .sbout_high_25(sb25_high_25[3]));
ml_s_b_hv_sw Iml_s_b_25_sw_2_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[2]),
     .sbout_hv(s_b_25[2]), .sbout_high_25(sb25_high_25[2]));
ml_s_b_hv_sw Iml_s_b_25_sw_1_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[1]),
     .sbout_hv(s_b_25[1]), .sbout_high_25(sb25_high_25[1]));
ml_s_b_hv_sw Iml_s_b_25_sw_0_ ( .vddp_tieh(vddp_tieh),
     .ssup_hv(sb25sup_25), .sbout_gnd_25(sb25_gnd_25[0]),
     .sbout_hv(s_b_25[0]), .sbout_high_25(sb25_high_25[0]));
ml_s_b_hv_sw Iml_s_b_hv_sw_3_ ( .sbout_high_25(sbhv_high_25[3]),
     .sbout_hv(s_b_hv[3]), .sbout_gnd_25(sbhv_gnd_25[3]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_2_ ( .sbout_high_25(sbhv_high_25[2]),
     .sbout_hv(s_b_hv[2]), .sbout_gnd_25(sbhv_gnd_25[2]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_1_ ( .sbout_high_25(sbhv_high_25[1]),
     .sbout_hv(s_b_hv[1]), .sbout_gnd_25(sbhv_gnd_25[1]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));
ml_s_b_hv_sw Iml_s_b_hv_sw_0_ ( .sbout_high_25(sbhv_high_25[0]),
     .sbout_hv(s_b_hv[0]), .sbout_gnd_25(sbhv_gnd_25[0]),
     .ssup_hv(sbhvsup_hv), .vddp_tieh(vddp_tieh));

endmodule
// Library - NVCM, Cell - ml_core_ctrl_top_8f, View - schematic
// LAST TIME SAVED: Sep 15 16:44:22 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_core_ctrl_top_8f ( gwl_b_gnden_25, nv_dataout, yp1, yp1_b_25,
     yp2, yp2_b_25, yp3_25, yp3_b_25, yp_test, yp_test_25,
     yp_test_b_25, bl_out, bl_pgm_glb, s_b_25, s_b_hv, sb25sup_25,
     sbhvsup_hv, vblinhi_pgm_25, vdd_tieh, vpxa, ysup_25, dec_ok_25_l,
     dec_ok_25_r, fsm_blkadd, fsm_coladd, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rowadd,
     fsm_rst_b, fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec,
     fsm_tm_trow, fsm_trim_rrefpgm, fsm_trim_rrefrd, fsm_vpxaset,
     fsm_wpen, fsm_ymuxdis, sa_ngate_25, sa_pgate_vpxa, saen_25,
     saen_b_vpxa, testdec_en_b_25, tm_allbank_sel, tm_allbl_h,
     tm_allbl_l, tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr
     );
output  gwl_b_gnden_25, nv_dataout;

inout  bl_out, bl_pgm_glb, sb25sup_25, sbhvsup_hv, vblinhi_pgm_25,
     vdd_tieh, vpxa, ysup_25;

input  dec_ok_25_l, dec_ok_25_r, fsm_gwlbdis_b_25, fsm_lshven,
     fsm_multibl_read, fsm_nv_rri_trim, fsm_nv_rrow, fsm_nv_sisi_ui,
     fsm_nvcmen, fsm_pgm, fsm_pgmien, fsm_pgmvfy, fsm_rd, fsm_rst_b,
     fsm_sample, fsm_tm_rd_mode, fsm_tm_testdec, fsm_tm_trow,
     fsm_vpxaset, fsm_wpen, fsm_ymuxdis, saen_25, saen_b_vpxa,
     testdec_en_b_25, tm_allbank_sel, tm_allbl_h, tm_allbl_l,
     tm_allwl_h, tm_allwl_l, tm_dma, tm_tcol, tm_testdec_wr;

output [7:0]  yp2_b_25;
output [7:0]  yp3_b_25;
output [7:0]  yp2;
output [10:0]  yp1_b_25;
output [1:0]  yp_test;
output [7:0]  yp3_25;
output [1:0]  yp_test_b_25;
output [1:0]  yp_test_25;
output [10:0]  yp1;

inout [3:0]  s_b_hv;
inout [3:0]  s_b_25;

input [9:0]  fsm_coladd;
input [4:1]  sa_ngate_25;
input [2:0]  fsm_trim_rrefpgm;
input [3:0]  fsm_blkadd;
input [1:0]  fsm_rowadd;
input [2:0]  fsm_trim_rrefrd;
input [4:1]  sa_pgate_vpxa;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  yp2_sel;

wire  [3:0]  sb25_gnd_25;

wire  [3:0]  sbhv_gnd_25;

wire  [3:0]  sbhv_high_25;

wire  [10:0]  yp1_sel;

wire  [3:0]  sb25_high_25;

wire  [7:5]  dec_trim;

wire  [7:0]  yp3_sel;



ml_mux2_25 I32 ( .sel_a_25(sel_dec_l_25), .in_b_25(dec_ok_25_r),
     .in_a_25(dec_ok_25_l), .out_25(data_ok_25));
ml_ymux_ctrl_8f Iml_ymux_ctrl_8f ( .yp1_b_25(yp1_b_25[10:0]),
     .yp1(yp1[10:0]), .yp1_sel(yp1_sel[10:0]), .yp2(yp2[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2_sel(yp2_sel[7:0]),
     .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .yp3_sel(yp3_sel[7:0]), .ysup_25(ysup_25),
     .yp_test_b_25(yp_test_b_25[1:0]), .yp_test_b_high_b(gnd_),
     .yp_test_b_low_b(gnd_), .yp_test(yp_test[1:0]),
     .yp2_b_low_b(yp21_b_low_b), .yp1_b_low_b(yp21_b_low_b),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .yp_test_25(yp_test_25[1:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25));
ml_core_ctrl_logic_8f Icore_ctrl_logic_8f (
     .tm_allbank_sel(tm_allbank_sel), .sel_dec_l_25(sel_dec_l_25),
     .yp1_sel(yp1_sel[10:0]), .fsm_coladd(fsm_coladd[9:0]),
     .yp2_sel(yp2_sel[7:0]), .fsm_tm_trow(fsm_tm_trow),
     .fsm_nv_sisi_ui(fsm_nv_sisi_ui),
     .fsm_nv_rri_trim(fsm_nv_rri_trim), .fsm_nv_rrow(fsm_nv_rrow),
     .fsm_rowadd(fsm_rowadd[1:0]), .fsm_tm_allwl_l(tm_allwl_l),
     .fsm_tm_allwl_h(tm_allwl_h), .ysup_25(ysup_25), .tm_tcol(tm_tcol),
     .fsm_ymuxdis(fsm_ymuxdis), .fsm_wpen(fsm_wpen),
     .fsm_vpxaset(fsm_vpxaset), .fsm_trim_rrefrd(fsm_trim_rrefrd[2:0]),
     .fsm_trim_rrefpgm(fsm_trim_rrefpgm[2:0]),
     .fsm_tm_testdec(fsm_tm_testdec), .fsm_tm_rd_mode(fsm_tm_rd_mode),
     .fsm_tm_allbl_l(tm_allbl_l), .fsm_pgm(fsm_pgm),
     .fsm_tm_allbl_h(tm_allbl_h), .fsm_rd(fsm_rd),
     .fsm_pgmvfy(fsm_pgmvfy), .fsm_pgmien(fsm_pgmien),
     .fsm_nvcmen(fsm_nvcmen), .fsm_multibl_read(fsm_multibl_read),
     .fsm_lshven(fsm_lshven), .fsm_blkadd(fsm_blkadd[3:0]),
     .yp_test(yp_test[1:0]), .yp21_b_low_b(yp21_b_low_b),
     .yp3_sel(yp3_sel[7:0]), .yp3_b_low_ysup_25(yp3_b_low_ysup_25),
     .yp3_b_high_odd_b_ysup_25(yp3_b_high_odd_b_ysup_25),
     .yp3_b_high_even_b_ysup_25(yp3_b_high_even_b_ysup_25),
     .sbhv_high_25(sbhv_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sb25_gnd_25(sb25_gnd_25[3:0]),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .en_blinhi_pgm_b_ysup_25(en_blinhi_pgm_b_25),
     .en_blinhi_pgm_b(en_blinhi_pgm_b), .dec_trim(dec_trim[7:5]));
inv_25 I38 ( .IN(net211), .OUT(gwl_b_gnden_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
inv_25 I30 ( .IN(fsm_gwlbdis_b_25), .OUT(net211), .P(vddp_),
     .Pb(vddp_), .G(gnd_), .Gb(gnd_));
vdd_tiehigh I117_9_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_8_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_7_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_6_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_5_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_4_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_3_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_2_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_1_ ( .vdd_tieh(vdd_tieh));
vdd_tiehigh I117_0_ ( .vdd_tieh(vdd_tieh));
ml_core_sa_top Icore_sa_top ( .tm_dma(tm_dma),
     .fsm_tm_testdec(fsm_tm_testdec), .tm_testdec_wr(tm_testdec_wr),
     .testdec_en_b_25(testdec_en_b_25), .dec_ok_25(data_ok_25),
     .sa_bl_to_blsa(sa_bl_to_blsa),
     .sa_bl_to_pgm_glb(sa_bl_to_pgm_glb), .saen_b_vpxa(saen_b_vpxa),
     .saen_25(saen_25), .sa_pgate_vpxa(sa_pgate_vpxa[4:1]),
     .sa_ngate_25(sa_ngate_25[4:1]), .fsm_sample(fsm_sample),
     .fsm_rst_b(fsm_rst_b), .dec_trim(dec_trim[7:5]),
     .nv_dataout(nv_dataout), .vpxa(vpxa), .bl_pgm_glb(bl_pgm_glb),
     .bl_out(bl_out));
ml_wp_ctrl Iml_wp_ctrl ( .sb25sup_25(sb25sup_25),
     .sbhvsup_hv(sbhvsup_hv), .sbhv_high_25(sbhv_high_25[3:0]),
     .sb25_high_25(sb25_high_25[3:0]), .sbhv_gnd_25(sbhv_gnd_25[3:0]),
     .sb25_gnd_25(sb25_gnd_25[3:0]), .s_b_25(s_b_25[3:0]),
     .s_b_hv(s_b_hv[3:0]));

endmodule
// Library - io, Cell - rgtbank_f, View - schematic
// LAST TIME SAVED: Jun  5 17:37:00 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module rgtbank_f ( Tdo, in, tck_int, tdi_int, tms_int, trstb_int, pad,
     TRSTb, Tck, Tdi, Tms, oen, out, ren, tdo_en, tdo_int );
output  Tdo, tck_int, tdi_int, tms_int, trstb_int;


input  TRSTb, Tck, Tdi, Tms, tdo_en, tdo_int;

output [54:0]  in;

inout [54:0]  pad;

input [54:0]  oen;
input [54:0]  out;
input [54:0]  ren;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



PDUW08DGZ I63_5_ ( .PAD(pad[5]), .C(in[5]), .OEN(oen[5]), .I(out[5]),
     .REN(ren[5]));
PDUW08DGZ I63_4_ ( .PAD(pad[4]), .C(in[4]), .OEN(oen[4]), .I(out[4]),
     .REN(ren[4]));
PDUW08DGZ I61_3_ ( .PAD(pad[3]), .C(in[3]), .OEN(oen[3]), .I(out[3]),
     .REN(ren[3]));
PDUW08DGZ I61_2_ ( .PAD(pad[2]), .C(in[2]), .OEN(oen[2]), .I(out[2]),
     .REN(ren[2]));
PDUW08DGZ I61_1_ ( .PAD(pad[1]), .C(in[1]), .OEN(oen[1]), .I(out[1]),
     .REN(ren[1]));
PDUW08DGZ I61_0_ ( .PAD(pad[0]), .C(in[0]), .OEN(oen[0]), .I(out[0]),
     .REN(ren[0]));
PDUW08DGZ I69_22_ ( .PAD(pad[22]), .C(in[22]), .OEN(oen[22]),
     .I(out[22]), .REN(ren[22]));
PDUW08DGZ I69_21_ ( .PAD(pad[21]), .C(in[21]), .OEN(oen[21]),
     .I(out[21]), .REN(ren[21]));
PDUW08DGZ I69_20_ ( .PAD(pad[20]), .C(in[20]), .OEN(oen[20]),
     .I(out[20]), .REN(ren[20]));
PDUW08DGZ I69_19_ ( .PAD(pad[19]), .C(in[19]), .OEN(oen[19]),
     .I(out[19]), .REN(ren[19]));
PDUW08DGZ I68_54_ ( .PAD(pad[54]), .C(in[54]), .OEN(oen[54]),
     .I(out[54]), .REN(ren[54]));
PDUW08DGZ I68_53_ ( .PAD(pad[53]), .C(in[53]), .OEN(oen[53]),
     .I(out[53]), .REN(ren[53]));
PDUW08DGZ I68_52_ ( .PAD(pad[52]), .C(in[52]), .OEN(oen[52]),
     .I(out[52]), .REN(ren[52]));
PDUW08DGZ I68_51_ ( .PAD(pad[51]), .C(in[51]), .OEN(oen[51]),
     .I(out[51]), .REN(ren[51]));
PDUW08DGZ I67_18_ ( .PAD(pad[18]), .C(in[18]), .OEN(oen[18]),
     .I(out[18]), .REN(ren[18]));
PDUW08DGZ I67_17_ ( .PAD(pad[17]), .C(in[17]), .OEN(oen[17]),
     .I(out[17]), .REN(ren[17]));
PDUW08DGZ I67_16_ ( .PAD(pad[16]), .C(in[16]), .OEN(oen[16]),
     .I(out[16]), .REN(ren[16]));
PDUW08DGZ I67_15_ ( .PAD(pad[15]), .C(in[15]), .OEN(oen[15]),
     .I(out[15]), .REN(ren[15]));
PDUW08DGZ I67_14_ ( .PAD(pad[14]), .C(in[14]), .OEN(oen[14]),
     .I(out[14]), .REN(ren[14]));
PDUW08DGZ I67_13_ ( .PAD(pad[13]), .C(in[13]), .OEN(oen[13]),
     .I(out[13]), .REN(ren[13]));
PDUW08DGZ I67_12_ ( .PAD(pad[12]), .C(in[12]), .OEN(oen[12]),
     .I(out[12]), .REN(ren[12]));
PDUW08DGZ I67_11_ ( .PAD(pad[11]), .C(in[11]), .OEN(oen[11]),
     .I(out[11]), .REN(ren[11]));
PDUW08DGZ I66_50_ ( .PAD(pad[50]), .C(in[50]), .OEN(oen[50]),
     .I(out[50]), .REN(ren[50]));
PDUW08DGZ I66_49_ ( .PAD(pad[49]), .C(in[49]), .OEN(oen[49]),
     .I(out[49]), .REN(ren[49]));
PDUW08DGZ I65_10_ ( .PAD(pad[10]), .C(in[10]), .OEN(oen[10]),
     .I(out[10]), .REN(ren[10]));
PDUW08DGZ I65_9_ ( .PAD(pad[9]), .C(in[9]), .OEN(oen[9]), .I(out[9]),
     .REN(ren[9]));
PDUW08DGZ I65_8_ ( .PAD(pad[8]), .C(in[8]), .OEN(oen[8]), .I(out[8]),
     .REN(ren[8]));
PDUW08DGZ I65_7_ ( .PAD(pad[7]), .C(in[7]), .OEN(oen[7]), .I(out[7]),
     .REN(ren[7]));
PDUW08DGZ I65_6_ ( .PAD(pad[6]), .C(in[6]), .OEN(oen[6]), .I(out[6]),
     .REN(ren[6]));
PDUW08DGZ I64_48_ ( .PAD(pad[48]), .C(in[48]), .OEN(oen[48]),
     .I(out[48]), .REN(ren[48]));
PDUW08DGZ I64_47_ ( .PAD(pad[47]), .C(in[47]), .OEN(oen[47]),
     .I(out[47]), .REN(ren[47]));
PDUW08DGZ I62_46_ ( .PAD(pad[46]), .C(in[46]), .OEN(oen[46]),
     .I(out[46]), .REN(ren[46]));
PDUW08DGZ I62_45_ ( .PAD(pad[45]), .C(in[45]), .OEN(oen[45]),
     .I(out[45]), .REN(ren[45]));
PDUW08DGZ I62_44_ ( .PAD(pad[44]), .C(in[44]), .OEN(oen[44]),
     .I(out[44]), .REN(ren[44]));
PDUW08DGZ I62_43_ ( .PAD(pad[43]), .C(in[43]), .OEN(oen[43]),
     .I(out[43]), .REN(ren[43]));
PDUW08DGZ I62_42_ ( .PAD(pad[42]), .C(in[42]), .OEN(oen[42]),
     .I(out[42]), .REN(ren[42]));
PDUW08DGZ I62_41_ ( .PAD(pad[41]), .C(in[41]), .OEN(oen[41]),
     .I(out[41]), .REN(ren[41]));
PDUW08DGZ I62_40_ ( .PAD(pad[40]), .C(in[40]), .OEN(oen[40]),
     .I(out[40]), .REN(ren[40]));
PDUW08DGZ I62_39_ ( .PAD(pad[39]), .C(in[39]), .OEN(oen[39]),
     .I(out[39]), .REN(ren[39]));
PDUW08DGZ I62_38_ ( .PAD(pad[38]), .C(in[38]), .OEN(oen[38]),
     .I(out[38]), .REN(ren[38]));
PDUW08DGZ I62_37_ ( .PAD(pad[37]), .C(in[37]), .OEN(oen[37]),
     .I(out[37]), .REN(ren[37]));
PDUW08DGZ I60_36_ ( .PAD(pad[36]), .C(in[36]), .OEN(oen[36]),
     .I(out[36]), .REN(ren[36]));
PDUW08DGZ I58_35_ ( .PAD(pad[35]), .C(in[35]), .OEN(oen[35]),
     .I(out[35]), .REN(ren[35]));
PDUW08DGZ I58_34_ ( .PAD(pad[34]), .C(in[34]), .OEN(oen[34]),
     .I(out[34]), .REN(ren[34]));
PDUW08DGZ I58_33_ ( .PAD(pad[33]), .C(in[33]), .OEN(oen[33]),
     .I(out[33]), .REN(ren[33]));
PDUW08DGZ I58_32_ ( .PAD(pad[32]), .C(in[32]), .OEN(oen[32]),
     .I(out[32]), .REN(ren[32]));
PDUW08DGZ I58_31_ ( .PAD(pad[31]), .C(in[31]), .OEN(oen[31]),
     .I(out[31]), .REN(ren[31]));
PDUW08DGZ I58_30_ ( .PAD(pad[30]), .C(in[30]), .OEN(oen[30]),
     .I(out[30]), .REN(ren[30]));
PDUW08DGZ I58_29_ ( .PAD(pad[29]), .C(in[29]), .OEN(oen[29]),
     .I(out[29]), .REN(ren[29]));
PDUW08DGZ I58_28_ ( .PAD(pad[28]), .C(in[28]), .OEN(oen[28]),
     .I(out[28]), .REN(ren[28]));
PDUW08DGZ I58_27_ ( .PAD(pad[27]), .C(in[27]), .OEN(oen[27]),
     .I(out[27]), .REN(ren[27]));
PDUW08DGZ I58_26_ ( .PAD(pad[26]), .C(in[26]), .OEN(oen[26]),
     .I(out[26]), .REN(ren[26]));
PDUW08DGZ I58_25_ ( .PAD(pad[25]), .C(in[25]), .OEN(oen[25]),
     .I(out[25]), .REN(ren[25]));
PDUW08DGZ I58_24_ ( .PAD(pad[24]), .C(in[24]), .OEN(oen[24]),
     .I(out[24]), .REN(ren[24]));
PDUW08DGZ I58_23_ ( .PAD(pad[23]), .C(in[23]), .OEN(oen[23]),
     .I(out[23]), .REN(ren[23]));
PDT08DGZ I42 ( .OEN(tdo_en), .I(tdo_int), .PAD(Tdo));
PDIDGZ I55 ( .PAD(Tdi), .C(tdi_int));
PDIDGZ I40 ( .C(tck_int), .PAD(Tck));
PDIDGZ I41 ( .C(trstb_int), .PAD(TRSTb));
PDIDGZ I39 ( .C(tms_int), .PAD(Tms));
PVSS3DGZ I70_1_ ( .VSS(gnd_));
PVSS3DGZ I70_0_ ( .VSS(gnd_));
PVSS3DGZ I73_1_ ( .VSS(gnd_));
PVSS3DGZ I73_0_ ( .VSS(gnd_));
PVSS3DGZ I75_1_ ( .VSS(gnd_));
PVSS3DGZ I75_0_ ( .VSS(gnd_));
PVSS3DGZ I80_1_ ( .VSS(gnd_));
PVSS3DGZ I80_0_ ( .VSS(gnd_));
PVDD1DGZ I72_1_ ( .VDD(vdd_));
PVDD1DGZ I72_0_ ( .VDD(vdd_));
PVDD1DGZ I77_1_ ( .VDD(vdd_));
PVDD1DGZ I77_0_ ( .VDD(vdd_));
PVDD2POC I82 ( .VDDPST(vddp_));
PVDD2POC I79 ( .VDDPST(vddio_rightbank));
PVDD2DGZ I71_1_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I71_0_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I78 ( .VDDPST(vddio_rightbank));
PVDD2DGZ I74_1_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I74_0_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I76_1_ ( .VDDPST(vddio_rightbank));
PVDD2DGZ I76_0_ ( .VDDPST(vddio_rightbank));

endmodule
// Library - NVCM, Cell - ml_testdec_columns, View - schematic
// LAST TIME SAVED: Feb 26 14:35:47 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_testdec_columns ( bl, dec_det_even_25, dec_det_odd_25 );

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M5 ( .D(vdd_), .B(gnd_), .G(dec_det_even_25), .S(bl[0]));
nch_25  M4 ( .D(vdd_), .B(gnd_), .G(dec_det_odd_25), .S(bl[1]));

endmodule
// Library - NVCM, Cell - ml_testdec_columnsx320, View - schematic
// LAST TIME SAVED: Jun 12 13:56:54 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_testdec_columnsx320 ( bl, bl_dummyl, bl_dummyr,
     dec_det_even_25, dec_det_odd_25 );

input  dec_det_even_25, dec_det_odd_25;

inout [1:0]  bl_dummyl;
inout [1:0]  bl_dummyr;
inout [319:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



ml_testdec_columns Itestdec_columns_dml (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyl[1:0]));
ml_testdec_columns Itestdec_columns_159_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[319:318]));
ml_testdec_columns Itestdec_columns_158_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[317:316]));
ml_testdec_columns Itestdec_columns_157_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[315:314]));
ml_testdec_columns Itestdec_columns_156_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[313:312]));
ml_testdec_columns Itestdec_columns_155_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[311:310]));
ml_testdec_columns Itestdec_columns_154_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[309:308]));
ml_testdec_columns Itestdec_columns_153_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[307:306]));
ml_testdec_columns Itestdec_columns_152_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[305:304]));
ml_testdec_columns Itestdec_columns_151_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[303:302]));
ml_testdec_columns Itestdec_columns_150_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[301:300]));
ml_testdec_columns Itestdec_columns_149_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[299:298]));
ml_testdec_columns Itestdec_columns_148_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[297:296]));
ml_testdec_columns Itestdec_columns_147_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[295:294]));
ml_testdec_columns Itestdec_columns_146_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[293:292]));
ml_testdec_columns Itestdec_columns_145_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[291:290]));
ml_testdec_columns Itestdec_columns_144_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[289:288]));
ml_testdec_columns Itestdec_columns_143_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[287:286]));
ml_testdec_columns Itestdec_columns_142_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[285:284]));
ml_testdec_columns Itestdec_columns_141_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[283:282]));
ml_testdec_columns Itestdec_columns_140_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[281:280]));
ml_testdec_columns Itestdec_columns_139_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[279:278]));
ml_testdec_columns Itestdec_columns_138_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[277:276]));
ml_testdec_columns Itestdec_columns_137_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[275:274]));
ml_testdec_columns Itestdec_columns_136_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[273:272]));
ml_testdec_columns Itestdec_columns_135_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[271:270]));
ml_testdec_columns Itestdec_columns_134_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[269:268]));
ml_testdec_columns Itestdec_columns_133_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[267:266]));
ml_testdec_columns Itestdec_columns_132_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[265:264]));
ml_testdec_columns Itestdec_columns_131_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[263:262]));
ml_testdec_columns Itestdec_columns_130_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[261:260]));
ml_testdec_columns Itestdec_columns_129_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[259:258]));
ml_testdec_columns Itestdec_columns_128_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[257:256]));
ml_testdec_columns Itestdec_columns_127_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[255:254]));
ml_testdec_columns Itestdec_columns_126_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[253:252]));
ml_testdec_columns Itestdec_columns_125_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[251:250]));
ml_testdec_columns Itestdec_columns_124_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[249:248]));
ml_testdec_columns Itestdec_columns_123_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[247:246]));
ml_testdec_columns Itestdec_columns_122_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[245:244]));
ml_testdec_columns Itestdec_columns_121_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[243:242]));
ml_testdec_columns Itestdec_columns_120_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[241:240]));
ml_testdec_columns Itestdec_columns_119_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[239:238]));
ml_testdec_columns Itestdec_columns_118_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[237:236]));
ml_testdec_columns Itestdec_columns_117_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[235:234]));
ml_testdec_columns Itestdec_columns_116_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[233:232]));
ml_testdec_columns Itestdec_columns_115_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[231:230]));
ml_testdec_columns Itestdec_columns_114_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[229:228]));
ml_testdec_columns Itestdec_columns_113_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[227:226]));
ml_testdec_columns Itestdec_columns_112_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[225:224]));
ml_testdec_columns Itestdec_columns_111_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[223:222]));
ml_testdec_columns Itestdec_columns_110_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[221:220]));
ml_testdec_columns Itestdec_columns_109_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[219:218]));
ml_testdec_columns Itestdec_columns_108_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[217:216]));
ml_testdec_columns Itestdec_columns_107_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[215:214]));
ml_testdec_columns Itestdec_columns_106_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[213:212]));
ml_testdec_columns Itestdec_columns_105_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[211:210]));
ml_testdec_columns Itestdec_columns_104_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[209:208]));
ml_testdec_columns Itestdec_columns_103_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[207:206]));
ml_testdec_columns Itestdec_columns_102_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[205:204]));
ml_testdec_columns Itestdec_columns_101_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[203:202]));
ml_testdec_columns Itestdec_columns_100_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[201:200]));
ml_testdec_columns Itestdec_columns_99_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[199:198]));
ml_testdec_columns Itestdec_columns_98_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[197:196]));
ml_testdec_columns Itestdec_columns_97_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[195:194]));
ml_testdec_columns Itestdec_columns_96_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[193:192]));
ml_testdec_columns Itestdec_columns_95_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[191:190]));
ml_testdec_columns Itestdec_columns_94_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[189:188]));
ml_testdec_columns Itestdec_columns_93_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[187:186]));
ml_testdec_columns Itestdec_columns_92_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[185:184]));
ml_testdec_columns Itestdec_columns_91_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[183:182]));
ml_testdec_columns Itestdec_columns_90_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[181:180]));
ml_testdec_columns Itestdec_columns_89_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[179:178]));
ml_testdec_columns Itestdec_columns_88_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[177:176]));
ml_testdec_columns Itestdec_columns_87_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[175:174]));
ml_testdec_columns Itestdec_columns_86_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[173:172]));
ml_testdec_columns Itestdec_columns_85_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[171:170]));
ml_testdec_columns Itestdec_columns_84_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[169:168]));
ml_testdec_columns Itestdec_columns_83_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[167:166]));
ml_testdec_columns Itestdec_columns_82_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[165:164]));
ml_testdec_columns Itestdec_columns_81_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[163:162]));
ml_testdec_columns Itestdec_columns_80_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[161:160]));
ml_testdec_columns Itestdec_columns_79_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[159:158]));
ml_testdec_columns Itestdec_columns_78_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[157:156]));
ml_testdec_columns Itestdec_columns_77_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[155:154]));
ml_testdec_columns Itestdec_columns_76_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[153:152]));
ml_testdec_columns Itestdec_columns_75_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[151:150]));
ml_testdec_columns Itestdec_columns_74_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[149:148]));
ml_testdec_columns Itestdec_columns_73_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[147:146]));
ml_testdec_columns Itestdec_columns_72_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[145:144]));
ml_testdec_columns Itestdec_columns_71_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[143:142]));
ml_testdec_columns Itestdec_columns_70_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[141:140]));
ml_testdec_columns Itestdec_columns_69_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[139:138]));
ml_testdec_columns Itestdec_columns_68_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[137:136]));
ml_testdec_columns Itestdec_columns_67_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[135:134]));
ml_testdec_columns Itestdec_columns_66_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[133:132]));
ml_testdec_columns Itestdec_columns_65_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[131:130]));
ml_testdec_columns Itestdec_columns_64_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[129:128]));
ml_testdec_columns Itestdec_columns_63_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[127:126]));
ml_testdec_columns Itestdec_columns_62_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[125:124]));
ml_testdec_columns Itestdec_columns_61_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[123:122]));
ml_testdec_columns Itestdec_columns_60_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[121:120]));
ml_testdec_columns Itestdec_columns_59_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[119:118]));
ml_testdec_columns Itestdec_columns_58_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[117:116]));
ml_testdec_columns Itestdec_columns_57_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[115:114]));
ml_testdec_columns Itestdec_columns_56_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[113:112]));
ml_testdec_columns Itestdec_columns_55_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[111:110]));
ml_testdec_columns Itestdec_columns_54_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[109:108]));
ml_testdec_columns Itestdec_columns_53_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[107:106]));
ml_testdec_columns Itestdec_columns_52_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[105:104]));
ml_testdec_columns Itestdec_columns_51_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[103:102]));
ml_testdec_columns Itestdec_columns_50_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[101:100]));
ml_testdec_columns Itestdec_columns_49_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[99:98]));
ml_testdec_columns Itestdec_columns_48_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[97:96]));
ml_testdec_columns Itestdec_columns_47_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[95:94]));
ml_testdec_columns Itestdec_columns_46_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[93:92]));
ml_testdec_columns Itestdec_columns_45_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[91:90]));
ml_testdec_columns Itestdec_columns_44_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[89:88]));
ml_testdec_columns Itestdec_columns_43_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[87:86]));
ml_testdec_columns Itestdec_columns_42_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[85:84]));
ml_testdec_columns Itestdec_columns_41_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[83:82]));
ml_testdec_columns Itestdec_columns_40_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[81:80]));
ml_testdec_columns Itestdec_columns_39_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[79:78]));
ml_testdec_columns Itestdec_columns_38_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[77:76]));
ml_testdec_columns Itestdec_columns_37_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[75:74]));
ml_testdec_columns Itestdec_columns_36_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[73:72]));
ml_testdec_columns Itestdec_columns_35_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[71:70]));
ml_testdec_columns Itestdec_columns_34_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[69:68]));
ml_testdec_columns Itestdec_columns_33_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[67:66]));
ml_testdec_columns Itestdec_columns_32_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[65:64]));
ml_testdec_columns Itestdec_columns_31_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[63:62]));
ml_testdec_columns Itestdec_columns_30_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[61:60]));
ml_testdec_columns Itestdec_columns_29_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[59:58]));
ml_testdec_columns Itestdec_columns_28_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[57:56]));
ml_testdec_columns Itestdec_columns_27_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[55:54]));
ml_testdec_columns Itestdec_columns_26_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[53:52]));
ml_testdec_columns Itestdec_columns_25_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[51:50]));
ml_testdec_columns Itestdec_columns_24_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[49:48]));
ml_testdec_columns Itestdec_columns_23_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[47:46]));
ml_testdec_columns Itestdec_columns_22_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[45:44]));
ml_testdec_columns Itestdec_columns_21_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[43:42]));
ml_testdec_columns Itestdec_columns_20_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[41:40]));
ml_testdec_columns Itestdec_columns_19_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[39:38]));
ml_testdec_columns Itestdec_columns_18_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[37:36]));
ml_testdec_columns Itestdec_columns_17_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[35:34]));
ml_testdec_columns Itestdec_columns_16_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[33:32]));
ml_testdec_columns Itestdec_columns_15_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[31:30]));
ml_testdec_columns Itestdec_columns_14_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[29:28]));
ml_testdec_columns Itestdec_columns_13_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[27:26]));
ml_testdec_columns Itestdec_columns_12_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[25:24]));
ml_testdec_columns Itestdec_columns_11_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[23:22]));
ml_testdec_columns Itestdec_columns_10_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[21:20]));
ml_testdec_columns Itestdec_columns_9_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[19:18]));
ml_testdec_columns Itestdec_columns_8_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[17:16]));
ml_testdec_columns Itestdec_columns_7_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[15:14]));
ml_testdec_columns Itestdec_columns_6_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[13:12]));
ml_testdec_columns Itestdec_columns_5_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[11:10]));
ml_testdec_columns Itestdec_columns_4_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[9:8]));
ml_testdec_columns Itestdec_columns_3_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[7:6]));
ml_testdec_columns Itestdec_columns_2_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[5:4]));
ml_testdec_columns Itestdec_columns_1_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[3:2]));
ml_testdec_columns Itestdec_columns_0_ (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl[1:0]));
ml_testdec_columns Itestdec_columns_dmr (
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25), .bl(bl_dummyr[1:0]));

endmodule
// Library - ROCK, Cell - nvcm_cell_1, View - schematic
// LAST TIME SAVED: May 13 16:00:35 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_1 ( bl, wp, wr );
inout  bl;

input  wp, wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nchx  NR ( .D(net1), .G(wr), .S(bl));
nchx  NP ( .D(net5), .G(wp), .S(net1));

endmodule
// Library - NVCM, Cell - nvcm_cell_2x1, View - schematic
// LAST TIME SAVED: Dec 10 15:56:30 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_2x1 ( bl, wp, wr );

input  wp, wr;

inout [1:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
nvcm_cell_1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));

endmodule
// Library - NVCM, Cell - nvcm_cell_2x8, View - schematic
// LAST TIME SAVED: Feb 26 14:36:29 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_2x8 ( bl, wp, wr );


inout [1:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x1 m7 ( .bl(bl[1:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_2x1 m6 ( .bl(bl[1:0]), .wr(wr[6]), .wp(wp[6]));
nvcm_cell_2x1 m5 ( .bl(bl[1:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_2x1 m4 ( .bl(bl[1:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_2x1 m3 ( .bl(bl[1:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_2x1 m2 ( .bl(bl[1:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_2x1 m1 ( .bl(bl[1:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_2x1 m0 ( .bl(bl[1:0]), .wr(wr[0]), .wp(wp[0]));

endmodule
// Library - NVCM, Cell - nvcm_cell_1x8, View - schematic
// LAST TIME SAVED: Jul  5 11:06:02 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_1x8 ( bl, wp, wr );

input  wp, wr;

inout [7:0]  bl;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1 m0 ( .wp(wp), .wr(wr), .bl(bl[0]));
nvcm_cell_1 m1 ( .wp(wp), .wr(wr), .bl(bl[1]));
nvcm_cell_1 m2 ( .wp(wp), .wr(wr), .bl(bl[2]));
nvcm_cell_1 m3 ( .wp(wp), .wr(wr), .bl(bl[3]));
nvcm_cell_1 m4 ( .wp(wp), .wr(wr), .bl(bl[4]));
nvcm_cell_1 m5 ( .wp(wp), .wr(wr), .bl(bl[5]));
nvcm_cell_1 m6 ( .wp(wp), .wr(wr), .bl(bl[6]));
nvcm_cell_1 m7 ( .wp(wp), .wr(wr), .bl(bl[7]));

endmodule
// Library - NVCM, Cell - nvcm_cell_8x8, View - schematic
// LAST TIME SAVED: Dec 10 15:35:50 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_8x8 ( bl, wp, wr );


inout [7:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_1x8 m0 ( .bl(bl[7:0]), .wr(wr[0]), .wp(wp[0]));
nvcm_cell_1x8 m1 ( .bl(bl[7:0]), .wr(wr[1]), .wp(wp[1]));
nvcm_cell_1x8 m2 ( .bl(bl[7:0]), .wr(wr[2]), .wp(wp[2]));
nvcm_cell_1x8 m3 ( .bl(bl[7:0]), .wr(wr[3]), .wp(wp[3]));
nvcm_cell_1x8 m7 ( .bl(bl[7:0]), .wr(wr[7]), .wp(wp[7]));
nvcm_cell_1x8 m4 ( .bl(bl[7:0]), .wr(wr[4]), .wp(wp[4]));
nvcm_cell_1x8 m5 ( .bl(bl[7:0]), .wr(wr[5]), .wp(wp[5]));
nvcm_cell_1x8 m6 ( .bl(bl[7:0]), .wr(wr[6]), .wp(wp[6]));

endmodule
// Library - NVCM, Cell - nvcm_cell_16x8, View - schematic
// LAST TIME SAVED: Dec 10 15:41:25 2007
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_16x8 ( bl, wp, wr );


inout [15:0]  bl;

input [7:0]  wr;
input [7:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_8x8 m0 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[7:0]));
nvcm_cell_8x8 m1 ( .wr(wr[7:0]), .wp(wp[7:0]), .bl(bl[15:8]));

endmodule
// Library - NVCM, Cell - nvcm_cell_320x8, View - schematic
// LAST TIME SAVED: Jun 12 13:50:20 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_320x8 ( bl, bl_dummyl, bl_dummyr, wp, wr );


inout [1:0]  bl_dummyl;
inout [319:0]  bl;
inout [1:0]  bl_dummyr;

input [7:0]  wp;
input [7:0]  wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x8 Invcm_cell_2x8_r ( .bl(bl_dummyr[1:0]), .wr(wr[7:0]),
     .wp(wp[7:0]));
nvcm_cell_2x8 Invcm_cell_2x8_l ( .wp(wp[7:0]), .wr(wr[7:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_16x8 Invcm_cell_16x8_19_ ( .wp(wp[7:0]), .bl(bl[319:304]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_18_ ( .wp(wp[7:0]), .bl(bl[303:288]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_17_ ( .wp(wp[7:0]), .bl(bl[287:272]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_16_ ( .wp(wp[7:0]), .bl(bl[271:256]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_15_ ( .wp(wp[7:0]), .bl(bl[255:240]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_14_ ( .wp(wp[7:0]), .bl(bl[239:224]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_13_ ( .wp(wp[7:0]), .bl(bl[223:208]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_12_ ( .wp(wp[7:0]), .bl(bl[207:192]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_11_ ( .wp(wp[7:0]), .bl(bl[191:176]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_10_ ( .wp(wp[7:0]), .bl(bl[175:160]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_9_ ( .wp(wp[7:0]), .bl(bl[159:144]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_8_ ( .wp(wp[7:0]), .bl(bl[143:128]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_7_ ( .wp(wp[7:0]), .bl(bl[127:112]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_6_ ( .wp(wp[7:0]), .bl(bl[111:96]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_5_ ( .wp(wp[7:0]), .bl(bl[95:80]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_4_ ( .wp(wp[7:0]), .bl(bl[79:64]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_3_ ( .wp(wp[7:0]), .bl(bl[63:48]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_2_ ( .wp(wp[7:0]), .bl(bl[47:32]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_1_ ( .wp(wp[7:0]), .bl(bl[31:16]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_0_ ( .wp(wp[7:0]), .bl(bl[15:0]),
     .wr(wr[7:0]));

endmodule
// Library - NVCM, Cell - nvcm_cell_320x232, View - schematic
// LAST TIME SAVED: Jun 12 13:51:46 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module nvcm_cell_320x232 ( bl, bl_dummyl, bl_dummyr, wp, wp_dummyb,
     wp_dummyt, wr, wr_dummyb, wr_dummyt );


inout [1:0]  bl_dummyr;
inout [319:0]  bl;
inout [1:0]  bl_dummyl;

input [1:0]  wp_dummyb;
input [1:0]  wr_dummyb;
input [1:0]  wp_dummyt;
input [227:0]  wp;
input [1:0]  wr_dummyt;
input [227:0]  wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_320x8 Invcm_cell_320x8_26_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[221:214]), .wp(wp[221:214]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_25_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[213:206]), .wp(wp[213:206]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_24_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[205:198]), .wp(wp[205:198]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_23_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[197:190]), .wp(wp[197:190]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_22_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[189:182]), .wp(wp[189:182]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_21_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[181:174]), .wp(wp[181:174]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_20_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[173:166]), .wp(wp[173:166]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_19_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[165:158]), .wp(wp[165:158]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_18_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[157:150]), .wp(wp[157:150]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_17_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[149:142]), .wp(wp[149:142]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_16_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[141:134]), .wp(wp[141:134]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_15_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[133:126]), .wp(wp[133:126]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_14_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[125:118]), .wp(wp[125:118]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_13_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[117:110]), .wp(wp[117:110]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_12_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[109:102]), .wp(wp[109:102]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_11_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[101:94]), .wp(wp[101:94]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_10_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[93:86]), .wp(wp[93:86]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_9_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[85:78]), .wp(wp[85:78]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_8_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[77:70]), .wp(wp[77:70]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_7_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[69:62]), .wp(wp[69:62]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_6_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[61:54]), .wp(wp[61:54]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_5_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[53:46]), .wp(wp[53:46]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_4_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[45:38]), .wp(wp[45:38]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_3_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[37:30]), .wp(wp[37:30]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_2_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[29:22]), .wp(wp[29:22]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_1_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[21:14]), .wp(wp[21:14]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_0_ ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr(wr[13:6]), .wp(wp[13:6]),
     .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_t ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr({wr[5:0], wr_dummyt[1:0]}), .wp({wp[5:0],
     wp_dummyt[1:0]}), .bl_dummyl(bl_dummyl[1:0]));
nvcm_cell_320x8 Invcm_cell_320x8_b ( .bl_dummyr(bl_dummyr[1:0]),
     .bl(bl[319:0]), .wr({wr_dummyb[1:0], wr[227:222]}),
     .wp({wp_dummyb[1:0], wp[227:222]}), .bl_dummyl(bl_dummyl[1:0]));

endmodule
// Library - sbtlibn65lp, Cell - vddp_tiehigh, View - schematic
// LAST TIME SAVED: May  8 16:23:22 2008
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module vddp_tiehigh ( vddp_tieh );
inout  vddp_tieh;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M8 ( .D(net9), .B(GND_), .G(net9), .S(gnd_));
pch_25  M9 ( .D(vddp_tieh), .B(vddp_), .G(net9), .S(vddp_));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_dummy, View - schematic
// LAST TIME SAVED: Feb 26 14:34:35 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_dummy ( bl_dummyr, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, pgminhi_dmmy_b_25, vdd_tieh );
inout  vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo;

input  pgminhi_dmmy_b_25, vdd_tieh;

inout [1:0]  bl_dummyr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M1 ( .D(bl_dummyr[1]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rdo));
nch_25  M18 ( .D(bl_dummyr[0]), .B(GND_), .G(pgminhi_dmmy_b_25),
     .S(vblinhi_rde));
pch_25  M8 ( .D(bl_dummyr[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M0 ( .D(bl_dummyr[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_yp2_8, View - schematic
// LAST TIME SAVED: Jan 16 10:38:35 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_yp2_8 ( bl, bl_out, vblinhi_rde, vblinhi_rdo, yp2,
     yp2_b_25 );
inout  bl_out, vblinhi_rde, vblinhi_rdo;


inout [7:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M17 ( .D(bl[7]), .B(GND_), .G(yp2_b_25[7]), .S(vblinhi_rdo));
nch_25  M16 ( .D(bl[6]), .B(GND_), .G(yp2_b_25[6]), .S(vblinhi_rde));
nch_25  M11 ( .D(bl[1]), .B(GND_), .G(yp2_b_25[1]), .S(vblinhi_rdo));
nch_25  M20 ( .D(bl[0]), .B(GND_), .G(yp2_b_25[0]), .S(vblinhi_rde));
nch_25  M15 ( .D(bl[5]), .B(GND_), .G(yp2_b_25[5]), .S(vblinhi_rdo));
nch_25  M14 ( .D(bl[4]), .B(GND_), .G(yp2_b_25[4]), .S(vblinhi_rde));
nch_25  M13 ( .D(bl[3]), .B(GND_), .G(yp2_b_25[3]), .S(vblinhi_rdo));
nch_25  M12 ( .D(bl[2]), .B(GND_), .G(yp2_b_25[2]), .S(vblinhi_rde));
nch_hvt  M3 ( .D(bl[3]), .B(GND_), .G(yp2[3]), .S(bl_out));
nch_hvt  M1 ( .D(bl[2]), .B(GND_), .G(yp2[2]), .S(bl_out));
nch_hvt  M0 ( .D(bl[1]), .B(GND_), .G(yp2[1]), .S(bl_out));
nch_hvt  M7 ( .D(bl[7]), .B(GND_), .G(yp2[7]), .S(bl_out));
nch_hvt  M6 ( .D(bl[6]), .B(GND_), .G(yp2[6]), .S(bl_out));
nch_hvt  M5 ( .D(bl[5]), .B(GND_), .G(yp2[5]), .S(bl_out));
nch_hvt  M2 ( .D(bl[0]), .B(GND_), .G(yp2[0]), .S(bl_out));
nch_hvt  M4 ( .D(bl[4]), .B(GND_), .G(yp2[4]), .S(bl_out));

endmodule
// Library - NVCM, Cell - ml_ymux_yp3_x8, View - schematic
// LAST TIME SAVED: Feb 26 14:33:55 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_yp3_x8 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [7:0]  bl;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



pch_25  M5_7_ ( .D(bl[7]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_6_ ( .D(bl[6]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_5_ ( .D(bl[5]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_4_ ( .D(bl[4]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_3_ ( .D(bl[3]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_2_ ( .D(bl[2]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_1_ ( .D(bl[1]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
pch_25  M5_0_ ( .D(bl[0]), .B(vblinhi_pgm_25), .G(vdd_tieh),
     .S(vblinhi_pgm_25));
nch_25  M22 ( .D(bl[6]), .B(GND_), .G(yp3_25[6]), .S(bl_out));
nch_25  M1 ( .D(bl[4]), .B(GND_), .G(yp3_25[4]), .S(bl_out));
nch_25  M24 ( .D(bl[2]), .B(GND_), .G(yp3_25[2]), .S(bl_out));
nch_25  M25 ( .D(bl[0]), .B(GND_), .G(yp3_25[0]), .S(bl_out));
nch_25  M26 ( .D(bl[0]), .B(GND_), .G(yp3_b_25[0]), .S(vblinhi_rde));
nch_25  M27 ( .D(bl[1]), .B(GND_), .G(yp3_b_25[1]), .S(vblinhi_rdo));
nch_25  M28 ( .D(bl[1]), .B(GND_), .G(yp3_25[1]), .S(bl_out));
nch_25  M29 ( .D(bl[3]), .B(GND_), .G(yp3_b_25[3]), .S(vblinhi_rdo));
nch_25  M30 ( .D(bl[3]), .B(GND_), .G(yp3_25[3]), .S(bl_out));
nch_25  M31 ( .D(bl[2]), .B(GND_), .G(yp3_b_25[2]), .S(vblinhi_rde));
nch_25  M20 ( .D(bl[4]), .B(GND_), .G(yp3_b_25[4]), .S(vblinhi_rde));
nch_25  M19 ( .D(bl[5]), .B(GND_), .G(yp3_b_25[5]), .S(vblinhi_rdo));
nch_25  M21 ( .D(bl[5]), .B(GND_), .G(yp3_25[5]), .S(bl_out));
nch_25  M13 ( .D(bl[7]), .B(GND_), .G(yp3_b_25[7]), .S(vblinhi_rdo));
nch_25  M23 ( .D(bl[7]), .B(GND_), .G(yp3_25[7]), .S(bl_out));
nch_25  M18 ( .D(bl[6]), .B(GND_), .G(yp3_b_25[6]), .S(vblinhi_rde));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x64, View - schematic
// LAST TIME SAVED: Feb 26 14:34:16 2008
// NETLIST TIME: Nov 14 16:17:11 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_x64 ( bl, bl_out, vblinhi_pgm_25, vblinhi_rde,
     vblinhi_rdo, vdd_tieh, yp2, yp2_b_25, yp3_25, yp3_b_25 );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;


inout [63:0]  bl;

input [7:0]  yp2;
input [7:0]  yp2_b_25;
input [7:0]  yp3_25;
input [7:0]  yp3_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [7:0]  bl_med;



ml_ymux_yp2_8 Iml_ymux_yp2_x8 ( .bl(bl_med[7:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]), .bl_out(bl_out),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_0 ( .vdd_tieh(vdd_tieh), .bl(bl[7:0]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[0]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_2 ( .vdd_tieh(vdd_tieh), .bl(bl[23:16]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[2]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_3 ( .vdd_tieh(vdd_tieh), .bl(bl[31:24]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[3]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_6 ( .vdd_tieh(vdd_tieh), .bl(bl[55:48]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[6]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_7 ( .vdd_tieh(vdd_tieh), .bl(bl[63:56]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[7]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_5 ( .vdd_tieh(vdd_tieh), .bl(bl[47:40]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[5]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_4 ( .vdd_tieh(vdd_tieh), .bl(bl[39:32]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[4]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));
ml_ymux_yp3_x8 Iml_ymux_yp3_x8_1 ( .vdd_tieh(vdd_tieh), .bl(bl[15:8]),
     .yp3_b_25(yp3_b_25[7:0]), .yp3_25(yp3_25[7:0]),
     .bl_out(bl_med[1]), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .vblinhi_pgm_25(vblinhi_pgm_25));

endmodule
// Library - NVCM, Cell - ml_ymux_bls_x320, View - schematic
// LAST TIME SAVED: Jun 12 13:41:19 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_ymux_bls_x320 ( bl, bl_dummyl, bl_dummyr, bl_out,
     vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh,
     pgminhi_dmmy_b_25, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25, yp3_b_25
     );
inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25;

inout [1:0]  bl_dummyl;
inout [319:0]  bl;
inout [1:0]  bl_dummyr;

input [7:0]  yp3_b_25;
input [7:0]  yp3_25;
input [7:0]  yp2_b_25;
input [7:0]  yp2;
input [4:0]  yp1_b_25;
input [4:0]  yp1;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [0:4]  blx64_out;



ml_ymux_bls_dummy Iymux_bls_dummy_r ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyr[1:0]));
ml_ymux_bls_dummy Iymux_bls_dummy_l ( .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_dummyr(bl_dummyl[1:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_0 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[0]), .bl(bl[63:0]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_2 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[2]), .bl(bl[191:128]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_x64_4 ( .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]), .bl(bl[319:256]),
     .yp2(yp2[7:0]), .yp2_b_25(yp2_b_25[7:0]), .bl_out(blx64_out[4]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo));
ml_ymux_bls_x64 Iml_ymux_bls_x64_1 ( .yp2(yp2[7:0]),
     .bl_out(blx64_out[1]), .bl(bl[127:64]),
     .vblinhi_pgm_25(vblinhi_pgm_25), .vblinhi_rde(vblinhi_rde),
     .vblinhi_rdo(vblinhi_rdo), .yp2_b_25(yp2_b_25[7:0]),
     .vdd_tieh(vdd_tieh), .yp3_25(yp3_25[7:0]),
     .yp3_b_25(yp3_b_25[7:0]));
ml_ymux_bls_x64 Iml_ymux_bls_3 ( .yp2(yp2[7:0]), .bl_out(blx64_out[3]),
     .bl(bl[255:192]), .vblinhi_pgm_25(vblinhi_pgm_25),
     .vblinhi_rde(vblinhi_rde), .vblinhi_rdo(vblinhi_rdo),
     .yp2_b_25(yp2_b_25[7:0]), .vdd_tieh(vdd_tieh),
     .yp3_25(yp3_25[7:0]), .yp3_b_25(yp3_b_25[7:0]));
nch_hvt  M0 ( .D(blx64_out[2]), .B(GND_), .G(yp1[2]), .S(bl_out));
nch_hvt  M24 ( .D(blx64_out[0]), .B(GND_), .G(yp1[0]), .S(bl_out));
nch_hvt  M3 ( .D(blx64_out[4]), .B(GND_), .G(yp1[4]), .S(bl_out));
nch_hvt  M4 ( .D(blx64_out[3]), .B(GND_), .G(yp1[3]), .S(bl_out));
nch_hvt  M2 ( .D(blx64_out[1]), .B(GND_), .G(yp1[1]), .S(bl_out));
nch_25  M27 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[0]),
     .S(blx64_out[0]));
nch_25  M1 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[2]),
     .S(blx64_out[2]));
nch_25  M20 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[1]),
     .S(blx64_out[1]));
nch_25  M5 ( .D(vblinhi_rdo), .B(GND_), .G(yp1_b_25[4]),
     .S(blx64_out[4]));
nch_25  M6 ( .D(vblinhi_rde), .B(GND_), .G(yp1_b_25[3]),
     .S(blx64_out[3]));

endmodule
// Library - NVCM, Cell - ml_testdec_bgen, View - schematic
// LAST TIME SAVED: Jan 21 10:19:00 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_testdec_bgen ( dec_ok_25, dec_bias_25, dec_det_25,
     testdec_en_b_25, testdec_prec_b_25 );
output  dec_ok_25;

inout  dec_bias_25, dec_det_25;

input  testdec_en_b_25, testdec_prec_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



inv_25 I38 ( .IN(dec_det_25), .OUT(dec_ok_25), .P(vddp_), .Pb(vddp_),
     .G(gnd_), .Gb(gnd_));
pch_25  M23 ( .D(dec_det_25), .B(vddp_), .G(testdec_prec_b_25),
     .S(vddp_));
pch_25  M18_1_ ( .D(dec_bias_sup), .B(vddp_), .G(testdec_en_b_25),
     .S(vddp_));
pch_25  M18_0_ ( .D(dec_bias_sup), .B(vddp_), .G(testdec_en_b_25),
     .S(vddp_));
pch_25  M16 ( .D(net049), .B(vddp_), .G(testdec_en_b_25), .S(vddp_));
pch_25  M19 ( .D(ngate), .B(vddp_), .G(dec_bias_25), .S(net049));
pch_25  M8 ( .D(dec_bias_p), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
pch_25  M9_1_ ( .D(dec_det_25), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
pch_25  M9_0_ ( .D(dec_det_25), .B(vddp_), .G(dec_bias_p),
     .S(dec_bias_sup));
nch_25  M14 ( .D(ngate), .B(GND_), .G(dec_bias_25), .S(gnd_));
nch_25  M15 ( .D(ngate), .B(GND_), .G(testdec_en_b_25), .S(gnd_));
nch_25  M10 ( .D(dec_bias_sup), .B(GND_), .G(ngate), .S(dec_bias_25));
nch_25  M13 ( .D(dec_bias_25), .B(GND_), .G(testdec_en_b_25),
     .S(gnd_));
nch_25  M4 ( .D(dec_det_25), .B(GND_), .G(testdec_en_b_25), .S(gnd_));
nch_25  M17 ( .D(dec_bias_25), .B(GND_), .G(dec_bias_25), .S(gnd_));
nch_25  M20 ( .D(dec_bias_p), .B(GND_), .G(dec_bias_25), .S(gnd_));

endmodule
// Library - NVCM, Cell - ml_testdec_rows, View - schematic
// LAST TIME SAVED: Feb 26 14:35:11 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_testdec_rows ( dec_bias, dec_det_25, vddp_tieh, wp, wr );
inout  dec_bias, dec_det_25;

input  vddp_tieh, wp, wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M3 ( .D(dec_det_25), .B(GND_), .G(wr), .S(gnd_));
nch_25  M12 ( .D(net20), .B(gnd_), .G(vddp_tieh), .S(wp));
nch_25  M2 ( .D(dec_det_25), .B(GND_), .G(net20), .S(gnd_));
nch_25  M0 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(net20));
nch_25  M1 ( .D(gnd_), .B(GND_), .G(dec_bias), .S(wr));

endmodule
// Library - NVCM, Cell - ml_testdec_rowsx228, View - schematic
// LAST TIME SAVED: Feb 26 14:34:58 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_testdec_rowsx228 ( dec_det_even_25, dec_det_odd_25,
     dec_bias_25, dec_det_25, testdec_even_b_25, testdec_odd_b_25, wp,
     wr );
output  dec_det_even_25, dec_det_odd_25;

inout  dec_bias_25, dec_det_25;

input  testdec_even_b_25, testdec_odd_b_25;

input [227:0]  wr;
input [227:0]  wp;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



vddp_tiehigh I25 ( .vddp_tieh(vddp_tiel));
nor2_25 I24 ( .A(testdec_odd_b_25), .Y(dec_det_odd_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
nor2_25 I59 ( .A(testdec_even_b_25), .Y(dec_det_even_25), .Gb(gnd_),
     .G(gnd_), .Pb(vddp_), .P(vddp_), .B(dec_det_25));
ml_testdec_rows Itestdec_rows_227_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[227]), .wp(wp[227]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_226_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[226]), .wp(wp[226]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_225_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[225]), .wp(wp[225]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_224_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[224]), .wp(wp[224]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_223_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[223]), .wp(wp[223]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_222_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[222]), .wp(wp[222]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_221_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[221]), .wp(wp[221]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_220_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[220]), .wp(wp[220]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_219_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[219]), .wp(wp[219]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_218_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[218]), .wp(wp[218]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_217_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[217]), .wp(wp[217]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_216_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[216]), .wp(wp[216]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_215_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[215]), .wp(wp[215]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_214_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[214]), .wp(wp[214]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_213_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[213]), .wp(wp[213]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_212_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[212]), .wp(wp[212]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_211_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[211]), .wp(wp[211]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_210_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[210]), .wp(wp[210]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_209_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[209]), .wp(wp[209]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_208_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[208]), .wp(wp[208]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_207_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[207]), .wp(wp[207]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_206_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[206]), .wp(wp[206]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_205_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[205]), .wp(wp[205]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_204_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[204]), .wp(wp[204]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_203_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[203]), .wp(wp[203]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_202_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[202]), .wp(wp[202]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_201_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[201]), .wp(wp[201]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_200_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[200]), .wp(wp[200]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_199_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[199]), .wp(wp[199]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_198_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[198]), .wp(wp[198]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_197_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[197]), .wp(wp[197]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_196_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[196]), .wp(wp[196]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_195_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[195]), .wp(wp[195]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_194_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[194]), .wp(wp[194]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_193_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[193]), .wp(wp[193]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_192_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[192]), .wp(wp[192]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_191_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[191]), .wp(wp[191]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_190_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[190]), .wp(wp[190]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_189_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[189]), .wp(wp[189]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_188_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[188]), .wp(wp[188]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_187_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[187]), .wp(wp[187]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_186_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[186]), .wp(wp[186]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_185_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[185]), .wp(wp[185]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_184_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[184]), .wp(wp[184]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_183_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[183]), .wp(wp[183]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_182_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[182]), .wp(wp[182]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_181_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[181]), .wp(wp[181]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_180_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[180]), .wp(wp[180]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_179_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[179]), .wp(wp[179]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_178_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[178]), .wp(wp[178]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_177_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[177]), .wp(wp[177]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_176_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[176]), .wp(wp[176]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_175_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[175]), .wp(wp[175]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_174_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[174]), .wp(wp[174]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_173_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[173]), .wp(wp[173]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_172_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[172]), .wp(wp[172]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_171_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[171]), .wp(wp[171]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_170_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[170]), .wp(wp[170]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_169_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[169]), .wp(wp[169]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_168_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[168]), .wp(wp[168]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_167_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[167]), .wp(wp[167]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_166_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[166]), .wp(wp[166]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_165_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[165]), .wp(wp[165]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_164_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[164]), .wp(wp[164]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_163_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[163]), .wp(wp[163]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_162_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[162]), .wp(wp[162]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_161_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[161]), .wp(wp[161]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_160_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[160]), .wp(wp[160]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_159_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[159]), .wp(wp[159]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_158_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[158]), .wp(wp[158]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_157_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[157]), .wp(wp[157]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_156_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[156]), .wp(wp[156]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_155_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[155]), .wp(wp[155]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_154_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[154]), .wp(wp[154]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_153_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[153]), .wp(wp[153]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_152_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[152]), .wp(wp[152]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_151_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[151]), .wp(wp[151]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_150_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[150]), .wp(wp[150]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_149_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[149]), .wp(wp[149]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_148_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[148]), .wp(wp[148]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_147_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[147]), .wp(wp[147]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_146_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[146]), .wp(wp[146]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_145_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[145]), .wp(wp[145]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_144_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[144]), .wp(wp[144]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_143_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[143]), .wp(wp[143]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_142_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[142]), .wp(wp[142]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_141_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[141]), .wp(wp[141]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_140_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[140]), .wp(wp[140]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_139_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[139]), .wp(wp[139]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_138_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[138]), .wp(wp[138]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_137_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[137]), .wp(wp[137]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_136_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[136]), .wp(wp[136]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_135_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[135]), .wp(wp[135]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_134_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[134]), .wp(wp[134]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_133_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[133]), .wp(wp[133]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_132_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[132]), .wp(wp[132]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_131_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[131]), .wp(wp[131]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_130_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[130]), .wp(wp[130]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_129_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[129]), .wp(wp[129]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_128_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[128]), .wp(wp[128]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_127_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[127]), .wp(wp[127]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_126_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[126]), .wp(wp[126]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_125_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[125]), .wp(wp[125]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_124_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[124]), .wp(wp[124]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_123_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[123]), .wp(wp[123]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_122_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[122]), .wp(wp[122]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_121_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[121]), .wp(wp[121]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_120_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[120]), .wp(wp[120]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_119_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[119]), .wp(wp[119]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_118_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[118]), .wp(wp[118]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_117_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[117]), .wp(wp[117]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_116_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[116]), .wp(wp[116]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_115_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[115]), .wp(wp[115]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_114_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[114]), .wp(wp[114]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_113_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[113]), .wp(wp[113]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_112_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[112]), .wp(wp[112]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_111_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[111]), .wp(wp[111]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_110_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[110]), .wp(wp[110]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_109_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[109]), .wp(wp[109]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_108_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[108]), .wp(wp[108]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_107_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[107]), .wp(wp[107]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_106_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[106]), .wp(wp[106]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_105_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[105]), .wp(wp[105]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_104_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[104]), .wp(wp[104]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_103_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[103]), .wp(wp[103]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_102_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[102]), .wp(wp[102]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_101_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[101]), .wp(wp[101]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_100_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[100]), .wp(wp[100]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_99_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[99]), .wp(wp[99]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_98_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[98]), .wp(wp[98]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_97_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[97]), .wp(wp[97]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_96_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[96]), .wp(wp[96]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_95_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[95]), .wp(wp[95]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_94_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[94]), .wp(wp[94]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_93_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[93]), .wp(wp[93]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_92_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[92]), .wp(wp[92]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_91_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[91]), .wp(wp[91]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_90_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[90]), .wp(wp[90]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_89_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[89]), .wp(wp[89]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_88_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[88]), .wp(wp[88]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_87_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[87]), .wp(wp[87]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_86_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[86]), .wp(wp[86]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_85_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[85]), .wp(wp[85]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_84_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[84]), .wp(wp[84]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_83_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[83]), .wp(wp[83]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_82_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[82]), .wp(wp[82]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_81_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[81]), .wp(wp[81]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_80_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[80]), .wp(wp[80]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_79_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[79]), .wp(wp[79]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_78_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[78]), .wp(wp[78]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_77_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[77]), .wp(wp[77]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_76_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[76]), .wp(wp[76]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_75_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[75]), .wp(wp[75]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_74_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[74]), .wp(wp[74]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_73_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[73]), .wp(wp[73]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_72_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[72]), .wp(wp[72]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_71_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[71]), .wp(wp[71]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_70_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[70]), .wp(wp[70]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_69_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[69]), .wp(wp[69]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_68_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[68]), .wp(wp[68]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_67_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[67]), .wp(wp[67]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_66_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[66]), .wp(wp[66]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_65_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[65]), .wp(wp[65]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_64_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[64]), .wp(wp[64]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_63_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[63]), .wp(wp[63]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_62_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[62]), .wp(wp[62]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_61_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[61]), .wp(wp[61]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_60_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[60]), .wp(wp[60]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_59_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[59]), .wp(wp[59]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_58_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[58]), .wp(wp[58]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_57_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[57]), .wp(wp[57]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_56_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[56]), .wp(wp[56]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_55_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[55]), .wp(wp[55]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_54_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[54]), .wp(wp[54]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_53_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[53]), .wp(wp[53]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_52_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[52]), .wp(wp[52]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_51_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[51]), .wp(wp[51]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_50_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[50]), .wp(wp[50]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_49_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[49]), .wp(wp[49]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_48_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[48]), .wp(wp[48]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_47_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[47]), .wp(wp[47]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_46_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[46]), .wp(wp[46]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_45_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[45]), .wp(wp[45]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_44_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[44]), .wp(wp[44]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_43_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[43]), .wp(wp[43]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_42_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[42]), .wp(wp[42]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_41_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[41]), .wp(wp[41]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_40_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[40]), .wp(wp[40]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_39_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[39]), .wp(wp[39]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_38_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[38]), .wp(wp[38]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_37_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[37]), .wp(wp[37]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_36_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[36]), .wp(wp[36]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_35_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[35]), .wp(wp[35]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_34_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[34]), .wp(wp[34]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_33_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[33]), .wp(wp[33]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_32_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[32]), .wp(wp[32]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_31_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[31]), .wp(wp[31]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_30_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[30]), .wp(wp[30]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_29_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[29]), .wp(wp[29]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_28_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[28]), .wp(wp[28]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_27_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[27]), .wp(wp[27]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_26_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[26]), .wp(wp[26]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_25_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[25]), .wp(wp[25]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_24_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[24]), .wp(wp[24]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_23_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[23]), .wp(wp[23]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_22_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[22]), .wp(wp[22]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_21_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[21]), .wp(wp[21]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_20_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[20]), .wp(wp[20]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_19_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[19]), .wp(wp[19]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_18_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[18]), .wp(wp[18]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_17_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[17]), .wp(wp[17]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_16_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[16]), .wp(wp[16]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_15_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[15]), .wp(wp[15]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_14_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[14]), .wp(wp[14]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_13_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[13]), .wp(wp[13]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_12_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[12]), .wp(wp[12]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_11_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[11]), .wp(wp[11]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_10_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[10]), .wp(wp[10]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_9_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[9]), .wp(wp[9]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_8_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[8]), .wp(wp[8]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_7_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[7]), .wp(wp[7]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_6_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[6]), .wp(wp[6]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_5_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[5]), .wp(wp[5]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_4_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[4]), .wp(wp[4]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_3_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[3]), .wp(wp[3]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_2_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[2]), .wp(wp[2]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_1_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[1]), .wp(wp[1]),
     .dec_bias(dec_bias_25));
ml_testdec_rows Itestdec_rows_0_ ( .vddp_tieh(vddp_tiel),
     .dec_det_25(dec_det_25), .wr(wr[0]), .wp(wp[0]),
     .dec_bias(dec_bias_25));

endmodule
// Library - NVCM, Cell - ml_core_320x232, View - schematic
// LAST TIME SAVED: Jun 12 15:18:58 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module ml_core_320x232 ( dec_ok_25, bl_out, vblinhi_pgm_25,
     vblinhi_rde, vblinhi_rdo, vdd_tieh, pgminhi_dmmy_b_25,
     testdec_en_b_25, testdec_even_b_25, testdec_odd_b_25,
     testdec_prec_b_25, wp, wr, yp1, yp1_b_25, yp2, yp2_b_25, yp3_25,
     yp3_b_25 );
output  dec_ok_25;

inout  bl_out, vblinhi_pgm_25, vblinhi_rde, vblinhi_rdo, vdd_tieh;

input  pgminhi_dmmy_b_25, testdec_en_b_25, testdec_even_b_25,
     testdec_odd_b_25, testdec_prec_b_25;

input [7:0]  yp3_25;
input [7:0]  yp2_b_25;
input [227:0]  wr;
input [7:0]  yp2;
input [227:0]  wp;
input [4:0]  yp1;
input [7:0]  yp3_b_25;
input [4:0]  yp1_b_25;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;

// Buses in the design

wire  [319:0]  bl;

wire  [1:0]  bl_dummyl;

wire  [1:0]  bl_dummyr;



ml_testdec_columnsx320 Itestdec_columnsx320 ( .bl(bl[319:0]),
     .bl_dummyr(bl_dummyr[1:0]), .bl_dummyl(bl_dummyl[1:0]),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25));
nvcm_cell_320x232 Invcm_cell_320x232 ( .bl(bl[319:0]),
     .bl_dummyr(bl_dummyr[1:0]), .wr_dummyt({net84, net84}),
     .wr_dummyb({net84, net84}), .wr(wr[227:0]), .wp_dummyt({net84,
     net84}), .wp_dummyb({net84, net84}), .wp(wp[227:0]),
     .bl_dummyl(bl_dummyl[1:0]));
ml_ymux_bls_x320 Iml_ymux_bls_x320 ( .yp1(yp1[4:0]),
     .yp1_b_25(yp1_b_25[4:0]), .bl(bl[319:0]),
     .yp2_b_25(yp2_b_25[7:0]), .yp2(yp2[7:0]), .vdd_tieh(vdd_tieh),
     .pgminhi_dmmy_b_25(pgminhi_dmmy_b_25), .bl_dummyl(bl_dummyl[1:0]),
     .bl_dummyr(bl_dummyr[1:0]), .yp3_b_25(yp3_b_25[7:0]),
     .yp3_25(yp3_25[7:0]), .vblinhi_rdo(vblinhi_rdo),
     .vblinhi_rde(vblinhi_rde), .vblinhi_pgm_25(vblinhi_pgm_25),
     .bl_out(bl_out));
vdd_tielow I47 ( .gnd_tiel(net84));
ml_testdec_bgen Itestdec_bgen ( .dec_ok_25(dec_ok_25),
     .testdec_prec_b_25(testdec_prec_b_25),
     .testdec_en_b_25(testdec_en_b_25), .dec_det_25(dec_det_25),
     .dec_bias_25(dec_bias));
ml_testdec_rowsx228 Itestdec_rowsx228 ( .dec_bias_25(dec_bias),
     .dec_det_25(dec_det_25), .wr(wr[227:0]), .wp(wp[227:0]),
     .testdec_odd_b_25(testdec_odd_b_25),
     .testdec_even_b_25(testdec_even_b_25),
     .dec_det_odd_25(dec_det_odd_25),
     .dec_det_even_25(dec_det_even_25));

endmodule
// Library - NVCM, Cell - nvcm_cell_336x8_8f, View - schematic
// LAST TIME SAVED: Jun 26 10:51:34 2008
// NETLIST TIME: Nov 14 16:17:12 2008
`timescale 1ns / 1ns 

module nvcm_cell_336x8_8f ( bl, bl_dummyl, bl_dummyr, wp, wr );


inout [1:0]  bl_dummyr;
inout [337:0]  bl;
inout [1:0]  bl_dummyl;

input [7:0]  wp;
input [7:0]  wr;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nvcm_cell_2x8 Invcm_cell_2x8 ( .wp(wp[7:0]), .wr(wr[7:0]),
     .bl(bl_dummyl[1:0]));
nvcm_cell_2x8 Invcm_cell_2x8_r ( .bl(bl_dummyr[1:0]), .wr(wr[7:0]),
     .wp(wp[7:0]));
nvcm_cell_2x8 I17 ( .bl(bl[337:336]), .wr(wr[7:0]), .wp(wp[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_20_ ( .wp(wp[7:0]), .bl(bl[335:320]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_19_ ( .wp(wp[7:0]), .bl(bl[319:304]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_18_ ( .wp(wp[7:0]), .bl(bl[303:288]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_17_ ( .wp(wp[7:0]), .bl(bl[287:272]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_16_ ( .wp(wp[7:0]), .bl(bl[271:256]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_15_ ( .wp(wp[7:0]), .bl(bl[255:240]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_14_ ( .wp(wp[7:0]), .bl(bl[239:224]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_13_ ( .wp(wp[7:0]), .bl(bl[223:208]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_12_ ( .wp(wp[7:0]), .bl(bl[207:192]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_11_ ( .wp(wp[7:0]), .bl(bl[191:176]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_10_ ( .wp(wp[7:0]), .bl(bl[175:160]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_9_ ( .wp(wp[7:0]), .bl(bl[159:144]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_8_ ( .wp(wp[7:0]), .bl(bl[143:128]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_7_ ( .wp(wp[7:0]), .bl(bl[127:112]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_6_ ( .wp(wp[7:0]), .bl(bl[111:96]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_5_ ( .wp(wp[7:0]), .bl(bl[95:80]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_4_ ( .wp(wp[7:0]), .bl(bl[79:64]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_3_ ( .wp(wp[7:0]), .bl(bl[63:48]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_2_ ( .wp(wp[7:0]), .bl(bl[47:32]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_1_ ( .wp(wp[7:0]), .bl(bl[31:16]),
     .wr(wr[7:0]));
nvcm_cell_16x8 Invcm_cell_16x8_0_ ( .wp(wp[7:0]), .bl(bl[15:0]),
     .wr(wr[7:0]));

endmodule
// Library - misc, Cell - vpp_clamp_finger, View - schematic
// LAST TIME SAVED: Jul 30 12:32:02 2007
// NETLIST TIME: Nov 14 16:17:10 2008
`timescale 1ns / 1ns 

module vpp_clamp_finger ( VDDIO, VPP, VSS );
input  VDDIO, VPP, VSS;
supply0 gnd_;
//wire vddp_ = test.cds_globalsInst.vddp_;
supply1 vdd_;
supply0 GND_;
supply1 VDD_;



nch_25  M0 ( .B(VSS), .D(net12), .G(VSS), .S(VSS));
nch_25  m1 ( .B(VSS), .D(VPP), .G(VDDIO), .S(net12));

endmodule
